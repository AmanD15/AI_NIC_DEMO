-- VHDL global package produced by vc2vhdl from virtual circuit (vc) description 
library ieee;
use ieee.std_logic_1164.all;
package rx_concat_global_package is -- 
  constant Eight : std_logic_vector(31 downto 0) := "00000000000000000000000000001000";
  -- 
end package rx_concat_global_package;

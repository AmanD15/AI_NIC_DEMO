

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
UTmxs0OkmJURXBOVdUGR7t0vPgcBU0oVnrXWTlGh9ogLy+aZVadnSNImcgn+4jLE3/0AXAxZXQ82
Xbw5u5ikwg==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
NDHq9z13OnSHCjB5ixLI6v+O9siiJNJuJRP5KO7VWFUgsdEdfLm2msHdSHMZWHSOwKZ3fpyDnmNx
BgNrMCYycBeI/rO2pKL2N4HQAMnhKOZtiPFF9n2RUplezsx3A1KtfrZPlHnD/UnZMT1dsl6klarx
WHWoOj2BdFWF78jqP/k=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
pd1c/MzUc/ohRsjBZ9c2FYMEVEx0/T+c02CO5nj1hjCkjBTD1iExW4b2fGAqq2hXvApptvjN3kao
diEYImrFYF0oK+4fJDQ0NDCFSHEPkV9IuYgpAy5fNfC1Dx9rVAZAI1tVIUXAIZsy7oaGc/ReA3s3
/Ev1+YSM6X62ouq0EXc=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
Ds2lszdMaBUWm49P9ovDqEJCNyznNiiJV1s10TsqQV85Goa2s6Y0q2oK0nkUurPC2r1U/lFQ6UkY
FyQj83Ie6eOpnawKkK55JF60SUgc/KJzJ7bDwIpaZjrpb+XlrqrzZU73J8jBBHKLoF1/Njgvn5Ad
h9N2MGH8gaas+uT9uDuZCA+ii46LQ3K2yd1YWXKK4uzoENDnOnWVcV9omYQiZt2WoMmuDtnHiiD6
BU9fNvTDJc2E+yqoRZLq/i7Vp6O2raEB1EabQzrK+1rVqoRBidd5D+df98jf+SVXW4uK81yOCvMA
LOV3/ZU0qCRQoJbwjKLC39h49ly0sWjEpfW/gQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
df0vCAvcFSWs5BffbtXlfaFIBd83+wey54D1uX3YAx267SlsUp8LU636/ulbSzkGShRGyHAsajTQ
lak4/g7ql/uNS4cPDTprvz1MsadnxOACDABIUOl7lg4w0zjMlnHliJydcn6lPMrRHgqJ6QJh1Ypj
8in4rFzqjprqSxw1d/10YsZZxkQoba/tmtftne+6yGg56W2Fvkku/OTLhJ4+2k81Et3P6Hl8rQs8
H3zDC5jgcWutFMz9ATChQpuoW1Bt6ol0u96wp5xiZl1ORv7DkneMNq66FiXR7uQAikRnfSIiT6/5
QAjuFDJ9beaONJ/7PX0YKv+VUGzRFq0ZFYEUEQ==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
nCZ8D9A90hmHjnYoY13nJu1ipj+rg1ZVc4+qcqLwK/I4sVkFzYXzOHfQZXQ7YKW8qcQwr7Ja8l+y
rmS/aej2Bl+/GBm2e8OPwXjYQfJZAcWrX3bukYUhs960X48k+oy8IM2fpLqIO5UjCHWUKDAmMH8s
veeZjDOkDvXS6zx4x9hZL9OB3MW0oK6L//tk4UtxPcVZEJmBR7mpHfQdetJlD12R2NEAOMEs9GYi
egJoRgy2DcxVo/qhMUxikMoNK8DRbPimHxnf/gi8Ss6Awc1pw8Haokg7dho4WvcGQs5jULvRh435
wbmLZ1FnvnxhHSbLJwY8aBTSiBsD5Jozey23DQ==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 504800)
`protect data_block
wS8+RLVd5I9wiDK+x+m/kUkD1kGFYV6Hbblpan1Ad9SkG4DzJ7262WD54UZiZ+sa1geIGLzL+w+G
BmepywO9W6XMyQ6Kdx9850d6HyryDUle0eePimUKi7MAUZa1YN41g1fXPIZgwAzGz54PYUETIt7o
IrPtcxmftMhw08u9SABRZ/aFSh2zSj7Tw7DOIjiZH9ZJJZHTIM7Geesyn8FpNE35Nl1p5cO6ITaw
/uq9SrTwwdxkW8L9fM8NmG9gEFwaVoMgTk5r1m4pTVqE0w038XvGTN8dtRrEnoUwZ+3PJTL3efKr
NPmQO4gmGYeLCHA8yKKu8r/YNKOJ7MnP25rGROCgwXSb20OvapzwPqHx5xnZV8cI8z9ETRmyw8KS
6CwpefxTY/LhTSXRdFhm/T0N0EAmK9M0ctCGzR+k+3/ewcFiO6RuKXv3uJEQYMVz7uNdfjploUww
WW3Zdyo4iyxFS17XmAYfsJMKsiT4CkaqOX145ZDcMd+7mAFJ+uGbDWHXkWk1h2beOfUrGEryLM7X
K1TxqcoSXnx6z7Lch2EPsAnXwtKAzJE5nKlXQOMc4cUm4ogDfm6gz2HpQis+KuLlVyC38RoLUAIC
K9C7614vW7wIdu2BxL4rLfT8d5DVzaut36DTOY6KLJI/Dx4psH9TxFa5AhdRVvDdHnCIgBs7429M
23dnko1JM9ZVNr6YlRzCYkPSQuE7oHxxLesZKO32wDxUbYFiI++4G91OZ8sFrSWsHQ+TPt2jEvcY
5AfDqDQwqEcEPv11VMe2Y/yud5PM1fbQRAwgR4uGJi10nE04fOuXCk6way5f6HN29chKgWtqT9Mc
BzJTjWbxBguhQmi0ZbNM/4G+bskk1aZDDLhRPKDWBLfdYBR/QRjvQ+3DZCKKjp5LYgfL5xloGobv
MPmn8c5d2BBXg23lK/zaZ8igvr/rgCKGM1pDklLJUcE+rH8gPzYSDML0w8gIJ7MvhO+zOs3JSjc5
HbWcemPbj4UJPRC81MLYf/svD/x6ybiIdCs2xX91fxcGGayjFHvHXGWF/LT8gMVn5nFm5cDNgWQS
oiQSY/aMBQ4w2PqqJzjH5l+0gZQKvGbukUcoXnkigP06SsfANOCQSEY3+K64Op+gLoQK2yPjM0Y1
FKmGRy+m0gOO/+4r3EGiQ/WqQQXQLzxi9YmE6lKp/NHx/tWf/Gg57PhEDS4ToiZtFG58+t1+7uEg
fPSL/p54sMN81icAE2d/aXoZt7lB6zzL7YucVxKpHpNLHwxiXxJVYkOpJ39GvkY08O8fQGUqbSmK
N7GkTuxrg1BnwW7PO+zXx8PPYKx9qEMl07sIec2jreiJJAuXQ4ZI47INDAyM7mfDJA6bETJei69a
AGHwT2nDXiT2PFvdjCKMCfhpv9wA5bEdaE5bRMaZkLl5NgtV3emjRFAg2ev54DbGW3kAlTpNDdMh
q76ayD65TACgmtm/MFnt/Sa8KgTUTQsRgjYuBgLB6DojdZrd196jU7UVNBCQqkBKQPqRN7E/X1Lp
Xv5vqAqhmuYj1A6lAHLoq8gcYqcjZxKXZhkuTy3OvzNFSvzXOUdVYZL1M1jn7kGRiC/hfre2u5Do
LeWiPWsz9xeQCihBFSF8bhbODKnitBok28DjgJOBuOZG11TZ0Ns208s2I/YBOVg8osL1Q7Sphrfl
XPPMz3gz43Th8y4OHmxLVC70VmLCBbOZix2J1IbQigdIIq+3yvEW7oILIRk7+4J5itJ2ipkR0zHB
vHUPWI8+6EXHfY0hxsMYBu/Uge0pE8d4SCQ7bWy+zkNEvo5ZC/thHunmox5RIhYN3pbPD3G0n1sK
6/xyvc/tnnGpG+XsVbMEVxYKElaYODvbPJkoEhcUKa3RWLK8nj8iLC+UHrwJ73Yq1bpYTg2zDR3j
fnS+POIEpwlZbZtPPmB2AUZ2t/x54VP6PwRnx1IP9NfZIt9W14hdUK1jPgvNxkpYCcFYxYT0uFej
FXBlzur0YpQJTD7sFrsJI2h+AzzrLwl3igu/W4nf3cZdAYDJEeRJ8ipmRo5qE6xZY5tY50kneeVB
gPBgmy5EP7GoTIWRIn8sIuab9QpVbWfaLXzrBrTFBbV2EozBP7tke/aeIhBKbHq7yKDz4IiXeSkZ
vI9+b5Fndi7+Tled01PWFi/X1PAAea3bkJcJnD7W1IEPm2ItFad+s4ZS0F7uH53873w0jbhS75xU
0iVqsOh0WnRiRhNT5OzyV4/pnbMhiO2/s45Vm1GC7MC2fLkMiabllZAH727tFV/T02CBGFmWF2d/
06uIs4wuGnO0r00K8cFcEDtnqx1Yj2Is6GEe40n5Srv6B1OlPul+3yYq4VYofrmN6HFfCeyY+g7+
RtIK36Zu4D+wj++JJHEhPiA97cBeeiT7slUsYrg4CEnXs4jlvIgwCx8eGxi2spZQr/oT7HSa0qj2
3YASpA5x+VMDzryycezZLeSm+5Enx2zmR6azjuCzouTQRofVUcKeGbZzBpIDq7JLXJW6M/WiZ96G
Tk1hJy2E89+6ZUxKZafVMeQuU4FtKtReKsOvchWDd8k/hvf1DHZQ/bTCZdwBvO3zKP5WE3BDi/Ym
U16p/TS3G7M+2TtnbNgmv/HpqVmGVLquGR4xo7wzgF+KobG2Uy5InlCpUxGmQY2TgDuingHEv2P/
tw1IFK6Swwtuk3cbzRtizcCS43uTxJxhVSOc1STEi1thL/r7VaZPuF6ebpryCXPJoIl3O/quTEbU
BNn3YZpSzEdxiU83m0gBSdhZnq/Ter5N0ykGroeXl03EoSwhJhY1Y3uSg9efgqGBw3JR7lXiKvei
IoAA42mn3DKZsDmzs9BSxLFcF1ZZNgJys2ortkmpcAoGQO8Bb03Ya6dEDY4JmEHX51p8d5x/zpL8
UUYJxTnbBWIWW6ZFAM/9Y8N1FWJmIWUIDd8gJVgaVmaezp+NvgVKsqGFvjdHygofRhnatNW17Qrr
sbGNHV6mLeXZ+WSf7dKDs6SQjgPWhbTYipVPHgqnPg4SOCD2f99+d8WYEaceu23omenaJY8qTDtT
3rRYOR7cqsngxjQ5NGsTv+4x/8qVPbXtWAHL8aj67LGqqu4cDZTZGXqWWzWFE9eAUtNBli9kDGOL
zoP2Id4YRBGRGnWCmVb0ddCHAecyIbGlnspcFE9PJoeZLOv4rybg2ONhamARWF4D33YJtTlXvdHr
m08m/PFUmQzf1N35Br7W/iX8ubz/VtXsO0zhTGHtgNQLdqvk4vIA/96jX7+M16JqmcoY2FjXu+bH
67ynPs/fmiTec23Z+ICHCHPJQIaXxh38QMNAW5S8LGblAHkX9uklAgBBeKV6DQT9J2et+7BKw28D
zxuLxmTc7fWbZXwMU41YopN6Bj6sAT1Dz6I+yaSF9kXo2ohGAZrFljrDcZ4WxTrF91hL0phm7i/9
EthPYz0giPOB2AyzvP5Nahrr+06XlEMEebebLaxSC7a6qj2eVFXpaUgepo+01hQ8je2qbfHGEQXK
SfOQ3hTi2pammxMj388VlukQ71p/xb/Jzw2IX8hRXdEUaqQuEqtbJ3aeX/el68A6IKUWv7G6E5jC
EZ54TlJmdfiS7ovidwMK3fFXH9p78bQCFWTg17huvDx8AaH6mNFurujUZo/XKngcJ5+pwV8QDlr1
z5s7LymZ5aF3Vo9Z/TGDpEzZ4vJfXVpa8ZSCTLWBoQPA9w0m4XhMwYgjBBHd4WD9QyIyutPnunrQ
PgnI+c8ASwG1Y05HHV+e8AUtMY2AfSZC1lMsJF1Xuo2+81TH9YVcKMlr+y+ygsb2zsP+pgNMMMBf
UnkZZv/q+vpjQv1wfrENw+uVLI3gZRz0s5czbz0onOmGlmj6af9bGhoGmNXe0Szu9UrppQucWJor
0+DKn+LRMJ7C2DJ4j+MRF8MLPw107yyvtxOC2n41NESZzJ8aGzmUj1WqmKFB0zRt34Z9Jgb5bq8y
ha7AEAFiVSqlqYIIZcZpm1wEOCmoxnViuut5hu1v5bDX4naoc9J/KBblNxpRi5uYDkHzmUJeXePn
JVS1V5N+XCvASVfaDC+Qqqs0xm+E62ja0RZX32dsSgQhkUbluvgpWUkONwCtoJhRi2foyz+xGMSO
KP8rayQNEwGWp5heWfYok/L7CdYBCLQwOYqzMhCQQBzDRp9gTiFl5ovfusOa0tYoYAAPsesG6rnB
2NqmNrGqNcruMPX+j7xkwZmQQJG3/DXOuZtduVzo+vrDWmGX4nxdeC07fJmXwA11E+6mhY4H1IdC
lNtolPYifv2nKzUmhykWSBDnPV4/MD3SSKXSK5ovQms9Fs4Adlz5MaYwSe7SmscUeSr+NJSaVCsc
ja7ts5W9Xtys3iYoyID8bvDbaMycprPkxr8MwgY8AfKVNi6D15Pz1krYBa7f3EmtIJmt6rV7wYQ9
OjPU+7NzEeQLQ5YnsDVIPKVBf0zsftYZ9sRXySnG6xQpfLBakk5wbmarDUIUUhzW8TatBF0JZ7Yq
I+oRGehtv1OWXXemtUDuBi9rqpAt+Yxicvk0wRClBLWqJngQ2/WokiCZlVMGhx+7sIn4meJDj3ZQ
CaJQjpupHESpy6lScCvvVYPTPSg+XH99hee4zzD84na3Kg+j3FZa6zYwVza3Zs2jLHBjpLG2Lsv8
x4ggYVcqxE45y9L0VhTIcOo5Ky/k2kfLr1Kmo1QqogdDKh7QvmBGEFQncw6IjU/VPuhsmqBxvGzs
8gk0qAaqefKzif4MQT7i+sSriYwPqhD2PlxBcjNL0yroCybROlH51i937s+PXo34zcgpV5gkhuK6
uT0XPvrTJI9EpuR2NzjkkFIF9T5DLnOOJfUWPPZHzsHvacBwnCqffqRSsg+XZzxrTxPsjR3pB8vB
diIZCFG+2p6lwq7Y1g8UE9hYcXCofky99QSs3szVuFw19XGXh9PT1ASuk9JfS1UA9tUty/9BOVo3
3tnUFM3JH1FPkcFr0MKQQGFZ4OY0KH4doQ3jezGFARg5KaCsm0z5lW1wQqk/YnnsHKZRpNubGbRY
UTWq01EVcL2x4OtAzeBGB9nVKClx5HOPEPJK/3qAe6kvh6mimCrIBd/A7bswFvJf26T6dSuBgiK2
s2acnItxUS9iFAnascT8xJGkWnmJL95WBiT5ft7mLDbUOW7cd6pIHZquU3tYRHWGwSOeexho0fNa
d7A+hyih5kzT/VZDZREKff0duDB1lQOjwsK6xSoZ+ZC9Qc8AhV6Kfy2flduILzOHoiXsBijUk6bC
hy1Q8s6Ol6LHJtFgLDcJNQgJfJwP/rgMGVE2M3uH++PjxGUvOHObFhPlh0mjtUcYmNyUme+rtMAe
wNwMmCXvaqfaVD5hiopm/wR3r2JpX87X6G7L+OyzvcMXz8vRCkDwRtKESGCMzauYnXFgXTmSOpxX
uESJ2VTdLC0d7da05drcrAcWTKTo1AUkMv5AkPdb5SMG1bmjoxkT9DmyeGFOOh0M/N2zpgAMLKcP
4r8xgvP/c327FRGd31DwK5oZGtFonra5LDrudHsUlyPlKiY+Yel1CicU6Bg7+Z/ReDQm7iClppQo
V8stJ5f4jDjBeLXUE3vx5Uws9KD144p/gnvon0+/eIiMDI6vwNzThQ5++xf/8SJlof7zESna/tXi
ijXKDsq7/NX3aAtYQByJISZeuKJcE0imyi1FfkfUIo5pE3rUTC0lOheXkpl5Gj5756lUypn9pNfR
P3HfbCZsdnU6/scW9FS8K7qQI7kPzCeTb6F3RHtcHlSbeYxb7xtxHFWqsGJSUCptjzMiOWg9VRBa
c7/tMxvMow5VRIGxCy3eCtYwOcAPUE8chCIt7o+TUm4pK8Gy4NgFq8hQhi5UK24SkAR1GCk0GkzR
g1fzMKCkWYvyJN40m478bkcGKnTltOJ5KuhIebSIROzuwKuHkiNj1scaRtWIGh7JQNqVzeMvkh/i
po/54pI64kaQajBX5It+Lu9qMWjkImxdadNSEWFRo5s7aJpIHBaUVoO+pjfOmm42vz1KltJKTb7/
oUh55bZFBjX8vGunUxSZpALEp5C89FpYWgoSXyo/Szyk/FmFBTKwt/GTGN/iRMfh+rIoGyBu3NMQ
teckDGKS2jZxXT6fwPZO2COhaNoqUPUBemQZP+Ss0MfY6qxeZ9QBeyaCkmAjF+1rQ4MlHUPzTkSM
+/ilouRFCquBBJhrm4Q0SSIsE8F82c6i1GsVVUw+sdtzlHbjwP4yd+Lzs02gk6som1NDiIKhLUnm
kuQcTN4+5xPXXTH7smMSIxls0Pi5SFcZLZCWx0qR7bATUY9NhPgPJ0oXkcAQTJG9pCcuNiEHE+F6
Eq8ZYDX3L7Rs5x7RUBZhqcKRyxiEssqwe0Kim227YfNmQ22L/yyjlB/p7yfX2Mw/72kfhRW5dk9y
mHXQvoZ+en5+ocamo5IDWZICBxZDBJwpIerimfacDZ79KOvmJC1IfkphWrbkCcaaQCpsluzq42dR
ZwdqsBEGJkJpbLGrFpCJe3MpY2JHfVIrWGDl1Y5viFJaxgbeIqdPluQf9texg0q58Yw3T/qt5FvC
K50kuMq+MF8sgqB6P3CGIPWyfoaUXqfC0U7Nk8WUDTlZFB4UK8u2m1JgvCMbxG7BV34b5O5WrdrY
CeZYjGtzqHdXjUZ47xykY+DMFCWiWrqDr26VRDjPrfZ1LQCfjPIOVKDXhDNTUxDwXDYW03C4TsAP
aQQmVI0tkIFqVvMYb+Y2leuesdDjFKOaYjw1cHEwmledlhaKbggSpceykX0VvGUYC9h2pfuk7fd9
bjGcV+dyuiOjk8NLwziPzaRSuTMkywk1+7gyLZdbDe6go7rND6q4dLLq9qBhl3j/2Izgk9UdGYWr
o0B7RX6RDJp1YU2RxBq4Nu3gXvta2L9KT1KWKqKvwgYX4HtocbKbYW2NYeiJVy6hqqEMheeHA20U
Ul16u/xP7sz9ne/IPSzGeDEllcJt7zMlmxsocOh53UOvK+7NR9waMGGiD6lbOpYchRadAswPKsjK
QlsuqA/OnjAEMboE6v/cE8W0TO/uUtEr/NgfdQy2mHS/dY+VkLzzd2+n1xsJnhcvaOyrwEgVi2Nr
vxHo/FhMnJZ2k7+MI0F2K92O73JOZgicIwzFelvWywfURmxgmxv0/ySp6rlUAx5bLODTjDDvL9me
fpaYXbpfz5/PRdnhJx6iwf16BK9kF+OSsGXkxiQPlb00A9I0ZbE375il2BsbMA1yRBoTjnPji30f
CBDWCo6PFSSnUyM2XGXu7DoYOQu1ClItfRMZMgvTtbv53Qosvg2SNQRYRfty+rFoXwlpV0yYudSm
MqOY/m9dpKMog3COJpC4DOPxu+UQTN1xyx9EwS8jB3tbmlrA2jby+Sl8Ylre0K6maItIFwgOI/Xm
hspNV94faR1jXd33XnPwu/bq00qoi/x/ZZbmLpQRD3WAs+ORf0eJWt4y+dL2dK76bDrXVTRuftJA
j9D7fzTftzZiAb7ml54Yhe1EYu1KanLcSfFPix/U06Z/UWehQVZKGUMHiOLB0jdFkZPWeUAIf8OZ
2qRvS7lfjiU62rZHXGUyyqPp2J72EcSfRdm97W8Bo8m1bVwfghdhZr2dSxEpPfOwni3t4UQvClK+
ZfthjFSyHxmH3ipQ4Ajy1cSp+hQ4hFAfOTMeUiQHBf2VECZEZHEO5mAvBvLI+cvSCypk4+LRjxaD
hfzriXxI6tTeO6zVNXc/GxdxjFw6CxqGrnbzMjxHLOEcn8eBXqIhprkJXVvHm5duSzdC2Gs16irn
FUBh6x+vKmsrEcc5wOxW1A8+hMkeYQEFhg788eDngM7xAnsKUYgsg6tlv995sQV8mrbeHrLAc3FF
Br9GOwkNSutbDXdbSqWdVsXzdAX+kmHbIZwUV02wqPzCnh5VjEh9HSR4UFAiJwbiC124K/523krC
ChuRA3UdHZhpSFRV0u6EPbl3G10kSaiwe8EuWRkG0k94/Ka+wcFd0BloNQ3ZJQmaVT7R/uGXfnuw
lj7Y2rPdGjCOzCJwSHs6OOHmtwcZj6XkNHiWudN6Hj81fNeCrF1VbQHfM5zmoF1JAGOtoh063CWn
f/iKlKyDeHuB9n8FqtNdgaTlCN9g1YZMMY9BLLrqHVLebh3rIlN4zkCMgOXFdwy7QSvwEpwwyLfR
Ikd1fMFEDFIuT4rSmXal+40Qct1gS1ZpxJIl+GxDvhlBo6vz54nIUhetzua9SzwTxfy43yhrTNud
F91vMvqLZOLvKSz622yLDmX6NL7togr2AP0+YFmDV/05aZJaSPcA8556pakS99KZEDhFNw7BiNWP
A/eHKYKBZ0U1jpm0/BimtadIJrBgLOkP28FmnrWEUyauscCgLxgGOmBC8TpGJZexUZtHTLqvrG/8
OTJ++ZqOGPsiySvpiXUaFfMyLl1yVGpHGE4u1nZ0L7x6jpPYi+xQP+J8R5b7X3z7F8n2fZb4+u89
2Iuna3jE/jzKhd47+kjmA4p9LnuhpBiq8/UGa7JAuaKOVSyhVvTHzJvx/6BrpIfX8zL+ohijC/w6
t1eVgsAreqAtpetTdnGw47aKI59upVbpzfugo3b9b34l3XKSui0ST2W2CJIDcOWBnG+zOmxJ5aMn
Ggz6nbDPzFh4DC7a2/fgS/vX8UplF0XdINnkY+FQDiVt2G6ZneevvaFOPtaiJF/1WilcxYIoCQLU
X5vICA558rHLZRFcwMM65MVBg1nbPheudCbhA7XC5lfq3UtJUkG3NO8OUHoxi3THAQH65c/0iqrd
4hXCLEJZ5fEncEYub6w/2xJji4dOe29KpXTtGz0KiyL0pAXzOI/XZ45YjO3txhWa0FrTQsYF7aR9
L0DwfQ34fXqWl5TOMSseAncN8aBKm1Ik0k66Cphk5ZuV8TNMTFbHCBLLLw7IHbUOcNberNcUTkYH
DW7R7xFLjPSeHnlc81xQUKm1LKxSPth/CfB5cpFzn6pH4lCq9t3x+BE7zepaE1+N2xGq6d54+Zgx
Agfj7a46TspzS05oXXNL/P9p/QVasQarePvF4dP1fMPti+obky0Gve+Wf/ofs3XYOCTMsy74CH2p
/lNofVUv6zKmG+Nt19PT4D2YwDTE3xVqgBspQgjOK/EHuXUh2XHaz0lx+LROBPeFg38ZLwICoyo6
f/cyE/lTH43UNngZDAQmObCwRWLzZwY95UjVQL23zLHdUlMTJ5nw1aiz6Dr2hlY8XPgL18h+UngF
ZrRmgQzRlXADWoh12H350foGuMZk+h+stTzrpVVZ8hfoFPL/qtXPc7fljBNhce143h+p+FVmflZn
OgAxLMlm8dbJUvISWPRVux4rVHd6u/JdTuKMweLQ4mto/GbjazoW4xXNHyuJZ+PAHFOQQMcRYOsi
fyo5RvYwgDB9bdo52T0049ZL6UYizDv0nYXdhkJZOjQANseid7qukHSVgAUxF3Z7dlOg7HQvG419
LjsLDH7I7Bmwca8Kl13VxE4flIgOf2qjBzKz5k0EbSFtMxZaBzc/aHNAJPObPmBk3WWfUH44CrEZ
a/3DQ+tY3tHRE95YUsYJWYf5Rz+xDQVkkSKrIl5ZDP+SbCAXfpOEojgEkeY7nXSjmIsgMDghUiP8
8nDyJc81hrksQRWImNfPJktVZXgbpA9Z6L6bY5yj1HvYEU+prpu9WJX7qVVocLepjpvERoFvHZqk
fIuk78jMm+tZSOfV/Hl71bP8INtU5QnrY3RNPxeqjoMS5qIkvwLmJ3TgTvDRVdHCVRS4g5+NA4v3
h/UT+AbK+z0EaJsw+ICZFhb+4/ewva+I7HVfWdFrUMSPswS+JQL+r5Fi1+iiVUKg0XuChO1dDHKR
F+/cacJUs4lVV+hnWfKuRDu66PDOsPpf/vj6AUtPJd/BmaWDoB4V2Y4x5p9/ACFZ6rJxG70yTsZK
nBEPdlmhY0R+X+kLRVlxpFmlc68D3c72LQEvlZcn55A2WrvnlJSYeaouUzGlyFkyLTRxZwLRccZ1
qk1tXPMxirYBt7O56GDtRndnSrdQnLKlFtRzJSLPyhs8cbykP64SlRaPPqMeoE/uFqe2fE1BVpiR
xcvMis0sfinw88161nWfnyfBsB6u1WxlYG0O+lSv7muYmIjT+tSKyruUtnYwNANI3Oy66M+2WNOy
UqVD1EyTcUDojusdL9yC/6ZzrVA5K4FCs2yd/C/a7p+9X0f8Ix89x8oeUIdR3flvGKjmVtM/bhzx
YGailbbPVeJPC5tgVDeD71geYbWIHXTP6bsLDu5BGnEd9cbrYs+JEo2+ExjmzClBzSG2DVeMa3ZE
Hyg1/0eZr+1feKfB/KWnSF4UpzRJ78xxmIjAlDCm2F2sc25PMdpgK1DyV17IdBjdN6ZDWEJXesjs
PwFYNS0dCV5vlV3Sr9EXf93jttAE66VIP6FvdJ974U1hmMF7muJxomfb83TnvoqrLTKjqb60rS0C
Wudb16DlkiMfoNujqhf3dLDLboi6QKtU0e2kpxmAY3MK8yhVwPLRj6v6cOdpQ9DLIgpbI0uaKS6z
ekgdwraCBGDSgOyQgn029KiV/GWDd1BnhmlKxfS5fUSysKj681ZZtZO3fimsVHvqQo44WPuh8Uc7
ZnQalLG4D4y6shTXsbSBiOrBEx0obb0gOZB7H7EIqW6UXfchvg+HtCSnR8wWk9t+ABnZsDRaZBzQ
gXcNHlWeJNu0RJT/teeI7Alzc3CQQnrrUyGWg10XAnk4kJNfr1K7p3WlgKvmqALARqMbWwuulDHi
FqH3+8aD4Hf1jwwfo2a1ieRV6FEzbwWa4PdoGFuQPWW1sSo8gRHZ/7+XQnfVMpDKB2NN67DNzCZ/
UT0PDKCgbw86/7bXa8HB7TpOvvB+0VDPkNTeJ+1ng2h3zU6IzQiPWZSMoHpqE6N3NUfUJLufx0U9
t5KrdiImovZTSnOdpYHDL30mtrZ8LFKcH9ykBcHJhUj019464eVIlfsvgX7E0+hizaJRMpgFc0cB
d7EurwF7zYZW1A24mvHpRKZX6V4J3cyvHcwmJONSE1Sb3nylnow5aYQJ2KGOvafYnfyWhUYPByH+
t4FN/ocZJ8rGZ6vV637aXcrV35p0ZBo+N0HqZpSf0l0AuAc6LmQslpxXjea3rW4o8fr8Oh/cMf7Q
hTpudGm82DJUdwvveLAj5fA1qBQO1ECW0IhpkKdbP6XeqAlms30D3Q861faDewicx7shJiOcFvfq
bYgpygvHShENMTiPbx6JTFlRQ3XW4xfehBlxI70KIow21ymIbBeOngVJ8SG8Okmmiyitdu8cIEpr
7vPd2zUqDBwwM2RxgT4e46r6cIAxjzIn7jLh+XCr3qk3TrBQfuGbw/ZuLg4oRo6+gNLoD0KN2PCo
CDMgckmIg/O7cMDJgOwdJHUgNpXWMbDKHKD4vJVQUGQzZpHDKPQMKo/uhDhYXLUSb+aMqVB6YTJJ
kNbbOq3ulMRcqe7qBmVgE4kfawWuK8nrurSgvN5D1ARXn8kvD/xsUPPSScURt0BJZJjVDJxkCQf2
yz2K/hDa0cDbUwMUkwCusls0eE3RjYJA5e25PIBsVlKP6cPB9AUtErjYwPoD8pAX4lnO4ib8cee/
w1z1ny/IPhlWKLc2tKvmxKzhuvVGIBl7b3AoBne79+KTbCUoo7+vK2CAf1RYXU7dc+ZClbL4nL+6
gW6fxxB4HGF2AwmANuDO2fZk+P7FIZtB4qKYW0SJWv+ggbsp1SfMsNMeIIxph29FqVzB2UHkmaPk
HtVwv6RS7EgTqXq7FONcnFToDB1B+GDYboaR2SfHi8GWYgOrHtcLc5SPqmNJmPrirV7R7Mwr/R0q
15OqqL0XL6Jn3UMPLTAWNOXkRDW5kBAVgqORYBuEQBu1SmGIy+TbHo2XkZsMDbUzt4Tf7KDxE0Vl
qmh2tk5QXbMVuSx/4HgiDezNyFbQF8Dya+Ush45LxUn+R4+75fM8LPluSxUuqrd3mv+PokjJu+VY
mqPznYt+yVptiiU09SHRKx3SdZrMZxsTtkKI9yD1loI3Ct8Ox7GKGrayB+qVqGQFpBmtC1iw/4Uu
kdhmwfat79TucpMOglqe5IAY564LM9ym/hCXRlM7QETVMn7+zalZmALtDUWPxaiqMxZ+rgwOuQIW
zwPb3h+BKjQHBsSRqskwQuFENy95q41/E/0TvyLNvpe6eH+Am3c5feqS56/MTBaq2tYuYqiNR1jD
XAD/xax23Ur6LYsuEfhRjynZot/Rfbhc5BpARIuuSxvvyRDsZEB/ndq4DokSu9zKSd2Yx/o29waA
+tN5acaTUAx61fCLUcl8o6AChFUrcFjn7oEym0cWJ78cgCwESzzAHozUU8iKOOTe0ZZEPpsLbJSS
7kaZpLdA498OX2HJZFwEMp7WfXSlt7LYb8QqioGB9ckc2eiulBMU3PurHb8juuyh50Or7J2vaGo3
0yj1pI11exlIEbE9MhNh/EmOdaqMaGJFuhrnvRz27NGJMjOR31cpcOl1tGWM/Me3qirXaE7Z07x7
RU7151i1tV/nFk+XEREKX5G7v+y3nO1xAxKOd1JSyTBc7L02tM461xY0Hh48Om1nukiHQPk+8pLe
G7d41/T75Uhv7tMVTh6wsCrlza7qnhHXBPphgNXPhs4EiiSNYxlPIzVuL3AsHF7lHuYOMQdS/hhk
ynuoq34qWidX1+O2F2Jm9is5CF1PFiNeXIatLh1PAVjygDGy/l7UdHnRohla1hMNpiVb2JqM+BpJ
DOR2xXkadyexukvXh/9CZShTTKz3PAUjjxQL5JDtpIZn0fCYe90sMsk2o9MQiWpl0amWLW7gDFre
VckDRplrb5LaM6SPT+2yPUuCPVGEqF8iyJICHPbJRWNiPJKbsSYv4J+gv62n7TU5dcZcRDfc8W/z
SnuMOKrP2rlkQ40FgmYf72IrfCtIqi9t9+BO1TdVNgxadKGxmEC/kEBi2gdSFJD2WO84a+MD1kgJ
vjOjPrX7OO2YTH05JNOfQe5WP2rjQ4FscgBvsJgqawdfblRE/JedpJQqDtASnhZ7sGNRqzwN2Jw1
Jrh3IDhMOXToAtzTpsCfr2NSt1VubJfPvur201K8GRWis8IBqDAZDxx17OH1Ad0ePun96hc+vSQn
93r7R4q0FfPrWRf6sCm24qhczMqwpzHn276Jf3jK+F/owc70no/jHxQvpxKjfjAX+5eomTYL6KYW
DbDUEOiDRfLD9SoHo9nAaI05Zm1EVV1OmvoaBCddEq3whJrI03XmfldaJpUDXQ9mYkn59mctM1xN
ZKWlUtLC8ukIS3EGOufek6AVARH19uipKcOB889497UZEcuIXLfoP3pUEGqOpotfoyRgMXRvFbOi
Bhq2AtDQ+oQi9iuUHMQCBjnh91a58UyDM9fyrhCk+ukg/Tj2DT5dHntMmhGTP5AHzGo17YQdpsoT
f+4dCm2SrUDd5Y7s7mPgmfHZp35npaxShykzNpUy61LTyX0fp2LGWHmKRUZZ6PtXDEl3P+HdXfIt
XT1nUW3wInSXJI77D1jyi9DvqVv/FyAucl00FpjsEplwFMevtlZCXpEshTR0CxVzWw3mtnyGd5tC
jjA9I5L1SVhge6NjjkOHkKF5lprpRGoHPxtfCjbH+f7flnV0nZzK8qS00duFCTAcxY824SUS7ap7
qN0Ho4fwAMwPA4duG0ZxTCleo2YWPeaCdq4sHQ0rdz6a4mTcwaK6Fj/I4JbXepUKtapS0v1sdRD5
QbHfaRKn2/IX/v6CAzUEfIJlhIYsNAxkgeR0Y1jrabq93q4jNGT7yRSOdMW9OBWyfsu4YRelxxQG
DiyA70aG00XAu4jA/S0NgshorzmPMjUPgX0XKVRQ69Br93BypkcB8mA7Fwl8qGry6qo2eO4P4bQZ
WKbLf1B03uJ9/msgkSade29Rj5kTphC2dPkAv3YIFq3kTNxx57579D3JkTMNceJwzFWaguOky0vQ
ussbmdzqaSgXfYFGtdM9gXY0Gv8mh9KaxiISOwMXSBnJ58s01EI4ev0Ea6i46kNReWJbeh/9VvlE
C5UzSBgc3o2LceLF8es9fjux/+2xqtdHL902dGYnPjGVBuSi8O49o337tqbqgBJdLt3rut6md/ya
nzzRGxFfvP2LPEWmc6PYd9tvCwvwuKtzuYj1wsSiX324UJ7wAGu3J6/hUqEETDZKJPl/Dptxz5TW
acOPqVKwr9FwLejr3mOhq3n9MHaM4RKRuXpSUHuxmiSsSHdhxpKxnIvVlgaAdV79tvBFgFvhNBp0
2lYlHDtOYezWwHfxbKecNPLe5c46R5E7KhkhPf5WX6yTdgHZcvvRFh/n8QD5i8fxx4/mSXnw7+ww
4xYLfzfukBxSNrFBnBiCNTe8EAOF7I4I0IFjDFsG0sVE6PCFrMN5oTqaytWeo+iw/THz535KKp6c
nTWlR8FmrjRd4szjmkQGy1ipV9QS9DKT4pPj3GPZrMhBdlE0WS9YdNiaONn0fmUtUX2RmQ1rHcx1
X9afbEV8IfaoJSFlT2oxH2gwsiDmqpGRb0kiYrhpAwxIutBsC0L+eRwdWXXhaN6+ULUw4zTFv6ev
2VtQiOjp2xruaGTUZCKCYvoWf40NjCIfoWBDKslfbGtzqwOyienHCa3ineKI3Nq6y9cSgY7mcLpp
G1Tc+pgGzobw7BvcD1X18ems8Q3cPXhAtT5JrgVY82uSfvZ309uMoRlUpQ0DYduajwSBTHNl/4oM
+xDOFjZHSZ2Dj/jNdqO82Ps/dQ4+qd5DGmGE0bM9L9IqqPEdjzLsOxcWn3d582uk9Ap+u4+2+Q8L
DcEAMmPNPuHZ5vifV2mmic17FzkR7fejoeqy6yTDn0uyorr4BRR0Y9pZJ238pqQR9B+/GmLWz+Am
xemsJ1+TF57khA6nHz73bM2IHYaEJzGxnMrTiqnPFH4l+8TDq81SJdAbidPzDNM697ZWyqdYkan4
almy+KFDFiQPBZTITTzTm/P/y3TOXW+o9+lmKXdCzFZZWF7dXewVoapsl17a63rsT55s/ZONh2Y/
7U4qD0QLTh30jAp0BREo8gnds4X4483es71VoI8+9GIqo3E3t+tXC+NAeyA05a1lOl3o4QGLq1gu
excSoajypETGTdN8zkYa1aMYuQIAmSr2f520eqGCHnIqEEcTbxYfD3vRJLzhskQ2tT3eNnNeGAeN
wwvhlB6ozjShi18WpP+GxC53CG8eyTntLiob3fGeheNkAlF4MrugCKGQM6qxj3uBOh8PqK2MoZJy
U+GEOE1p5mUX+cJ4VRafdSgVmBa1Cjk9BEE2X8ETZHZMajRgoGwV7TSQ+pk2J/dLb0WoHxjzfyTx
DK7cQ1ICPR6UDJ/IylrczcL+YJdXj0XAOU4npI9zfxVBlFUGHL445tfiL8xbL8VlJTT1MgWF3CvL
+8LloviKo6FK9WGY9mzPd6Oktfx4M3KlBBO59UTGNiRNCt2HIlYt/4K2q5/MjdepkEmw3jGWQFpb
w+J4MsmPVCg3w5gXKRPY4rsMRCQT5S/tJQQ8cA8AZ8juMS7P6GnROBzkkdgZoe7wed+49I/qZXWq
te7BAsiSFptC4BpXFjVWVNMpWPQyIokr8HuFwExOLsvMMEULcTGXaW3olYrc7a9QPZh57qACgI6m
/sdvZdvihrqJu6AxvWVwAXeQ5ljGFoac8y9zb8zPgGRntlHJ0s43m5lOA67fIeWpIbfnT676pnc+
rCxNkZkCJnVCU2brUlxnQ6VyflzaE1cjb1bAqJPbS6FbuPLRBG3M0h/ygFva3ajLemNvDe7QVZmG
zc0x/llSDp4+f0Ad1Mg/ujApwL0Q49eN5tsztsNh9pdVRqmeD2iihyqzTggEH7ckPQtplobwrwsX
2jzHrJ4tAeSg2W/sfiDzj9p20ZKK2pfunZzPpEHqvP2mySQ2Hey8FU93IJpY0RXglNb87FdzWWv7
ZbJLQ8tpYj+l5XNAFjVDtBLJJKegd4C4LO/OpWoH1Rfm64UJ6Q0jKsN3+bM95Qe0/e4usMT8Wnf3
DgbTBRamRB70LRFG4BRPdLWtoU1i/Vu6bnMaU75rFzvaSuqoa7/QLYFCd9OeqQekch4bPKKL4d0v
IXCFLRb+FWM7TxwPkZb3bDaram5kC2f8qmfD6pXN9RzL+HFOAYs2CyDdtfFozGsM6YYDJ2Qxg2d/
NvVJ9Uihfqjg7KKdQWLxlA7391XcmkmJ7UltOCu85/k2oM6rqG+7Y6jL8AKuMKknZu6iSoNj2r5U
gQwXZ5TV/FEJskHCj4IOzsDx075Ro1sKAXCoaPyxhHqgUl1XNGsuh/BE4/+E+0t6IfHA55BGtSi0
CXSE82V9De1xqTC/yfh8L08TpYWw71VtSsUCDwXyDJl7h/64ElJey9Ef3GhFS1JnaKy+uY09b9gY
m8VuynOkrdNW1D2U+9kWkx1ao4m5WzAm7AUzhg3mDSTDzg9XLlUsQ8EpERUPDecCFpgQ030HVbRl
ZivnjxhkGGDaKNFxWY1tdAti30BdLNiaHjMJ+S9ne2Q4MOHCuXfcycLBU09M+pt7u7eVv3/FsIxc
QZNnd4XAfEOUKAtXeokLmFwvLascVL7OzVSMzW5leeBIj+h8NdxJwq1WZOuzLuYfJs3QQuoya8yD
xaqrPo6h3kyXHvHhWkTUHVc8kwky/t1r7XV2JA15UshSg2A/nND9GsorrLKdVXJl1ZfoTLGYcv05
EQdEoiQBdiuIpmBj+m0tzKi11Ay7ViTy5ic0+UIcpiqXWY3IrS3VW5yAehNz6cz7NEVO6WchFv8u
H6TD2rAdr9oS3kGQmzYfuoqXlnvGvATlSquYll7JFz1flD0vi8PVKPzNeEsPgMyFqu4DYZGKRENh
sDj+Sh+XOtXTlqhcEHewrLqNq8TnbaZtNd9qtA6Iwjy5tGtEz4LV8/6A6R3rtv9iIXU7adWQSvgm
GFbBx262EAQkV+d5TfNees3qjnJuursSA5t91Rdowuu0K22Q+qAPpmD4Ss30/1YFhqAwXhKwnVsT
Ih6TCpWhPw7r99YLCK/hhg9hXfbX7bsa4jfXh+T4VxWS8m+DkAfD5T3igKHeYwRD/tkRPAafZtlQ
GqhVDw04Z4eW6/sTzCa1XTiIBk2mVS8ME/3A7yGXbmL62ZXcFnWrtMS3bi9j+HGXCtspHlSb8lSP
UxaxCaFbWS3Jt7RvqItTqsGX3yZ+RxKKXej6+l62WuCVCojQWGwqLxR2RvMNmexeB3+Eb4L6OHtl
mea/cgzBtZhTleXB7oUy1OliB6VMUafYe3Y+iR1HkR0EaPYMK0Ss6pQOe7Ni678kFnosOSWL5Ece
xJ7c2GXGqtreMJl9DvJZ3IyxfO9sHvtPs3vtSY5Q/8MBV0KApBzTKG3hplm3eqFodP6Surtt+ChG
BXidzBpfimwyftLAxe4MqNIuqeTxoiKww6U3AJJirowD0MYJmWdsfIfOX+Qh/M3K7cJ38LZT4Vxx
StI8HSlZMBUKXNmmlQOtWo4CgoIMMocjK9OHZF/1yYX3j9fDDMYi4JkFp/GwRpRBeo1Od4V4wUEa
yaIAzz0g0X+R7U78fnu7tqPfPsmG39HsKEtz8l4Z7Tb0yK/pPdZG4EP2aBCcX+VZ4dc9VLUlCx/z
NWznkIAFO+E1dTh8Q9Wk5VcqI4X+KkxU/u7dXTwIJV6I8Yz/4lV+y9Kz2NEAl9Rqe+sXritb/v2d
Kg5ua+v33yyoGXw+FVlw/6SLVPcXsCw7PpqlBA8aiieccCPdy7y0/83gOxYW6uN3PV8r4P4Ft9IF
Z8CIDY7ZKTVOyZB6U1hMb6YsX/kXdHC4h7JFZKi1w4DX2aRZguhrO6QuWftL2jbHxQtFewrS/6or
vR7paqSwfP60d49zDznOhsg5dKkjm+xodsFc5WWEYl8lONvjRDV50m+ax+80WPiu+sSfuQ2C/75Q
g3a6Zo1CUBRJ0jaeuxGowgCznzed6zz6BiwGdJuPG0G8m5aCBrt0rgBVuomit7CxZdTnbrEdfVQa
3jE/qYcQ3VLJ5SFIlrw4MV8cQMLqXE2iyJbsjGkV1+KAfvapFNS0xv+j54nB0J/3VAy0STTX4Vw0
1hSXWFjgA9tu2Vmt+q86IiqdgTAz5M4ft5jWp7rKtcfg2xar95HnzloOyz/BMN4jli8LkNWk6HE2
YtsW1bMJWJlDDfi4fqSgRR80eAHtNXWc7Fc0Yixybh/KLRfkGCMJBijShOjHoznXGf0oEL4oMWl7
PIJUcga4A79+qWQOp6ntIIfE+rIfxOsGNragkjHQwl3WC0EpT7hgvoEId69YXJrsNZ1IGUoDPthZ
DVoGZeHGDmVgP7+y7g6yA7n5VJzTdehHr6oUkm8ISaSVt2kl6f12on4SN4Ywz6oi4WAf044yssN1
ktiLwGfxDMdulmz1mxAcrrGEma697OJ2+8pwAF4fgeLIH1ANdUiMCzkTiPXdeFlZGU5jta41cFdI
xXsTQzsaqz6HHv/oj/hzWOoKD0p2wFKcELpVr6NdkY0OWCI6QswXC+YfDKDVo4WoMQ5hSv3M60dk
zqYchMJU2i1QCXT8bApV2bmLX+qBRgoRGZ7AbL7h715X+4Uu0bL9yd2OMNnnSOWM4QepNi3upNkm
SShrCI4ihPKRhXhCIGvPzhDFB/XiEWiEigFnTnbt9Y3qpm54PtPpK+8oQpZ1IeFhhk0GtnTCQ4T9
qnM4Trmy3RZubCLjY5lf5pj1ENZC3n4B8dLIG0EWxKFfh68+FEbEmTsli+wnAlEGVqknZEqK6Gfz
B2PhP/w49Brfh+tTwOlReSTKO9VJ/jAufOnhd3yqwVwhtkHa0bCt8Mg4r9qYer5c++yEcfi4hgVS
eoS3x07k8OaHNBp8HM3H7E//849WP/fuWGxoeHL2o+rggMDvUJ3WIGpytFxDyDJ3uW26K/+2WMey
RMDfoSHjk9+a2u2XbHNSChIhpdtdcYFKZcwA0iwa+NspW+EFyACk/7xqQw9xdICcJKS9rF6WOG/X
AB0GmydW0srApe+zgUvhhuJOqS3EsCKgIAh0sxhFlpWCmCOQnEJcrcESAoeccTw6Iy+dqNNPuxLI
6cUxoFovGsNgoi0Jw3cHRfFpNNFoKttCYUHaHoneZ7edmj2te4qVDwI3WIx52Z5IHsjnooMNlCh+
fcDoXvZyTmwnDnVDqOoFpA8ccWby28A2St/51PzMitjxbtLmgm0XOZlHY+ceYdE4k4N9mCgB5t5y
sMBFzX0hK+ZbsWoNjw48xkJnAz7Pdk3hDqUROAG7ZW8h3VAAOBl5a8J0/kp9W4zjf539C3okDTLO
FftEKvzadcMbBPwC+ov5+wtSdmow9cO4eMd0GZEaDuy2eVpxLMIZtWwzASLzfjTqt7GfopwTz7oH
N9xE79eH7NofowsFef8OZ0UOmhgYLc11MhseZ5UWuyuY/p4XWd0TD1u9ygik3lDsziyjCO+v45ea
BQWDoDPiHc9m2Q205A1IaXDGrXsR79cDT+M7Cicjgq15qByBZDy2dDAG1Yp5NmoM3AP/gh0wEp7G
xA/UaLmiSIAYUP2XehaJ2Omz1W6s3j5Dzu0IqmYajxllD3RRVFE5zMcgbSmBaeVxOFr0GO9njZ0Q
WHZW8z6Yt4q8TKFJxh52z+yjxLaqyiuSWSk4MDAAomO92wy1HNiHCcqxoP/d58wcPsua9cCt4ZoE
UJYiJVUOqdXfonSaXE8s99VtZj/A0xW59jsEWPOUxvqyn0/02qBMsYhXy826babzQquVejILLqmS
8YC5N5Eaw90PvViQbpdRMqsSQC4ELANUGL42qpHpwcf21ZPVdSRGEu6X/j4aSwBxqJlm1grOBinf
PJ1SVgN8D+Gia1WbPzJGvdaq7r+Ym7jwtqzHyGpi6//NOORbch8laZsVNYNs1aBh97Zgc0M7SnLE
qRgX6McYuFtipKLlk2xciQSHEZHoKWvPTksuRam6UoGFkmxf6rZjotbY4tSo3R2GmG4n5k2Ils3u
hl9+aBDkZqOiqwhs9ZhlO0fI4JGZNopiw+h3pfMsGr7kJaEVBRjWuunFeEm5lKD8ixEWO9bWoStS
AmfE++RtlLy0AcQQ9TeP/v+/KHUslNp38P/8jEMypDwAuuNvxRM/P+Elvp+uQUekzk0apg7F3bb+
cw4oA4JXpyTg86NdttVMzBl+5uFL4F/qHeBVV005aSB7l5sMFxYddDdnlevLhKumO91QmSXc7F6k
Z1kKRVA/0KWydS+wNT3RFD5b33tY6ymCW+mBCT5BLGV869mdGw6YuYFX4Sr5V5xbPG2SOvI/3Dfr
T/lgH4AoQiLqbRHRWr6OGU88jFHql0yUn9n0yM41+TkkHhss7sJL6999CSiyf4tQpqHILNNPnVBU
yaMY9kcby00yIg+FfxIgvYEXBddBn5UCS2eJ1dGnWFONhAGXuzyzawEMIk/OsauNUCqA9gXrJdSt
KuEu6rO2vrx559mdUolnHWGFOqITrE8++NT7OMBIn9vg1VudTaqFMlY5bZlNvw+tPF3pmXoJYGlA
aVk6Zj017GaFyxCXb3fCa+Y//JyUf6EUCPBnT51WKr56VgWUw0+/55I/NFhcGbOkfRlLrxiRF54j
MLBf9yjPGJVB59n6UxCytUH4LFWX10JNAIozvrnhgT1swJjlCHRUNUQEFGPp+RRFo5tcHsKNg37y
YK2A7HpjV/FBEVL99brmmwrvrgJp0VPngSmcymiGUjjslHdBnPak4KZfiPGPVwL0q3D/w7k0ZCDZ
BsHJKhdpIIVu/KdAmkAcyuMkmTpKKcAfY5abIcyrveaqbEPj8+ax/cj9P7O3G3k57Abm60axxMvH
R5a+3k69ShqR4C9XvT8xbiYInxP0/JlkhUJ1CvCEizPncaMwJaeDO53doGZP7ACHiZLWw8g2PimQ
kkVCZeZu+yiUcy+ZVDa1u6bHBbcbJfITiE1NZug+NEa4f9J3jrvdWiC5OZREJLXuBNL0kZZrqYRP
hsxOzaZVk+yVgAlB68wu5/Ka9NkBZcLGvtkrUhk2Tn++55B+uKyc1ErjrzJu6f2skMrunLVgelPG
rRG6Alr20FShwNKwaaWVYogUe7XIqXWZog2SBc5X0HXuyoK1fpvDL8YoV2KrzJqnNUs/Dj7V2JjF
Te2gX7w0QA5MuUnzL5FOHk03sYYAyoS1s3AlhajZxXNjr+/R1dMUVbP3mlXXD6+3du4DsVX6S7zl
OfyFTy45UurNJuxpIqgBXvE5i4SLwR3cdbzOVBituXlCAlOOy5j8Fopnxpclja7vQtv8tZmhCgk6
HdrYNiEOWznVXqWSGCqwCIMv/3/DxhN/8yD2DyuMHXBKQjqvh+HWhYYXx+kb5aL1sazTeTHA8XDp
BK7yOIZMlVM8YWh5OHRNmwVLhUhgvdBKQld7crHFqdyU+udjmg9XHxg6aye5SKtURmCLKwxvKcsW
BaSoiVNT+m9AXFjUjsoX2B0vW8QiUWMQzku/thqCoYyA0YRziJ5LJZrxyOv/egbcFcKCh16/5hAX
h79SXFoRDk7sc75Bg1H6ZaGAnhY7w5HSss40aMOj3y63kdtDuvANTnSETYfWoA12p1Jqp45n+qQN
rN+SkyNRlm2bdTB6liSXEBzZmLxYFMhkxT85gSGQC8ijcYb6tXQCa20YAdVX67y2LYgR711csZlu
9A4cubq45tcudohRt/qfz7wHmQKeI73VG4ygS/LHhbKjjHf9M65zRIyOd/cZPUp52yJeF411K5fT
ZE6bmTgD4VQVRFajfEDP2bk/ck4kIgqd0vrHyFpsS9Bteqt5wuwLwZJ2yIfanSpxrJWOE0oHlnxQ
pcNqbpT0+vtc2m3zcV5o6kqC9NyJFbu5fK2ZOMTluxxUmMl2QPMx8czuxj8zRrPCK9nY5zW3/0sk
RqH2L5bFDq5H5yIcPFhv8/Nd+fkdrBMpyAxlQySUObSgbyfWci5vmcWVqXUQbuFUGyi0Dey7DKVP
wJZ3tLX5HoP6tjLfU6k70XCEbjx4oiNcudJLrokL45XVF1DjzKYBxr+cY92Eu/iHT4AOvG3EqcR+
+VFjyubCRlw6A/foRlHPP+FhvE6KFXYOv6Eqlm7io+l4nYfnrJxsHCYIzp130xc/yZDCvTdHO8pO
RzXdd21CmIs/8oBrJcE1t6+lPIzQZYz3rS8hF0d1uP33J5WL34xvfhqWeWYgqSUk2ljOp3vN1hc/
nwAb6ScN/S/2k+Iua+goVbYYSFmwYhK/TTCkUxzIRYaEwGQiqRuR9AWgUIfu3BQg3ig1H8IlXz9/
sg1a9QLzH/OA1D+NzgxO+Id/BoSjNMg7Y12wHW1FaDnxcV64Q0QoFrlSz1Fjyjuz2UnXJ9JKkpsE
mDGwfcjpWYkoHxgIYeTJKFw4HAs1dxHibCcQ+A9pRGKgjVb69PuVV6prqON3+JblZnFFf83xca0h
HBzmoN3xM7pbrh0b1F1QNq5rLVvZVb4JblXelr3QLV2SKoT3QUo9ElGUD2EUMLKsxEZhu6FSgktk
MuEOP7WItRD5eHYGXJqpvjP8oDmnINl0x1n5M4auh/PLNnb6Zq/mfSLxzfUtHSAyqzJZa05sJzWK
5vHPfwdt2+AfAHWJwgcOqa8Og6KDzrgm2f3btpU1zJbz0SkZ0bIB0ELETYH/ubH7jqgU0Vxo3CFQ
CWxA0OQSeK8lAPBt4O0JZ/IMavK5g2sL2r8kLNAug2MBNbWaHjpU2zeYBDeLNqe+4vlkxcBLCDkv
2qbDJ/J97P1xtEQ05gV5z1x7Us4ewrdE7kVWLuz0hOoGSWJRMpqhYW8fDtty0fL0hXS6wErto3ZA
wYqFebowx/Vp4JkJtDrXNrTYCw/F9ULxO7rgtLa15NasTnXCdIgVftRXHv105KemhhyDXRGb0DC6
INduaUYvX6PPDJ3tDH7ZQXEs6tT5kWW4TC+YSWpJ+VkD1IF0Yw3PW33Qe6qBLS+inE3AOLDtFWdn
GnL5lhmpw03Zmh7MbCkc0B/nqPeoqkXxkiHSSecLrMt9IQrXoUszggiQhyPToMQTy1TJ1CNB4TrY
Af1Zr/PRUpEme2ckjbb9n4E9QROilC4Z4CexT16TXIgl/PszSzqloLR2QGlKYkH5mbUnvnoy2clw
B7+fdE+jP0B1xOPM/ZxqPKX9upwf5lldxoZ2+uBbN1SUtfBN0PWHwTmBYhvqHmuiMyVS4GjORIpW
C1e5ZMQjacqwa/BqheDQ7y2rM0BfkEWTBwKFlf0/GC5ZJQ1qu08Abudc/IxcO02tQ4zt7HhQeRbw
+YhhyFbKYGP45/by5ggO1M4MGd2ZoDfCwYudsF25MN3I2HE6HDHTtxVxZv24mbIStwedTKpM8B0t
sCy7BlNchzYzFeHqSCl5C+IB0meZTRSLcqh6M3e850nRFEAyBbSSrDM/cTrwkHszhHl0au170uAM
Ja7LjxXqI411mdp0F9v/f1fS9ZDXPYKPla0WTIX4Dkz1g4HoL5zP0cwfgmtW9SQE+QAJlI6TpyhV
T6qkgXnbm04khAp0bvoaHrNHqYRAk5IY66faNkcFxbaKjvLw18ks7PVMJS495DX9YLxb1O2hgUea
k8VLG+21L7TzzOVyg1u1cxfiFrWvYZhJ7ePHusi4ucidU+ZihsOlFJO7I7/usxPSIjVjGkTHregj
VgbxETU1Q6ZnN1h9X5CijkE5Zp4sVh0oNXG6eOFosUUB6OGFd1YIEzfZLIxHva5WNSA0diUJLS8X
WwfbiAGJHJHO7l31DG+D0zKSKfbAGivzcnpVI+iyPzNRY0RkvXkyimSkpM2LdVIWbjSzlBjjPh3v
KVmDO/hdWOcmL2lhZPWCOla8PNAuVpY4j+2ugyAzM6uFQF0op419FbQG8QXqW1Nc9ysDhQdlAz/o
PL0nIX/vkNMk/xA/vBSkoix5gFv/uKZH8wUFRw38Okv6mMIL9uttiUrd8ZZmc9XopQyo7L/EEEGz
B7N1X0AqGTBisUszmf0DLQS8tiri9Cb3d7KvHriVbyzW78qdLPyMnj8S1sVt8YfbjkkETY4w1Ynk
cNR6bDGeEFDNG8PG4eOAVnTnPAN+zWwt5dfhefWxULwYN6sBtK3qaHm7ZYBW7AfCkALte4t/Uiqk
yhHeEXB2iqPNxVkQyeEnAYS6TTMmYx/YvcqK7mxvQ1sqENXXKSPc7kzZwd4s/yICY0pkzzu8J2Hi
j86HG/hJwE4cESVUNT0Uo7/0+FV09snuL5ANp2arilYyPx69H6kdntlJfCxAkEz9dahF+NWWv7lz
zjlcyD6YuAEB2TG4xzb4yitSHH8gePr2x9XH/dSyds5l3I33GiCWgOURG+QNLUBj1eA7f60Z5DkE
tcMEZihirYfwTby6C+Tli1eIDeS3bPeyGhtq3hJ2DxcS4CWGX8hPCWkUknheejDb94bkoUJLEuIS
3VDUjYdZA08wokmp5biUDggbCdKq/lqGghr/BYx8OgxDOn0U6McxRojNwPm/+FPsc67y9oK0SZqz
Do1BOikD2YsLjx7G4K2GBYlrBEbgyo4DpcjKM6vyfqv0gr5g5Caavv9rYEaF6p7YY1AulAgzJcxT
fTDP0wGQ8wqLWaqHIhZ8HFAKKEm9VYGU6xo3DNC/h/Y49YZA6qIy3Sr2IVXBLUBx9h2lvM+i8gtP
zp0zNp+qOr/AeYzM+uN0/LRKIuVee2P77GCMPH8r/aAcaFdq9PH05oFAXsEMImxze9dTNECAEmcZ
vJ42JHtWYdudAlVrLuVP2PXOkBPPDFBRVVEzAPJ7q0WrJLKgUgh/iPyAzICaKNYO1GoM90c7bclT
poYQCV2uJdiNTo3qc/SvTDWgP/9SMhFIGJ/XhI7oA3fZPzRfi5NRYZXaZYsn1tAxjx4bTtN6cDOM
QCZGi25RrbfIF7w2uxIM5xR3PPpxonlDytoih+XU7e6YC1pU3TG5M2SLbAyWARkc9NYwePdXkIP/
E8syxdBowXArIqF7AuSRJUdDepK1MwRQKWqonQbC9UH9GfK3JcrTBq7gRfLfqIl0V7k4QG0FESh6
z1E/fA1QXZtgcuZpasiRgyJzFssAMSRp5DH0ILPhU7G2IeO/SisymTSbnI9f5xoQTW1h8qP8NBE+
JdrccwlMjHMUTEhsx5GBxMt+aNrgAfD/NReuBOzvAPNoE93uF6sn4U8KblVtb3pXcszzO3Hm2FWV
KO9X1NDi06LKyd39OtyQogYy9gHS7Av9XzBZ2X82VSA1P+hJO4ZVxasPlM9dOwMXIjhpL06ZyFQk
twMh+y2s2g1x+2S31QOs/v316wHmYa43wDVt/keRogqc9cPFd/1to+K4ZUHSyXiDbpF6+vr3hz4l
yI1U3gwhYpKwHHMCCtS3CIg/S03eGcFXWDCI0n/pl27Xequ2umj9rWPEnYp4KhFasGPBmrvnJ4O8
98bSWEqnoVvtiRa40Un4WpnMeEkhDpPUXSbsfVGXNIqWPU4MDvvikI60dvh6bfqExS6J36etvM0f
qOuKvAqcjkMj1F4qmzy7zddEujg7ujL91b+G6LUfFlqgq0lUyhptLDm8VqN8R5iHoaoZJBGleAvi
I4h8Oj3Arl8Vf0tFioPpV3Xjq5rUioOCSIUf7zid/fFDsRytdxiLQDm1YZguDQQg0yBy+AuxAeAM
C6V2aqMsWkAoWqfFEDOS4lPreW72XLGRH6+20PbGBHiFohsqo+CqIpwq1dxsNq5qzjFbC48kE6/E
UYk0RLTCrjhSr/mDhfaaiWhJh4CPxO8Vnw3ReYQ54FKzZihR9LrBF0pGwSdG+chVYmDaSpQYtHmP
lg8H2tOZWC2YscMsPejeYkEvDTbftIKB+zaZU3MrWsjJIP/dJ3829XYBCyj0URY+b4uERADxp1bn
iW6goBHINqpsKFu/qjsPpwbRKKdW6x52RjTV7gCuF5jhGBGoJPPsqTOsrgb/TYtquO0ZcGUywBIX
vh9JERt14mLcpB8ft9HOkBOSf38Dbbcba5oFHrXjaQZqn1Y/yFNBMjIpTUIcveQUC3HYfWVXjfyS
wEjNXkVMDCOHxejcWINrosjLQxwF88N1F36N+VjFig2dyUbJK9x/AXs1qU/bBmhGlZZeM1xyuXpY
3u1Yo/OylmGDGl1mO/BhHE2S53+frtZieESjUGdVeU/uzOlXMoIbb48dT2AO1OvDjLkm1xwn/bbE
n+iqGNZKuHSt5ktlCHgx3sHIg3S+DghKTnT7AXtxXnFiNE1Eod7yU+5KYqVRZF9pctKXp8jAZFSD
IUwuzV9/GUovWBIsXCtjIGhXCGv5FOxm0LKv/R4HyooNBDDANIFCnyjL58hE/dSF1Esc9lLpdDpk
tx/cvUTMCIQRbzzUjsVfh/K/3nRlTRN+DXZA7ePG8HWBJiz74ieY9Rm5g5Ge092lORa/Ax6C26/+
r2Wm6Rq6SHMoZ/mfiJBEhmsYRSZo4++vLn/C1IQjyr6SCWoy66hFiP1rsRb/Z7JRQV4UoJloJYwX
vrOMEdgew4qpH4uS2U5RrLx+tucFpvQaFbL+iluaEIroRQlHMQfWSGqHKS96bfw35u9t0lS6tDy+
Ue4jily/+SMuggH/4DgVmiifYZoG3pEogfz6QmfIleTUH/aEzoWr5OqpFIyZAQ/Dqk5vjgLCgEei
H8s0TALUJwJoxSv/YJHGF2Wr/83aDUckwXyG6Y6OR8ArIV2HLNq5+PUg90OtwJaD22Sff21k3DZ9
rEsR93XPuGNriFjBU07G1B0pnuBES/Fg0tNtQnyhwNIRwZCAmdbGfTC+Uio9f5YqBSnFOQoD7SIJ
blymwkDEDfgRehhFWb5J4DHc7BEd8ZDKak/jKP+rDiWKe2FfES9g2+MHVROX5pqRP4oQgrB3+M69
wilvyjGGqiLxIrnKappva2OkktbvF5ywEsH5Rha4ZoljIsOg/4gahJT7ZqeA2urlnxUKRX498Bnw
p29OaUopuxFCDPSozOf6ZJuz19WSOAMzDo1+IiV8owNg97ezAasuSZByf8fmsJvgou8BkwUHyKCz
WtoAEc9tuhwqfug7kwHKaK86J6OdI2dEccZjvB3Vbouyg0WDX2tRDKvHwEOsOPLCleovRKnQ9q6V
VwBAWKjAgvDMmxOiVFNQHdcl3K52kSNWADh/Y67QKE1BCS0kpZOb3Pxb+MSxAuRW/KemoHTpr65w
RRW4+uj4TatpkoNHMriWkhU1d8tIJUhGc9uDi2Lbil4dORVIruteHd7TGzcDOgtX1MZvVQHstcVo
xbIbVdMYpqvWrfZ7jmQL3SxgUeD0UA32zqi9958t4hxOekwqWX7XhgT8cFKFk78N1GOsyyjGnXvL
Dc8FQ+57UhRoFVtbj/oLy2hMZG/6L7fMXJ2n/kHV2vD1YrybmuPIQNE90lNBM73CWsIzXfBMWJ2G
iyt/xJOxb9irjNig77Ufru9QtHzi0KuPZdMCv/II8ehIleDW/KtK1oGyDsSSMnDIN7vSwDl8ROn7
5T6ywyMFglR5oXi4UHglSChuugymR1WjDfBXrxKU2O332urPq2hSYo2n3/ohNB01cTZ+Tbyds7bQ
K2O6WCmWZeWimy5sMyBDjQbK7UHpUOJr2axIX5fmWAh2RLKnlq30E44L0F+xAlsXvOnvtxPL6knC
yCMhP/vu4ukXnEfDX1wNn2gL+YFP3id6yt8M1YMpwJgOW2QfI+f8GmLl+GGr+ebNtNP0Fao3Wtbs
WvsZGmYY7abvcdUCacCVPmL8b0Mwcsrn0IHIQoPXr3eW7tm50R8NcLuo7MDxNwhNQH4VaF7RIhQE
dAv7nr/Up+GwoR8GV6queN1D0AS6FotUprXs9uvfvRDd61VtnaH8whjxvunr+zBKzY8GFvgT/lNI
MyMay/84My8ToQi+We2kEmcsjP2wz8BHTsPDnCvzzktgYaYwG6tI/gSWsrL8oXI3RcPVnxm1TnSQ
oUPFYVzvUF3Xtv8OLU8zqJRrykpZV0NBczj4pLUsAk6jzYX+smAbQvYMOIfWq7y57kLtU1er/xL7
/G8EfO8+QmB3WPTUwAhSf1t633DCZGyZpet0+f3nBw0H2TcPkwYuhVMKL5iIjJ9zGUDxtjNdaO/7
l7fq22xdsM75GTZJLazuchEn9Q+C3ojCRtJPUWZsPyigOqIhcUU0SsMxGt3m99wHQ2Uwq1AyHdT0
LRl6kJnka/mRM2hCcAGumKqboGhOX5tTfp7V+IjUGJEsV2dxHE5zzm5f1ppk5u+gp4c+P0os2S8R
4HQiJOHFILGcoCTDgwM0L2hmYhwlF1H+hx3tFUy2Nq5NVEc5TlwUBDFUkqacazVt3+Ry6wj+fStc
r0KsU5WoPvakcVLpezW5nhATAAZAScYIuuAhkoI5I2vLmdlR2EHZxf6t5NY4z9C/NzBZgaOgvw1P
aFDs4dKB1aeflnDaBDncKZ6ASLF/FH5mrFHm8FWExBXSGW20l1zPkUyko41udADxVFnk2sB3BZ/b
ZcpyDS+R4VPB1e9WKppz1BsocjPRmF8ooJR0LnS8bLYtwk/GYgRBLApqvh4JX2293QX4n4tlyyqm
03KwYElbha5/d+y2eb9Gd4WQGYRWtxJZuHc2f2jPh3yx3u/WFl/C/8h5frv5X7GFLqpspS9POiMt
+90TCsI/36R+MFDdXbNMxW8OoCG5GFPNCGILEwuCLVkgUGtdYicnczoY9LN0NKBXldHgj7GBlsUB
soRNN37+Q+iuXvvS1adrE89+IrbbyyoMqJfQmJRVg/xBtt7TR5aty67ps+Z+WfRFqy7iwu/JF0RJ
B35EyLkUgvkJGp3oypfEe37X9NAvnbCrjJxITPG1wKt/7f+h0hpydShDsozEiDMFBZmWTJ/DNzqB
splBcmjb+sDMYrSmZkuIwX4qSWr1XrCCjAyql2ysSd1qU5tad51Cr+yxhUOp2Y8gIEywRGqriUF4
TOGTECOrIorc4LQwna5omV9frgdaBpQtgBElEoyca/LxwZN+gj1eFe3cvZIq0xRE+LWCh5dj5g1t
UBiseSiZJ8bydyS3yx3BUAG/CcV9XSj5qHjpHAQcDlJYvahE3oA3KQ4E/jk6yMrY/DP/lnVrSUS+
gJ2NChFB+Wrr229eiYnlL+E10VggaDhVpEIa4RIruxq1prqxwzJaiKpf5ZHZit9qJ6Jk1hgT+Qtg
tiXQbmPtWYKcgMB+k5vn04DAyLOyhDNNLp2EfjIe51U6HHJ5dYOXsPaKye/szQlXjKSm1Gc4DYxb
l13tRRdwPFe8Qi7kAKePLasBIPGd1VErMQ/cL7tVWpB4qTkFNsZC8lHsD5T8pcUGpxj5kj64OnFj
U8j6mCWfFy1tca6k1DyB7nbssBab/nxl6LLYsrgHhureWQ0iUkbjxmrUXF8n+Uh/RkjoPcLmsYzK
FYvBsBZDCLuWZPvTjp1gC0MxuEHJ+llK1bb3WjLSbm7NDW8J9iFWHoeikZB82pcjhpZuRjkERy0u
EpYHYwg61eQQuIXpbxbHRZIuhZdmSQpEIXrVAY5aYQFwXNOWSP+tP95J/OU0xYtg28mxPXQ0u6rs
bjGCzeStW8GRCAxc5GiT06EgBvRFLeSk4DpkrnNMw6uXun3dWuSpPUfjluSUtXM4GgsVX/+arPOA
mToGKofsY9JKwN/Lh8XrSlxKSWscGGa7uAGYE9mRfq1PWq+5g0UJB92rYhcvY4K1NcZzW5LuB78T
as3GCQC6LQiOol6gCzFhr7iU/xtjCZ8TVGPa3A2VoDH651N42/tNZPpbpOXUdDI52LUPNeKoDEhI
RHM/klc8cGMpBc7dd6DImJn6WmkGHQeS/EmyGMdhM2UTSJZPxLvA0qBZQycDrQVkyqYTVS1u1Zzz
RTstCFoc3Xtoi+oc+mAr0HnjQEj0etyF4VHkKwJAe1hoZaXAFnPo8Q7gosxjZG/OSnlZj4wE3pv4
Hbw9GtvdpOxJ1QzetDwZEZCX96Z6fBxliVO0hOzKsfHkvyxtmiKyH7PfIGjwqqvO9sf5Rpvc/NZg
vbo1nmlHHzyjjmd6Sw+hkWfHoJnoqm0BH5G23zr9F4/aWajLuyGW+vNbE1JXFJlNL5glYrRQmVBZ
yG4BKvR878s3SANKy99iIRVpSDAErJuQ/dZtRZMvAXcS/Yqq1Ku15aYZodBhfx/kPId4MNxHsOrA
PuqS32grueaj806ZPD1m9mAh9LpO5o5iBTl8a1Cfo/Vbbl9LGUb78sMvJI5PR4FK2UDZSmjraNQ5
WaOt9ADI+cHLhLXshYc+RBIEq7hB7OttC9KhieCtquN5MZp0BhVLR87V46NHD8d4c3dkCDROdUZh
j/AMgRIyBnnIHtgQJhwgwjDyyHmUDCOWHawX7nhaqI5zUeiZl+S9K/qaeS05jQMcxJ5FLqGSoDFO
AHy/zs69rYMCzv8Yi98d3f4EqSE3kZfX3D982h9/S4TakchPpIObH/VahP4mT4zhj6qVClfJwygp
JAV9+GSYBA8PO0l0/fTSmPUSArzi6wxDOfiI0L9oZoO+Xghc6VIW3hd5oq3CNawD+jNUyydNF66k
1KSYA5u9xInydDyGfTS9KYtU5akCd0C1t4WPWGiQv3Ikemqpdo9L1eOhdX57vOkSyL88Us247F6k
mSArNxYwIfDHsFdbQB9rVkhn+EIsufdW3SbJm0WrPZJ5rDrHiyXJKQ59L75JO3rpsbNlkGr0eiAt
SPwzi+BPutWSXj20DU6thD5QiC2DQ+VwbsQsnmdbYIWKAcmqaRO2I1pBl81eBzIMUgnl96wKW+hJ
u514Gjxa/IqOt+nCbUB8mdEISLuXSQc/SyJyiSFnMv1TdS/CL0GRL8tRMOKJFU73gS4Xn26bErF7
M0e0OUdFSKYrZ+TmiAzVFItgOyeIvmEKmIx7mNI51jCngjOKe9AMcAcj3qe5EDwsbgB12HxgYtxC
/cHmS7aMtr0ffiZg59CyyjdsqdTZuIb0h7SRLxl0keDrzaV9IaUzjTCB7PMCO9wnfacuUdsXjg7B
+1L+PqBHUWN8fz7MIhiJWjfq4NuKGXp6LujHj7dwVhwVdKWQEF1v+wCvTk2e9vN4IBpyjZlZQjAq
h+TtA7o79qWLRgZJComyIHNSsZ4u1CD595FiOE0mYAJ97OLek5DfOEM68ds0amxtF9JLz2FKTPar
DP3KSVWvnCpk7+4FZPkPZCJaxFpx09jj1+3+bxZkMQyXzz4PqeFYU6ojL6HxnRn3gtC2ebaGrBjP
C7VM/xwdQpS6K1zIGtmmEOJESrK43s4ok6pTWxXtFcJ5GKh553k6WvuBcOwxhV+1jWKORLIRoVHz
OK92oVXL1sAvxOKxtOYvMNgvSAJrPM/Jo6fOz81KZUh7rEc9VsDIGMul3TwyNttY1iZwyA3ZyLkN
A9lDJbe1t4P0DnQ2rSR9jgIsRKfLmzjUsWrIdnfyZ0B0I0zyE/EJ1F5zpzo3G10MBt6MMZNny+BM
C2bHu+uoKpkj0JotWT0ZbBQJI/tEdZ8EyeuA16+aUJIqtzy8DCbzP5luN6Fy36tJBmuzvbjkAQ0L
AeLsM4HBSTSNNKGseuNNETLJLa6gC/qMsKwTlsZASkxJp81UgWXWe3r6khpvggMn9RWW1uJdn3qy
HVA7NcxxZtFh2xWoWR79CqtLjhhOSDXUax5BI3Bfj8qbJrCF3HXyMxjHt23f6r2sExP7edMrEa6L
2bxWR6++s89SsCwlA3PDQsnU01mZAua6Y3PpL8Mw5qN7qftS5btcfgPZWVSYuSrgQ+Dzrcty3ymi
Vlmb52wwXCebiLTN6YLAuAXntj3Mh5eZX4M0dBH98D1vCWkGh7tVLmJidq0WFj59/6n2bAlK+uUH
5CF/1AkSBSdJoPFVqNROQ1h2EB9LsAKZeXvFGMadR+YHEuKM36EL+X8FZbDq0JOGah2WlgZifySX
iGCzOfnT5VOyT08a5/XtBZLdBR5qrLMZXFrIqY1fIFqZAJ5Cy+87ylRK+KXqKFobQP5T54NE9AZV
uqVWcjaf3iKNHxJgFjoLFR2w80eHvXdnWuTyL4T9bpLD81B16T8qtttfR9ZStSxwtOifX5QUvl0l
ITCzZ4y/0Xs0FZBMKG9Xf9NWFmyqZO/IRP/6OZkB/lpEmdIuNgbETuKezoCmzKSQ7+uVym7Cx+ON
hwnkHg0LSg60hjsO9IIIx1tIlRdjkFjTjAIzllpk22XxBx/UDHqPG10qLyWwH/XVIrCQySxeAkoH
moXC7eLsi0TFrOjyQLHnZ2Xc6rA/T3RopoqOphohh1BpJI0Du9i18Qj46qlOTC1SLkCDe5b97Yb5
bfJs/vzU4qNk5Mx39c8Nw321YwM3RF0q19ZFXSgCyIZ8SSbgUde2HSYCt2j67AgOpcQ/6Uugiw48
2Zmk4iRNCRfOPmU2IkzVXllD8wxSw/bqNmBBXtWnHhbgiOFqYDHTz5vvP6t2r3Lw6J/8h35b+FL+
KgRCvghmLf2o60fYjivCx9yB7FoYEdiOtGgRt250518n0G4kho2jb3sJZh/tW6O5EuJ7RgheVWZe
E5wlmUeE4c2xMiF1wR09JRruO3mH34y/JfJavYbV1OC5lnJOGahOobaeWK5ktq3r6j5KhVrWO+ad
OnUChae0lA9NFd94zx54fvMay8dU44PZLbCBxMkBrS+MiTdzQ+PsdbPjQzSogQY42CnZ/XRVJs+v
n9vHv/7eRb5bsiM1H7WB5IdRtNywKUencEtF7bgWswC2v9UT6DQHdS3KLD0jzmkOZIqpCfW0Izb7
cmsk35hRvwu4KGZkyccHqFyVNaiRqQIg6yY8oiGF0e5TjGynHHpEBKRKi7HY29w+WDUWCHlcMkOO
SNlIZP0B7hZD2veHCTf9H2lqXxfZnsHK2hu7FqQGFNPwGHqpbZ/Zk7AWQYQKA/HZtIhTASdXZGFX
l3LFFFEw/6aygzQJU1t7IWmX1nf51HLu77ezN/mvk1m86fsbER0FZIYXEC+KMQubkP5jtse+9lUv
3wsvPRnyg06ZU6LwAwfA3/3YA6zzskkBTmhuzXHra9nCTS67o4EMDjrvMd+gU+twasEUcDA30f+0
gbHIgzlDO0AcvGqS92lomxZCGFbko142hIQrcC/UChsS1tpKl0vBxk/UPgmp1KSmSu5rxiE3uGa4
Ws+GNq0tUneoDx1LnFa+RBN+n9Fw9KkaJlfOn7Y5ZGeCsiH78Tx2ZQLXCsjQXSl5ciAAcXY2sIu3
lNGrXnz3eAsIHzzlGDhSlWLWQEsH0NisING7ii9UsWJUrnjEJvDiL1kOUBJK6EIq9dXeITgvW/0X
sk1rJF4W7h4A3D0rNSG6g1soROPHZHbhyiO1erBZc/OQ15ewta6fm76XOgiRm/cnhTdyzVvTrZ3O
d0d5wZgcPBTNNAHA+hCjv9ePfizuEcrdEPkHnqoXBDW7q5GoeItJ10QyUFpRcnm7zE6uD2MbKlvj
Zv1RAmCAwZDH9I7Uf7NveE5UGsW+Q2tDMOkaM6aF8DzxhKFYXh6z+o3YRGI7pp9T1Y163EIWHhYb
v1cZb1pdn6Fd976KXrTKS54klv/g4xlT2QVaq5C1ol24puyqlF1G2/MfyXE0mI5v910EcJQECwCv
iyUZH4zOXh8pewQe0tEwSEpDP0VrswfK5yDDY0qtpbNISqbgzXsN2gmQAQAqGTxFd2Xk4A+3xsCE
U+oCMZj2KouPs02ptR1xg41zbupM6vFelHstU++/9Tp+ax7PfG/pyGZJqgIfXtAdfisvkjwP1u54
18RRvzg5iq7JHt2T2v16QznCpRinw+jKU2aYGPaYzn6lqCH06clCncP8GOOnWvMWufA3O8oNW4Rp
3RebrIZ2gPeI2xXFLU3I+HWpenxmPJQh6vyX2XCJow+cNZBb0Ua/0IyNr2h5fl8q4/cNP8OufWVl
WERwq9zPq9pyeI6qxDQxClWhlP5Ec2RAw/BZmdOV20Xfz3mheR8pF0d4eWuZMz3K9SWNaaHI8P8i
pjUIyI+/mcrk26wcZ314axj38JMuY68S0FIzLsihwBfg/iBuNT1ihcYDoaeZFdhh+W4QHmdCcn0l
tcrE7OGSimuL16+IQoWj6MltqkIKOfg49SztykJ76t+heYoTdWmuxFodEgsBsrNuk8t7kv9QcBtu
/z/frsTZEdyvQHtMWl2CZKG5+mCqKVV3uX96H9GANZe98ltntQmhYNGIq4JLd/Um3ewLd3lY6H9Y
aHTdCPBS9UQ9cY2O9c0aZUu7COZK7oKIFA2oDXY5Dxb/gW2tCtTrGniT72B3/66L4uk8QuklYInW
hY6U3EqJX+N64G44IJiPI4b1SHwEFlFJM7gMpmR3GbUNIlBYVLPzagmEVUDrz4Jd3U8/47lR3njr
MzKEXzzbzCZx4AZ8nSaG4f/01DWsHbetsUd8yy34y5NBmAvCsjKNqU0VXefeGcI7VtikVFokQiUt
RhJVYQg43NGYCSsLHHTnU/VAPgIM1QS81nDy9H+AwqwQb+90690JnNJM7H91lu0TaLefjcyU9psj
fY+S2dnPJesJFO2U4ZPY3vR+tw/wROZ8DQ4ULcVMK40WwXXdFmuOZMhhNAqYqrXr5viHuy37oLoZ
mnyYWaw3tyN+Gw5dDp5BcA0Nkr4FCxTCGmmAe97wdrIziC4qCGj1GWts5h+hjZLfMF5tQ1mbNDI0
Xr4vCDHJWzXMn4u85ETl3DxpIACha3zrNbaprHZpUWuacEHUP+j8ZKNSLMp3dukj0W2FO77M/ewW
pDpmdLCXGVFWPkPzRmV1mBWep6hSwCr5Y5hED1Bi5ti7kxzzVfLW3bRih6Dpp4qWdbas3+ypBSqz
9uPZjUHl9Jv7Fnrrn8WiZb6APwShR5fRs7mi78njPgOdkbDqGOKl+Ortf1c1cBpjm1hbyoiV9Y7+
RYCLAQvTdSSN5SkWiUKRNQiXJRKUkxS10VySiIxouCm9tLiWBCTNs/9aMqvWlSJ6+rZKx22vcuE9
+u5HARXyZ5hyTbksY8aEkqpM7geOH3BlGcRUs2KLySZXOy1VrsByStpfdN/c9FlKa93ShWj8K1P5
l5Lsyv9dn0KNAFNBAMVL+vMbJvJhfChmExpMVJ87H2GdSQWBcuTuBqpyvhfSKwcrMPBpdnAr7kgN
7nyWvyHwHO4FdpFbfH54eefj7LAJ71UmLjUpdBHhqRbSD0VY7fWteNZI4NMWHjrxeorBa5oajUnu
P6ldYE6vet3LZnCFs5SYwETuDWgvaaRH7FCcoboY9zUFsp0j0Qis/Tzikj9w2/XPBEkLBYnLtdQM
xYbwjKcxQaKZsG0hAZhdPm7iIRG6J17phBKwl1NAiYYn5Zxm0Zi9o4Wdae4xU3K1eCq+Ht/QIX4h
civJGOttzcZPtdPwRiw/I4IkNSk1MRzL6hcvk+U7IOhDVzfRnYjLy9hjnfP7ugnpfeMMcM0Ukmh7
R/MQiWxMrQiHNJX5Utc7TcEDheHvWykzZ/Ek62+myAuu7wgsxiu3fot5cmNYd7zEsYYzYRdwAXkv
fYB2wYV8H4ODYo/Z4kngRAoY7ce9oKr98Bnut6PP/nzpTrR8H23c6fDd9hUxRDwfsZQXPPmvfjnc
wPKzDNYN8spTCLdOpsAVGo1pK5MOtcn5GdhlkMja4TPrxZg2Ij3xnz1/1l+n07BGt9Wjn2mLgnZt
pK9HRwduhFjhrggqUDCFljHtWEHNwpf5eEAa9NyxoLggWWe2a4ZgR60vKplQp9KLdtTh523YQOz1
fekijjvkBaQZj8cMRE8tP681EnUxe+qNgg2G99trRV2vd2JF8vhkkxbZTqYNyiO/B+0QR6LAKAWp
PIX1xDcIUKFEcM/sGcAOpO4IrS3mjN5u4ONqS6xRmAyzuAw3T/sC7r7O1OWnGiGoeXchKuMgd5FC
Y4vcDAXjEYlD0Ipd5WUtLYwFbhEfBsmKllu76IS0g+nnHoSbR6R70A02RLUmsHR+NNrH+AHMU0AY
eZyeSLaGhbz5QIz47Q12+lW2jZvuRKPxypyz0OxAsxM9GE5oqfT8etI10FOfndQpmSQWnto00Iz3
UTENABwbIZWEuzZoaRwuqUMqDaYRiJ989sEbgq2Ekt+6ucCltNeIAHz3tUzwk0JIg7JsqTEkj/ql
NIADGqY1mYBVZARCH2toFH5DoZOQjxxTKzqUYO5wIOP4WXrfkAYmzPV3wiibptVmufbMGAWYu39l
ZbSd/MXDLW1dwx7eSxFcuaHrJnJPDhNlHj27a/UYf/msm8FxmWLwnjlOAUL0+IODRlcyFNiFwvU0
ptSf1YcZNoXn9zm5f6d3Hdb1OBzZj/jc+aiubwcxvCkwCcI27X3Adza/TTjGxAt9YwRYPqmxzq3P
PVfVNioxVYaMUIkc7R9DRRCDE1i4tfWpZAkmjfMuzih4p6rHBhnu57vVMHehfDFP6s7pmj7cj7dX
G5LFNpABety/usncRMf2XjHmLt1VobCOQQ6aIr//PpTYgeKZ60POrUP63oRRQWTY5RRYMIiV0QT5
wDpxwHV3IHhtCsiq+wrIiJiMdPXSvey/ADljCfOfqzyQ4Cl/EUpG9jGd0Zpzsov5HDjEhtfxq3yA
w85akmP8vYq7BRJASQVLdNy7Ds5LGiI0HOPYhsLjHrFPEPO2VB8mZtjC56WmGSjJTlRZ9QWWvW5h
hKtHaSCSNSK45bvV/lB2xdBwEPlvaTHnrXmPRCikVi91PO6pA5lM6Gif+6Ivxdr6+Bn3L7kBEXWB
y5JlDvXqMsWEe+/Vq5i3mC5FeTJMMC/xZJJNhBfWdHkNTUhvGjaaQ2E/F9DRtiTg/vGs+mpC2D5v
3Ll/2AIMt1MAvepYUqO4k2VKPfiDo2RpEgQQT7JvhUrN0Gw4kqCxoTQiPi3dljm8VNW3MW5P9dqX
2CoXE69tmVqFWzHjbDqP2f2r78qJb8xy6eSLcXelVYWdL0x+i4xHPGgHOnoGubEB+PjWN4281lrv
DNF9mTUsXf6kPnwX9fF96AZ99YtBO0QQKvcdzF56o7ywEIrqy39ea41Jd+laJ7+tWtKOg4Dli8JZ
KDZMsjgOzu/ERN9xQohihhxlu/tedU50IQnptJ2ZAKCcO6RDXsR6rDjHPNsQezWP7uc2c2ZnApw0
mSf4bY0JEUGsuK0CSn7X3iVPUzaHghiDpgN02eE1G5Yj0v1SlEuK9Me4uSF4Ue02vG2hPU+eEWAI
fvDpw0I9FAsbwCgQEQvhyiVK0FQehx4fWrO3C2UQMzwtlDoPnib8IvCh5QuMu0KUBk7HHCz4i/a6
eBCP7V3RZif5F9Dh2LZ216AAg6LZPKD56mZRbu3KSg0/rsGIU9nD2v7XsrSvnzHqfc/l5qLkypL6
UeWF2dxfcgg1sQi+uyvhbQJQmal7RtIPkQmXMIKm6w1Vc1piEUAJXj8DpjDbA2JF2/4Ap718iUDn
2u80ZLpSt053h9MUsVvGFOAW+QuBvFmksDdPT0R16ITUfUNotl+nGmPeNUXrxN+x+jdgEwovwd9E
l2a5hrdeV18XzoB6H1IkVeV8W6oK4vpbW8ACp8tfwrfE6Q5oYSx5FWoCgKsk0hNAY1FjBG24ulE4
k5SrbyC5SrXhcNeBF2/5nfelpTjvp2nWtYzHWl87SuTZnFYSDSGE1/9xdGc8fS0Lem0tQaPE6LXJ
b3AAtrX8qwcLliOtnzY03fYRZwOvZL7NpPf/3By/s2kgSepqXBVr+vKUSBIJstAVrZ4QLBhIFQOl
5IHaKhqh7lNUtz3cvwe9rVVsr+K6/vrEkP5QqAqX3gDxCxmE3hfiYdBDeaUGnBW8BkQG+h4cpRTS
wwgr8iW8V4C5rSntROFCKswI+ClC3ex1JvhwyVK3K+KjIWCB447fN2hbouDg8JLg0Aam2xxKloZI
fbuR2Na6hxTQYbLpQtHUkoG6sxaezFqOU+nQXuQmQiVM8wxoYXreoN2f5bTtMFf8fyHt/4r90AcB
SH+5saZfcspQLuFAoeJRxvCHAscdDqS49V5+v4HHVIev0OgF9xCnPny9TkLLtbFvOSG5MBlly/UN
WOT80iVTgvT1kCYfh4LCr9rbjZSv2hebK+IVhlphPO0ZAfHIitQISxSKUQEr/9t3gi+klAoBHDcU
St07ttuK0diE7FpufXyWJbjBApCuJCmk1GGJEY7q5ldoXhJQIFPLInJUbJ6gYPYEprG4EqIdjT3x
l7tslRp3XY35SUCdLGUSyN3P5yGh7nTjD1RP5qceXPkTPHZAZq9XxQXsGNoUMLXs+9IMUCxBNO2s
zn3nCzNqL/AAZUafImaHkd0UN9F1sRjTlkOEXzqir/g8ZOupB1XomkDTWJmHs7wQqJ00jmyqvX80
yIGnN5GBaaGmjbO3zqK1BJZWVE5hCl6GxbCbA9zrshggCiCylbCKAvyDrzWA8qptTlNJxiPIH+l+
Hk0pemPvHHg1xLWVJ5NlaKYNn6xrkrFuXBEvD1E/lT8Am1XA61QAN6eJ4Ump4OXOK8TpXS6gdbvN
bwETNQWkzT+nH66OJOTZaQYqTQkQzXd9qqn/7zTLnszHbLPcbjrMSguyXpbKJI9G/HDvzl6NFqxC
eocvqAKGjlC60vq+lrFgeDNI+Rk5glzdNuz+k9Wu87m+cQYme3hbM2smL2xl4/6rU11j74W0kf4W
kAPIbK3vx1NFkB57xURN5qxpJsfIVzflfYPTGJg/lZJXym9NQXD4FCwc62+4XMwbz+59zE/KVJzt
d97CCgaCeoHchsWS38ldhSk2lvzO3wpMTHkNXn/ZJm3i9lrOPJxFCOrmKHVzd+joPSwxyaynBjC5
dNvTUlGoEAoPqZXg4n+MSvlja3uxz57K2TP5DR2hoTxBqfjN5/PSNGHT+OW7azWjR8iDvbttb46O
UH4desRWJc14AeoQmvXsN1+IIzJiHwBMmnZSXWhgWRvUfJ8rINeC9H7O6C2XnZpGvdlsi6mkfCkq
Y7m5WSYCKZyHejfsnKCUvHq6wshW8eQcaZsafLMHUsSdYmJhYJGY5qcSlTk/ySIoAyZ+A0OJu6se
q164AgKcg+JQKV44FF8598/uqNXdNU0Y3ahWwpSAdH3cENilsjda19JPUbP46MpmjqUTAmPTlAZ6
HedYVsmUn58r/wM+m1DtAf8i3rSNcb4QGmSsJ7SVErwrVZeMNjgt6MAmm2J+/xUUzRBrI1xUzQCi
ytHwWJmjeQoBQ0pzryn1u4kYo3h/5eVLQ1sHXIYxFABkIF8exfiaF85NcTvM2RlTmJMPSHyupE/w
DUWf7M0jWOzT93ja9t9gNJrmmwRfijMNbAmssQ8UjEZYMRzaYGADao39gIAp3D/CGasOItbvIneA
aWt3HDv0UZcEfj6wvetokWEEjyO1r6FjlG+JzHW378HknlrqS4/JnrRTufeoO4X5FlJZAnu0L8KR
qskGgAKICNVYojF3msW/8CpkwfOxP3e9GpZ2D2B2ut+sph4SZ9Af70lR+6C/64eYR757du1xnATX
KbbZDk28jcha41hsbsC6fH6RCzq5+fA95x/oCxtlR8NtrR8H0YHzdFwGUtiFZbhf/HKUktbddYoi
AOx9nplmXRuUYtj/1kOqhFuoLpKeIizacumV+CTGzLf60O4O97ytFGAEZGapm2qbYmvKZMqGV8ak
8eV4f2pCAz/M/7ZapG7+nKfZUzfZ3ci/iaZ3Yxmu9J5EWTzIweiOA8cPKUwsDGhTkJj6H+KPu+Kw
GPqVSBBJ70WX/Sd8ZHg+6HWt2ix5P3RVT4Yp+jQ0KB4Mnog/cmGvhltMh7ivjHV73SeytVld0XFC
efik4y4OHJDUiQbAI3cT0XGOGUvPlflRgdk2wTUYsIzJHzny0qlv04/kGdhqB5OZsRYZ4/8RIU8a
FHcqTo/X5gjsKqyXOQhcBjiQKtE92+wLTIU4SxZ/z1koxkAwm7oiWsMKppcbkGH0UR6YzbAwiIF+
jxia42IFPTXhRVZl/flR7PDsMz/NulaL3KD3etnIPODIhNY2lbQi8pElK4jQtZEoc8cEtV//0SPh
5oyxADE6Ad2H3sQ1Ida2zh2T1owF3EATO2GpPu1BKV6jhy3CB5Vjom9cjrfaOTmWqIhKr6LzCPWF
8RkhEamuNQWJ9Z+jhbv3z1BBO+jfaz5J5r+/GOU1pHB9hMctENUg/npBlLdo5c8moE3hGQMB2Lgo
KUzudy7SKML8nC4zkSQxUthHPHNxn2xlnVJ66kdaqowpa9jnW1XahcoC5n1DNrrTPLCB6Wj2J7d5
ZLTteBiAfnTSwpfr6FLksmp8akfE0bQDfSLIkqNWzp+1+KLuKQDGZJLmYMAgpnlz/jguXKZFmrHx
p4V7Q307vH/rOLpnoH8XUwz/sXOePeq/hFgKsZd7WfkL3oWq37FzRESiDX/Gs2+y0cR8qJDc5T6t
JdlCeOOSbnIQKpnOB87te00eKHDfaLxNKnxgckhFFtsfYNboYOvpC9BIAlyNZfdoEUwHZgE0UTBQ
OufUzBWxq/wTWlmEd+JnSXM1AkZqkt4TXr13NPS7/QkYKqSkc8QQpj6krsSLfriI3Pd6h49VB6C2
TkMocEvdLnFvvlRecaut/QoEpNLXiIbUDyY2NPtjjwuD9xg/mOHOXed2wgnO44qR9/52wdRW9Hb8
PUwownIXGXe83/kw1yWbH8eH9Jr8t/eZkTbjIJjw6jkvgFm/vcaXD0c2vD+BHzjK0TfYLhn8QIdr
3zcEf7XQnV5MMX5MJnaWQt7KLN0xsfm1c8Mkf0geARHAlv3koARHZu8IfJ133hAzhX8EguwFBatB
rMWQJYP3qrZFW98zjblU+Mcy4+GbWGkgAhr9Ruc2PtCW7PL+PbvmP9uLsQVzIJUHF2jU81E0vLy+
f7hhCNIAiidohJrY2C55JvQnoYihlXa+nCXwCEe8Z/HgvFFom3sKWUkZvYppzVPESMxMvBmIlcyh
4hOr26eHdqOzyS10d3luEnDNKF0SH1+/UdvKL4fZ9JW/sHYXlNqhsS8g3fqtfAIZW8V6htnlQU1f
jrTAgLuLNWyd1n/kARoL123bq5HwvDaUDDw4RtwzoMCJp+nWS8IXU0WD28kMNnbe2fyNrAT5muLa
MVjMWJn4JDcpClljjDdrNjzdvrvaxMH39qk9oSjhWgfm58WGdNdKq1bsIvCHbGFr4bdo/fD402kB
O4gTAF+u4phi0tpIhW21fzGnUgYg5OhcvNJ/NXdnd2mVgp7vNr1z6+cplgpikhy1zPrWXcWsO+8q
mpuSwV15xRyG1u9pvQbXM2hACeinyxb5PNuQ8k+FSEdf6ByZ6uaebGxztQBXjF5EyPdgsuqLcHWZ
QN+AggjClgafX46vYh0MKD28erpy7wmn9iJ9par1QFRjWcjxzr5XCRvrf/bZO3zsGc3bg5a+gQjT
EppMT2KGvM5Kk/el45zhrYpwUrgZbBsz1pYevy8vrHDtXT74SWJNPest/UwMTwwRuTJbJAy2y4fq
Zi1BqS05QoymyFdWwrhe12MOxT5IkW1v1HVHW83oobFv2xF//iwQHAH5QuPaMr9HH/3ryOVI0rCs
jmPR/qrAxTrYPbhL+9NPdhI06S68NlyWvfvKA9lLFL6yQM5itczNeeZcTYnbTWH/BsVAbkmNaKlE
GpEbo86jKkpPJeoe0imX0w0a0et1WIWzMNI9th/1UnrGQfPpFciuIDj0c/BBRPM16tB6rtOcFeHJ
87EEk/1jB2pFVB7M2k3X9ul/XOZMxh42FKlMCe9Jen0b5kM/azlqo3+BQ+KjsZlCoMsNxC7zYFXw
nRsPOTF7ivsDOMHXBUruj4nfTywsTzJRb9EsilOeQCHksAEy+03KAHRbhEabeHarTaJBlZtThF89
5alNqSWw4tjqcAZzzMuqnprRdzWREaEVm2OKR/0dhcrq5A2ehnZKL0VoYoQcuuFI/Q84R3IR1sTt
ZfY8iGPHqv5HrKHEF7KYy1sWZOnnTwY8SPxCqF+1FpUeViWlyhY0YoaggfzobqARKgi/Ra3LKTVZ
rIWQcLCLFMR0PMJCydF6VIXXIDuTcttdosm0fuUj1QTVXdX7Ju7xJcqZp4YoFvycAqpoBhnSOJqJ
OcRII2DvnTJ5Sa9Egt5uYF/GyPh5hRE5RrDjsUqXD392EHW8Im+TqVNWdcUk1OARLCU/qNOxj1oX
eDeL3TqT4weXnIvYsHs0KOgw+3VP0pN/8QfWW4ALp4Sa7F8BeicRdcRcqzGlv25IiONnAfX1Evy8
0DQdgPsXuA/V9WKqOXgb5mbGlur6igZkE43n8ci44jWoMFXvLdM0zGBKRHU5n20qVEqgfJ84g834
tm2jWg+QZC0wywy96BLXstwSJCEbfFGUU1vWsSEoeP+4Ro4z5zj7D87XPs/Olsdx6vsHjZs/tYTR
uyazmL/V6/ZlgT6njf5YTvRFCNRK5/2XVJJ8sj17LyTI2BXoVw4sPs1xVGJjckwStF+iDGGMDjso
H99meoo0hyltV9fPGPDC+eZleJJNXs1+QVDplC7qoXp4LISJOB9ebs0YH2v5BlIGQd+g9NmGtUSO
4QkTW/XHh/7xEq2Nt1ULXi6cI9EZcAxYWIIcoWWJ+Gv1NuHe2QXFNdF+g6xvbcVVCQJbQIy1rr0z
RS0/tP7u6uNZV7acsW23J8tJ2fO03lo27UWdejNKRPyVHmcFs4lNbIhQqgsAsrGngKsYgjT1qyAh
b0jmlYdCw6qp/OAg39Cn/7rX0enxfTsworJF4sRzdrwPjYhZ9WFxrAlZ15LmLBEHgjGw2vRF0p3U
6yY+/oIRNtYc4MdvuygJEqW1NtBXAd6Vj89dmXUPBGr3UP386hc7L6RfnhGSfcb2XfNL3tPBq5vd
sxPYYNVL80Y7e6gB84h09sOFf4pMhfjdQayWzhiQ9gDBYwbeBPNvMK3L7r9ypept9lVRrkZp9Emv
ctR+OOr3p0behk1lKOIq/aru4nfCYY37tEMyj1GmDGkJtwGGEnFdmlUKnMSWTbrTLDqIpe+OF3/T
l81ZpLfqkOl5zYo40htjhH9qLaTaDSvtU+GXKY/N0IUXL+cE8naE7f22Fi4fXFpBYUuDfK+dbClA
HeqEHdLQ7smyKcwK9dmJvhd36m7HdkaoUho8zMnHZbzM9GW3AddK6IgwwIrL0tvNEEx8lO17xTfP
EnPXbcPfVsTredkydIEnlMcaPTyZFkHcKa/b3wEKcBF9IejT/8E7SToaqJIChgKyVS8GxNWPW7TA
bycg8T+OGowHw/AwhaDxklcC8PUcsgqQZ5+g0dIlX9dbKOwETdYqtf260N5RgpfrLONb+8LPYxi1
NqW7BNWgZtoq7V6h1/dSo1gLUi2xoYmtXfnG4jkWiqBBGVLexsUjW2rM+7v0m4Ad9kJp3ExIavgF
PpN7WSQCE8vBrDoeCkwFOjvkIFIrCo9FXA7cbBqzra4cAIa/j96AI/lMzzI9sWB4OTbNRkzWscoJ
txgWjMz8QjI9NkZ65349SD4U+K7oCE5edu5oZN2KPc+8+ET8oi4K1GkxhYWXNm1ZYftOzgQ+G9iW
6RvtiPaSiFMvl8zaQU09E13ieVDJUN8yzO6E7vMlS7Ay13ZsqTMv48S8MBjWH5MYeRbtzLxiLb7q
qA9b1mUZtxmGxEv8cdctI8Bf/4//hukSIgprTF89cHgAT1W60T48JxUyyWUX/eONpMRULvjIfg+1
nq9NP9xgHXCYcwYeYUVt9OWeOC4yW9k+K1CDK87mTqQ2kIdZscfuztIc0ljvBzzP5zRFgZWfz2ag
NkFDu/48h51N6Q2mfSfxTQnwAXWxcNTZ348QG7AVoXaapDGEumvlC2/egYqtdOWJRWGEsRuG9nko
LRynbPYfhf2AMKpJ+n4l7oPqKhtrP1hFh3TRoeMkmUtr89C4DNQ/K4yboNu69KnPDl52jpx4ubTr
shroQA05x4zpI/J6MoZP5fuNbdKVqfbWUaUIx3k9wAwI2y06QXhwp3g4oaX85Vg8+2bmTBHjCz1W
VOIP4FefqJ7KASjXZM08MUnOBphDqLHhTuYtLLZRftdx+0dONi3PVW+etFZ8jsGmh7TAFfeL2Gtq
hfSTFRnrniGUx4et3CmLE1r15zY2B3qFZyPCZ15G5fOxviju6BcAlG1DBBaOyN2K27S14WnF+K18
bMr3iKf8iYwcaAaqeTVlBc4iUvbLgor1Huu0KSVW2WRA1FpGShWn+UNgcP/NHz7HtNlYix0iTPo3
JmqC/H7hK2Erut3AO2dVskBE+FzEbXyxFuLKYqJB5dCl8tcfSaLinpDyF2g/xAIJEZQ4UNvEDDxo
Q6T8txSBHAeqGvEO1u7MVZoKj1hUv19tdUy1hp8uAtDfPTnVhD1bE9odeP25a5lx3nz7yvtOVQbX
10jKFWymJHwCDIQdUYlmjDdM/e0/cKc/dOu24eDY92sWXvjVMVYYYfczkllmXbvAeldEyiKt5w98
8IZZdqseKGx8XaYuUB39aJQqU3z05DP6Y1lKB6U73aC267fHiiAlj6Uhg7ODLSsTAGMY2CzxVEQN
fTfXH2zFvBmg+866DrAD3X2NlrK+fHuMmexjF8mIlRd8zkKWTWLdzHnF6CI7taJ7PD+Ly1Ktxp4T
I1x9GMSZ/pIH3meS6L6QLmZASqseX/wosQ02aL4jxy+QbCpz7sdrfw1YDBetkxSgTYMyxKkZV8aZ
5fS98bymdByyVJI12KtGzVJ00z5vgR7k0q4t+MIkYy4Ova1hsvFEpigRqtpWJtwMvaOj4+alsPDr
uCnBqM+A5mWruRlDgZSEar9yE4qhNcz2PgEMx41Q+ixqfrc7zI6vYc5XOdFhPpNCtjp8qf8SLzeE
XvMPUls1llLFf72porZNJw/uSMxbkp/syYWdX6BH77V9YScgqonC1a3K5Qux1AjKcztwFTuyH6un
kVkW1X1M2DRsou4uYusy/xmMLVrn7LEJE0wXQwA53Zvebs0/kNS6APIk35VmfZeJWvHPX45XTsyk
z1woerYS1y76R4ktc/rEt5VtLi+OKczVRi4quHqZYH5+io3Yvd26SBd+WKrcyAhzjg15R1jPjEEZ
uat2+gGhjxawzBfzrj82P6l68trs+pjX1+pmmAzAN2J3xVMyKrlW6fJkUKtxIGDKvcToldoMDk9t
bhCBQ6bKM7eeEZVTk/d9hyTOpFDPwuaG94WE/c0WfMFtK/GWv8v5GMUTKkYSezGm9qN6vTVgIvZx
qW1S4KE820YlkAwjc0/zX54jFT3jFCOUs3/rZCIA1Yend5eMP8Ijiv564djVjBf+nbACU6L/Iyog
pktfMLMSc7SSvkEDLk7IFdbpQwAnqNa31ZdkmIuuRdo9/q5ypIcNKn+/XqMD5OXVOjfM6z581QU1
LL1y/zPl0ObA/imq1sqAhULZNMoh04xiMsUvslhEJDEAUyhNSoSKT/Km83ToU++hX/ldBtr5erGn
dgFbSBhkQLhv8Y2kommRfhRJafbKzMaq5yY13Nuj0NvMSs8X32pSLW574JhV33+cynisBySS3lqC
Yuv/EI0BN6VLbxZkYxOs42dEtbKVXLfchhqtnobexm1m3rgFJviwnoJsUImfGzQIydRVsogbrJAH
7BYgWVSNhODGKsxJikGHyO66tPy3Slg1MWhnEudof038IwNj0+LvCq+5r4Vs0Si4ZyTDZPp6aQl1
X/tfSMisIpLpFNxWja3q0OedzX3h9NlBhZxPh+zcwf0Lq8xIrVL5JSMgzsWIhDt28ZF9EoFOv8hh
chIZscCIzDH8tCUepWPWJVQF00CW2zWPnJSKyxoJ3VhqHMQtaKPyko2srA8nUwBNHuMJuSVlqvYy
BERZcKBB6Jsw99Kzpvygq+2CFXIgb9ubsNNI43ddK30qv90s1401F/9N+5h3aX5uznGm+pW70tPy
LTOVP6pHJ0MHlOl20xSFHfc1htFfdRU/qsKGahL/DsrN6VFg+d5AFt5zb0BF4b6dd6FiXA2c+E0S
++9rXQNNhuYldxUFlhzxiGm1lh75xAwW145FxK9zNefWeGdi4LsEl1rETDV9QcN/8ZDmkWtgKzBr
SlnsQO1tFZCImsgln3UDn1DS1eRI/4VPi4R0CbZcEdZd5pi1vuqWIxunqJb8JKFdrogztp7Lrwkm
YZmlgVKh9uTWE0VOeuMhc5Yt4ePZzzIeyaxBkt29DHSwqmPeX2Lt7baaiTZqYUpmnz4aCMc0eezt
co8fFcZK0TX2b9ROMXsck8OnbryW6qKwiFm/p7fkvgCkiNti7OEb1k5a8A8Nlw5MsqXJPM4enXLp
ia1PHaGvbVxA8hu41vU6YRpOu1NYmoUaPv4pjEURoMBYdmnwAte0b1czHe4YWq3A5TXQiykNS9qC
gLNsIrRKGgW+zg6Wt3RnsyvYpsBTU9Ygyx+DRYRXnPMVPagG2GQBvM9uBd6RU5hGnLIGKfKJteHf
SxQ9XnH/6H7s8qgQuihRjWNECTgp3adnhO8c50PUV7Bbun7WvgWa2vvm4eULQrjcBq0LFsKN1SNu
AG740kdbn5Vf9FC/Vt9dKIQ/nb8dW/mbWUBcWVtBczCMoiDlJTh+AaY6UdU0TlB4rMvL0KPkczJW
m+656hwPD03xshJfrkhtpIiGvk28AZCM9j9WtVWBNhblb/aVGv7mR02XugvEPlhoqeOOfce579jX
ZSdHI0ZoAapCid0jqBrp7UUpe18a4bh7F68EIHaAh57kw9ZqWLqAUeOBIvwc699fGi44F9xtJWM8
WezcZLDWj6MKe/0lkFUuw+w9fmy+1OQ+IAS6wagizvSeJLBHEBzG24mw7Qw+GZst5tzlP5KyDGPt
rTnAoPtnz5fBynzReTvX9E3g606/uY61a1lKXU+/4/fd7eD0gfnIoXuMS5IlZrEQ8TqsW5ZK9M7s
Bdlt+i04KQBNkNBHRA+ruwG1x5L89+B/iSdrIRr4W6ktIy9KUMz+P7bvcm9d21f8I0Bku9TtAPsL
0HJVh6Rw9I0pEsUGR2qTuBolY2dlWYxdVkw2AhPHvpCYkdfZsSMRAUX/2yPUAoa/WjVFBPkaEX9f
x0deZQkw2fceysogtQBVa/174XfJVyX9EjQIuJC6RXSi7i4ygRsUvyZ+RFiY0W4fMGxjVC5EwwHn
70AihGrVCvV7l1sMLx2GiuP80MLeD4s5aURMKZJTs+M5mmzUbSgt88uelWhOc/+J2KRA3e+OJyNn
hNLt5KAP8NMQePz+FCnS62hHLKE+G8+eC3PZxmPknN7BTt0PQS9N3YySxhwLvV+q9qnKwYWo4LAJ
SWco7KUZbMcb3y07Fs+gx95c8NXSSsZbARndZBwcjy8ij8+/yYyd8m2qWUZkr2IY8ASTHIUSuffk
CtQ6XOzOsVbuiDJB08udsehd6Sj1PYK1L+AzHfgg6FMZqMu1RXeBelOSC3RV2c6AFh9d2vK5TVi2
YEI/F375Nud2ANXmbqn7xZ2anzJBYg3Pahu7xg6E++d21PSWzlWqjfRPx1rKW/pvGHyI92dXjYEe
9zJAKwx0CeM5oJOo1QR0H19DyzspmsRWPuKeg7ugqIY945i3YXV1Ca7AgwO9LXJs08yXidh7qMZ5
yqlGDAUBZzHF4/Frou0BgoeOPqxfx/24g2BS0K1CcZsn/CKTgJs/ypSxSKiA20akPHzeZVWXtmm1
coQaXzYw1FKTYgxEtSCb4SmaVPs+0KDU4XFNjSc4CMGYhvZGce2TWxrO2AqFcSRcTg90qOnnXhtE
8iDFPG/V1OUolgg69j/enX4wSkfcR0pInKLGIEMAkRirQ69PND0ZydZvV/TGm8HuQZ5kKCjjQe0T
GLjSunv47tXTvarEaDWSfY5PyoNDk5vLPSQ6z58V+NY9hiJRZ2Ki6oGSj5W6HLCYhsuyZdEF5c1w
+Y0uwGpnbdbt9aW6GZAU3W8twkBKlEMh6Bj44atFWEIU/jamotXyV+lGEMZypSgkCh3g3gdX2cUc
EweCW6YWXs4F1mzbuB5nuoQ3ZM6No7+L9FAph/waqZZos0TMCxngSFfnqb6gDtHva2wcOXV41H5Q
YV5F3tMFYv/drcuvt6qmfX78PV9Ay/CWGVWbXJLo4oTbDUhX8ZuxooOMQK3Wv9si1/U6kkKBYbf1
d+yvB+pc8xqV5V5Sx8KF6rDQC/+a7Z7pIS9FNguz9lAE5efv6QLNlpP+n40Y26O6S+a6QCoVVZ/g
ttf1l6o6Wc3c+1pyTDSV4E12tgPorP4+wSLe3bqVP+5S/3+SDcRBnMcVVJw66WtYHOI72ivGoSKb
ivVg6k0e2EIwR7EqbpUUT2Fs9bYDCdzlbdMOO/S2a9ZoDzM/SB10n4DOyAC39AVhAAQK95g/BZFg
MiHwHNjPeQLMkMrbL064cGHOHYeAc0XDl7lG4SjSCeAchVaAupy0tpj5jOlAXIynr7mHjqJQsGiD
t0EUrbNNqRXvpBAsu6iQPXVLn4624W11CtVWmz7Ly9aSF5NAAqMGt5rRmco27ywaLCLW1oHygNFu
VAN7Ngq3Xit4KcbvDP0hJ4XMCZXrfvbpIo7JMXt3C2P7C5n4oDy11CzcThBnmoMh9X1q1kCaljZ5
vqaVU1IodLW7wqSf+qOAFq2GuSQT+85SLr/aflsvoSex1Q9tMojnvYw7rprPF+J6Ks1FgD0LbV71
Qdgrp6ozbFE1hMDxhGAyrHaEoW3dlzxHw/tcxVQVrY0Ik9Ii/lh8TRFtkgLZQUZNJht6RiqK+/l0
aJyDQpoZLva9oOilE3Jnu8je6PLKglCffG2rnAr+y51KomolVH5REL4t83kY6NH8+5/NZ916Xac7
oxUgLD/5m6T8RoU2DKjw0B1mS9Cohvkb78CdulwyEWUv0FsLvJZ0L/024kMbzNmzcX5yKGv/MqYH
E1ol+zX6RjovhYnCKiYGrIQN7bZrKcE5TmBNPCEe/vmniN5vx1rVIFdIioIfTiPDl/BX5VfDag2B
sfvqv5vq1/lmBbU7vxxkOIaMoioeBOH36sFqPH2vW+/aoqk+V5wqDkCtYSFtfjizMulGzhCCOlHe
RRO7UvuyCDPSA8TdNUdxS86O7uiDLVw5YLHLKMWtJ8RJTbUaqrxAfsh+49/ItgF/3634E8PVHHOC
joC95PngGFZtwnhy2eHrZKytKCtz6bZJgAIqNEYcIlv339D5weCveutI/tfWgzoiXhbmR72dUoM1
NLYw/W278qdIWhSwrr78FHWc7XXWduPTxGjCKJ+OiNsOHBadS6aMGPV2vU9A4pb4vDnRI07nd79C
Q+uZ/XSj0glNpm8toDJcfVebL7pW9n/+QR/MefkAAQb+kIxv1r/XmU++Hxt1PELz+vfeIt3Ky1rf
buw8gVSkKuyv0P67r2RUvolllTQFWV29YvYlM4hzd7iXrTRRIkSkGwuIytiAq5pYwMiQHECamEOA
j4vfiRehKUhrV7aL5DfIDC21qlHFh9bckLiyUvcnpW71K4XG0aCxZM+ZLokpcbKYXShyCf0ilu6/
FbrqgWBAroFO0F+tLtUV6SkAqP/ku8YshGUbFmHEUhzbuHciV3GtYRdLE5WkED50KsmuYBNrrM1T
vOvMLOUCQN/vyKKpLmMxYql9Rs7OKuVHwr1XTkNn9eKJosO5dkusKypXDSOs9f0STvXQHq3cY8Wk
YOhIRnJFnbKOd0OgxYmhXijy5HGMcLlRXmCE6v3Vs8mqs6E7zP81nqsNbZwASEnxRxqI66DbZ8jr
j5pPLKqysdpzdb4HRv9ZuZiYxyyf9+ySuAOsjkRWFymYpKZuDdDmgPREmNMZrXj7zwV0sdL96wlZ
IqUE82e+0chEkCndHeg+vyMJDj6UvRr2YIN0Udtx4z5yE253YniJf26qPAJ7Epot6T2fv3O9DPH6
i6W/SIhrgOzXU8ZpMmTRXaSfK82eq9nyRdKN26E/QmFwWsFkSRWKd3vUy4ThE2NXJUKfDZlkLJq/
gH3zXRbDz5b119Sr3H+9vswTgtBBPmPy15A2PcI+YsRsxFtQauphvxJVlXpfbOpWjzNl/zu7VbEv
9vAAiEyFJLen6B2OaQk2wJKxQfCVERdMhcLEgqLOyVHqoUWbt9CdEdROGDfga3r7y965qdqG6xH3
QP83Dh7TNz+gOQGZAv70u+oKyK84/cxrGiovQWfcKFIbO/iugnUqJx+NOI1OuE3hbaEtTSBPAnPW
FZ7HqhgH9OAJqWFFNKtUwzjc1Os6SM5HlpawfPdXnO71Xcoe8rKw5AwKZa673npkg3hm7TLlU6h+
SKgVlWDqYO95b3xl9audIbtzfgfoCOjfw9pm265SgZZmJRtCPnCjmmNzYWuyQuKs6tLdXByoQfmq
mwkRhw4UkEaawLwK0QDHMlj+m+B42IEwD3CS81ffgXVAqKX/mUrvWcPE0aYd78+fRIuq8ytmbVp3
6Ssh6tnAW66JuP14scW94G4M4fHwSxDRHPzgGOSggere3+UwsoUAEYu4iocEZ0qXn1m5D8sPAVp1
PbL8YRbCkCaO0FM8tnpudJ2ZoViU8XOC41xx+VlXnDspjSCds0wzd7f//qbEgKBst2pUMJ6WT1w7
18c/uYNO1Lu2KnXOuKTki7iJJySrNtoOt1rBzQx1pHrd6wSCJAwG8Uq4ZaXM/2PjZ1dsNQI0kHfT
oSeiQc63flI0gyNIST3XKETMBknEV9bzCNQQzqzkxLO0KsDPxdsMrKO0MegLaEgbCU8F4ZitAmHZ
PqT2rAjFAZPz1z9g+Ynpl4CyNHQWRCf1xHokKo4yXVc7srVO5tNRO8iX2LI1eIRltPPrc2ll47C0
XuxrLngk7aSAlk0V78pPrX6X+Ra2cRp1rrqptFK0CjjQbrVoq97s5+/PdKpf10JcG4XHNZCCNGBt
78F+xu3Vs0PPrEdhIZBo6yT89YhJ7eR3d7wYXGXpo7YeJciVVhujTo/0U23/7jrvmq6ysw779hbB
/9cPYwAzQIC4Os25+Q7i11yRe3z88U8Ix69vUBAXEMzjM8cTW4/J8Ue/n0jNYV+WrVdDXA008L0A
h9G03U+13shIHsyOgmNKxUsayCBjTl4BZCeJ79U10yHuKzsepNR+9d2/CORrBAQJ/mr8iSWJYOU7
jR5bTt3tgl8pz/cxZxuZ1MoczDGaJILQ5Fh5O/4E39Okb/I0oD6jXEfMiqp5wp3lNlrXxkBUflIO
Eiwa6fR+XPC0EDgnWrh3dE3+wZ0jOo6xC5EEt6vFBYLoekdbCfvKoMqS0lD3VqYFFXQZyBj7sT7M
O63mPwt+PB/EFn2YUw8w0kS1t82+/P+PEHadCQqaShGgCMAUnjhUWUwd1u9oVInikyfIELnYXe24
dgiRs8SnhwRaEmXctfynsEP2mz5848Bv2jM8UnG8BomozAOPJh/tg8aADf9Cz/kjwq0nEIfX8n/r
TOOsBIHTbh6CqAlmbdoJ+H1tr9fV4jRfFVBF3zcVgiLl+U6aOfpU9Xiu2cuOmHta6eqxusoO9lIs
9kcllBwzk3jG+AYghANSQNogf4HkIeFLkEgWSTQYLJkdmmWSifVx545sKMYMbJeY8jdqqpzzRDR/
+Fy//8IzRKvNW8CXaxztbgcYU3E6pIdY/983nokKBV6L1/5SLzTd7utFoZYJ31yCy5CJmJkzF7xZ
ZMTdkptQkG+wUjHbf1vxNketJjkVfcHnJCdLop42/miE/gldbvUo+5XKlU6l3FwtZU/LEj3oHUco
nSKQ3fKsB5J2gchkOLZSXW7Ngrp//I7NkZS7pyk+q9putNTNTGZm4EEvwsnXfwMSoAtdq1C3tovA
yjxXL0c4Yu+kPkioecNG03OFIOZd0/kn9jKnbfacXkDyTdBHPcFtLw9u0EPaBJ+RYdP6YZCPsZRd
iwJN2k/ziCtpM22IqMJxZyhvjz+Ql/jcOYXYHCn2dxAaSUzvzrb0RtaUhigL0CoGhTyxyJgnbzS1
oxC1d/HzHVnWECKMDAT01T9DpLGnX5t/wIgaASKCPvWqBXu+CehKqF4K6EjA7nrTLSlyEFX3KtqI
dC9Gs/EpzAr+jqxh3tFi9E053ebrRECIcDHLi/g5XGFgRmZ7d1AYlU4+B0jQv0Nf+gxgWex6+rDW
o2JmGhoFTrMypGMJuMkdh/yyJPtWNc+ofHWwQdNudPMr72iq61/8lS4Nz89BAMqjE0ANUSfkhd68
Ao428fh+IzsWtH461G0ZmHPb/TySS5b+hdbuDnSoZhdp21Ju0MyIGrSGljpnTTOgrSbv81bU/+vc
IXFImYC26Hud70Aj1K1TrybsKS57O1sUVMvw5Lb5mMwYJ601pVEAsng933eMd/HQgtiaK1EfK/jK
HqmkdiBZtV709puks0T8u4vAjZSC8wSzbJIGh8m0arsNoDlHEzTums5ouiQsXk0uwlptKh3tubWk
KSoNT2jOXwGW/HSlqdMcu2Z68W5yHbpy1iW9d25+kV78mljygA1tsrWTXbjSi5YpKOE8t17KNW7+
UaJwxAAFNsn4cCGaAc/LMr7sU98aasjVo7CIvAc1nQoqobq4SK3hkwkd4eZtmoDGd5/LGD1h9zhG
XBrNr4RZAVPZ4f5rwNfpE0QJdmMA9CD1TEK1vbW9PcKWqLRmAQiDGbIDpkPVs6dJjY5X4v8lvNy8
GuZU/SKhDw79eiEZvDghQ7HUZ1FNjWogAxv1Mp58TAuSkWUqL9/3kn0QTOvwMmiBwdrAfVhRtPbH
exGztgaGRxwGJsRloYtZ3ecuVhHR1WhQI+u5Y9F7W4BQ9I6TqXoAm3GFFCBnER49VaI5v6Q+UKWH
8aRha0cixQRf3MJN6r49FA5mZOj+OO5XmWt8vrDcY7Qj5ylytM//PfPAeVAtHPswhYJYJ9h2tcF4
LyKdxOrXb2m7aZUfQ6NPzcv9QZJMnXSFp5GgCoZ0jrIy/riX4j8GIb1186ekXYPj67VJNf9BpE7/
kATcaKvAeT6/xFvyQImDJWfe2B8E9npka+NKh3SNnNe/6XdwY0QkZC+inddMTO9TsE1eehuhpFa2
kZ0QE0mfNkZGx0ZOsfa1sA8advO4GzYzlMp5RhU7mSSNYpkze9NZo8VdV3Q+r63J0Fu7eQthao3e
YZZ3J/thW3B6c/rnZ+gMWdh46986ucqxbYtEguKggBCPP45PRNKB3SymxeRAdECeubN3htapfva6
1CA1+dwpuB0Y3K1aUyXv+fkhdApPqfxrA4iS36j7z4kpTDim7PJzapoCcTrfrZpS29eDnZVYdx1W
V2MA8OQnvD1mSrkCG0J5COeusw2YyM2O+yksA02idVdpVE71E1h241cxdK1s3hyyVBkO65BNka00
YA3FXyVxLoVoS4XMvJS1KnvtKRAY9UQVadQUwoiXq6t3MXnNYnxAOR81IqgbbuU93IAJIPeGlbjo
WQOZaxedE5KaVd4+/QSydxNqxyVD70/KGllfm8HuKHqJhapPWMRzgjzXgZlOyHUyU5vcmsChrjGH
ywcdjfKg4RsC4UjNCd7rBY7VVq8aACfBwB2XqVDTpnd/6deM2iPpuFSxc84E2k9jI5Sk39AMf/4o
b94R2p71ELe1bvzq3KbKwBjSdEjmRpRGRxNW1QBfEAsKIzKXkXKOlJDmvsmZwDQmANHs3eDJlqHo
yUsO7BHhszn7IhFfrM5aYIdthg2jIoj03XBtZP1vakOz6mAgU0165OqZ4Ijgb4fzen1OnD9ZUD8K
VYVcsMl1uHlq8pBTRMZZtXDaBjaradqNgJUcmogv7XjCVIDOELbhsIVomPOXragXvLAjSI+apXcK
lOJpYpJWUtoImJs0tCuLsDfaKNj5lsOoZmCaCO6yL5jMYZR4WYAEmpJ6/Yl+/Wax3xW/xez1lhBl
HRBKY234qmkotVl2IqqB0K0Sp62rOkvUS0yYIBTFzODBpngcoiNwSKzSVgML2yz9x66/XbxqbS3M
xx96kNsM29hO2/NxOivmxFxcqWsUNX+V/9vlE5jMY433zx5o9O0XSonZhETEZVnSeeu5ov/QUaFM
fK+pZ5cqlNdnwi85A5giosCO1+xsXrJcTFeInZwneYDFqm53xSiQrwBYL6VYgeyvicB4z5TLVM+f
S2kL6qi1ZTEKxZt/aKIisEJ+orF1e5jpf09Dqt5m+jxQpaYqdHbczDm7Cs6KjkwdgZ9D5m3PkSww
F3e6GWye97tYwY5CMU8pfj/AMg+hnX9HakmzwHVntc5ZimC89O/lUUP+cDz0O3jtpSULM1AatRyj
5sqnm5z9maH6jWPgLYALniGNoL396sYxNcDWo7i+h2q5Wd3EQ/3Uz3/C1dCdMfEUZh10tPdhizEW
lcGnAnSOot3izjPzttjXinDTAMv1rvq7D/KLnb6jgSeTUVenKs78KUbF5deJXXmVQjy3qjEPCcHP
S3jjlzNttI5wGDt02Ly5j/Efe7PN2ZbPKByuoa2lVKXD7lnYMqNvCtE9DeZ1F6/d7oIC+mY/V+52
s0twoMOlDIVBf/J/DqmJu5LBRL+oOsasFYqZ5SnMIOfxmWCw8DHGaetz6GSmSD6U/CdhbgoWURzH
U8sY6eWJFmN8ONl88ZA3ueFM7KGkY9W5qz+qAvd447Ft/EvDA4BQQzeLNfCNJyCMIFn6EVhRJlxa
Ux34UpCWOu0upSFqbGKap12MGYRJZNiLWRt4Lnj4H5JgPGwafy8zd99Y+//IKjum8Z9NvdvzwHQc
ODFtaNihIA7LviPY3GZgIWtK0LLmwY/blUZFpArQS5ri+x93pk+YKg+RkNteuPtzkH1VGwIjk3/H
XkJ5xn1hgV2SjtcIpZvZPqg6PtL0vVUzUdjEzgVzoPfl6ASmK4uRmsww8EdJnMWoReq+7a9Zh5BZ
alBah4A7GEdNdhQ8l4nq0etguQ3FEFShItCBqZyA4bYJr78FfIuFwVjj/BsifRAMVlOw5oi541gD
tEgeRWX9YD6IHboX06u1QHD1WBC7AMlpqjIiBzn0tKvzfbl83az732OU71ymyvlP0VxirvWOMxKh
WD7cq12e3GArO+ItKjrlTcG4RCiegI0HkejB312A94YP1X+TrrCG9Pw+oy5VRRPNhlXdCxAZ1ETg
CoXZdoaW0ZAeQ4V1vn+jRL6gzQJw2mFwAtKZAPQRIimWGWp8Qaf8wRriims+r/aXe2olV7jAHj0P
BDKoQnV6CZovsfYZcUWtXmHKJcJQmPXV6kcMdMAOwSvxJCm7y2f8NIUicYbh2PA9rwQ8Pm4TtaXO
I2P+m7k010bz20wgFzHMgdI/OkePHObWkQoT1f3MH6a1LhqIW47UP9noUgT3W/ESkvN/jnY3RjGV
oQflixEHPygAEMjS7f2z2CjDCOlXhUHVoRrYQc/lb2Ah6tSkthUG8O9Q0TYnEHeD6gLJ0FBu/O2T
HIqmCKuABnaCHLdE9C/ldZpgdSDgIwfeD8p6T59/d6CJYQhNz4MvKHeb/xkV3PC0DORaUiLWeDTZ
0VdXGIdULgurdZAKP7xdnbh0NcHTZw4/u7VkK/Z7Nw31TlUN+dTyQ6BZj63oR4ANDXie2NOx1Nrz
f4Mkiro8hRIMDHvg0HNxrObOyW0oqHTLncPlPl4MvziJ0u2QkQ7YPJFXQzUdGIru3c5sE+KIHWQI
tdh5V+4bnIRTyFCNF157K/5VhLuNVlXxbY037WpLNWocllvGcn/kLNGaGAIigr6Nwow8RRwlslGR
Qclx4dpfiW6UIwG21Gp96IhDvn3IhLFDx6IogqXBKg41uaK0BXNn4PJYL8zTsYiTPQ/cuUq2PEht
lluXn2vGQUvUwqqj4A6bUiQxNEjnhvfMaicnie8fZXBE2W6uyyvBeGxa9wYRSX8RIaaRSKcmsL1u
X2+LeZVu7+17UBh4gXA1arDfmAdfRfpUcRINSnCx1X4DeW63Nqa8zkHpWZT9QWdhoFboo8zcl4Jx
LreUAYZXxLx1+2blZos//lh0KXs57K8KBisCzEgb+ojXPOfg0hUGMY20mpzbiEC9EKko3jo2GDSv
hwcIBEnzCCg7UmYidYB1iuuyJRqEZaXNfqObDQgoppn63uWMESWcaP8EydPp60EP2wQYDDGTs59m
fhAIUMXLzIWaqqKnIdqVMeACro2m9JI2RK43MvlQ48txoQvmZN5LJB+4vD4xGEuM11cyBSrwA8Cw
f0ar+FmscGL1yPGYcfCbe3kAvD6rCtwNmfbbUPr9MBw2T+EnUyp5BIw48TdoN20nUurHG3S2ZQiJ
cYeRL/4FB5y+pLh31z2LptZet+BnnKYej4lC03ucwFNAD9Lnl8PEbibjCUJHIGi8IpOaR4TGr7SL
Jh6Zm1xIRVOgVd73bf8y6QN0u9SwNWR36hXXPeqfyLgTBJCP5WnU+CsCHGnHhwNaRm46IDC/u4PR
hV5JQQz1xLKoYAbTeljLRAY9PVDnR4sya0lypBxyiFTpiVap+5f1B83MoIGYgB9gknNnoLX6BaP0
EH68BKmDScupJjjQ2wAEWoRfw032fq4ungkmd8dUbgqpwJ6csQ+kjVd/ozfcogos+c2yyNlj83Y/
wjC+x1VraAaJ1Mf5dO+xoCf5sbD8TZxm9c4KyTOAq1N6hzuJkq4n9opd0YxKxUefExV/18i4v0+x
cudjwqaJ7O+NynnawU7ue06lCmQhTDzWaWtk8uszsBfKChpCKAahaeduiVPOTQrGSxBMK7vXTIdr
+KtVXkNc7J2WH7N3FtX7nSpQUDVYXhrdFEZd2NiHDhQn+NMEM2TCOxVTCNCPeTmnZ1ZJwqHz/i6w
Q/8zihSJZymsKQi2jhKLUv17SpUCO8a8j0UhZ+Bkd0LAC0d1vXADsr2h4XmAswpswEZ0i1r3gbga
QK1O+NaVPqyYD7u2QZAcNLGeOhPVgXopB2XYCYpq2Lcbek+kMhdPBIv6xjr2yug58UGTwjn5YwC0
GNf5hBRoiJ+t1SU9TGmW3tvdj6R6urae1gd55yFvhlxDgDcqo3BmJm/7AaXEe+/C1qFFzayBC79C
P82HwYnlQipUdmHof1MNM8u/JRuzfMW2WXMI2JE2DvI5hSVW5IXiI6BbnWI1gHdz5xa2AlcXZWz0
UoOoJCtOUfpSdhUFgpTGrLGrv0Rb31OhIbaXk7dWkhGUWFFVS3S06tiPZ2a/rsvqCxfivUayZBCv
YKW8v567aKxyKzEp1/3+W5sK+1SvluFRe6NGdfXAEBI6lyoWSK2Z/GpQhPz1qtOsoe/nVmG2qPet
Y8l5nv+oRtWyJMXzXVG6aBQcZGtLQrahK/JC4DfD9vJJ5Kiu8zYO+Ms0sNB3hQkgNl6fMl+4kgCJ
D+2RUaWz8y/DpIYxtk+G8VOk2vcVsqxDycSurG907xSEyNx+5MIoN1psxVl4+GSF+gFpsqT3K7Ij
gq6itGzyxPPuIyX4pLJsayw4eHqcWzGiaHqg1G1wkEDBoAbK58j1CIFY1Mk4Nht9+6zWH4tXLbUK
2E6oX3UfxmPr/G0g9+Q/IDNd9aU81AG7ZxLwaW+0o3hOOvpHSq1jfjigIAbbIQ5m75QRPel6bHYs
5UbS7NyU2147z/b/DGqeL4iP5hpDpDpabL5MGfC5kNp+20egIaf9CFXNwqEI7NmB906SLPk2fBeA
KjZHQX2/U1Do2ItzkUdyn9Cu7SagvFSUYYu4WwcuEVEplx8GExkhfHYcEpdy6dJPgD9qgKPcKq9J
mVCVxLyqrEOMPxsIcrKrOPF2TKVgK1QEhgwpbYvPoI4//3f5oLw2qxIln0ovvGFmEth9FZFXcCg7
ezH9NPhdaz28Cbrc2E/3DiUlPV8kClDy4tNAbE5pGL1Y8pByrpOyjqNuKhemt4zQHYFX81v3oUTk
RCf1c78BnZI1m02XZ6jLY25xbfKW9OYkgxj6jcF/snz3DltJMpD7jiHob6MFkcuYdm0cFTKvsik4
Sr7jIFL5o+6snJ8u5iUduxZOf9BE9WkH8q46FKFANVh8JDfTf7qATIM+x2qulb7WVeGy3TKVOwIg
h3yOaZmtSQnaTIn7AOLBSv1zjHou9NCbtdfRKInRYJGBsxFSDSuFUcsJzd5cf01VDHpeIHsTh01n
p+4A1v2pX5ekVvCKxy1RqsHLwPbiQFz6YddLXyB2gZyNVtqSsnkl/tZmJDZ8OkU63+RNQogbsToK
qt81W/X3rv7IjtwP601tihqKp6CSirKWg+RAt/BGW3rQAa24oSzVyPywsIvj61gNwKtrVvLycXOO
ILumk890ssTKiWVTZWrOrNjTmbCTfKZuvpNGR/bqw4nWw7GCzrjynISNSTCyYXb5ZAPRm8DTevAO
6xgUt4sInDT7kzd0JMm0Gtp/GaLrG/MMNd2WpFbbktliqJU77r0E/5apXQDtyHfgiHdsoleLqytP
bc+2653HkhLYIqLRFm3w8rNmgypeBdFZvkz0z6yEimzZ29IN4cZOLKa0KnBH4DQGTMnYtuezRbnW
PwPodMx2pUDy4xuue8GGVsvbVYyy8Uqpnh4LCxRqxx3/R2bkJScTHlAd2kJh4dAf7fasWDYL7lU8
zfhUbuvxNZKfx3JoPfZil7TGYcR9tlXA5yoGw2+orIl/BfqtYvl+Pwi62qK8aNMNFrIygDcPURdt
YPtJTe2/dSuSOwAU5qcWBL/EbQ2wsCic8scsex2mRfzwC1LF7Llv8VJEliq4cb43I32WF+x1OFZU
ONjSk3piGCMb/V3X1DTciDh4dRwF/W+ioPnI7DCXVOQG9YksxE1L/d7QivkEWz8SV1yehnQS6xsk
qilkLg3xhr9uGNe9KTbeO3xVQcRQ37u580XQVoK2m4iEp8T69SW29bTtozvaaqp5rZW1ZY/as/iu
JbX0I9JallRVgWw7FHQ20kuvsMWOw9L9LY3KTYlHDjNCcr2/uJ2ZFZ+J2feeJfAgr9e/NoSybmzP
WB5LuLZBmeFJMTdLbg5QomXcJQFGgIuN+0HCo5yQ7eduwEMIKVGtUIH+lx/0VXKwNDl2ydytR6wX
gh98jzHLDvj60y3Bpq2RJlFhrM550Dvv7gIhiKDo136Nosaqy69HoVtAWvT1vfjLtyfq71BragK5
3wMvUCItG1C1pC7gLgEclknlfUKC6gkF9q6HB23dxsU6SFJXn0zYLgrywBQ94rXpeKrYBjtoxPA8
QSjjamWHLUZBB24uYcB5hIEFVvXqVoGV0IVT+tBjc0B/d/zgoIsYmcctsspcuoz8icFRranhf21k
vLhfOkik0oHsjDVSduLNjeWk/E5Bzyr3GDRpKkfykEpn2Z9YI0yhLeIzCUgDIBmSZPLWH0Vq22V9
rBmkSafiBMYIBJJID2YV4YlUu0jrk9fzNbEdvS8Ys4v1n2HqL4Jd+VwKIQacHC/zRqJfUbFn29y2
6VsGG5e+fqwPLhs/n3QzUoWygqF/qlBGU24qMOpfs9qjzZkO798VVADualoafSXyVQM9RmD1VYhO
KoUx9lojsMa7+LQVmMRLPca0S4tW/0pT5sbaMUOzA1Z23slm+qSiYavfS62+lQbMj732bCWtgZKQ
kVnMx/deQ1dB5J5/i78W+spzd1Xey7Lb0JJXxeAHHY694D9IkuGFgNdkwiw03Lj9Uff4tK8zPNlW
UJ2rEE95VIscR1MiK+cE+asrcsDII4xVAxRWXhzvFdp5pitxO9cbR//R+4+nJhc3b8F/6wlf0Kbo
8O84wk870pTA9UmKZVmyoBebUSKkp4BC8dDNMC1gNl1oKaeab8GdFYYXTU+itOKoc4IplQM0JrDh
xK1yMsOk+zNN68TCidWszDNQh2ptICJEyUnpPxbsgFPG0UVzjZ/X4XipU+Z9prtYqvNPIWhgjOc5
W8DNs4WuxBfgelxVzL+3I56iSiNsaaGWLclltXejBwi3x1apdsRXUE2vXofNKd8yjEMQzQ4PZEM4
oQ65cSplauTsRMXI7fTWQhij/tJU6vnCElKltdS+Zx6+CSq91MA11C+AWRkDKo1FCzEdrEYcJw5P
iXXeTjk+ksTfWyF2p3s+Fei7KSFn53N9sQ169qVTOiKVikeJbn81RBvXDGpxlRt0tv/YbVyBaToS
y6+zRlPWmK/oQs8//apmrwUYA5zRMftUr14fapC/Sz+0tnr/1ZXHCyVUZrX8AcoeKLDWUBmJKxek
kNPOApEIkyDZ06offXvsRudvUbhntPRkNWWuMv2XwEGHX40qABY+dpeEO0wuGI0KY8qfWObMYX1i
/FrFza8414OEnTRNeokim4YY6LTESX36/Ba+xFrKCMbqXfWY3424/0VQ+pxXryaYhvW5iWBl4/ZH
fAGpjPvR1u8aY/g+2VL3jfq8mKSwbL6c9kklXqrFuFBfocIZGWagP0AK6J+49GYCsLhPGRunUG08
a5ShXa+XmCpy5u9u0Xsqm8nd0nLrnZuoqHB3YW4RlEnnuzccobvE2Jj/EUyC3KftwetSNkSpn3q4
9kNgBx2DG7oXtnQ32+P2NNWV4z5PJ13ZG8DOJj/Fy//O6sb3a6ka5Q+wHLnVw3jnZ4L4xzIM0/Y+
977s/u1vjeEH9OTEezRCECpyBr+uYoyVGsRIvznNQZ2Fre2CabGsVEUkarxkDVCSMrDwaWTz2FHc
PlSJyijSpNWfj9OSE/xzo6z0/sQ+iCj1LKhfLfoO2xLqmOGvlVDd/8VT928yQchbfC2S6XzqMOZD
0huglp4vHdYCpIqY+qTXoQIEExZGROv7ZmQxg7mf3HEFsZDo6/1jDhpW+8NBLdI7/FKMoi6C0up1
1tPN90GqlWpNNBIyV9SYjgEMsqttBWeOBU3WRgnFRECp1ZW8HdEjs8pIxnwTlUh3vEdvtK9MZD8w
DmYeMeqBv1oxLfWaXZw790gBa4U03UGKVn9XN/8xWJE/L6SNYLW1F8jr//ffMxQAF+vXtWQhcENT
uFOqODqM9BrnPPXBXCLfhJOgO64KlDzH4AKnQwS1Xog4RGs9R2vhSqhYdknOgQcHWACrxOP0nbY+
21VOVgaBeLm67ZSjeY2wW3eU09VIzkcfv1RDpJCDK8IWnKGw5IZ3TsW/EXXbym3Oos5sscQ+P5DA
3rjGddcIJT0qur09UidGvKcfaV2ZRA5H6HemHZAFlHwQP8wWT+81ETu8i+1sYt42KzYWCstwHtxx
Dj+q3qgi6P/ltDJC/rRpIhRDI0LgH3rdKA4P6wJdxqdKQsIE+drwUQVjrpSAoq/br9ByNnKWoNY3
7/uSKGpl2DaWJBzSqDZ6z8whaW4Myikh/BC5yYeoocFj+QOaH6kuWEnYxDSCYqU5GBFSxy7sy90y
1OjgLdZ1H0ilh/LrniLgon3NCTN5w84NqxX2psnGj0GZ8K3YLpuf+tzqPxmTQwCBnjslFPM+RfiA
21Mj2qs3NyyEtl4lmuwZT1eJ92ZaR2OedrPJc+OLEdVTtlv2UcgZFdwBC0mdVsWHaXFR+QBidvaG
SZ/0/YesaSbj/FMI7mm7D/9EEof4OpxuO7EPRTH5YyEFD0wW0tM+oKdbvmoDiH7ewuY+OFRu10J5
3Ate5UTCESAQYIiBZOElZzHLZVyXd9VM5NbS1qjOAou4XYJDeDbq2s7GTAA0+G7JEl9AwLKQQYYb
MQ84E2meRqT/6+9bT0v1UCvp8rnPzrH+KWbQQalNFN0fZKZL54o+mOFiXGOZ1Yet9zd3WCr8qkyE
AHbNS1Atn2cKGfsqBph3/POqrqqtzQt+cOQDQlOYbJI4wYkzcBUxKg1uQeOV1NMpwJUDMKnrg0Gc
1tL/f5ADCUgrMNw4g6yqaAtYeczn1jN4XJgLHHzQsQfKJT2BQk2hTPPYHR0ydJkKpfKdk1FbvAKN
heQi3uTHKvS1aR3QW6QVtKIoruiYFiQf0pTeNsfjXcrxpzQvR9CnbDF7KH1wZuYm+Ff4lD0PkKcH
xMAqplYwC11bvzW7S4mu45sGrmd+DDmKLWDNiFcWeBDGI1Fo/EEhBcuTVYyiii/eEsxll0Y9SmJO
ki0wQfNhVSXHenPQJKaTK/nmUjrx+iZwyC6LX80olE2e1A5dBQGB+s+L/t/Bkmf78cR9PfKobeyy
5b70SJ4XbJ3ejbw9jt5NJ/IwE91Umfmus803ELg+FnmLg5E9ObZ4OyYM56Ei9arcsrnn+oE8aWW5
+h5dixY7SeDabCyCbv+DpRz53TmO80jhw9Qn5xNd4wsla7/CjMOStjUknfgH0r6Y+PXAQyOfQa+j
fzgUQ1bpDE0UTj+nAhZl1N9jGlU+T3jlJOnbiTUjou2sxpcgNUuMR8am1GPTSOGHRhoVzCQIDzew
30EL9cfYSRXN1tJennVuQdGO08Vlklwe5G5M5sXAijann98b26E6lLdl+ivyRSOwgKqV+mhP3tmJ
lvc+qTq8mGjXCKPfx5EnDXb+YFAzNdKAIOAW9pSMRYS/RqvgVsjfI2vWnUThG+a5d7+px59PzodP
SOMF90EvNqqecIXE5P1vtKigfNPoKx7pVerViazcLpLAKse+kbHgW/Wy/KVnVkqTIwYxj8aWmpFk
lzeqwd581pN5zMJMmjYxmZCx8I3hJ9Fre+KneVXZ9o4/EBUIIogP0pbOR3503u3TTmPDWUJNGphp
RCJ5DztQY6bwyimQ+zG4jTeVwc4L8RKsfr03Pnuie+RSJFzQzHfc0om4SdvemX8D4yUmywgf+ziW
cYKOXAan/IGKylS1FQRN3GVlBku+hrPLLVDxre1zgebZGzzWzpyehd7DHYZPJWRSfqWii/OspdNu
OU4czLQ6knuvpfLumyH1PynWoPIkhxF1cNwkDzdKJQwtsixCaKNwI0EgtROzraL4HSEByt+bYn5Y
gyM95U0B1q8UDZqNNJjrHfpbIvrsrZw+tcO+GOelY2f8yxL5RDmumRid1bAuatUoCImDM1n3TP+z
ipJ+0YYmAa1nbOJYeXkXqpa1rMopTQE24ofQn7Gz9x26eQsxtUdWMlrIuud1k2UBBmhdONfKYJWB
0aKNW3uGTwdIEd9N/1xe4Cf2Tc9VG4Vt5f/FFC6hECFx77O55hPNkz/0kvKjzI7UZFVrgUkUMkji
nSbRT+xc6YHZyTZvP6q/z3fR9x546YXoFdEzKeBSaAUoyL4WzRukiPU3TBL/H13brnDyI3mIv28/
IqBeKXmyeAv02UZo2ygpKMl4Kk9svssCEY+uExacVIQk7yxkl0idzSHzHtEUVv3B/gLSiaheB/6s
Jf5CWuS3m+uSLZSF9xkWgxDA7HRNxY4XCEHG9i9IRB9Z/2jkB5lZ27dNCE77nRKkHxpzOt4BVL1G
5MkCFdDpTBTZP5MwL3dyFFrL0JpTBPvOTHSSQV0fAh6v6cO3t5FadnbMVqxlrPDihKj3XjgNoqn3
OLBmVXbhGJbWA/rJfiSmSzou2MjI+KwgouNBOdIBKQEBHsEFZgcEQCwOSNh1092RUshXKEPSw3FO
YNv2ApHZ4Bu7mBrzC/jIH6DEG5r2Rw9+Dr2glCAYUhgrXdZGDB260JrURzhzOJUb31TPqn7Jxca1
YCzz0Er4HxYn28HsLtPOygPjZUzU9NliOzYxQPpAaSpKX1TeS1h5IMvcQgiOeWO9EfdIqdPhy+Uf
ssLBInwL7tsgnJigT1XpPdOrOFVvVuN3bR5fI3/UW9JfmsP4o7pfo8OClwrmfKHz0/dzbQXqu/s+
LZ7/nlYmf46JH3/IxsApD7/lIpdaxUh1grOWbPOVGmrTgZtkOEVpofmSxL/1Tq+M2+dWOSdzLaPP
vgK7MuWJrOJkex8jEc5Eimpo/zzJqNInoEa3s4A7akXIyIBt+nAVZOPLWW5Ig5MuLOpzqxLp4PfE
79vfo7MpkOJWSZWcnMhN+f/ZOn7+MDDPT6KMLFy3C5boRBesBO82F+gs37+A9qfnGmmRCzPccmRc
Lc4mD/TXN8C/MxlGOsyuSODw4EkdTZ6PgFuxYIf4LkW2KiVSHyr1kPUAOcBYbi6a3+a7tv/VbfXk
qKmkQjxq5UJ8zah+kh76D6v3d2cGFVFo6mkZwNxHMm8hcGCRHfHjjaHH8w9Ea9/zDQkXKiPfbGRT
6gz+GkQZ53ZRQVZ1KM+xlvJsm7Y6JtvmYpIAXzmqVTFtQDmX0lerEN9N8uaOfXBzEKPZNZz5+xP5
qnq+LqPcLEAJ/WFP6cj9syw/m5/1drtVdY83x5xMkYzZnpvC4JTZNf3QQYIpTyi1WNiRrx2nB1zl
LybSINETojcZvLG1VX0ycnvcqRD9osvB6RSI4Yoff3EaCdaBU0Ft4DbOdEEYiPj73GA53Jn+QcGj
NVSu/S1UZqLFd5DyeHME2dxpK9HXKFq7msUCrlkTfK3SM/ENC7IHxZ/LinXnpjXeqGuZYL56SExc
BnnlOXm6KF+jlOx445VfCSga9bRtTYfdpddjK/ZgsUa0POOpc2vI0gyM0V+VEYNE+RC6RONB2N80
C7P4IUDgyCrHmw5x7/SrFVSn40nbX8qLJcivBntDysDZEcakCX/Odtl4XP+8qO08s2++hCWDwtE4
VRbQRnybgnYmatPEVNEfGOd9S6b9C2Rd5EIUbNp46bfEI0nufhZDO0YfcP2OZ5+PrguuUIwvRR2g
q2wR9Rmsw3ROz+vvf0OOwQAHczEsCentD1FNwZnDOAr6F3cI0CVjEMAMvYR+vaqyKiNdZlCiNJeV
d+rCOa4F2dgZy9T15KdHXRn4llWtU7ewgtTJLC+gqS1tNqJnn+u0l1NJLa1xWeJMVbgatJyNmknE
mN7wI/GmqPw1G3jatl2KvbPQ87nXUHdZ28+9ne1E9KZ6ZNHBelWkY5YlvkRBOGnVZwpqXyDV1W34
Q4Gh94btpLN9g1XhnwUm44A0U9dyH5G/KumdEPaeploYURZtJqWTHawAVpg8uAssbXamMoHbyhwI
ljgGYEfQ4YG6Zltv7zLef0ziUaHIxfdXpE62Gnq3JA+xe3EEJaQo1zyPwiVZCoU8QHtLjdNtHT2s
vXn+yNe8sVqofx0qOTy5ElKwXCjTBEV76t33eMKLVfMb05Auc1ghnkI6tlszz43omY49+QupkwwI
oJIImVKvlSzF6YtOO/Rcbhq++fCKwGi2ksChOAKIZbIvidFbrc5fSr+8PpD8i7ms5V/90sPoxvDf
mjml7le786UVEDJUfe/nHx59++UVGmyCN3EEl2Q9MRfsGGky+bviJVl+28ZA67YE9s8gBifzL1bg
BR4fRvybRHzsKXiV/OAy8MYE1pdeoJbyLXMBd8rJe79DhszK6I5Fzkeq+0eswwy9YjrEkTG2p0Rs
A3uKYLzC5qyukIAyCojSdGMEW9HYSV/3LtFBt12OrLNn4bT+MT1XqPYI4Kq7nQHOYZucJye35iGs
nQLNxc6OzT4+OH0eYKLTeqFvHMNYgcEKEbPPcckgSFv/kFbcJkuGYoi3ZlRCHIpAuV7AzEh2fhPE
xa8dhpMCOCwsIjNWrlM4rKulLeRxtDjdShuBmrJsrG9qN3b0y/0wfUf5Twu1GgANHXObjF7KvjGp
Be+LX2cD2MwfojvbBMHEeh55u3Nu6/6PQm+L3YxBMU+pe2dJJkBotW5dxsl6iaQdha0A5CaVLAvT
evyLtHOvyJhYoiIGBVYvV815l4una4OYqD9mF6szYK8IApEo4750nyI/cL05s3XKeUdpZGt1r1N0
N+WqArWWcJdRgZYJHeGEh3A70v/NdL6hEyvXdoG+utd+IVg0QjBz+8lJq9VYR+DORfOy+bQObCGA
Vahdgx5Y+xHdczPSTzqc2zrkmdJ9Rv7LK4SWA4ptHbxTPArsme8/Wq0S8dGsMq+d1smwTV9iZ9Yk
Cawxj5x6jto/sSJKjWBFHLUGKtJe/qTb5+PftJBCG1fW1OXaxC1ci4KKQN2Wy0HA/0NpCyUU/a3x
cDdueLtr0vAd4CrTIqYiHY/Xk1BDlPyCnS55o0pKhhQUNlZOCdVqRrPhbEh+GxSlhUJncU1SV9mK
lap6M+15SeJHPGjqQUtAt5jUU8BvOaci/JYt/aD3HAjaaiditYe8IezhTu4tIfGhcqX5Pmq1+tBq
eIW1iJDYatzyHmNsdNXwp/He8fOz13vXkV17AnhhrxU7jjacVgzgpnmBT2PJpc9jQrpBqdUueb+e
CckO2QBmxO8spr3v95Z5XqvPZZP5Z41ql7oktxz4x5PolBhZo0dhTl527YA6Y0Qs6YRtaCUMg3xm
K4SEIDz+1bEW+0nc/R6AZfvYQCiKV/f8r5w6TDyE6KQIPQJLsstNErxpwCX4+fGl77UWnra6gHAo
MEIMCzosdnGGPq4zviGxGwI1aSYTF0G0kjNWm4GgrTZJhWoMQwuI4j0MxyFyPDRjidsBJsq72vzX
HMpZSeIC/4fXHshKbkknWCTRYr3g4Hk9uEnwcC0ALgz0mHkxZ0IYgUuJNx9F1L8b8YpxP76BNV/a
CNve7DC9vQRaSYpMlrVIcVCUrDkDc4/Qg3EvohRSrEfn7/8ZuaXsGsqWkFQUZ+iBZD2p7+ILoY1w
qtGBPZK4k1wsn0Wvs8ya+On6LCZRgXYDbnOfKQ8T+HPkMGuCzm6ixjJp906l3vAtcPZA9IhESb9n
bnuSFPzY4PtWU6ZjumLJeDVv2DTN8HXeh938WlOSWR1EmMo+cK7qVo86YoqF70GyZwSM61Tzt4Lg
oXReFcgrMW5htWwfaVs9ouuxqLmC7qhmLQiNMJhQteVvX0ZNusZ9O6PdaEBY5HNpOxemqMRUVWoL
JEM+W20dBMV0kSHMlst/YW8sQC5v/HizSGAOJmXQHqR5ldOh1b4uNVrS8m6sB99WNIWgHXkgRPTa
GdfpNE6iscnsc2Wkq+k1YZHnOtp9L5lLdBQmO+AGIuLd5YhRnQZIKGb6hztG/eXNGou0Wrxqvij0
zpBEr57jtNMaIpgeLAAkfW+t1hJPMASBgdug5sp+exSYptqVVhMo+qgDi1e6E6JTztWRARqgDKbN
BLDGlBMBV0nUHm4i8F4hNHT+7Gh8x0/rpjCqU3KaT1vU7YVU/7fnhoPx5ccfFhAoRt+7UPaYuuZ9
/P5d3C4MiAuoXHV79oEX61M4Z3tueSH1aoNFKtrgn1WxAdPo9WSxDCV/sJDLyi1wSP2FeNGFGpai
qCsYh7JH+6P+Ie7ZxfQlC0vmTNVROTYPQdHF4nCnG8r/GrXPe0Cp+6UZghs6+RRJL8UFlV0J6rC7
+8lMWyieTXG2dZaGWPihrB5pVIMV/e+OpGVx4cAssbkIPrZn3/AhmtJv4En6rRr40SJerzzig8TY
cQ3Dsv/gMc57rEt8JFKgYlxexpG1C+wfeVffk6QH7AfNNvcItS+aMPZP3MB1YRc0j+3qI7zuwuoY
eZ4nwR41z8NtjOZoV27SEL0mWsSRXv2wdM/sthRpfR6vo4x7+FSVqvKalzckAFZwzfDgoi/dLTa8
PDM5NGUGns74mP+gB2gdBUihEoPzhU8Cl1gNt9iz/YvlQ6M2i/EIPi/iZ4jNVbkqOZfXPwRf4he3
cYUimu3LsSgrgd5UUPcB3DPI+x5gWEL3MPmj4XXoggOUdCLLjUZkUMGLd8+AfqFI9sLxMYIzx/+g
OZ4XhhfHqqBKUk2/7mvOi956k+KtNclR4R+yBmcxwfsemhKPZ2eQJbISgbj9V/jJ7mWMIsEOIVFH
/85fPzbXdZK/0MNpTc2GbijKxp8vzwnYwqCi7MRpB7iRvsWpEnVXiaeQHN1x0IiKOqTHblr4ppnk
5y1bLCUmcPrLYLxkGfPUfmevsMoBty1T+bFX7d53vDUnfx+Tw9fnfZfUvX34RmhWIibRh580iH7x
Nml5wQRi0mhzwoD4UvV6iGE7jRWxQadWdfTl1I+zUqLVK9ju+hRs99CkV5cqB8ob8ixAJ4pthGBq
Ra04g9qjgyOy2IFdhKoBTPqoj82f35SGBPsbEy3l9TRojhFLkdUM/H4QXz4ZyWsPmggrHH1fEQ6Q
chpxRVRP/Pm7b91DYJcRQU3OL7PuSVBVkoqwao9G9u2UtC9et6t1whPzFxmfia1YLkrsCWyR9QuL
0ASBPjiCiTzCNklBzm1lYUmXWnMO6wbqNTILTZZUqDuSOTR4JD8EWXWuoOE/yPyzwIzZfzuxOsGl
hShit1IQeK7vAxOVQmTa0SsjLigcrDJcwZAuT/LCU84DdI01PKxRk/p9qDr2lR2V0jBY90tjyay2
yLI8Vw9WygM64ts1ge+ObLBjz73KNqWt1pKOa++ziUZNKAGuT+Akh06oLtm709/bDbir+ofErLfP
p7xXjrckwbarZhTlzEiBK4hq9GuzIIqFliR7I/VFtF4wf9Zhpv3nxK/9AVFKuzBrIdkfX6rfpeJq
DQ7BarRVmjW1it8KtWl8jfjq9IWR8mZFIi3IlfNuXJzr2rB83RCWazrQ9eVJG6EG5/3roiso6PhM
OD0UQc9LFRXFqcxhlPiIZCnATguL2MkjjfNDGDFRxy7Qha/fkQ9VKikjYRmU6lFlIWM30Dnq03B6
Oyj7oI2Hbq9K+kMZyzn9utXX2F/5fsAivX69OPGKU59Zy7B20EEwUwofVPKJdEYPzKA2BgKXAZrb
KEFfX6iSCMS3hAAakRsSRwW0CApgTiebkc4wUTgRQn+Jlfz9QAGJe99hBMBfVDxqFrrGRSAHf4o0
kJ7hz8lzMwdpFDsOKegXNFYWPCRBj7e5oLcrvE9zxE333+lOIK8Z+TtYOUr3fHKpiWw3dPCULvYD
zyto/jIHQOrShBKu0nrefqkQmTq7I9HyUJqPiHgghgoCqcX4wbCmQizOxtxIQhUJMTylhWOfx0jz
GUVvUO0ExmKUKPqGjsA6UdLiWSXoWo+/oaLqz8comixNq/O400xeMGlYulUGrQ1E6LPRwENfcq7F
wpv9EhxqyhAdTL1mSjbFD3r+8pD9yVuXYGJGDgfUWgI/qJdnOpzh/BMckI05Tb+MCumabWHsm7bp
LP2O2riOaIarNXd6FqZEfrY842lkpJMENaJg46v4eh2m0J+rF68cDip2d+xjihrj3C4j+iN5//qy
mYn9SfMz6f8DhBQ5VUCpn+MDGl8tpm3WRg61Qk2c2G1bJTNM8EWz48q23Lf05LdCLssbNDWJhs0m
yiVW3wV9bmNm2S9tgSXHHAGm0pSz+btvjo47EdbPTuGK8o2NGy5obV4vMdotGI62l0k6iqJexA4t
9AzK9Wkhic2x/Y+ga4NsFPcXR6s+/E2qljZfYNWuGNn1xNAciLOzvUgO3+wLl3axd2VeE9dVrIKP
nZzjoRWbLlajPy4jjWI9NM/8/oO3YuB2ASSjdbO9m96LdhEO3N8Uj2Zaf9nORKTZfKln4xMdYKH/
mUP1/uAKLBpVpxb1e82I3a7HlSAxknxi/1/gvPc+pXVOeZ4RI06OHzvqKIl9u+XIyIXfRBkJ9HRi
S+Rjxhvj43VLZXDk36PCUMPnudrF5Z6dILZngqiml7j3yUKfUdwtPEX+NSxNP+uyvO9qFAARqUbb
mZTVX7N4n5/VefSVzIA6C0ZUSKsqMxFNt69RoG/qvsi/0Kf3WRQVxfPn6biOMIsALXfcUNS11GT6
cSPaLsXqmh/eYVeTGQ56mSiwwQK6QODcoU/LcML8wbdq0XjbYJASWr07U6bOe2Cf+I0komW1hxmu
BxT4rFxMk2mOyh94GWh0g2qhdO1Rx4GUELwLkorFzI5tXHEjxvmxyzufHXvvHYuLmuBsnkg/+r+7
mUigfISABu5Q5NpJU28/S0jT5w7ebQpVB9sHAJ5ZOej4DcCXn2EIeSSdkHUgG/Xs+o0Nd2Dg6zP/
s0yTW/A3FWNtokEuRuhfO2fFqxYOheHT5rQ+jR/87dpAxWspIA1KXWnPXtjznaTYMIaW23Dyl8Xb
UhUH0B+bINWZrFbn9hnllVnePvklpWTFQ5Qmd5US9oXN9c5eUAVNTONVugld/shuSGqfEzXMdPPo
WL9XCKdJ+kCg43GqPvsZwqGcIdazupIyNXcSSMLFgL2ZkP1ADf0lHQwMg0itv0ouL4TA5hUnQn8r
9iFAxHX4UExCBmzp1w+tH23dJc1VKhXnulGsBXrB1uaPymwrpJ0L9BAKYOziSOLVA99bFmxqlsZG
m3Lkr3gC4txMZLHnEQoeLgS8mj4ZYhuHFpbQfe61cs3Mhktns3kJ+Jn+wdp3yHv1ROg1g177Ib9n
EuKyvNioRTKvDs9SoYsh4q4OlGm8rM29qf/Sg2KfeOa4SoCiCvrpFVDH90aKfNjPlcwAyyxcGGWn
7WTxaeeyKRoZ2PzUEGeVQCBjwaDYwB4dbNQh98YmYbjz7sLoJkWgvJ6Ay85MXfilqgZ79jhBakcc
lfgcvywJIiM+4v5OuDdYxFjYd6jtImfS+LLnEL9rt0DRIeoxUpvKJ93FfNRpMr7ZwGh9kr9hcjNr
flr55gl8LKiK80anmeUaWNTRfIE/7X4emaGdGS9ZBdTmDm80YuiAVmkltcCIoUE2CBv8K/f+xrEv
mOpF96w6AsC7xnf4Ww9Rx5vXAxoB7DbUpB9GrV5cjLb5PgQDJV+//KCgFvy2ZrFXTnmnfmGwtV6D
FPzMKrBeBXtRlM0WempsTRua6P++7fM0a5xbzAqQX9t/qmX+lIXZJbRpcSJWq3jBhUxEsMtkbuG0
3goarwGtI59QK86AGq+Y8BmV5/RwOmBqj8Co/X0/8doK0CF0Lt0klDUu2UD98a5TDD/813crm4pF
lU8dmcEl4B0REYMpjBG5bex/vO/dN1HU4Uc0Y4t0HqDeTsTqOZ+XqD3OtDzj9W0p8/YxjgqclpEf
fGsVhToBhZxPeUsTNZJWnXUDY5u2/5CdnfikaXW4ZC3K+g87mL+duP7GaRsVXEUjtPFO1i2ZWeV3
vfEzBocib09g3devrQxCzjFaeZ7BMphS2FsKlt4s+Bb9mI+uIqksDbL/Da9KUcH050yiL6B8WnHm
5dBFevG/eOA9u6sw5Glv8nHqwM+KbzFDq+xkqqCO8wlhvqr9ay7N02MusHraKob1vt/7fR3IFf2R
a816iadkXSSEYZf66KGp7+ED0fYDI8WZO7likrgGXmc0WTu8PuHgbR6e9B7F+E8TjSLQYEVHliY+
6baM8KrBz4RtuuhcYGE8LydhQsNhyGi+FCEmeyhbJJvtHNVwDpwZhftsYPiAyBZAIb4m+98c3w31
GxtWV9vmlePN7E84uyZrBtTmfgTpINWTCsHas5K+Pp2xXRee3IMub2KX0qZ19knCRs5CE3aZIeZ2
t7ACBQXb21hGLcQ15dR8wgDMv5cENGIOpTLTVXaJYlEQCQMvXgUQfBA/L9sPaA6Lig29c2f17Hkj
eoaAZ++IM/KyHSDBnmCh4/xS2OOqPJDgeCVxHJTDhZ/73w6X8xeTUjaN8/tI9ZlwdGKIHmoKuK/l
+gUzNmtFqq5qTS33BnVQkLDT/aKcC/rh5hg1Z9f4VxD/PE4aij13PvaWOOGBcO07Kld4Drq5fPHD
pjk6pGMpiKgq052t8kGKjxxKJE3ZX4uw+pTt/7+jrb5JimtguDYwtaOQe6wxEQ3ztiOGjjKbWPKl
xOw4hfQeoU1kq59XvlUBUt62E/Xzg8e9kMQwWSv2UVp+6zn78ygVmHJVrOl0JUSbwAIm5AMB2ReU
vpVxXzMoFUPch/vK8GHNyVqzNB5rEhDtx8JDQrOABWaH/y8qJcoVYJkCuaCMDDck/9wFb2/4o2i7
FiYovxR3uGApQXb8KffiijGXmJPgv2Y6N6/QV39TcfHwKiC0oawe3A39VlvDZCDh2h4+7yqPPJHR
8V5Rz6RVFnfrEEs2teXuvBQt8so2xjvWPHRYsIa5cupQ2vFEiLFaISApLE+U4woJlFxtBiU0jDHu
9nM64RagaWeoPInX0LPrwSHrNNt4PQjuTz9WEEu83G3TbFtsvGazs6UhQ6CPa3PWQfqAWz0FfGle
fjO/pwYS5o66slLqHSSI/CX1pnVtYj/C45W4sL3eDlpay6hhQgf5crw0Awg8JewjQ0uCkGRA3kOi
6N2vzlPlr4wWBFZFD6S8AM4sytP6rBscYIK/qrXsrc/J8F1cg7m88T9wmNA7EyNQTgIfJQOgQFzD
d9FJfkX2FHrVrSr9Jq6Kg5OqdSUdiJ/4LZHOLGCm58p3G42y9S14yGInUsMUpc7uygoQQRbpbiWJ
BphL41WFhBH1RuuKhYPtxHuQpoSOnoy7VjQTM0FL8Yz/SulYJ17gEq/XcjIfZSyDHWyuJf/PDlEm
pAjADaRlxRqtMi872twK5en6Ulnvdy28ZMJKHzzy3fUnTAFGcr7+SY0UD+Fs51sB3R+gmhxp8wh/
jUx9oz7o/hHKnHShi9UMN99sm1q0unoIBuaWfnFsJrt/hMEQ8XGONJ3PV+IelDYovgOgLkUJ/i8a
2Q3vKRNtEN/d8QZnhFJINKvvM1uF0p/s85Lq9RA5UUS1iu0RApqVJWK/2elSqPMysLCbqDyVp4Jk
aXupEq/50YGoM08roy2fzyv1bVDeCW+nlSIy7nhxKJvbuD0hQ7Ojm9slBmMsG9dZ50uxmD6JEYlO
iNWws8pk7BO2ZiaXaZ0WLv+7IBZvjIYGnERpg1G+30rbM2kajscVfYJgyyMP/UiyX71XmLoaHvhj
Q51wmngOzWwP38FI7bVbde3SktpabSxJZl4H4/nvCKfHzRrXBHDTrutvPRLCQ8wB4FATIP3QrSgD
Mf0z9bHlvgghM/VNfUAZQKyRPBaC1uRucrSVW3vSn3BtwSWnj7qBNlcwXFZFItzCObu4E2QYUrzQ
YdXsDI+CHSUgBO8rDGl4QGb9E4eMq9W/IuS5oEnIqjPNfVSQcen+75onXZIUcHiM51L/I8WmdXeZ
2wJlf3hD/d4VbhzG54Q5gGiYJKc1O67AUHQU+hyT5FJcVHgPpQn0kXrD7JeHBnwwzRqT6uhBN7iV
0O2Wsccpn87i2h9EngCgSYMdqt/8ZyzzOa/Vp2ZY54CCqpYfwZ3ZU5kS+x290bJx5kH8IwiUbQq8
/VVBSROzOflsTaGGwy54n3ELPUDfHFpHRwKyoQQ//bn2GjGld++iKaI0iSmLBpAodXjURZTToC0y
rFGd0kYh7wJe4JL0AGP4dHzzvyIH1GpEVuKNYQ1oG0sH9XDiV/Ngju9B5WTfDEaYkWFGdn9M5lLp
Jupfik9muVLse15zemu+vr6KqsYkjrLxdTmaEgzA1IiCagyMYiNJ0WPHXfPuwzmyCvDpTTB4Ezhy
hyMBvhGxC2haTCoe22gl1C/db63PcETkchrCd7kvSp1xucmhdXcobKBdKLDy0et8io0/yL4U6CNF
kkqh4dBLoIx2gMzv2CCEn+WEzmmHxdXeoDyVpw0pCh+ej7bnMZcozse57LCglMN6vHMkWtgBYA5V
ZS3dpNzssWj4Y/a90x6wjo4HgRXegBoKq50NUsMuf2KbJXkgJRgiau2e0FrFjc97vMRX+FPl2Nax
bdw8RtJtahqJgMUIASHe0b/K2nkn1+apAHYozzGQIii0wjg7wsQHEhdwEQczTxC307K2skAxPk9y
Z3TRifEqiDtkPTBpX1pgck4tDReS8+1sQKpJ0IuMKnp1YwqhAEld/JB/Yc6oI9PcYVJ8VofzC4xf
N1JdQw8WZcecqXUURPz9Su530YngOGiomj9+fPRrKMGtsBf7nEB0+THRuGYBe2PPZOK11KvAAfPN
5NJHx20RBqztEGgtEEfuWI2dF+Ki7E+KRJ+3NqQKJVkrJ7GM4XIxjo4P2Qpkkfxj4wO978WhQmgk
4xASu7MKFGgSWQ4xRLO9G4VirDxWRhlEq04GNeFE3YK3lGMqz4Dlx8qUT+6+Pn3FNOjq2JiuRTi+
cCfSFBfBXMEkwEIACnLPfuhvwapkU05j/gbx4ungofdUpvURkNSvGV/G57blL2t2kcPoPcyhgI/R
6oqeLeht08u2et7aljDzPlJgvh/UmW/nP0KODiA93fKEESZ+l4IOzNiW0KMeU+54BfMKN13LlCnH
+n6UzH+d9YQEn4eKLscXIQJJ+fQe6KwQH2VughpLXnzw+nlZsGUhjDPDWTjgOOHO4Li5DSBeeqDS
CDEyrbuyVsbou3nAtrJi87vdQxWeDGLFlvFUmBDaEjod4C98npjrj8pvwCWAl5nGJFBuD854TRnG
EdwXFMETWWd3XX7S0Heath2T/mMG/kDdR48yVniVnoagTqbUB0o8iw2uea1EVmHO28y3QdJ2k0v+
7jDlYD1C9loiuIHGQax9dKAVYk97TxWWX2+smHYRCRxMWZ/4G2NCN0T90v6z/QBm6RaCfUuy6wA9
iAwVJMjeW5flWoUfv+6Qg86/WWBBLKeYjc/b6Q398YZ8r4SAbC+LLXsWOz2qYKI5RBTAn4aJK8q5
5bhfISHQz43TPgGewd/mSzPiLpe705f8QtROJgg/QqCFDzL5D1ccptQe2uhAEM8hsZpO60gZ23ax
gx+mr7l5clsAG0Ysxl8vOoGlvwezV250ywtqvR17pAA4tW7cjkpNhqzdQlMnbTHBhAxekQ12ONSi
+o4EC5sCG78Y1Cz4uxFYbJeVW8Jwx9olrtVhn9Ldpcf/uKVng0TMJIO5p7SZfO2N8YVSj/Vuk/ka
5tV34wtNoYjrWi65u+zrB29tJ1TdZsFVJkd4/rKzyEMlvUVPxwR2FzE8QV4uHGkwPPK3r16GFFWo
+mYLsLLJCLPf0/uv2R0dsw6bO3jsIFTmPaxJ3bpgM0x2K5YOZ81nYLChjdp1eUGhlkqij6nk7V+3
ud22Qc5Mrg84A4Be9YQBE5YEwj3dZRNcgPSe+CbgtW9VSATncsAtT9b3uu4ZhDLhH//KFXPAFSIs
bazZpbNFFPHBvYHGc1FxxE0ZkHoavgX6Ng3zXUh6vPo0L+/f4Pbhpeu4Ba3Q7dRUHw5162vgNqvg
60Q0cH0f47r8lGbSQ0dADf3s+lf8d+ud4G/TKH9jjS7Qm6jBYGM//KJH1hfb0ObCX5ohqrA6ZU4B
ua9aCpUP3lMhVKYfHS8gwi/9OcR/8ptRcSzFmplyMwKbbyHRe9xwUJw2DrAzpP66gfvhTovHbRHh
RygGwfb45mMPUXHeghbKndQg9PuX7GuxLacBvzb/OZzMCTk9WY+1a7+j/ThfM9y+h+J2b1oCIWKR
vc5ifdjcHE5ypmQ6TY/Yhw2LLQ791mTzITXK4SfRrAXeCgUFgG+iUtG02LXfU2jWTFsL7Db5rpkU
g14+aJxPhGwGppOocT3DhT3ekT9DkwstqkK+jPj4S6kj9Uwzf5NqOkrKjb5P5cEy3B11U1hMyIhk
WGBYosDJguozxrYbX8q+JSfx9EEyN4C3Fy9scCCvUpGkzVartKryQyMBmVhYLpf0rIUh3c3VVZ24
pR+uKNzm7GSaeJ/Xrne6pjQjYPCSvNn5kGj4eeplQVkQSseFlckk7poLwcjpBTrAiZHxXM2j8LWn
Q91gsiWQyRWoib1QFxqNDk2FPAgMOWxLqVflAd2Y+NVOJJaAhT9xo1tqTH0BW++JblGvblhWCk2n
1ucmCWFffu/flI4EvE6l2lg3AhQI9kZVw6JCYt3375kqZ38WxLpRM3w8u0ZIKlNRaAlC2Ym8sYiK
KlJkm6I/EDanCeyCZAxoQDOcUSVEa84eqC1wZkmomQtv3Pt4ZroqWAO7IXusvb+1kgpZmplenDWs
5q2JLeUDRKTFcKo9HgnvJM4sr65njFSz4t9FGrrEKRxsb9259NOELzVKPJMNWqtJoNHll/Y2BFjI
mqGTQvuMkGhpO/rg7nXe2fQNiYxBVjSTeh9oZVtCPWqL/kYZB60DN26DUb/yBqOmVeN1ZiOvXa+K
mRgkWJBQ++cgCs6OTywkjARp5t5yh6TSgNGXj9spKbHDwOPn6HmvulzkN2EiXX5+EuME/cVsMBrZ
XACvJ4oNBAvJSt/1rFnlH1kQn39NbVwE/G69QXLsacPej4b3PAYzlImG1NHuY5vtsbkicDD2bp3s
eulX3n0lEevOTZY783MAVT+BWc7ZmnifT2LdtJgzkkYYvb44VlIyuNcA+cfDgXfkLTOTRchjBB7+
wYigbZly2acQvX/57Rh3yisTJprxfjYX0ZeMjrBTaNkIiOFPfZBZQyeTUDImDdBQF47P1TiRWGxD
fG56o9r4FJMb6EjxhlaJREr3Q248DVTtP/SikEf/h+PteI1I2psHcalieP+Bydey/rv4FP+F7kwE
47MtdHr0m2l+rzbcY06eD+TYYFtiYJw5jeKhOMEjya9Z2xWGchgrxcLvCw759NBMcZsgqvKn6o1S
e4PxUPs4WMg5Mlgfruv66K8M1/ZnudumlkhM7qon8JL6QVeKttkZqLIiR8mVch/DUJyJL0jE6WY1
DKv9ltdx0O7vZOl3lfmElw/Qrew8Ut8UWYU0q4zKJonnX/wkPtxYkcs+dEyfqr2Vh752PI7c+U4b
3oNhJLH8zZmTW7S/HYasScB8R6CF4cx897oX2KPix7ocrkKlZuy0tc8IvmoNIScel32IuFcAOVpR
7vovP0t38hmpxDHFYG6WWhSLXFIfiEL8boDKaP7PjP6gydxHHMd4qgI7cj9uu5VeFiQ42ZZPEbvw
4CLz6L/GkhqMSTcJVbWvL/dP8YmbUWJ5gP/JUFovzkQUVJAOGq1wTZWfdroqJ7qRdzR8foCPS/Mx
DawO3RcbwMWF5DHlv/bglV7XD8P3wzfCUcdJsnRqXXqFgDjMoXdLt4PAR3x9nxcxn200uwRUxsos
nY04OmcB6TnpF5ZxL0ofv81C0qdXur0qpGQGiRz1z9RCdBy5Vl50FxizMep/s9N+pwlF1EOOTqzb
pdTeIH293o2B+BkKvbNIgU1SO4SPuV45fNrcNq+OxhGcpDV1MwZBGUaxG3sSzqS+sXicAmNu9Amh
p5pWawJzFT57DHVgySvg3cotOmSS94PbUe9ZNaMfmUW4Sg0Sh7O5HtSso2/i7rguVokPkVqVRSso
vhhy/8PwE2+QjAvX90XVA6NBlO7kjGy/7Fk71baxIlgYjxNV6X8GU5Rm2GhUwNBM+Jt8XEQt1UrI
U2MtwhjK1AMb79Ta4oj7B6ZmA0c2OjOGxVPDdBXl8hHSUeRjvzzufEEJSbF7NGSoWIlxu+sNiCfs
gU+K+unGtuc6ZenaJBsq5rgIBUyrvgq5NWEEsSXetejLKpgWwXqwLYWMr2mOGF1RhGHnQqE991K2
xUKZkYYID/L1ZImd+wkAu8klNuFrDf5cK1IMqLIKx20RRNS/fzLAVzBppefskwHTz4mb9magpvpU
KIy/fAAenvec3ci5uNTBPoGEawov2M+arzqOGpB/gZ3nzL6zrvV1yBQ9I2TjOX3X6vb3iCKJDSlA
0XPz2pugDfUg7q/H0/kCxZ3utFiTDw40+X+qhkV09fCJ/EzDMhrZthPVzAbbtkeBMwusUw5XNLuA
BNiaJNAitgBOemKvfX7FWLQ9EOGJBfAhenjr5LQ9x9G1y0aK3bVauHKUSMeW+P1DoUSvjXjs4FmH
TCQW4OunacF7SfAc3XpCkrmI1m/bA/CbjsE+NWNtzrlD+D8l3S6HMCU4PEbM+bUK4UJgqB89tv2o
XLWhK5NC+WFKLITSrZsbIxyHU39uJbvDX7ZSQM+nPlmf0JXYRPkHAR9nIzqecsjCDNuXe8fAOYkN
OBTIlQbWxrF1vtJJVtWGxg/7jtgilX/9eU/lJOUBpOffJlFVvoKRkHRT3ZFTfjOPPfZdMOu/O+DJ
jfvblF5lPUsmLwQaNw/25dDq6gfG3XQXFXZWjEfZ8Nyo7k1fXHBjv5PXGU5Te6NdWbP2tGj6DUQQ
zcpnEoKuUpB55aLwBxv9wyj8D9U8D4LmARkXWn3YzOs0urx5+EJa48YfIizOryEHfKp8ZBpfOfsT
HtSVboDDFFOegorUzqkLKFLrNNbAyU6aUaOp1MOWUg/jCNhVuY+eU6O+ux5rzNnr/Am5XwkdbBPH
8+EMdWn56BAA5WhCkzsSujtj4M4HEdE6yraUjQDvWFPF5jbu8ve/e0xbkqO/MjYQbFcOlZayfAWS
i4Vm538lTUBMW+8l62YD+mR+rM6YTvOAC/+PLeDSaVa+PV4e0jKJhm0ydCQTaGjQmP6HBCTz6IL2
V9tTnYeIwAheCcAStvh8vBpVSjAxdMalJVWA9NphERFqICVd7nOwfag7aD8A+slyJffX8buNpClD
cINpLwo/Ej9pDkmOfE4IfwKW+ybBincPt05Kr712I8NL079y4Y/rpi/RsHYz8JhufBlq3Zbgl7Un
rO1f0JBad7rU4l+AK1t8NtdXOV7KFT9mNvPgw3AUVhfiWSqk2CHJys9t43ufwmSP5NkBA3mqcutF
0oMJI8stY2vItr0j9eyZS5aqAqrwg0TGiNkjPTlk/f5FTfjS5xvetgxiJZmluBltVoJMrPl9v+QL
PNbqnyyLcK+06SCidkuhvlYLFv/iq3dLcPI0b8h+reGr1RktNCHt8xICimUaBKyqRCS35QE54ANb
dCUVl7mnr15TmfHzF83k/2Rw5kG0pgAWkYrnpyghucXDgxMyASwIABClp3bVHlSdoFF93kNYig+C
y/gc9UrrMr6UayL5KVewOT2qHIYYrb8nMZxoK5gfnNqL6iaRDmoleii8NDrWFm7lKBQWk+/TPdaN
uucH1ZiKON/WbkShGzUqJkx2cQDQqTILvrYOoDqefFv1BxM2utCVEt/nsdBaxuN/TCWQfaj+wgAK
FH8gySe9WT9Clz2fkKkPqUhbG8SGhOLkQyqG0HgKsbYv0oSFPkApqD+9JVq98D8tj3g00H3RHsP4
/DujcJTiFwK+1AW+csf1bkP3CN1H3y9Crjby6x19JKRoJxau+iQei5pVxNNkkQz1R7HPuqpjT0Gb
hLyw/TO2z18VDkjezRkd3JrNwJoKG76NZ2cWsE3CNRitap5WvQb959b1ZGq0tUlLUWIC2f/hSNX6
1MMbc/q7n69i+NCWVSH4hwakWdpQwjy7hrZdWCSklfV6IVDH9JFhO9wTyle3MQ579pUBxBv84fUP
gwOzfx5XD9fzutHzNUmjzCfUe3OEid85hi6ec6ZQQ8VcXEQwG57qXZhFOs51LELyDATx2/yNADa9
f0OCWlqk18Ck4D4wX0WX1cI3+0NmdZY5mul/sRIs57ZBfaSIRNqDBQ4gWONUdJG/s88LSiJCyXTS
9/PEE9xI66Iygrbeo/FMiMZlQxKRBRD7y0mmAJDgZJZg1+UC8OBdhDlzyk1mnxR0zYvG6Yaw57at
MmLvymw9J38OuqavuCfvd6CHnIwkkPt5YxjlUDUGiP0Hv//kn8ngbBtvYbiFeARcNkpym0CDQdZZ
OMSQO/pa9yjh6vOEtd58yC2K3fCh3krMqs0WIhMOEdmpQkUb1Z6SUXzrUC8Z1vRni6sCltjvGYt6
g8efJP9lf0bjFOrJ2sNbhcBmAKtN3sWa/q94tKp9p7cYUR3Xsk8nm9MOdXO1D7jHSmkNip/ezGXs
ceP8urZAy6kGjhy728j1EBosCQfYLA2TAF44v3ezuQWlzNks3Kc7I1Ak01v6jW6IBMWiTr5lgkwI
rk5ClIuH8XSVfmWIiV+Rl10I+dbUVQAIWx38My5AqLugYB6s3JS7MIBh4h0wUda01KSBldoRSJ6r
xqTT7KVgajuSCs+LqsWaxcL2Zd3gNwHIl1G4UPzqot85VoNFr/iSxP+gPG2zCCWkQ0CntDop6y5M
zvPJqZPM3d+6BCwspl73R1IhMVMhPltynm8x8QUZQRAlr5LotF2VPmgYr6VfgJxGhHjNRtKM8eW8
zPURKl8Y5gmiWeV1/zoUyyuaPTL/ctVn/bQFKp9U3LNvmvcwUEVTs1y/TxQmwhdzS/y9IyS49xbS
iBL/s7Cc/Jj69YHDd9wqf5apF4+PR5XIiFDY8LfFMWDeZ5XziAqsDrr0iudMpOmSUvQ+pRM3zMGw
AQti3NebsHLrt2jvGCgx/BXb3sSUAbc675IzHMs0JFnfP/Oos/JseS6lB5t2Gd07+5UaospUV7z5
Yj6njkpuNPl0ceACyyZ4xSLozjXhAIY6pQk5tyGdUFAdrNanmGWRGqJOghqq5slLzVQSREwL9+a2
D7HzKc59cy96LWG97IFbpyuoNcsQOFaRaPjri0yruMAC+/6kN3n7REmbfwF0h9wbxEAiYuILCnNX
sv54ASVP9U39gxyLNH4VHaOs1+IVGz+RafL0opAsv2QJK68aDi/jYkhTDRwXPVNwhHGdGGt95OSE
HJ8sjHUVJgd/uJMzUtDHDrMjt+KOxN/0wjEoDDdvJBlIyo7HgmcJLSPtEVYEsezw1hW3Dd8/I+UI
362DZzq8lcjwqyVG1Bg9usb49XrpJR0jX2+YXX+JRVx43LKXmGa0ngG/Ya3bgpGGKv7nwne9AnT1
gCafXVlX+bQNvUr7pjQXXn9+JaV5rkMGkbj4R+Krw6EV2Z+7SbbMQ51mwNJOjG6VuO3VIUzH6H0t
P8iZS4F3L/ES8ihVvYnAS1F/DOOPFOaZNvFiKXhDZu35iSH7KHt3FlGXxz+DZzPQGOn/gYXhiWzm
pxoab9NPmQZA/x2Z2XMCn2FUEE9neAKHNeSOVwRYIa3YviUK8e28VbJENVwymT86I82ZbO/Hslji
VRqH7TCdbMEbohN7s7k+m+czMHJib5GzqDPW0gu0TZUiz4u7sBxQ5ZAkAfyuDBGIHzlyF9Wndtwf
bGO9mGUtoEonkUCpaeRgrsPr/U5LXwIviRdfTMwb4HrVMX7UQTVKYcXVGGMg0ZOp8M96pWbEXw0A
/mHXByg+qJkZLpP+9MrCwrGC65RaK7GQE+vmjzwkzjTAabHweQOAlTf+mYH83+68JylaD0PAy8rg
UFGcNzjXFk5Tg7gWJM/H+vD/E6D74Cb7gMB3I0qE8Z5jeL8sstQ9JVQtOfUZsqPo/WzckuYfEbEe
kzZY80x3AF2JCcHeLJR+H3Z6wrdvV7KIzM8hFbKpBIbWdGooRv2Xux9V5E4z+KRQth3O3aC7s7kh
RPiwNCCly5KjmwnDASfj5CG2b2wYWNic8/CBsJnHTspNsMivMUszD+TF92l1Thc6HiVJUpUzgpik
b4QF15Aw+1MQCK66fdFriAuFPu+ow4LmO+FCO5y1WFkndtfeea6ZrTIvpXER1gkiF3J5ST09l3Ph
SO9MPhXr3kQiXibPo4/2zvTXcdiGTfOgrpdn1Sdwrj1o0sZNrZP71BvNWO+npw8/TLsVD7Xua2qB
eIKX+VUZOlCVpMy1DCh3PYCyqwiSywrC8+F9N1FV6MvaqwAoigeK0IATQVpfQ6FFnHHPjR4qspFP
IdG64uV9Hu69e0L3Cw3uq0B+KobvX6j4jQnfIJzPpk/V/3u2agr1jATN/e3GEg0Zg+xmRLRCNcvj
/QMapmTiCmOyaDhNwattZ87LlAlRZZsI+xX3xtM/W+HEBV1cfXNC9+kEhThhBMLOUgDWE6VnEQgI
sbs7V4xChB/VVp/C/J9FBRO/Tvmzz4iC7NPTNtyz3zaW5rtN63LesJBIe8YqXDolXIB/Gms67SoA
DL9+SikGVabObzxXuZ1ZfcbGIEMvF1AJStbie8xdDq/ZjM/lETYt+Uf74EPYlqgnRn2UoLBKZiQS
PTwrnY6DixoUKTIaOcct4FYurMUwbEozkY+vzfR1Xl23eCTfIP+f7nSBTUYdYyETcKmMuDv2vuJf
QayIpgomcIoyN8TLeyHluYwnqgQhHL6MY0V8HPZrHYet9ica20ewyv3ehFpedVWHEY3munjqaEmi
i5YPWhYUtj7qLUvXIk3A4UR8V1YTlDSgbinlFUu7RJg7AKrJfE96+tWQZ+YgmRHfsEqKg5hcHVr6
ZxUH3bDLYzRayCwPJR2zFwUibLiaTi52b9jSZtA2+9AglDYE8iRCwezCuvJuUNPqYyzLKJ7wh47+
ODxuU4mzIFu4n14zB3GIE7NiXd+DnOEgcYFBBscRu4H02XXwJVYZicnag2rc94XuIAeSNLddYRBh
yUVBGUKGcD6a/ReTcN/Gtx9k2iBRSJCBVel4E+tY4LYoVXNejBPKnuLsFGS30qmA3Bxg0RYgLkGS
eeWYW8LzQWBVtIxmhOOMefXDJY2oaV++btnEWIk0nm4EmFMbnHODQSSJU16aQIe57u7ob4Tzd2pP
SC2e0Fzqn4ksDLqaNIYQxwuJc2Cww1AqJXroPC+S5g7Oj06V8o3XK8DlfBYUBVIRJ5uAaCYTQDB5
DoOkjrDcYLjYKFEgCvI/NpF4dBlDwa1PqcMSjw5AKqKa1Zytr+/X0qAahDusyrGXmtWjJiv20SmB
BJz2OkAMfWDrWvSsG5nBetcOPcCr/1vved22r/DznYcp4zGpgwddC0Z40qs+oYBolCVtTK3fdiEt
h9YGWLltZ674N2iDEyA3o9gpxCVXvoVpSyjmTsqiS5Jp6031dc/gRnjn+POq8h6ZG8CB1S8Zzsxr
0L8bBxEWzR8UYhWzsQlGCMI8qTui6kmHozxmkNBA+w/NDI7vUaJTfZmmxWHE6nDSyLMpKm83EG52
dV4a0AR6Y6dfct6EPJf/CFG/1tJIT8WZp9/KtC8DuodiViO0+bk1ESRPcR3eW382tsmX5b8443Ks
B39NdTbC9Pw9rxZT3d7NaKz9+dK68zOIY5/tGgVpo7cbEqNZ93OyKBI0tVTzvh1F7nBUH9U7iYHC
H30u3m83hoEOigo4CuFWq+6z/RWI5PlxBQY/s5dhrU5d7dL0CLWpHSXgGwmRGdah1B98prDInxjj
zbAYWNSmzmMYRhiGekE0K3UErcJpbbeKjOq1gtX0oUlH0HUGWoaWnDVWe+kIDBtBdQmCOgOEbOsE
nEOBD6gkCRdSnV7tRfa2vzhM0TVJxUPHoZtD8K0+zbtRmepTA5grHXmc7LszPM6+upIVXOI3CiBr
K1pGwHuCKo6CTAafEKIU7I05QahBz1hnNfcZpoN8LuYBnj2iAhnsHrts1zGfZqW+M1dyFPA2bmmI
SR20DrYPA9RM07u+8ps9YxFIrlmRYSgb65tMhAHOnPvYth9JLV0yRON//U6ph/Q0Qc6+p6z4ck/v
1OTX/dRE1yxPiQtyR/2tid+Za0vmardfknS3u8lX5kaX1uUZtxrRvmt4RpTQBzxK8Ep5L1rZ8Mbz
HEDPP9S36Djo/CzvZ5JxSQovR5OSRqwESTlSqixPSBBBDuWcnUU1msT49IZTM2HIRI4J/7pbelOL
hHfVVFpTDiLOP48bA43Dpit5zTaOEpvX00y2LA83zL/1uUNli1RO4k9A3Gsu7PMtOisRhzeis5Ex
6JVLIDOgZi1xA5cu9gxqkclTH2L0v87pVAe/LnA9GOM6Re0vuwpizR/oX2fcb3ZGHdV6zTFMCFHH
sRFa7JgcNbLQIbi5568aw72kkb4eAx+duuHElMpX2dFFin+nV3eO4OJSYsXvaurDAcgF7nF90M+u
pHKKOyI6JYLMPpYp+jPeq0PxGoQEwptaK07E/13foPAZuelQAbji92R6ba5qFrn8yEHViIQNCfQV
7zNCxTOm7j4GM/u6+W4Ai9k4vPfR5vZXeeNznAAe8sKIAP/TKqNB1CeurRsFL3JMlBA7zP96+bB3
nnkrdrB8bLRoAR8ZhyFA0WIbM5/vhVdHDTSluYPwtO57mPBNKOwQDOt3sNMZnslaNjorYiuqVCd6
GYc+lf6ls6qW4g57f1yCcxaORl9WKg6tGFR0+NOdXaT3ZEmKzp1QlWeeyhSgLc9dYvPo10Ao72QG
71o/kwYITIN1ea8FYyvxzfI+m9MtFzlKvzelsNSmbUMMIaR0fDc6hmQ0vO0TugJ0BbViSpOSlFli
y8HmfM/4HB4UBAE/IXDs54qjcxC0iBK3q1aSuBUil/dcz0SrQe1XI7cHVy5ldRHeeZxIxl0alVeX
ouweTFEDVnMALIOBR/Tp4BeQkryOj9AoD///aZGwfQM1KhK7dxE5YMkGN6jDjzVNJaNTpSgTO9ue
QGIccngk3VYGoIt0zwXqmJrNaCnojTFh4gqa57pCMSVnEh5K6fgZnh91RBiF8B8jkmvp9G2Fp0Gv
ySyEp4gMgxizqGjzGeaa/OnK5ot4fXUQqRgUVQgBbLmnw1mru8wxEm5ceeVkSueK9igwbVlrqxdQ
A6iWHi5BiH6/tQrOvS4CjZo9EsOX3q/EF7wpIUHFqdqkgtf2+GAjpkAXACJrYqWVcHNruGwEA2Jc
NhzfFSBxnbDHuW7Q9h/IvuIRH66MT6gUOcN2tJY5A/YQAZgbxaUlgWUbWXzovKVwYbIR4WcuuLJU
z6ypjDB8pHxLTeCENmpCs6O9mrS+3+4L9lnVn2aaec1mRSg/k4pg9hwYWzZZsbAQ6Oc9tI9NQNIu
rOYvexAkk1hvRv+Lm1b7nH/F5/rtVPSIgOW8xAM5Il695vZcL77IxauiFm/NsBpoop1ErC7b/psN
Z03FPv3YmnEKkCcAL5WVc5+BRg5sUVPmBwYIgUws/APkusNRtwjvadgDfn+j/vLtHnTgh864U4JO
VWLHs/8LXz2IrJMXyCOrIK7jC4d+bvnurB20WrMKZbOlCIk7R2sPh9J1PKhl1wZ2rfrr2c3y3OQY
3xd4/RZJTHiunAwpklxx28OhlUsIGfjNofy5s5xp04GozhZDfXgsqGYfEaZIvDiYIIzTQwM6IrTc
28tTHNX49DlU3/P8jIEQ2tqVmEsP351sNruuELTP1d5xEbhGfdL8CN8i6YZeNXHo15D7hxgXuvsZ
RZSpAYHKjsNV55N0qxKjwuflj3IucYDyodImhgSck50F5/fJ6Q+MP9wLoKUb93sXnkBwLSUMMP5r
aIymxFC4tfPxphsmCJwYei7u+xYiZ/lF9I0w00WL48A9qkhVweoHmVJYCFOom/oAE20uQxcF6tzx
B8zsYImUY7ZvzlRtztUBfOFmQAObt60lLpxEXlCrB6VT/GbT9LWi8Mmbp0m0HKRZfUsjirqEPG3K
3oqn68xGHdtZThxeuIme3TyPCo4hauSSBLpJuayXw7Byp9mNAVgc6YbhqwWBEIpdKR4CWX9/nk6b
b0DtZNJFI62cF6IV8ZC6DgVyF4/0IFdENKblAaV39e624PLBy8fMploHtIxadF0a4QRE+dLbm78m
eQckcF0sEkjba4DtykvnT9ert4KRmNGCX4+Dn9BCE9adDxfMN04GsF86GkKKn+LMHPrpWfiCyQ0G
PZzKaqBYs4TV5TxKyiG5T86Sv+utu2VbG/Jl/uKC2FpPiSLgKNW9DTKoRd0pYiFVbiXkno2RIw8r
TsIrnbAV1C9LEFjo7WAB3sCuT6gIAzz4/TcL3tRcXOtDDJpurE2SDY0sBb6CBeOqWJ65sapskq/5
0yFeHIeGdk7Nx6XclVAKJj+OtoZJHmDpM7g8ZDzA+X2UY5GsNqIF6Y8Q+dF8NTuBlu9iYdIZXzh9
LCerfCVCTcyNSyAFgpWUsLPLJVLG7w4RKGgmRh4XmOi7WD3sLR1lQrISNrgGmm8f4lSLm1IzUrNi
SdNJ9kxtvUSqPkh41UiouJMn/iTrAqj9SOEf/Kn29pU/9tja/Eq7vrwRVOpq1jsV2yepjVRwSNgw
IdFCULp/NWNWlBCqzaBbZ4WVsD0cAJGdXb1TV1aANhBFBDVDek6aKI5gtkk5UBSRyTOmHgjiM/j6
4npUHsdDbHnPTcTSFriJNQvr46SPvc528l9rKgnl/+ilGrPPTyRzmfhmepq2a1+sFyRprdTH4XjJ
CpfJzyMgaZFz1Wq/ROTnYtI5883lbH6nF3Pm7NeccNNa361cykW8vIct8cociO/WdGpYFUf6kicy
BIq1yLOrLqM7js54GY9UiHqI+hSk0HPLl3KkwI62CBH71QuNUjXfbXSU3Zz/cBQtpqs+32PT0t+X
gdnzHTgcBtg/iJMVN3F6wX+L4HnfDmqd2nL0mOC7uGfMa2YMbGL3kh5HDZB94JLaCWy6+/Q6qmRq
2KWIpMneEw7/78V2lsjS6Hlury93Srnleja3BZy88ze7YGAzg0IfqXNALzGUG/Nr7IDTsGhuO4i9
0V3fSsgdfAWCjaEpKyv27eQb72NBYMN1mVD0uaZ5QWxcOku3/rdT5rwgM8f445jYLQAoZqlaxZ8B
i6UyHdAP7YOdrUiP6Oq5G2/Pku5o7nW3U6YWkhMRCRJkmuj2bK2g5ObxsDNwt4Py5/g6ggZrYimA
t7dbaEAX3gYmW9a6AHuGMjNEiH8QfDbr09DdT9FpXiW3g8Oyg3BJiwnXLgvMMJBjnLE4fyCa2UzH
HDaCeuN+CRkj6IHtExjWrBss6ubI+kN4XFVlSlNpld/+PXE8xH7fCI2AkH9jB5E9x4jnYW3yrWk2
lX71H8WqNiLQ2y07s0JFxSjkB5TRvUQK65LXOKD6AVW6JaS2SDy5Ry5jVc3/+HzjAx4hxdfCNAsM
ROaiNLWp5fIg6tigEFjsQGIXRl+RQQuIQHdlmUzwNEHibgevTufx78pzyOVQBd34q4x/QLb4nghq
xaajup/c7eS2AN+X3bTjhFM0cnD5c6LCUqQ6o+1V162c45WRsOSHGMOAOmNuK6iKRGdH4Vtl9/wl
EVj+zs5ql6tOQ6iacfqKMukd6rzAEHSwfMYCQ7yUoM8ibjV0YkkC87UVwEUjr0o+YG3ZtvRQ0HQX
j1qEq+bbZEa4DbVh46HiFFohFcCLzy9v2HtFK1scO2PVvJSbRd9jwdwyadkmDRt1jN94fg3ZOVlt
KB9KdG6w46ORU1gM6A63vUOOdmF26TJoOYRWDAQ0yIw5Nd/EWFARL9CopoUVPhvPvH+OQgP+gdBl
ZEOfO/dmRyQ2ducMLqfcblBly4lS1DskvH0CCC7c7g0jxn/juvUstOcVA2ZGUdTNiiBfjuMv5daY
LjNR7XHeNC351lAXFJE7paicRu4M1ZhQZ3Ry4DUmFo8jr/OiKS69waYgGKbkrouoBTvZgcLPkfDe
yYN1GUQkjUq5+QOXX/OxC9OW78iO9+cHfVXK9TUOPPWGN1HFmw+nErOExF/B2kU4Gp5wQ2NmbfUH
DRILIV3ukjaj4z/zGogVT4BEgSw6KajteL4kLh4ZApWK+n4zKrrfuOn9ZzM7YfVFWNV3eg48tnHr
8XFf/Lbsof/l9UNz2BiO2VE7thnn/u5QYbOsUFrlU06BqUdP9dr1QbV7wuN/B95nVAJ04iKsGwPv
/jspZllXuk7jd4OQV5H322qJsvA/exMur+DNijLAC4QC5fYsx+BSgk93VDd6yD7imfZN14HTYVjA
PqE/WalTd9/H4QK5KHrM35lpwcMgxT+OWkSVO2sK14Wm8nLYG2jswFIOFJ6nkY28wa1yn9H2s8UX
TcUVZbB3eIBcZyou2J2Y4hFnocJtvozpZV/aab3v02EN/3l7wNls3fDeuubn81g577Xtqsl5QThV
/V/zncyl7ExsptoSzE3/cg7m4lYetd7ocPqCPecn3qfI1uVOt2QFl0RiwxUppTCBrZRjUioBatFu
AgtE8NF/b/+hDVHd9dAIBxF5sNyxNHsFp64w3lvQNYRECfNYy9rhqq/FNiAEoF/ZtppxrDD/zgIw
/NlG2KRN7A34POZtUiR8kdR9gGC+aO5+TDWBsDNZfp7v0KRmlDKb/58gScYmEt2a6yoSgvNMMIvA
X9xzbRlZ9H9WUrnOHHukvG0gLpYzkkSZUl7UvlRfohAu+eLiOqgHtHoI6y5+CYjZnrsAaXtX8tPN
TomY6eUMGLCLtyHFvCtIY/+KvZlE+tn6qI7AVAdFMAXLYpoevJax/XaIzoPgVfaRx1E9TNwC2E/2
Ms8afWbjIOMI6B/ejH3cWqxR3/TNln9x7tALORKlN60oVtYZTnJ1rBDUkoBMPiQFu+He11cWkqX9
eZ7/6u94patdEfu9y5kxXy1T4HdxEL8WbBsoFqWKLVtNX7RVkeg+lKMTKbDuCaKJJq+DrU73Y7BL
TrvuX3IZ32lfc7LqTqhOrbOAjTKVrUrxuf5bocRAP9T5EzmH3hgaqBNGWGs87JKzbH4Xj3u9zydk
87vAPJfSzL4jhzIdjkrBul2VItRHu1+gM820ITepOX8d28plLNUC4AJjalGUPi++qMkasZvo6FW7
zGIq7XFlWvxn62kxt5sc6VE/FG9/ww9PwBoLHVgI6nn2mzz0+m2naauAdbFy7dtJfApL8akmosXZ
mzBeSD3pL3dKOpoqdxBuJUR5B0IVap3ETRtCYD4R1UJ/jkrrVWRDZzFILOapdw2m6iuIOYUm/nsK
79uxYcdyNsRhzg6H1EQC4WN1RYrb/+rxJcy4KTsGp15x939bt4gF4LF+C7GTgVv1eQl4vdRstSwY
PPai3g/RY9lxhsa02g00cuhIo76gpMQGil0pKw2JTUZN+ZbevrgXVnR6fxEXYvvRj/Ft3SdfmpUO
DfMggAQhSuZJMmD5nrDv8xYRErZjC3hOu++Cdbq3pZx6YRxYvxD9WpmwAn9WQWmW0c/snX3mhBCw
LyizZZHYktEoSMRwRre4COqmD3sXpob1J5Bt5CFQyRY5+dQKr3TjCbHPFYy30fnGnmJb5VOgU7wj
6cCPJT8xKArVxaDM8W50wz4yE9xB3s0mFBCV7Csho59J4plAhdrS7bnhxMCeO0L3e/fMHiuPpFUD
9oJr59jgHnKKcKtC8bTF1fap/s6UoexPRLXss/V3vjkkdbhCZZPuJ6k13JlrG4VOCGilkCyxLC9Y
NyyqdePc8u0x+BzY5cPHFOhvZAsaOBQnpzdMo95SQg8y3Xo58RH6s1gIWeYNlQ63zRISy1F4nAdC
HOP56cHIvYD34Yc2rUsnwxLj7c6TCgRqOoMx0U0fg0WpZrNL3N+OFEQdxxdZd1N8u9JxS031+eSG
jLusEkrT5t92ODVGQN8ImgsSvvTlGobThYOW7/B76Fy/0p90BYPGmq/CmR1xH91rFJVSU5cEz3FG
NE/+iaapPms4C+/9fjarBHPsU897eWuEuVKHv0HS6pRXHJDYCq3UtzarFBeK6eyBBbcbbJ7ni9m4
LicRe16/eEOrFqxPmfHCTBWRFkty3MSE7EhLaYPGJ1pvlriIN/66SoHKyhH6hD9Hu2NV04OWzXdo
ptUUHeUc57S99fUHiP8w2b9RVQ/DXBHyGKCFnnxByLZZFgR8a7b3krM1Oe2Zbc8sceCWa8xID+Sn
2aDNUVqVhDYlsx+wbyTHba2FsVY0Dl89/3/a3x5/7kIGPcxh07kFUYrbQaKYaMVobDvkUZCcawo6
+UOr6O+DoOxccwEyWGtOea63gMuUKMnq1Thkzhxm06MhVf9CwG7G/RAwmxjC1Q+cWZOwZ3226APf
AgUN+pP1xIImjuFcuqCpl+Oxy9gNawCfG3ET13URbJ5qICuEtbnCKACRFvcmX+7ZMDnzNE5wH39o
PemAS63I92AJlluhoG2KGaQ5P5//9kDuXDymYeLegzfB/h4zpvUGvD/1VStpcdKUa0YB3RjnGhb0
sGgtDY5Ab+gEM5t7u8vLdZVW4VL4jd5m9TV6uS6BuBDpl+fSqEqMVunNsn8YjWxEao1gXpXpSF4/
uwyc3+kxu+EpCoxfuEBDowWJF4AI1SZzjiLy+6nIiI+ELE9T69bbwqM7+0YPgITwie6TzTSjmMYS
OjE84EsBTFbT7Rbcp9XyAVKCy3wp9p4frX0xZ3STQeRKdSHOUOLIT+O24P30eGnm4W0Q/+zWpeCU
qucsQxZZOmedz68C2C14mBOHyOZwDjLHy8EfedTrNktYs88UWT3+hsFJN6v5eMupRa8WyxKdyu2Q
EtLNEkHA4VxDzWcKCmQ4GUikNPYeHsmnqvhpiT1Huui2u6Zmsr2VE5n+H/qMlaCatiUtnlEQPFoL
y+oDQdl2jtTACQDYDNO1qfeHn9ocNdYMyiG63rzW5LF1ZI3HWZlzACylrkk4UtUfTFthW/q9LtjW
efncs97pK24jkVMKfO2ZzEYimZ2Dx4YWtPON5HDhlqyRrZJe/lWQQq2M1xmxFzg6ekT+ffUM93gO
OF4+dG3L7BDgINvBL/JIwqmfoCJb2I/pe6Ru43nInUE6T3HKyeg6WPr90guRYSvsFwxf0lZsYL3v
fLbTLsXZwPFGfZVFOcp1A3KKx1h9Jxb+/Vr9IsfyAVoUKRc5DdAJnd5+D4JLIdqLcS6UndJvYsLU
jo3HwHObrYrg6gW5sl7tgw8xvFTfgtLKTh5bDqqaGQQMoY8twTb8cuHYTJgq7ap/3xPwoq7v159U
o7q/vAAW8nAqQnfldPJmO22p1g7Ix7EPgfmhdIa5/23suerpMcWe3SeT1DDaMVXlNce38H4C7gFf
e0aF2T1GeO29xz5c3llPs2L6SUOKuHCNI++Z1h68w5DuS8L4haECdeshOz8ZhuF/9iK+OxFX7Y28
VoDo8ifSNPb/SDP43eWwum07m5KmfZd5GJrXps+5TAh0ayEfJhhGVpPf9LxwdLk6NZf7L09XkwLm
UNMPt3P1EslfE7sSZCHV8co39MxxZZC5ls6GckciHCVhNAUe9Y//vxUi4L91RTRcxIY9G8UEmWjY
jgl71yu+CXgJ5+WCZq9c5abi644B+SIlwCIoBHfN2Zt5olwYtGc/UNJYwfWydVbIaSmoIotmwFFM
m9FxWToZ/90JN365Z/WKD2rLuiMkAgbXFJagzuHf2osMV6sBm1E00kibK1VkRuTzzS8xlXoHDJUl
h0nnh+/mC9TOnma/L7tzJM5KJjv7HYa8llgQyqNo30tre2FJPjEwDFOXNl6ikWJUkywGvUVj5041
NKUcNxAD0cDz88W0Pjx/HldJsyxTvY8/fpdqCEdkS569G5OUb5FuBDDKM3V6Rw6xL0o/rSiikkso
aJffYEEsUm4h0Yo9gUp410YWFd+RKlHU59SZ1zMt5fdWvIO014hClu5c55M/xJet4HeI6WqiOobN
53ILeOCAky1ww1eVffmW0N915aCbi/1KfjfJfNhWO3g/AGaoHEXQHyi35+R1jIM4wdBf449ZCAsW
qWIAlTu5A4PihabaqVwDDgRVYUJu8aA9NRlRJCyIkkO9eSm+Dq2cummPJ85c9A+Up6V2dT4RvERw
SlLcIt9wB25HOhdczSNmIjjq/BoOiFAiUdr1vFUymGNNne+4TreUK919JjziknnYIWorNn/8PSsN
Ep6ks8OxmoJmOVUrOKN/BD2iz60uKdiSQXWtPLWtCRmI+PFx2dquWBIlpwba39ci+M/sf3xHvIBp
4+K9Z8Y2rRkIzinfWNnz22WGYpIylov8gyB8rFsSiPsbwQT6RiUW0f42+rqlw9yO5HtKihqri6Kp
MOZU3hY8zyiL3LFHKWSYWu3IkYbsX2Nf1+f3PEP1AhvDFKNRDWKLc/uQkFZu4r6hEojpiQ/wAVQk
cZGQlCpWC1YF/Ckozs1HoZHe5Ju1s6gHDXPWS5hX8Zp/KcCHSZb3vxwz5Df/VkzzSOMJeYLViXV0
S8CYle9a8r6mcrcUHrG42CMwDezZy18OVKPnRGPWcw+6qpNZk62m9rpbDZpSm/n1znaQejxXeZ95
zNxcSlADuprmK3rqVatIUF/0LJY3fWniktcosK2JfGsh/aq65thI8MFWPyXuHD2bor8F1BfZlvI3
2cY7j+UvJoIn44hHF/vxEBj45Y8tqs1YZ0Jse/cCmGG+fG9ZIuqpetcZWsqcaVb+LXKyI6Zvf3Gs
0onrqjLkucqNZxDxX6nMwQ6ppdie34jB8XKAZVwkPWsy8IoGssS802TikafcFAZuqXdAB8OP6PdB
9muL2eFuh0yiV2exOv9JuPqr9N945fClvZ4mHOYduq6oH0GjGU7yrKCLGA1SZRwdF0gk0FjNvGU6
adLRoa6NZN98ThX2F0UdxmTcIEYhkiSk1DS07tcX/cvVmM1w+r+T75QUsXty/JxUX8CXBMcz8UeC
NR+kzJMoTHarDSYWDsnjt1zUIGIgCzur4otMcCqcszkQ+d8JlWIXupXc0i3ZmeUe9iaQ+61iMncB
R+RX72oJtdFqBUqo1V9HBHGdHaFBZu3VMuT7yEGOcSeiaDh2Y9IKmBB+87eKb1hqCIoSGVYKGhsB
TupXZqLArmj/Sxj6Gvu9RPgGrQmLVrzuZ97jQ+FftVKgPGIf+6wNgVEyJHEZQIXIDzD+ItUDReil
84iMyTgrzQsZvb3028Lnt0p/O2wemgTLGAmRxQVvXXCTGy9jKXkRYAq6pgVgKwPqPAMi6AN0dzwo
m9S7OwRbbQZl1BGZI+OyGZyGsmneBVE9G5CWZLqKy/KFTK4M6SHYcgelZ7C76LGg+tOpwblA4Njd
+DXNh55xqrBKuXPmfhNkh6znY1sVOMugG+P5H1rZOfbiuXzLH0NEARQcv3u1G3vChWP5Pr0EOhBj
l2zGf2TrXclF22fH21UehJ81rVthHvyPWkqrWDa7wf8J2xEKnIiialteGW/1nSTWLOzGwkRqt3Da
Dghfn+DDT0RXTVxHo8MjC0Zf+4zFhoZnbzp7fXLuHv7E8MQW0SiASVnIOCdelUtE2oV1cB4L2Dnq
f6dabOboEgkf6rbRinyW3T7Cr4OSLghhT6KusqwkX266oumgOhP4H+PD4wE/sAYMjxJPIKko9Y8p
+49CW8Ug+sMIoyX+JQFccns5/MK3eay4JYy2Y41G/RSh1h4Tz3m5n5InxqHivDl6Ut3GmoiOG2zA
M0wWIwl5xrd7Ye1k8U4F5m2MO9PHAon8fugzx1TrDI5pA1CggNpVqPibZPQhxeBMe2wX7RbW6Uck
H/DaeYzPtRWsGUFgmE8KAFZlxOK64NFGbSDvUmGKWXm0RzS5VrcFO5AbPi/9wU5qTlt6MXOUQni1
Z4c/Q7p1NSAnW5bidW9tuXHStZILy6CZsthi8jwUEjWFFYQbVK8V0t56fsmybGNG8de0+gbLSqvL
MpxbjqCtD8xFb85U+43/Y8ac1SYcDYNnT+I0EmjzkUVIPVvDBsy4v6e5BAHNrleIU/uTA0Mc0Y6m
oPdML/PIvfbe+kzLPXCzlQZtbBaY82u81ChnzqLusJtUk5YMMaahu4iKoJ++KxACB6o0CVF9LNje
L3hauOAm68nTomRo2BD0uW0DqHtezSe+TTNHYe1LZ4dtDZesid/3blSsCq0w70y5nH8VVlp66Myp
L8r3nfpGSNcQX9x7EJrkDPcbvU/JBvV+R31YpMuSw3ivOAHPUssDL/awS2RB34j9WqyDkQNiH+cV
OcpXoHE3/qbSJVObUOmOz1Z5My2p6g4oawULtZQ7QvPYHG4md8pJsfdb+TLCm1aeptBZDbs/TRWI
wxFZN9WvzuqCWzspiJSYTpkho5WFueFUAS4tfbcW/S/Tuj3SiRwN4IPtQbYwugBd5oohdm+L/xQQ
lcKgQNQgpuwBhpLSGKbZ/nJOntmtsboHg8UyWqsYE6xOPGU7CK79TcYa+hrcrnAizs73onXLM/sP
SI+umDD6BDcRPD95xm2UQJommcaRyddYA9bCZe0ViNvKXmUS35Vpla1x6SrfpcOSLgd0gQTIW9je
OekEs1jgDu4GsFPiIwqwQqDzKo2TyJQm7P7X37glnrpEJyqxyUrN/zPyU90K3zGEq2VzSkebBSCn
MGn5lwe5+55du8kLJjG0bd36Kp5/kC7yuA6Xi7rZ2UTkFNK6u4vbYA1w/AagpSrLyncpWpgXMYN/
x3xQVrSlY4jwg5j2DGeA8UnXQu0SOkq/Z/626Jz6HjUVOXR6891NflUuHWLkVsdRyq7p5VOMNCNT
ARyBIpelCC3MDljZ6S3bMCKsDVGs8fx2F+ZkSIUmb6U/0vXxAcjqt8T/iv1GwM6T21LydVIHp8e1
t5QdEusuuyQsCKXaClLczwbTfI9n8tFW4ZTV1r/xRQj1KEFukMpzjUOJR2+hpPMLdOSLGMVNTjn/
O9DP+C8b64AXO0fOgQ5zhf4pKQr3lI6lcePHOcMHKQcYYrvTtOEfjlqJoYtQifhcqroirIfwkfFA
FtQbAkiGSdBWT8oJUz7x075KexOf9aKMKiVcveEJZqkGK5qqS9M4OEmJ4hjA3aOCNlDXSMewoPMT
DaiqLBJDBB1qC+mvmKNMhTjfxelvrgbTMbMxoBIEURdFTZdwOERW3cYtsplhq4IwjXK2i5OLQn3Y
y1SmgRbxdtre1/IIrKKNzJ0yACQGMduBrH5LzrqUxsyrdKN0/FC4ZjqYxJJZnaO3y29GS/Q7z1c3
DQuXhZtE8iVmdNVSl7nHzswCyHa8S3gQzmETTys0UZ1rTRN/28S0DG/zH/PHtdLjK01PodKp0M/p
om3UpVdS9AgVltsHAqUDMNc7L1GYQxz0uoFu4p/zuQPsIP721WAPwXUTbEF21NEQZK4KhUF0Xx2P
6UsaV64Aqk4S/52fho+87+wfI5OyENbiC0PGYDPGdIDl1byHvZavS/LH1kAqUA8mqamPQfPRZaYm
Q8NO/s/g4DEFEDUGGKFwj/HMM+nTyencd2lRbqj9L3JeNIGOgeFHVzwbqM6AbcvPbAXl10I/gq8r
daL+VTmLr8Yrk4Wc2DTCpVACQ8bDioN3vNKn1VE8oyV2ValhPwCHjxganSxQBSuA/zgzFfZdYCIE
yeIrti/v6WnKmG0Bc6599ljBvXxK0v6yrgjsLqlJgrf5grpzNjcTS01JD5/0gN0VDbzFgEF6xL//
gTTtANZgZyuOYUF8H+gcLP/hIPyWQYaAcQq25W91qgwX3c1rfXsWSD7fkbDvpemRBSqTbJrgt0pj
XaWK7fflXQRnwqKofXqfkkkkUC3CKnSntNULpT/tZQwXtL9/DLN9bjYGY3BpA9ze7DS2Jx1x+GeL
fS+5H1wMUSqvxu+Zy6lOk2+qTPbuqlx3XNQ75POp6Yi7uUuwIUDQcOGXnrSqNVma1nzWxTEIx8rm
+nu2c1IrzKzrmE3BDpygzbWLHKfKEmkSMpR5ZDDGJEzRzlpTe6RqM/xVUNWWq6qzhmE4JvBXXEet
1yvPR0a8SfHmATkIzKGqrCXOQKEsTH9ik4njUAQPncwKoQA83CEhu1ziDUF2ZND94oFWc8FjSWTZ
2NxHMwUe2gGN/5AN8dLHnG4X5r9Ljmp/L5sHsO+RKvlf+fsKOUdc/iM51k4vKBazT7nT4wDb0Y/6
ghGqTrHTvpqh9Hbg2t7prgUCepXbmw8WYbSp5NVhcRKJ0rLqT+YRC8wy3ERoVCZgY6oqBMhLqQOt
pHJxfM3eIUAJyXYFZNpq8OVjLPpGjRUyQ3az0rLaGRQsBQSTEMGj2+hg6vINJ+wn7m3PH5gsQ7SD
VJ+0PSIefOCfYHC9M2oHQrQi7p9U9UDms5TghSGwhBjJ4vF+GcQTH+AlrEzx4cz/ixdR6q8wGTrc
K6vkfdUSdi8wJcXmUE8ROzRxLe91v3diPOh65VsPwDhpRl9RprdsH//+Lhk//vxD4tNVpkUnukxt
NqtofUSLEWmDL00x5Iz84SGilJ91UlpKvMXbjtL01aTU01haz/266GGFG6Q7hs28tB6sNanBz/mj
+UZzeRZc40AsdYAkh6M9oCdpXUF6FdzDjzPpMMkVDIVLBqVslf+IQZOF7rSAStvfOIWpofHWHbI1
0M73bu4HUPuP9fmjFBjJCAXt7kmkgmyvVv0Ou+5JEcOcy/ZSsoBl7c3GvXdNPAkuhoJHcR+Igp98
mlMi7ZbnlNHBaAXEpJyGk4N36Cn+HNRAzDrQCXNWfvI8L5a5Z/cRD2Xg/ejF44nu6Zsr5TWdutR9
en6uic0oOkJJyJpcRJL1kw4JWfBBkCgXzdal+C5uugQYCBtJ+9n7M9ZqOWrveC+9kbO2bW/qrCSe
L5nfEdJN5f5kxlRQ1AuyRHAET3GmlllRUBQPYgOW/2YUQ1ErSFmr/wcLh7YcceEDhSTxw9pdktUN
bIhRUyLon9NQjCmSHtIM2Uj6dq7DUjHss83apNEzVLKCzuURxUW6bYA4pbySK+43ruEUUWV3a0SE
VjjB4WLrp6NYRnkkR4SbzGKLm/BRsmdio4PfDzaArguoAkVNty8tJUQLHW7k8HhTkHZ+C91aHCXi
86Y/KfxoBx3MRsQbx95SDysn+8cUMeKqTp8bkqSfGzqoDXk6a4FJnpRo2hVkJ77XVZC9l+VVoTdi
cxAjI15CrpLhohXLFHaQbvKCDpkcuyEA4x65nS5KmpOk9VcCu5xPVCTmCUcjqjgYUwxrRbuPiasN
NwA7PKJ7oWG9XLMhV9w+MsyWH/civj4fk/5SE8iaC7riz0ddBGC6yy/B+lZctSBeg4bT71GG5RW2
C5MJ4qBwFS+ntQi/o5xODyBX5kJKVmzZX7F3SoWAcs8U/nS7VJCH409yXs3eEXp/kVwtrhNvkKoD
wND490ajuZL5OfF0RjZ056C0mV8va/IYlYVf5lgn7JMEe5jCssMfQLAmOQfS2oKmmwI4zcracBJ0
KjrCWGlCwqQJKsAXDTEmVRjnZ+TSoYRSkCiQ6WQyPFZVUDGcD8KG0IXOezamNimELm/QmHAtwj+j
NRX+hDz3gxFc/uORlKCttSYrpFTawQcx7M0qcm+bxYapvQOhD0hL4Jd45N4wcscISkZvEU/Wlluz
pENwce5jgmJjxRO54ixbf3mbOuh1LkW+oMj9feg4mS058OYFcPLFiRSXsVB9wxHEH4lnQwS/WGFA
SbjnsM15+w5NKNkDttwqEAoLqBMPFVArP6RdcDmxI1x7ZajHB0QWmKYpXXjXTssmCdhNzDe2kMIp
6S0nT4/AkVYdpKyOaoefG+B/G9q4XU2kuw+TEbYxGW4yOb1f9RGQZHDHNeFMw9ZdnC9rWakDXiFg
sYDi067G8KrD1OwqU8HsI55dvetqm68UcyRRwdk4BnAWiCGy3vEJ/m7/ppjAbKtGUTttSr96Wi5r
pio6o3AQblQv7rhEU9TP/SdjZK8a78e+iDqRnaXOXc8OhsKFEU7uKojEQ5T72eS2FAcokl4yTVDN
L9MYNPt/0ZZF6jqPDsNjDWLMxpnWmTCRtqH/dZ53KtGe32lmgZ4ClK9P3fUlrb3fqdcv7Q2pFB0k
yEmybrKbdHaii3U9ojU4r/pqbAONytG1NnllhIDonYQYqI9gE6ipvfYXJ3Y0S4NyguJr9+cTuAQA
vbObiZdBygKRbnHDp4r6UhNgI69Hp4B9BRTi5WkP/TBnqmv63cx/a/fbcvKOvnjEnV2OpaaZpzS4
Ttr8xvArgXhWCewSzMx+oGWcYqDdamD+5D94WiVzOov8jNU5kALstQ60R81qp9zKLZ9KJ/FhTso7
SZcK4RLKuisdS0+jLYL01YetgaesDVNQPMFqqMRrHD5J/p59MqIZ0bj74O1sVhhY4U9r4qtf3Wru
qAzzuQl4n2o8QNV5rFfGQOyW43h86byXK5U/HVN4r/Ymw7Spojv3SIvltJ1zxOY6AIqdcF96zt7l
pPh5yLScZLaPHnXj1bEezL7hWSuzOsjVJD0nOyDeQ2SmlUGdTjPO8vfMgeiy6/KLz/w7M9EnSBER
pH7WFA/63kliSEdwJP/Si2IruLfMZpYRNmL6pMZvD3biZpcVDQIR381A8gDk7gpAeFgn8PUBUWff
InQcV3YUal5MD8WdHP7OL2z/K5Yj/NHeFS7Pb5Bpdj4w22zeFVcT73cwjY5CmUtOoAI+0nGzw3uD
ORs6aFL24lsNWiPSKRDYIj0QybmqVXBsNXEaX4mAL5R5OJa47IZodF20zjjpSgW/mxrStN8KznVJ
1wcV+YQvmoA0M4qNZgi3IFj1B8lLD7t64QFWBZMWm+aSEwHVjXTGHHad2QWeF5cst6EG/Pd9EASl
nXhkT+M3BYD/EfkiIV39DlxQOS9B/2HlPf4yoBDk7CLP4RKGE/zMP7iSNH2eiGddCVKpRxAsyE8K
Yn4AJCHj00LWiBaA9hFz9uzwDmsPMmyzD3ARiMfnRsp3HSsPczuHm+5GoqK5dwR5P3lEX3LXyr35
vF80gbfgiYZGaO+hA+F2B5mCdFA3tokdFl8BF9O3VZQ9eicuIErArOUbqFEllotS7YsRHb7ihq6n
FyQNgd7VfoMY62pyY7gjmsVyC5iXY2+VqXMmMAFGqml48DkOHYcEi7WdjBoVlRsz5jP2g8n7RP1N
xMHIkp9M9YrcTokbpXER11mzY9GyfITqzMcHM/W06rgwnWGnp4A2TT6XGV+AI7VtzNtGOCLLy4sz
OjCReTCvBigN2b2rjaHC9EoCRa7gH0tdShmMtoozUnBJWtSZzq2zNHOxROlv4tK0dZNCQgnPn0Bj
dz6/Um/OvlIpPxrRIH9Kf/02SJIhIFrmLB37iD1ge0Y40Dz9+cxL8b4lwqijRN00qn0Z21NW39Bb
FrrRsCTvS0fSZUNe/zItm2QKBqMiKiRXY/qnK7p9i+E3vU0SAOwe5/LeNg85dZ5xlhjRXX1iH0V7
YgQ14LtO9RFHJNZx6/upbLslaGqtuepZS6WxsfFZmqATJFy3yyjsdBGoriaZX5LZMuIVTEcP4jJi
Wt2cPLepaZ1SgQ3cFF+ORp87YKtTBasTaVqbDzgsbkw+uNWf67n2XIywa4RtV019HU6ZtqHbWjmk
eV8rTdFcyW4kPHJkZ/k2dyoKVWErYMGWV3AO0hdo+34fdaj52lPuosUmIvsjfoa7AZXRm0u1xml+
CR9pi/GRv7W8CJBBzx1kPT3JPistvSzoQ00gqRbbG4KGC99nwdjd5CGprO/g5Ql4SWJWml5KsQb+
gHJfDr+XHWM6Muu33rI73sJJigRPyvZ0I6TN8D3pPjOknZZflZt3wyGVVT7+hZ5pHSeU1BpEKpGP
cpelor/KRhN+2AQfzbFUX/fh8Yvp3F3yugtLXZtz4v/zX5VeEaTYwT/BECyFSb/26ps3yfTzPP3y
uq23cpMkuR9OtQtwvAXLqRHtZuBSj3tzNgvjl9EbmhwRQiTJCex7FrBAxF7iz2OLbSRyMsJxLZ/b
y5/VTL2PxZ+zH+BS55HFNpHPEmxULsZF3Z5kwN4YBkE9rypZwqQsIx1SrTQnUhSTC2H7aAjyR0Ad
qjRYLhyDb8L5YtanWfZAdAmEOOpXmZKnjVd1XBF+MrTYkanUO2eN5nyAGp+5+24hnM4GP+u8bQzU
gAs286ZEcfT1hy9LMjwpTTtsaISbsHYbLtXmBEOhR3Xw0e9/WjhEThue2Gl62XtaAsr0U6p0jSE0
kfu/eRCbuypkOoux8C0tuV4Ra0xoA1bj49G2BX20uLLfwQOD0H094bWSzGrkpk/9vwYa7vDjlW4L
6msIE73bagKBW6KH2XpSRxiiA4V+bBvLjYMDMEPKb8mx59t9eHxjsH1iYn+d23WfCCaVb4JueDO+
payrJBrPWdQ5RAxLrk8UemlvQ5/6l8Nnnt5YphUchuradlOvC6ffnynAbVfE3Tj6Lx83Gti64mn2
Xw6GtEZdJvlnIDmUt75jJGpiN7ua6eE0mr/E8ct2Is+AZzMOCGrEyZ0Ijvcmuujtvwf5keT008bN
In0Uu11KFczP5nA8kgHnZedRbChR6jLPLZIQhPUo4YlGXtHH3+r1nI0a1r1S5IbfcooOj5QCMwu3
TG8zTQH+MU2SCgK/Rp3aIVwNmObTmKxhGrm1R5zly6V8MTzjnqqeiLq1dYSKVZA+mkkxQfjCidEp
pMpzh/cu+wQgI2BDrhgnwzxmUNOXxhnzBF5IWWY7FOMJutfXHP6/ENRCGJWWoGvgV/JVhZ5KlJzi
c0mnlTwwudyS3hbnBq7mY+KLCG3iIHKBp0Az/u6Cx0sLpeOiQM8M4E0YJX/3PaPVwNFUOASp/TNx
nKMBWfe6YgnwlZYefBuUsVJ8ofR29tvNoSySSnrbCYLDSwWMQSzLIIO9u1J6bvfzB7l8GHdoST92
P3VgqbkSY1VwPgb7K6NxRvLoml2q8FAJ4HodvC8D+wXe0LMDlifYWbFZLwleMBAiqP+DZeH4Zsl4
YUBhLL8wHRVHXqFhpFlPs82g2dHTO+9ArHU1epkoqkcIy5gfqGK+j3uTsPSRUDqb3QxI9QItBX61
EfnkOvzmH1grahx8DeaLVmcDVsMXXwCjlXmAD07MrjZJYgZ6sC96p/Og/5t6eYM0+6c2HiOhmAhA
tXkgUoDi+lnQmYsycYtGVzA9kI8vcghnPr+dhzXmMxGt/N8umwBGX7GyqF5dq7pJzpj/ygVAgAtx
xWB2MyLUWCH90ap7eSWYKeWPDTPjb/C8sqyrLPHLpUgfMyfrmG340UsLsRQ45DURT5rzNXvyWZFC
7AX/CpMXEguNpBk8qB0SuchmXxhaiLRPnvGzmKM+TqblY5EoRax6gbiRZqlB5yIWNl/0unxD2g/t
f5FgMKLhd9y07MNFVVLAxf3fxwS9vsr7dJXEb2btXAxJm2X/A4FmyyWodNxKv3E1hu0mQnas4MoY
j6uMoqh1WsJP+mSJs5xyZ6qzdKPrVS+eoOxKAdDJ/uMBSiIZCcmZz8YQqnNqmlCISQmHwFIxpku3
CjRgp6W8m1IlcNAKe4LKY2uifTmr56vM65K9Jrv1+MPitb76rzjfU/tDi16xVNMjbqHcl2zR6Ike
dcfZ0ZrTAtlZvh+am/L3Agif5veLbGdG0cNjPLt7VW/8r3Bzp33fi17cASatd2CblKFUIrsPNN6/
ykcrM/qDGXDDUh2fEyZ5EkyU44mDICw35zHFLoR6xyvzKvcCoGskv+b2cEB8R8sAbaL6xeDDH4eM
gRblzvbcFjw+aUh8jAtI2kdhUlQbaysnNRy8jsD8ALQgYtXYOf575hMwCP+iMwDxfNlNHjnob1N+
4PqoqVsmWInTkKMfCrdvlVO4ZP3Fn6EudsC1mSO29xhEWOk8cHX3zESck4BCOAL8CZso+2VU7CDy
+mRVetkZwh16AORdRri8dMmVHIlojxaXf/+dA8DSTmzbJVeolI8gEjxzXPotL7v/C34X7o22P+zF
2wkww9X1Ze8luL7LTUpTaYGiKzvd19pH+7YtVV2GMWBYGyQnP7Qgge/Uk177TTcdE8A1+Uj+CJ7p
U/r5H8UDLmD6GgNDKQN7djuTxHyiaCieddci7LzlPHZpH3LuDuIpBVzaO5M/KgJIWX87q9/wiQXy
maA/opT9c91SA9phtA08F+OMyu+TbyLA94sh3cySOzHiU5MeLBtHkVJDpcmUcDvteV1K9nAlLTli
vuRa2q0Z4r5rDe0641ehhpucvJzzZElrHX+PkRG2WormKZbDHY5lPlLLt63/4i0yBkJF/p8gcnTj
aEKm3wW0JzpQG14c958z7spXV4JTp37dKMb1KWe57PdPZfBJFvWQ7DfHow8/UAWIVzGT1D/59ML6
ltnrmjcUg0bstzWbR2/eUyiq/7kPs8Mu/Dj1oWzyFxxjWR9VTYrh6ZqmpAhFDmhdrE8JGAVlPtub
MKiD5OhFPNEzQ0jFoMkKh6fWxIx6imORX+kVzEO62G6tGtpF12S84KQWRwDiS+oeKfmTtv0dI4/F
GiSmyZK9KZpLFCcPSkdp4n62b4HrjFlmaM4l08Dd50MYBCz8apSuJYyg0k5HgHsYLcGkmRCBPR1V
46g7Vt1Rwb1L/WYXjWVMq1oLw4pw84CtVMuvkoP05a1uYGxjj7UDLpP1I9T1ZkDQkun5pBBaTFsI
CGQ84ozL+gXZxkBHx8Fn0CeakKVTZZArtK3B//9e0byvL9VoOZz3Jv6ianv2RNrWBFgsIwLkzn7D
RsrcTK/9k0SGA0armrIzkTGbuP10H+P/yZtE0dq7fYZhimPCP32tbAe5vza49B+Z8RaTq9GP1YlZ
V1+NaNCbsz/M0OfAN1E49PtqncnfXzkcTm4jUCP/oM8VmZnUKrWTk+PJPKkTl6c72a3BT2Ue0LSU
5l6xYjrvtyDswqoXoKm8yI7HOj2+yopqdgdnyu8JkYapWxYUMX5FIc4tRtvsK2KhR1e9ghGwDWf4
ACeIKg+flT8DUI5TIbbBt7IH0aqObEkAkKueCXIleDUijRfzmNw6+gkfm67r47Vq11Yq7rXwczs/
fSx8XsR6ySr+BsA8PfofimQrRubhI7WA954iciuvefL0qHD1PYKVyWL9E0waBxQVFzvOvp4gBNEm
unWi4qK/Zpng/Xz/KwWENN2kPo6ETJSx6tYBlWkatbU2G3QwcE16I8vwdKk2x975/2gyHFuJw1fg
wEtIMjJHaF53DLOMqgPSl9qaVSYk0tEfUqgrCJJoz+f3JaAB5ojHThSXvL0d8uwoBtrWVD/Icp+g
tvYrpm4CC3SiQ5wGMRLtoj7O14VuKbKxvZsSsmM4VkQH7+iZvwH0T2aZVXUwXEdJF2/K29EVJcAn
gavu9uuXwhwg0Jxv6pV3FKi/lyOKS5G5chGamCZs86wB4zNWsVnzy8Zha6JuIKSma7hafzB8yBiS
p9/7KyPVmBqPa+7VEFp47o6wtUFBhJEWeNscWikWZUcUcg7DjTZUptshZY0YnS0tNuU/YPL6022z
KR3pfx+LuKQ93bnTrMsQBbRitaDEMLZoR+svBQZ2JNnnmSCOqKnJj1twNMBsmuJ1EciMkYGUOYQD
p5ZefErBHDZDIlf7vZJVU/aA0DFMnrd14tK7349ngfeHK4HDdlFAzTJU8Rln9lTatNjIyl4EX0rw
9FHJiuQ1gCRSB7QE1DQCNfkTvuJLIME2JBpvyqUrFAJ3+23wvElZPhJzDcH8CMgK8USzuqK9NGdE
KqDP+cGGpDgl1WBKrQWxTv8CAUNavpBLGDI7uXBfs1sE9/1r/eUVMulCJVjlpRX6Plx7gzkgcgfa
xTcsqy11+Rx+o/Yp6i67M7QkvQBarqvKGo7kYOC/YMtXIVqU5/g/eQvtNPX2BIIf5lA2JPuCIOZ6
ovSUNsrZOUyN/713qcQnPQEc8cpo0baIv4utqUAselFpxP7MHbxa/XRWLeuD7zzyPbOBoX2bw1m1
/B933XT5/GZBt9JNmlX79w8v0bhFjm+XEXpYjqo9NumGhvKr8xZG4K4tPrSP9ixW/IeY1EonXGZm
WlzI3oe4k0vHHvNiMT+cXGR9BtnpuwZlkcrtQrZ8H8k5z+D5Ec7L5J+LoLbN+hnshFKhz+a/Zvv1
+5wt2NRizUvEH+R+j2kCmXXON4DoV11+jQADBotw0CLKMbeKr1w2mwKQuAKZ6VoA36pLxSoCDTTX
h4tI6sZLKkMKmEeBocMKea1xPEeY0jlbwl0eFQT4bwS+GX+x4V8GjBevW/+MoPiTP+ziaaKh03ri
MdgSV8kTm2kCidC5P2o/UP0e03qxtRbAWnfA4JTeXDaMZ6ZjiZuLsV0qUPqacESYeMIqjzU5OU+6
5n4Ej34qX6jYwk6AZY3wA8JCWzi0SKZSCGZRTlGBys8ixnztTDI28oOcRwMbXwkkrYAnywukLs8O
61zyflvywrUu0LeSHJ9zXaNsk79M2MxjHh1FGcMEUWG+DNuXrI3pc0JUv+CGdSbsP9161eTSDZGs
vhAWMmhWnI9LcsjLTXI3TY+SoUW4umSbeVSbNuj1qNzSywKN1D9IQ5F4SIzr46FMjmRGZr6NbIVj
3Z6uRBFDuf3YPSFcazO6+Uh9MEool2Oc8OIJH4cxqi9T6vK8eYrUDMjplVP602JJA0+habfhCwmI
3+lHZ4LYiMGGSzvOU4Gj3GX4x4LyQTv1FC9z4iQc2DQWndDcQtWpCs+hTzy5SGAOvIgHUkGtxmfO
7L2cT3qzbxtapncPzLBj0hc8owKcgxr0fEzEg+bEHF2zef4eB8kpx4RspEnYIbsVUsOknOSJyDDy
OfXxMbTwrS4rJ7QoNXt4gcwEsCDCu4cIKbSM730/XRHaaXyXYVCfZnZvjFxh+4leHGVSSMkWayQk
6uKpfrECQ/VaM75YiOCfdg40PIt23QbVgQromlxxOas2iIfl6qH0XzU7hmWeAujZYDFgueqtNNDg
9jPW/Ub03pNwDeryya5aycdTDmubErf5OpLwoAoX+SdBCE1g/TG344pQw2roaCUMVDL2c8ns9lVv
LkteVqkiJXIy2YR7OHX92Wr4xyHcojw0WU4kORMIn9s53WzGGmcYTDvXAtf3Nlqz2xeBU+riObxd
Cak0Xb8F3lIEWw9z37dvJXB6OgW0qsZBV/BMrRJSiA0+gqnkkCngLH8G5d2Tg6o7/jkp7rwZUmzG
Un/3TLgyi8GtUPr9L+60oE5PpPdD+b+1gGZ0xWf99y5FMYuQsKLY0Zwi3jgarIgy2l2pwu0X9VE5
ANyY8YsgUWTSzXYIAtOSjDm+l9n1PneVflXxo1aIstbzUItoBiHF6a+Q4pwqrHITo0fSTiHVUO6/
ZiHYemWKM5mxqKyJT96o+I/7DbijRK0088b1kf5bNqpHDSen59EV8MJO8/iM/G43GQET1O0+k1nR
J/UUA9LYc4PphJFuxBDgVnP/91QhwzokDR86UoF7BUtvhuq4iB14nT/1QGrli9wSieSvlF4BW2/a
bZoDUjT+mpcWH8KZoDnXv6SFivPMkjmU07GDdz38iaJ9S4CI7xKRdcXNvGCtoPCU82iprJv1iwwL
ZKrlBkkDpiJ7CBs37UEYom9FDkbnPyThJF7hyLvB6Wt8oB1tCHwgHvLLLOP4sSsj3PWSR/BhbdV2
d5sUVgt/z1VTlBpf+wbybSb13CgND9KCNed8UD77tDTqvRu/3daLVkKtq6IywQ/MQ4rIYhA+3XSg
saoJgac+H1rCVAsct4Px7FyPpLYsK+61xjx2WpcsacZkLhf2r0PXlDTlNldW5IKRXgKG8l8Ccn07
9GQbPLYXwOdvjcsax6NK/q8D+0wVKoE2pUgmQ54sbMhW9/cpaidVir6SEM6hbaE5VEj9z0AcRy2q
PSw70z9fpOon+FkvfjfM2FVcYREgjevl0VT3vTQO2/netPTGQNi2apvX4CoYrpWSUq2HS0rn0LGL
IgOb5zxiHV26RqUnW3b/Hkx4vfdjSDiTWgnOrTSTFYx19COjsjFtDdd0gvOK0nXKKN+So9RF6TT6
iAMfX3oVgK1CYv7UCiDJqb3xfGZS/Cye71BFcobfcQQWu3rS8XX/YePiGctfdFux6kJ0pzZXkhW9
ejQe+21xzJJ4Tv5s/VAT7CTtA443LUHk0H+UrYkTHbJf7pD2q5GvJk6NcfOV+iEcA2u2dMemLQfD
Q0h1IV+oCXDomytJB0SsBiRD4mNxNwUAfVaWLxsVzNget9SYbl4L0WowV+FJ9NMMoI7mkbIh4gEC
5n9NTqX1W+gqxNpJ2raiqdOvNHd+okIm3B9Ekw26i0/CV+3p/SDj5pnwUdlxLL8JmOeRU/Ihp71l
6+pqbHlGr5v+FjeVYMtCdIPqpUGwpIVzBl7zjz9XcqPFtDAVCeAVil+cvxSNes0SKIEgT8Vs6Jxg
+gUksv6SHHrOl7/gVuuu/gKVEW7cgbnGN3RDph91DW7++GhCbuwPEuO8wsQ89zZ7cC9cmPYr8vm9
RAIM2g6c8Are0lQbBhqtAQ2sdvJt6hiOn/jl5FxFy/BcDtA0eIKAw1FTYBQGAiqYkLQwJSiG/Mbw
Xdwd2LHh0tQ59qngSDAqBSLPL4/eW/ebGAoBtYY68mQpp4Q9bXJoYx1CggkOh4BcNaD/aos7l+/f
CvgZ6YAAzlW4SVSMNFEnwY3NVI+1F5chOKnlTcAjAecn4GPhh60vuvgzChlRu4GKBZIXooiUp1Kf
D4FqzPG3GWNdThaJ+cfmT/SmjuSAkLIGFCqq7+0rSnf5gY7EH3u2gonMm2Li+T4+07tKdF96wGri
ic2Bm4YQ1J7ZN5ho9vXyTbBfRN2wFL9pPb5J/Zn+7ofV5O6UR0JM+qPZPcArDkPAPKzK4rzjKAv8
KM1pBwTJjXYOyn6DuhSoVFSm6/vh8Y42gJ9WxZVBmDZIi+hLSrHPM2ggJFHm8NvzVEV2TVDW9sl+
NjPjNVT7KCte1a4Jrz6TtcBOXHen53D2WkCHrZIQBfapfFLTjkvJSv7OzkU1HKNA7AzoRFhIUrfa
/28OznpDHEPXMHqPR6kEr3+qAZAKiNhUBWCyZd6E0rKf7xwIy9/inxP6mXiEAt2jBKNUtV0Ba8nF
JLz/wKjTplnkdOs7cPxZ0FqrdlFuhUHHVzgJOGxviRuhPufHxU6OJdF9I2znqMuJ0DXxwWv97QbA
EJ51aDNfa3n5R4TcF5huDo+5d6xzK+AmXt5JQSf2WUrdDYRNi1d6Od8p4LllNoiA6vagYiTKPfyn
VJ/h/9d0bBoB4vlVv6yzvWozIuf0yglgDCV/xglTvuzkIFRsqmlAafZ3sTTONpGVkMJHX1Mr7iFl
syGrszu38N/DY+GCm8NUKXslxz3u1U+T3bcLJZqpx6my7lhbEcIjmOGs0ebJ/QBUIt5ex5vzwupf
s2N2cKdWlqYChz22uPoGQqRX0eADZkNkimkx8BIXeg9P2Sqw5gt1zFWe5SAjEG0rHGwOEo5Wq1ca
QpTKUrWZbJVTsF/xth5Lt/AHlNigjM2qvKjKnn2UQBKCq6pU8kHtSWI1SgNwA15ySTEs6ZB45oMP
KGN3xHjte+/W4vuTZzv/nWixPh0rMlu4A1PXdGIqOwa+As8YzitAaFgnF8dmDs3SOOLKn+BygFiO
Ru/3wX6PhjztKwxriPlyVi3g+x8Wv9w7yeQR4n8e91+DK0NIy6eB5/ukfp6f89EeOGJDfY1piL8r
GRSztg7hFyFX9td82FWNAJzmh5FhdDmBWgXeZ/xRHc93bQX6zsH4W3ORQ5us8H5alvlvON71IIfQ
gWc8RizV2Yf4UnCu9Ya/5f4wR9z9fwetaVjGocyoFsn5Dp4py4wFuAfyIRSxxAM0ssVFLxL3rxSm
kFZEIUzx9GLrwYFcuKQsXBp2qKGyj/nATEbjHpzFaxLzc8XyqEy6zMm81q7DD5Gg5S0pZBdK97E6
XjXR80d9MwCjKgYxBH6Vm0Kp/Ay/+evkK+XUyFCCVBnGYjITDQ7lsiLOonzAXMlaXec8xliMdxtY
/YLjxEMK6Zqz4gFlDmhwmBCkO7/De6slew7qKaT2LRtCNFu3QOInqGotPrfjnauUmcKG0Quo7EwQ
sWCn5Uqox3UqxvA1UgaQDiH+d0yWxsWIapgKMsXtimMD1QW8NYC9mFU4Hb62WjvNkktD0qcGGFom
ddLkPtRkN+UiW2QKp8GCDJxwDRdcl+TeSovE5QIHX7Zr9x37WwDYR2RbK2IW0AEL5fYvOaygGtzJ
da4H4zoVDFY9PAQNTA/7cPPfwQJZj17M/I/5qbo0HQ3gDnKIWtGYJS+kW+f/VOXD/GqajjyqX+iA
XHIveNgdES97Yo5W4ZxiXHOpfkVuoYUg1aQXrIB7kS8ZA+A7fAY6Q1i9KvQJEq+6swiHzlSwcLRx
SR9hXKH5qcF+Z7rbz4xZo/HZJUbjekDQ1hjOOrnkZAdCmNsCuRmtT2340Qv0vYORsw3MrC07wCFw
9qJUaglaDa4KuwNgQ2ccUnZMCxPf1A3VRB6vRdncTOvkOF1aAY36hbuj/KLiMYhJWSt7Ga4Ysfoh
vT6oEollQbXCcKSS8uaxGRR8zguMkn0PWpDw5BMwwAZ8xwWsM46xieViYNZ6YdpllECkLmOJgo7f
9ROo4bVZKghanCFEVIy4Hfmhs0W6U3tm0pQN6DLcNH1Gn64w3bgR9jduJ0k+dkHk72BB6VXkk9uV
qrGyWbzG9ESX+58RkAIIjg1SnHBSnuZYYq/91687S5FZUsjL0iUwoVfYzzal5R0++1d88hbaj7jL
7q7xeZJqNohEcSp0xgLJqdXuGXen9hKNk2l0h+JwXyY4a852jP04XXU8nni1e26+nYjoK5Z4sxND
m2pSPMByTPKF5hZcwyAI7jvjbcpRgFMjRqGvBoYS2SvcrDuIGwErYe7UpwOmpmD8HAV04Q/AyOxy
m/dLiwr1az0Seca93/C3bk1GbFJJBfSaZr6fLOoekfLvPBqp5NFWtLQtLhztdqCe3FZ7FeYPIYMr
DickdcphmHEkdW5JglDOxmlHvaWy1UIrvxQNlA87bhBkqTSnaHwPNx3WlMUYHoZpb3+YQuB72xuY
L3J1PgAzplittknxLlWmUR/Ah9uUAvcYJ6ya41OT0AMvguwPWJYy4DYKS/gJ8gcq62t5raNwLNs/
Y+5tY9hOOgcH46G3dsu2LExd4lv6byADCjuij+l7gBoeTymI6AN6bfuxDLnZDfGqgUmHLgSOD7b1
/o+JOv5pkEk9CmyjXzp4WmWMwslhkjB2JtEhgHaelWoKB31mIJZc+g7TICllLwCHV7NYoiUmJhAO
jzR+3Fo1Iik6iTN0YUtpt0Awh34EpR8/S9FEuDp+sKJRycGE/Drd0enLWD3dVBKxQX1lsovfFqNu
ubp5u6ddIyyJ+PHIp+36e+Gfzal81TNv9SVSlqtcRL2l6JsKiX6Ox9I0Vi9QkVFP6prsS4bMW1Js
ixKpSIAy/SRCCP51Y+MPm/KbLO54TT1jvHdqk9Pt2Rt7/Jc8JoKb3u9orJ6Qcnz8Mb+9liMdP2nQ
ndfgtTdIpsWYWfWaDpM6GjT5DVsjOR9Mz07XvuGwrIaCLvzj/TcZnYStO3f05EQckMvynl72TRxl
1LqtMLqlJvWLHRyL+s1iSA6i4AJoQ1ECxxcBd5dq4Te1VfBQv8Y3PGQCIzZzMROKIdIA4zvrSAqr
AB10EyF/oUjx7RjwDjlYm5ViHVpU/RLR/vnLWBTB4rEQlJeRn8QI5oiybixty1OwTno1LF/sLIfk
ZFXDxm2GyHksz2WzymAoSdf7Mm0WOGbfbaplut2KkrHBEPuMvkSIu3tX/AH6Z96mgR56VeCl7iGo
KWP8+8jJfZFHqQlklBhhWKxg/DbyH0Yy4AjCWX/enc4KpKeyRRXAch1Zj3cUNbRMNrb6434mkisx
eU9xVmutReswnBm3wKArqvgVVD+1lu36QHd0YaW+iiYf2RF7bDYWnoBeUChZIxQ9sLcgAQiYpxTJ
AaYBbU+8GdHr8ASlxgpGnfv1QagfnR1acL5OOsuS1f4AxEA0iC4QnCFxKqEpLMlap2UVbZUiXtgW
sFsj4vKbfKXS9mdxFG/PE6STjLoWc04lB0Wn6zSbC9lz6FczwQP7F/k+Cm/P7N9c+iZqdAs4M/JK
ULPXrqCIgMzOCMmD7GIyk3Z5t48zjIbQpxN6g5bEKOm0GmzODDxibNrmTOQ6SK4s4VjYZ7IFTB1n
U2lOYv5cQHCV4SATvQH9bOmkHm9YSClK4wydHece7IXCWqiAEuQxYGx8xUV+BM2y0YzHT0J1OMVn
/QJHN7H8M9ER55on5CAkxa9h2NiVvbVHwmGM3swwt1uXTM1ZTi9IBd80Ckry6DYQq90tIhKMxvtK
AqzS3hGjd7BCoO1uRRu4AIxUcnJL4eaV0KYcsk2kboKftoRarHZ2OFOvQBSznh3ndCiRgF0DpmR2
a95KppIyxP/ASB085+F7BpGVWbWYwe6MEG1/b1Z9qNAmYAsv+pmOwMNBl+OpamWFrBg1V6KgABiQ
H4ROXCm1KMWfI9q2+FwGkhslE1ceZ1zx+Opqbbh/kqXCgJu3IYNd+lghl0+hTBLKOM+4KoaulZFZ
4VGJsB3fywVQaoJOpJDssguIiD/CIYUYeBlogwVXzzT7x9ydjpR+OZeqpJiB6484ThUw/ylSXdAo
hMLH/00i9MBeaemBfvrq/VyaEsRIdQzd4rjlWP/abFSsOC0gD5kWBSHMwTnA4RO4hSy7twgFTH8l
7oNqNwaz+j4kcIyXgRRp8mjXA19iNLu7f11pRBt9sovprCga12yJk/86Qcnt/dISruE2Dg0HdHgV
KgrPrU8AihTZ7DszpACJFFeMRBe0ut/N374xf/9RSgRI5nmF2bNEiVpX6kwq5iPb+C1Oo5NxIjUg
CXA1+L4ymu8cLXMBJzwgHtUoJv2O9XghxzpdcPf28L/rRUbxxCHZbbQMcje70Bn15EB0AJCAaSru
hdUKdH1s5IVp2HCB/t16tVTYZRjstHbeYIijxcEvMhkG/A1Suy3xwHrSPhULHx7t0IIG8JoNY4tb
5jgfTep7UabqgaymnVsn5sczUVWBUITRq99pLCgCMTqNjl1v4huEH0TaDf+yTC4xMuMweObxxAJA
wZgahlVQ3U70uy7LC+BogeIWmSIdK2cUpt1DnZvUqPhYC5MuaVxkGQUXhPxw++6TBetTjlmnAMeG
GJQFLgfs4uXnRWN42NPbOsvBeR4eyf7Np4UdM+upJYqDQ7db0YUnVQck8jU527s+nLjZx6Jt6Jeh
Ww0K1tA8NC2HUKX0mAf9OTP58zu1+QUEp+nBFqwpcbxYY+KN1P/Eut9ZST3hOd9eQbNNguD78Jr8
G+uVBFtTpljsrqXppiGSn007WIBZ/VIdITE8NLoUbyWGeBAEyKwW1wkVyLqlUxC+8FS8nqRmFLTg
RLoubDQBufhwyH8Yzd/t70Kd0dvBEZFj6tMae+d54x+IRCcdG/nmMImsZH9VYOmREGibNaVg1AVH
sYmKPcHe3fUqpnWra6bgmcKD0a8wWGYmTeYaPpdovmnXW6IwgV2AUsoBKkybCOouaQ9Po36LyvyE
mC9Xf7BzK80u0v48xJs/JnYMHAUpeU1PhKVwJEE0Pnx6ihbvp63qbANFZDE6wyMkUN/d6ko3+c7p
CRrhpiYVj4XZv49KJryj4Vz869znw4qoYnpKohfygbLn3JC0lFjwM9cxw+MrOvB+u7NJUDJ/GkeO
egpHiKKjaRFWY2ydClcmUxeIEkCxoU8nOMS+le8EDNI2orgHCbHW5/MiPL5b6eitbHVx185d4mNi
lYeqvfePW0Kxkl7U2k71c5avLteTGXaeOBgvo5OZQITMjDJvvImosZjayLJHPvtq5JH6b3uBCG73
xyodfE656dQs5F1jkAWcHnAVSxx/Ux1OAxiFyBnLEHZde7XewCC49weod9cLSdlMg19F0ZOR7XbK
+hbDu2SMimAmNSo70oIBIH793rygNQ3yyZXYuEPsnnoLP4uxE48T9CgDhCpAIWrFpRvjQxzqSFjM
fxO2B14+nqQ4h/1aMUXmDhBqfxjeF6CQvHXjRV5a9sMTkgxvK1uv9JMWsTwE54GFbcq+WrlOPPaW
g417arR35AIrcJwG4mBV/GcuCkNQ8xeGW6qGaGkJj4Er9AskXeNaVgLM1ozFJL22rY4q9fghoh9y
7umyqLVOzvbBwQoWvQP85195sWkw6I31PyVrNybu9Si+1zoPzHsW2wB4OhaXgFgIB9ZfZwIBf8ZU
Me++1Xq8Jg5zZv9EaYDxTCk3DiyCbLtxsEtL+iwNcNnKioCZEqlr5Y6bQUs9+mWgXsCJlRYFmD3C
BnM1nQ2zufOv/5ydvf1coc9lI4xTy3cu+3b1mBEHdO8tV33wiFOiT1l7lheqmI85wNm8nyBpL5sw
2mlfIBdtP/HPqpEALVguSnKbsvO9QkUKXGv3ZIZ//9U9nfwh9zf+bh3ihlgHXG6pNCp+juBqVxVT
kSLvzfG3OkezIf7gNQu1HxEoCeGbHlDmBpEKkT90mLCdMCHKUJChAB83zjKrWNVei9jnKy60Gj+2
WYEeB6+L1Ic0ynq0mHpbkMiHwTX2tIhbrUeKCcGYYilrTZp84AVMGaMR0ZzInRPAGBWYkADPXXAb
fbDNHBugf6JJGZ+ZQmA7ScdGvNYhjiVvjo8DAU+guhLAhzR9lgVB08A7Axnwd5e21dq4dy0TAsMe
qMKUuxPvwWx81Uct8MWgyBnnpfAs5E4NNDKIc/kImNhRno68ZzSlrSRNcf270kHIS2Sy+mT6O0hO
Uxvelto7TS3398gL2xlrXcnE/+oCNDeXOA5vdQ0CVCUj9BDxb6y7d2e4Gj9Ur4nlby/9hcl2ojuN
rwCYRy39bd8iXQnZQREX8ZfrPl2ymP4OFRPIJyiJGtnUpCdoIviDjzNa5X8lJQGUOZCAAH/06P2L
4d/uyEVVIjIq3UXfirJz2QIBajA5MA3Oc4nLtJj4YKS1c9gGQbYk/p2Bx3Gg3N/fNiFJnm27Q63R
WLPyz2rdWHrdEisAymi0DMzvootFNKWr3uvGsPJMQ3q0PwRhQ7HRJIVqjJ4+5Y3Dcgck8MoQpEHf
90ez56NET5aRq1euk3qokDOMsk2FQDhR434dIwei0wRuZy/FoiplclQgzNOZRbiB22zTiqcy60/T
vzNPtLpcgy1s4OFOJGsyJujumhjFTtvbhJ5emHP6UrqSSvAGghTSi1Ai+swbvVxb4FGSifJDJe1G
MMBpANhbDVHP7FauEgTzWvwxxdTCKEj1Z6pQYYzekQBX9TpmEr0o/1Tk0Zpck2stoGAMMj8WKXEm
TIfKv9+jB0o83A5d6LMR5kzSOyYCgQt1CTBQg0HtwYZoB2at2XzXA2GtH2QDO0R1borUNy3+b+Au
K9jThPkKYBn1yDfY01XFgwb7DqozE4vD3fKi+F/WBz6whQwkzJ8KkjHNk2PlNjjTmi6axMWUIsKZ
xqAzgBJegPOKK3gvz1UYKKcAWlPy0Zd/VsV3wJGVUJzLMaSYjrOI88V096c9y2Mfzjpf5eOJtPCW
GpYqSPIOraLd/dnJbbP0YY1wqSjnTs/AH7Nr7kjnfLmJ+9VWyBZVXirzyFNcpbSLXBmGo8sAiuUW
njg15mGG1uF9y9XFkzT8A67fmldtIwDroDP6qo0wMiwaQQthzRARvhaUoJ71KFrVvvszxdNEKAE4
w9XdDvuFn7F7loHlyYbmvnV0lOC1GdmEvZE+98urwO9Au1u9/cJnKZRsX8aERDYX5tsRISR8ee5N
MSbt+6XogAvJjJbZUeSrIe0yOaQ7SmON//HrVoL82+usiXVIvZk8IO9jkVk7D/QiswqyjIP4bJx4
w4BKDB6kS8KY8BLpEmM1IKdsZYAd6ANrZqd7hmo1x4QLtPDo6Lok1L9j5QE5sh7AS2v497RgEUY3
otI3ATnVyvNOGy1maveL4H0IATjUKIcd+Pt8H7GmjVp36mxA8H9tktM7jUZ4xMWhKPZ3obtpaLPH
+XyeJGSU1SapGmvtWAQ5oMcxBm7BmJzCRH1wppAUtsE/Y9FMC5XjT0020+XpVZzAh6gjxj+spqdI
dFjBUu7QjyZF9s1XxI5KcInKrwTN3ODVdD56Ke4R3LnBXuTsefOnwg9dEb/yh76EVrJBuVVPIysX
Nnt0r+7M9JaRfvc5ON1/9I2beHqquakpkuYwVLjYAE2Acoqev0bS+V8AoKajh5rWGmjkKxqJCyv1
Ui0KvuNZqWk3VT9IzWxEculYwVDUdeMBmNRrR1EycuLR7S4lqSjXjcPVdTa4fGvS0D328fQ4irTD
ZZ9wYnnc+fMrucIXV5K7sNBrRZke6KOlYM0uMHAKHJkkKEgLF2pKcyWW4hujCPDOHKrNaYoUy9qt
5PtQglIEyaakd4JghbDMdzYpxNbKW5nuLsNuQvuzTPZjgFMFxrwGfRtdZmV3n1wZ1LOk5yCNkPXx
se7awz85HI0aq9+I+ZKDaUxmfloB2nILbq4ulbLvNPFrwe1yjsj2I7MwdXt7hETTRPPGtJQjpkM0
u+Z6WNQVOHmj2iJD/0mtEoWfrCFundu6oehBCz6Xa+PniFIWC4OlmQg6ov/cZfEyv3oeiIMGWUpU
PC/LuWB2Ox2vmlLsmoZIXWC6nVk0tRzx4fAqfwwPHlzZA6LmVDroOFVigOm7xw7+FobkBweg6ehe
LO6g5cfdsrWv7Vnibh9ukhCAkfAKIzNghlDT+9rhOxYqo07h3Da+piDuiqRhAmJyLuAGFRNVYEcH
QWoFcS+RuI5eYPu9XXiLZkGMyrjDglqqllcaQbCHwEyl08Xm3NftuRayWwOI+OGP8yMZY66bqTVH
PAkb6lX7WhEaVu5hHylUNPs/1JGdZ7Ec4+G6W/8VV6jZmac2uSHJMYqVTrTVKLHy0CcObBaikkRc
MsvomrO8PykIqbhfTax6nBnru/BpKLybGEHsJocT29ZWebaI8fkepTd4M75e/HdEUyQfVWbz/FX0
BOnNFNQJtSs+cXxMqW+JYXC723qB93mH0Y/9zPcKegR0Af2zyBvbGbdx7GkXD+dBByPwZ0YwkN+q
eE9khNTZErIICeIbvPYsSnoJZuwjudkZvx2ZrmRuXwb6aVuNH3CxrS9tEtP6kuwnXCkUORoe+m5z
/0j3eAR+wOs6efzi2+8SWznNzjafJ0DDhQvDQ2rkZ9mTXxpn+frk/pGnEDl8dm00omkHXiyoOkNB
JNibM28Sr9o79SWID2rI7+buSmYXYwHmD5vZUABE2a85cSOtkjvZU9spCFdNsnYfvK6O2YbC7beq
0EYzE+i3nnPvIfFUHtTMFxL7jEmlb6t8/z1RyEj4vkICYI9YTTWI/ZBv8EfuN3sTVmAtC8EFcuZC
YkAB+EWAe9idlkpaA3tJi1xtm1cLIxJWt2KuM1B1c3Pfu1gRm7pfRIUPmgfhvdFoTQB5icS0l2Yb
xx14gP+p8dLK0k6TNCyFquCHrm83yiwmn7m6MlLJS0bB41NxII+JHfxmKGoHvRxr8+HkfRSboxf1
LehLTqnrgvEEEhhWS7//2bU3we9xOQkHAbCIi1dCYhKRy/V48D66Ir6JJQO+py0UALObhykZMHZM
5Zc+9CVo+tknPpSBIOj/DdeGbNohtupA5rbiBCUr5mUxlrWtuH1bRY8MKm6CnWX1bjnMQs1txrtW
Ne88HClYsfbCTrbdCNPDkJ6YVhe/xMWX6x3kQ/ArVHRGDLJiXwDm9UP+SG1Ob2bRRgCRDIj+uBwX
V1vjAvQ/4/F6Pi1pKfESjVQVjaHaMX5zNYA53BvRnyhMvqMq3pE3HIS9GBQv5sjtdUC/uetZijTL
EtAlOeltreIkJio0SEzd1EQsek+41UtXcDRM4rKR+9AI+Ra5lOHgBU5MKau2postA23bHuCqRIsC
Lfl1elwoa51BWEGD4s1ekvTcnX+yCW3BblvueflnuCoz8rgEXJ6OG7zoeh4bI1GzG1uTwyqsm07D
lFI0Ya9+rgFuh9RQRb/hrOpFp1aLKqwKVuMLD26Bvnxn+D8lWSpWCbXsfvg07+FxgF5tsKSekg1S
fV1RhsHoSlukfCHEh+x/Xq0IYSF/U78VUS2Z+2r8bEW55OgZstcnbsuFG77Aj/wQzLOsS9n2MNpz
XxtmqaRB6rWFqlSpEL3LuWaN4XQ3OrNhP4OnejwmJmzLTJJzOWDoSlID3uHwdD7yxtke69H8x4hR
4bPoKTRf1agdwkDISMpYgSJSQnpTXBI2/vjtzZH3ToEqaTWhqMUKGLl4kx7x0FJhajzlf3jwnRDh
xelFO2AmuEdrlkI/3KZhBeiz84XLf9Elst7yMhJoc0B2slqG0joDMZk+Hcfsqtvn3DTip9y2Eqbb
kXtaMKouwJVnFQGpQ8We3wK175ya+cB9qtax2yf3T+zdDnA9JskHSAxLBqGSmSzRu4I1psgMAefK
PpcjQNzIoe64SCmheNCekfIj74nTWREEvWR/Ruq+f9Wr6KghAxLMz5G2JVAKIzMVkHdGH/oNOBp3
fu2kiAN+uBPzvRUzQjPpYQLBuqCzWN9R+YN2k80WXepo/lbzyiOBe7EeeEJuCEcDPSWPbh6L33Ye
aU2Cy/3L1CM0GF1ddoUyjD04Riow90mdP8Ms+3TSsZmjVV9gY/YXZ7fqbvfLQoPsSRf6wlQkvoAN
h/XhmmIff7cNoggm6GgvNED0P3LB8ivkrBSuSOmIxxU/0pTJM56IOcnFUubuRwEPL1iwtYtBKH1u
yOq3uAo8hiPb4AowiPox65N8X/dYreVf5SOIB5eygr6HiKs6ZY/pjJm+DF/m0RYiJfRcUwEnXdJF
g6c3PjpChoJXvYHy45vSkuto6ZW+0/yKzjkZPhmN52ZbxN9C/y+/DuDO9OR5jkU7T90s0YPLT1QF
Uw1FxVz1vB4aAPNStKV8aaAKPK65DY0wzjNHktV2REPrBqldiGqccqHSTcj/hpaxRM7kOQzqPM/u
/gdow4M3kLCAcehxgMNWKdubR5yFl1gV5IgXXT+2TfUfjhyNTiAE/22g2moE4tS6edYdzNG5rixP
xV0ng/WuKOQZTRpvl+aRr4Rk4DyPfis1xUCwlyRTPxfaxreCMq7WdfF8A5be/Nn7BCe4Hc8d1T6x
emp29fD5j/GSYYAxrREdx5nTi4MqZdGBaAxZKzy1CBL6wERJXeUtzTqMRfE6g6niToUIyynDa90k
Paiy3gyV8NvT85htBOGqzz2GPmUJWtfXAIMlRnOPMmVkM5E4YS0u73MlBDAjaFOD08sta+mWa2Gp
x+pgGwISgwNcrNItPrQhKpbYu+V6MfvbW3LFjXBIho7x00YNz6utGIkjwDzSoL0rFLQhWTokfEv7
KxS1pBIgs+719ORdxPu3djPHOqXz9RAygThVwigV1WaGVyWwa9d9Gcrl+CKgX1E24pmqIOScGvK4
pUENVMNPb04bgcK7hfxHHx0t1aCTg6n3IhdXAmD5YSLieVAMTubq1+MdIxYTVPfyrqoPcXyQGHaE
AZwVS6btcT1InlcXtFatFBMzy4ag/brS+vj83ZXIYG2yj3eFUJd7VXszFpvV7RKVDP9NXWbop2IW
j4ko1Q/r4RDMAUOlf3brHLXVKuLwQPn93Z4+xEhQFyj1AQg2vBhcvvoTvHoTYfiG/pUAl5NyWqK/
5p14hOz+I791BkOdeYuqQOK0rJQ2tuT4irXnXRWaprNW43wEl/6IkYiXyITrHdGKAFQgSclcY0bl
8I5nyrcva+/LBg03dlMaacy/e+/QYUQtKrUOI6c8ekA1d/tFbSuwGWboDddNm8CzSHOcRRhtP3FJ
+C3MA90JMvrksGo9zd3LuxEAjozrI48mjV5MvNnzrmrCRB+j3YnLgCY3Izn8sX6YHM1l0zzwVEG1
6QEPCvH9nQ5kJ1bhUsf/fRzg+vrJfCPLRMM3ExZFos5VBR77plDZoITa57dTD2bDpothbLMUhknZ
7PuKmJNrZznYGomjceR56wdJWsBZpoasbAlakWxFO+urH0zT8hqlgD89/SFBqsup+zMHBJEYxz9f
SWuzBlRPH+OoKZqHUgacoOIYh5NpShmZgqi4InonyMwFfCg5XFXGAORPG0ragx0RI8uNWHuXK1xg
y/01IhyUS/XDGJp9YDpyd2dXZbhE7XFTD/HL/kLuR8ZoMPkY8bpHn5zCrPyWT5qavRoPROMV7jSf
yhv/povc1cQ9j5+bhIcsIQV7d3Q371uMAtVhGkMSmrmZT/DH38Kztv2f9aY6xmrFh1L1pVUaiBBG
9dhF0AsvFiwSUBeMlWulU2DUa2enwvz1sbvgToe3Z/gVPxknu6QZm4INRnouLwqym88Ryfcyhx7q
rXLROO9yAezVbZ/k37ch7yETrhMB2A5oFvJD3OCO8zW6c7argS+quTDUoZG2v0Cr1eADZRz0jVD4
NxJNfB9FhpO9GecBXoHweWalMkxZ3nRlSYWFfVLN6QYSwcs8EjYmZ0X1urRZdqZTZQkQPwjD3lsU
Opk7K8dC07u+I8yaaLsmnCh/dfs8qAK7xFTEvDfhLdnL6317ktu+H59/BFrFEXC1uW1GxrizcOqG
LL6wxRXCoS6yoiEviQAEQ6yxkQzNZbAyVJ648q4Sa527FUZKFhrnsm3haIhpg83U86jc9i/2+UTT
/RKLk5wQ8qpCR903VsSuicO8wzPeDGPsPBUgCLFV/uY9vEftSi0a/eXpESvMb6gvcXF92psyTsPM
uqdXszNXKAjcSga4DmPzvdJCUXQDu8qGfBPr6To3X7dUv+gWIg6jDu7hDz+DRQLZTMISuJ1NXQRs
CAoQ6xB6qeLB9iyv2gjg9iD1py2uT/nBbLDILNY1EEoNdoi/eXEcUZ+jIzChsb/vY8ShGH4eVlBp
amqHmqC/JLg8I+247RirpWIXeOGYkIg9io787KEQRRN8pw6LuMiXH6c6xqMI0dw9upoL5VtE2wvv
reKTnEjArCi6rrZoQOVSV5eT+AnBkhZjrL0AfNTKftMkBnlWVKt1dLa11RTAsAwq+kwh9fvtpDO/
sAqv9CBr9S+TttYF4qHz6h6AedVJTPu7RcllsGOqVawH8tx1WdzrIiMmdQpT85HwoUkdTGo0u7Nb
yYAGzBQcSU/p1eIIIyC9kf5Z/gUclJPR8kKfmn+xUkcUnoDcbp9SMekDtOdndOpzN4Hf9SLCt7Wo
BLcNuldit2nf9B6Mqe50tx0QY+YiuXvg2F8RifVQUOnSIZP3aYvO+qvh2ElJfmglXMGw0dY1gM9m
77BDI/odfesAmGLfa6uxIAOyXdU/oBW9ZgE4OyxsWihRyQgNFXgvHRYZREEoihn0BiGMjHCO9PE1
/TgKa4G5tvFO/ir3fd6XJ3aR2GzN+jgBzxo9D5Yk5jeHxxref6m+F6WagxYFKCDkiZGh5ZtI6OdS
whfZ1zh7WfE3IsgJEEHoyZzByR86IMU0k5ERBs8XvBKyS2P2gqjqO5MdPJIAcLsMEmvsZhEMoEEc
v6WLonPQTR3TS5XamytsXo5a68xFePr/qYSxvHbnmKGPI7UJDlUBg+2eLr+K86bAbTynrbK2nVJb
kheaEyKa0m+qELPM8hYu8lM8Tv+qGXE8vowO6oUpujnkThr3ilb5GD1QuryHDZdN66WaxBjQisp6
glFXaDfJ5Ttb4mC32paK82h4by7KcHC40XFFH2QS+jrJW+Xz7NoOVNCLJLhxRTvlfjIvj4z8JWhA
Oan4nUOBOzM0bZZExWXq+6ngrla/LG2o/M42bgNmOUiIz3nXkV/1eRFeRGB7ZThal6BNSapeFiVg
t67st+bZ71m9F2054NFpwxHJomoPMTAAP0Da6fhNlXzAOhvRTJkAs910ExGBVD5mD3DOVQq6zVVE
fKWf+iO5xPSH8etGLVLGTKenDcJVmP9VejgxGqCIthkaqmtM8fBt+t7Wn4CfVDNMq2LX5LcQLu9d
aguLxnbL9bzBhGFbj5JnHjaetbUB/GB2+ncKybes5bX84tCH0KDBQ7c6CAj8s8BwzQP7cIltU+DT
1K+ivfunDN/zyXzRihObRTaQnWIVKPuB+ijrlUVe065rWKD1PbqNJfsxQMwHN6I7l7vwsl6ZXwkJ
hO+1uMboYABOFe03UIG3TyZBF/kMVj6Tg0SvY7Ipb7Pqyh7NPE8QmlN4zgFQuzaFc+p2qQA1JPAV
cJQAH5r4G9JkWPrEMH1j9Pjm+U9LJ/S4R7Pa35oyilDEms7XtljREr3QZlIOVkLcw6pPKTvKjeGC
zkaoIxY15E0XYBP1XHOYxgd+gFYWwm9bx5EymX8LBL05RtmIv+e4ADWP6ka8FtPu0NrHyXqqqlen
khUSyjzIZ83EU7Ugs+Sf0czujhm5AVtHKCZun/aAOO20Ym+Q+Q2Qyi1v0ZK4Mu7U1qPVut+dYWaf
D09dM4WzZuJk3Xbgvvs1v9nL9nbQf6bbxj6tOiiXApVo4sTDcd8zhCShpSVMZD9XIgCDajU6zGGb
oX0Wke2zy7QZFdrNuGRYwoHwiTKXwunvVYTCWsYJBFXRsUjK7YZ/WiV2crFqJmX2cQhmgGpkRv1K
2y8gFysQDzql0XGhK0CcHVqxLSbS8DLFhEZCOkhg8gavv8bxlQb8DeWjn3nqmbuOPjbAl+B+X8++
1ldkjeZGOBcA6dGuSoKjdEKVRQNPqOPvMtaIG7dVPPCFzL0JPReuOWLHlXGaXrulmEHfSUKEZr4+
nwH3WCaRJG9LIt+F9Z7Eazatm+i9kwtw63XTAKvaK6x1lENRIvTL6dSBaOMgFuOsc5ehWD9uUQzn
wGZUNF9VyVOdKkpUrP/awUpGSBnYoAgeYjEZOfALD37mzyxvlTPb2f/NvThyluk8V1jc5TC6TSqs
PKs+JVoDYBUBbJn8urDE01qABCBFdyHVVLFFVUMqOCXlPSUBziag62yK4p5Y58HoPXqJdyJyJcyN
mqmup6IdaRtC2iwkNX8TT5SFb6NtlOCgEQX0yOuDyTRih0wz2mehgfyPbL0O5lUpvKB/Dk6BPCTf
wrXhStgxVltv4gDtwrupc7fyTvtqB0Zk0dDuQO1SUZw+k5frOhjKBc64O4xxvPZxtnqa93R/80rz
xy57Ta0psr13Ioq9k7x/5eQbcamsBTe2vWtia/GYs0VpRLX8r5ugM7zNuRzBzM9wyiJbg248kxK5
ucz2me7m4IZqzLV2E8G9gYfaQ8tnAe7FwXRZHIuGladdd05Pda65ymUGmxcAA6pbzvqrqdfUlQpd
aUg3RMNAM8Qd58UNo8V4FWsP2k85MrfXihGAw5myBJb8Kx/Tei3mQjDjfNtEkp3/clB6TQ24WzDz
MPHjbKhtJm5VLd/hhbUVLNRccRVoYMd17F/F6lOHXDwsrG76sLlUFEacq8gO/1x5JUd7XefB2MB2
CaZJpdLao+iDIGJ+xUza50fo/cMaHalufvuIek+YEQ+rcS1PMK5aMcX4pUE8r8R4mA0J0x0fpK1p
w4zDu4nDDwybpZi5NzBNkA9uIkeu9dFdKP63z+5Vxi4dBKwsHwBeb53s/yGX2+kitTXRTbwLmDBZ
SyTkRd7pRxZw3Qyp74eHa0qqgrvpX4oI77d/Co5fQYQJYnRHE2lVBid505Oq/L2CfcXS8v5UsVLb
nb3gJkc6VzlikdGZRE6DSfCrTGXtyQMeNis+J1EdRUj5zKT/Wau+ICK5DMCixW76OzVvk2MdDBLu
ZHgaLInXGEiKiPRANr7EkMl7tl6b+0UwfeSkm9s8d2m2+j98xslv6gaGDzlLb7IkJliv1QHKrK2Z
w4rdircZYqlLzxAQo3pqtqJJv8r/ENofgwQvcJWNps0yoJZV12pLgYKxH7HCPBGeLysaAaKvmh1l
dJ94CU3g+xxHSzKKcZfZ5VsQp6hUCMXcGTSHlNJnxOU+0FDG3BtT5Rfiejqj7iESrCFPfFyWDaNf
eiBvbC2l8P5m2ReOblB4XTB3eO8duvfaHddvBbyMk0xfrUOkvYeUgzS+SN4icwXeXLvvIaLi63Hg
/IUXswHspsCWhKzOuhWtyzNCEhZ7cljsc7Q9uzHhT0iGKBnEP0Ai8Hvan65PE+kSWbJ8pwVHO/Qq
htkdDy/zx56YuhAuwuOQEvQNN9F5+dQRE/FqTzws2RqZGNqkMNDZLYfFwBXpb1isK2q1ozv/Pr8O
n+6vb8qoeYUCk5HBeO8mww2dJ+YH1y7UeEmx3rQbPh4+bfaWYsja/UxNFS8Pll2YM301C5PMfBPD
GVxty0MjSS3UsEJ7iMmYbOHw9bv0tmVYlg7Dv+VkIKAGkAGHspDtrk9zz4x95D77aVO7M7qOOQhF
cpi+fKNWENyxZQh2EUMGV0w5cI59qjoq2EEt5zWx6S5/PMCpBqd8fhOX/U+3INASwMHRGqliIo36
hz5q7kvKeRIhdZpuR3/rS0T6KeRomUKj0wEdG7CIf3XKNV7Pmw3Zox+aSkMoe1y54yBmOooLX/gr
csMBwj8Simkww2umW9wAx8zn22TqlK15K8RI2ayvciI07X3Pn+zL3En3F4j9a+VoFb+4C1PDH3zI
whRsZ1USxiLXxMRMqi92RB/QBm/g907ryLPqtROh/4TbqSLeHRwWDZjQP9b8WqpGY1m9syIQURf0
wkfz+3BQzC/7Z0x5UC+81vH/WHR8p/3QYJAHzEeVNm2Yu1BxxILl8zqv8+z4cXosQOzUj4zNSp32
CUxWnmsXJeeQow3UaWDboiNeiYQOnuGst6AyegPvRDnURSJsNrI1l7mu8cTH6clR594gVAw6zNBR
CuTPPOoOTQXjjkVtl0He43MtXTQU14kahtXGVBuLOfouXB9nTmcsWIDuo+9OGYgLzgd0uzn6nibA
4oRpfGuBJVt6MH5hUUDGwYYt7cRQ49KpBzYIIBVF0TX+3Zo2eDbohiUhJgtysVL40q3shYboTxol
XVBoxyr5Q/0uyTx60pdkKQ+YwZcRzI5/SIBDWqSgcipt1YAg21/PTRC98dHgEuogrmP05/JSPl9J
MWX6eUKWFMXyo8G5g2EghaQGvHcNAgO3m3+oBhHWZQ75gvV8G4ASzJgmVn803oKB762lYXqiyIn4
N34YmRyHIlGp4LqCqCxqWHU1LBKitPYDJ2StfTXF5hmPrV00Bu5X/GtSEARWvGobqhg6kqoxDyJ/
TBRwzULC+IL51xX3iLI0GasQLsqEQqiWHGHpkxck6wLWdBMxtaVV3GNeGari9S9MThNYCQW3nA7M
laU9dzBVflhWhP5hlP0sf45XaiI3jA0deFoJ3xS6saIr7XoWmMn7aaDSbs/ggEQwZKHRYFqpluEl
U7vn/XndaTwtjX8Zdxi0wHye7LxGKCnrVjYsZ9TzUoi7PX7s9XuoJheeSA/0b9YuCDkpVhBrULW2
6V9LSgghB2PJ9PtNTne8mojCe/QgmugHW3/1BI92vnUDnf8W9OhmpldxhxFGXWJxk6cJdiIXoujt
4TGxep06QHkc1c8Co+S8tI6UGAkDmrUVhHMhAowRxB8Mp7QDGje71vragKiJ0IQdQ36aiDC59Tv0
4z2dXN5LA9HBlDi2pQhlZ0+xha0k2eREXYrAL9usAzl0v/3Fs+1C5cpaCW4dCDUiW9AC9HcJObiR
x8umrK/42LrzsujJ+MJFNReG41ke4dVJindTq92NRe4tfj2mx4Ad0nTbtV1KvEKBuuK5fGtwRD5d
3qB+lrarX2bkrmbUTTk2zlhlc3Ha/dUOdYB2tk6w6XlWlekmO/AyEfK6ktHT2NRE6EwQFYvBs0lJ
gLuiokecDUfb3NmKU6LsOebIi/AWGWcSXM6sNkU7R6EbTPTUo05ptyflxqg4PFuvutjbFpYYpOHz
LMsV9JbXwrk1ZvsWSvuJPjy63Aqx4O5AUS04kOTS1yv0M7uccQI4BHpe8c0TpRaw+dL1yce7Lz4n
zc73gPkoa6BjeK9lrPOd+NO1u/PL+hGbKswg0fd2yeO8o9eSzIxMEtPbKngiNYcJYGxIYf48xz0n
+fYqPqF8R4GWLnvmgc3faHr0C8Q1SVIE89qRNwUSPScuprMuQYQnN/MzT7o3rFr2kYFO2sZxQxnq
XwfOe/rf44YeiFeT77y/SPTJQlZaQ/B8t01Dxx6WN1Wi1NWWjTVohP8fptCR3PUESnSHVCIWkFut
B0PD6mpoUHad3HyLTFIIkdphyctIxC3cdDMaPG5wj94ivgHxx8ItgVJpE90AtJri3h6X4cwn0xoT
dpKe4pbjQ/Yx3QqbWC8yELmFUP4wDmOVGpNlrF6XQnNcPGVC13Vh8lL5KWBQHwGZ9JEgcDrthgxC
KIHnobgVFessmvi+jw5cN8ZLskGUpR8ly2DbQ34mpgyxqPgnep299DUwNJSXpf4PHq+tUBiDBzuZ
Yhho7huMDgrxiFwSkA35AT8V2H41dmK6MopGmM4g8VeEHKxyizP58zny1d+8efJumU7houkjs9+b
pV7XM1e6EXXaX1SRgN6+dLmcmkJIzwifzw4JcZPfeyLpmLtw3X/AxdWxMTx7XciEmiN7oEpzFtb1
mZVXU+RPUJ5Aa57LWj2VCo8c0Y325sZGck3deUJTwQYZVxL/wSsAYuuWPqDe1VzhiPsnMKX1pGlz
wShrmnZzXuXugZAGSoXb2hu9KKuM4OKs8J7fO131/tYh5BDlKtPHwSd2J6Zz2ZOLyM7wm6CtrGN9
ERvg4GTnN/5p+cEWFVj37nazo0juBPq3Vc6QywzMXdrsV5pzaMAwtZZ4s1HAoK/E1g8od4GbeWJy
J6vnN/gEDRkI1xVSWKdQNFCWQg3ucXPkZyy+xbPzOgCC58wFyUdI6qL4lsfaiYXjURLX1OgQz+Sg
RCU2qNwG8JtVUGOr/oOEfCwZzFKuPTmq4EaUrX+0PBcdhzZRQs/pMoUfnUhB1XmIkNZZ4+Yns35g
0AlP4yESYGq4W2K9iy3Lks/d3oMnMJzsyz4zO88P2PWfi4IoQ3s+s4EMyQIS3hgxG1N78nG18skW
NsYD7EEgmCqZt4/ENRwAOEk954634X0CwVgg25c8QyOmLXSD01sxcBjJPuE57qu8iQItiAFrpqQd
8SvT9NtLYXVRxjGtpaOuBTN2ZOL7DKeQO3xUklL4qbRZSghKziBEd6b3ch+XOR0HETOUXbMlHnu4
Kv/Faz5pD2RBE5Xrqs8ivPxG6PxiCHAQGqnU2P08gISjVtZRgZy2lqtdvIRTPM/r2AI6gZwGGjYf
iv+lRPl3/+iig+CBRB2fn9a2iskcTP2x4awy1PHWxlrzLqJKnmGNQEWIaFwpuRf01aZkRzbLyVgw
jiA74U0H20ASkUJZ518rU2WegXNOfuIhTU/A4r6cK+xJ1Z+ff1DJsdZ4FKro61HstXjitL9vSSco
dbIcY4YSsDYb48tdBfrQ9La0dBGzMtFwITMkMSGCx7MwV3IKjyBIBBmJ1YOkbyel22uHaHith6WR
hr2PfwWscbut3dGc8klsdBcSm+cYEpoI7ZHi01HtdwBGWGnUygRAH2Ad3Ls4aSb2YHAJ+2/a3JLj
yJT9qvADxFGRsOIEo6O+mtSPC7/piScfoPXbZBa8tTF2Fkoxp42k68yY6Ju9ySXq9ZVuJ3hjHxcf
KA5ATRYzWXp1g3yg4QGpaeUR7PsYNA+vptBql64G2xNFJSDZamOalD0CB71R8OB0AiUVZWFpcPhV
mWwmPYq+SsEusIWhJZyUy/hYyyP8kGWWDbHyaO+Ty4feM3ie6u2fhO096IPP6/I1qLrLbJ9QhGYa
ReRANcnhyCYiMjPnjKtEBb6zMmMxGcajR9e7lJ7s/OWvrezdTrTLlQURRMu9tF9s+SHOfQ830lzM
C5kjg8ibnQIH48XdJizszOooP15FptKarEeTFQjsgq31V9fVhZYR7eg7Mbb1IFEyhL5x61s/pnpE
it7hwPzpHM/kBlcc/e1P3llDNY42NeneXjSL7/848yhEG07/pustOh7AMLY6QGKpk3Hi1wruz0sn
0LiWDDiM55qXsNMEGa32hHFKZr+yU2VosGPqQ5P083YC1D++I+OVghl/Cj3U23ug0BGjkcKufmyL
eha4p77ER1TgTlcKXYfpJgVUWCAkuyii1yVUcrUeXu4g9Rhg4+sEdY+1WlbDqm0Z5Bt1zPnw4Roy
Jkt3nNokuKpGXBa+o0F8sn4+JsqJaUMTG1EdjtkM3pjJy+VQBFEINnp8qBdRl9uC70v+jqBJ8Nde
Nf44FKepEpYAqzpvgkEo0c0GQ1+KSQN4ZDuoyJWSdY3AMkBCfBNwJ8HjTR1YjGGdzm3yLN5BguwA
WTZ0j+cxQXevhF6HchVrgpZqINFtpqVn5fBrNk/Ipmq68o6N6AcY3l4VSFnRIdDumuaclAyRubb5
wDi0vT2lyBmFlTN0fXeQ32I4WKZgEytMlQYByhMUYSnsg0HQppt6qqdUeKzv7kUNjJYJ0NdhSOou
eDNgNv3t+S6jRqr27xxHlPfaglNEUdEcGyW3iT7QkroztVitSom7yiVFKPb7kwiD/dW0nNgqlD3g
Htqmkx54J722d0HJw5y0G6WLLRUFv1B9Lk7oTPbp4euRtNGuE91V7IM86yC+DcbQw6e7VB+RcQ+T
SbjJVhDm9sVmDq2+mlFYHESVTmra3W9NVDmMtCEzlweN2eS4sbMRD/UTx0bt+iO02eE6Ci9oIKx4
8b3NsbmhTzS3U38NTpTW9xjEJdekfptq/zPyDbaDrPFCpJ01MbNLV7tId3GZDYdceWo6zvWykZ9I
xk3UqWFdeMs7yAde5tUJmSb+bHB+2+XGpGx6nE1DOsEcG0NiqPMY3KL8OzMyz9zTfbHu5uLNMjct
qeLp6OvHj9MN6+xXFlskVxNTh7YnqW6vGxhTfCxYTMP8p46+Hv3YNODWEkoJVGG8n2wDX2ml9TBn
dPHIKWXjBwp07LXaGUn2NOxXHT9GqUPBWP7d7uy2kcxTvPKILnBUH77CF5sdY9+ga45KxiyDFccR
EEmhdFgIEXpoP2GPkbY+0qVeGYwJtWq/M8KpZx5jXoTTL/26LqMQJmykksvHCdtf1D1LNJwnQT3G
vNc71A39mVMNefffansr8Ncdkaj9L3ag50m8/yE7qyd3K9jNJhER+YtN/AJ56buoPyaHJfB8IV/6
riymye5eP8sXNgHsMSmCqCARwtqTI+Si1yBKg7OHypjvW3qtnodge6XY8pmwqzrqYZ76C0PmhLg0
AjGXUZqM5VddK7LKGfURA8/Ewd3CNXEMgD+t++7GWitHH2FQiS5nh9XguEiR/Ff+HZjeUterh2On
L0f6vDZ4auwcnBl1njvnpYboZPfQFoTrZZcpkA+Kvg54UgaKhSaanB96hGhF9gTb6u/KzcKYrxQz
veP600lXvwit1D5dYydh+ug2PIr0NAGA1jI9hPh3nhyVQ3LO4LFGbuwkAN/krBC7es3LQXK1AwMe
j50KpbtXPJvTELUgK2zqcsx8MO8lNx/hZXJlz/MIeCb3xrVFDlS9jGwMfHJ3weHyE+ywM7sDXg4S
n6tAOxugCGWkAQSLPwExE6U3znv7UiRxBdYPEaffg7aqqoUVT1Lq/u6JIxheolXc3kq9W+mWBILt
IZAq8JYsDiRRLz2rLNxdgd8ym5AB3fylUKSFkUa8a5m1ZzSyK/9LCCEH3U6vMceZ+z07YOdgoDId
QgBXwbyvKc3LHDEgPMMIS/ugkXzs8U3KiImCDsn/3VvLj0FmpITInkWkzjVRTh5kBsSN4W8hvCBb
mcQBfAf/E4QG6tqQYrR7yccjAHXxfEfHJ50Cv6uz5BhBEn8UvkuAC/GfGGWyHkNB48vzMEeJM6xB
Na0stCFwyv8yB/DLRR1/vUVwzNCh3DrFA+PB3XK8em3tXAH0MxjLTNUNiCR+AZf8tLb0v3f7EVen
JWBlTJw+2L4UJOqTjLpmci4aIK3f9YgKFbT/s0WqTFpGe08iWQORjYkgJici37XamZuzB+sk0c7V
vjJ9rRCDNvBoJCrTphxRpQE4P/J5WSISgoqdAXz+KDPKbvainutPe/DVff/WgjICFO6UfWyF5Tom
kepocvB5Y08tzNpoeBbHL7KvNBp6kSiknznhQRJ8g4HZiSgDzgj3DkIpxlCNjbrTNA21gV6wnvWD
oit2Mv7J4DMdaRVBPpPPT0yuv8G7ynf0wA+o5Q4yMP6Owi/XFShcVu/J7QWxCrYt7eOlpH0I2IJ3
w66jzC9LXAkFLRLBpGbJD4nYdcnAHulpeevZ9q9hm10vncbgGbxdwqmC46hThtKYnFJz80tAB57W
1PdKsPwuLrcxK2ch4WwoLohpeQ0lfLpht45C+xAomnHpN5LCvmanQTy7KeiCKU3MggtCFVeSu5Px
bQzzVM5v77bozTAhYdfvrnwKwqyGFgxJg5Jo52wIHJ1UYXxl+D0yibhDCfUa1wvvLUI9hAMSTAGC
CE8Klq2rWkE6uNvBtCT9jnnxpXWnHvTyxvIUfKPFcj+8i7w9NDV9QxZRf3xE/X94QCXc2iljnfA0
INzfL33182RyWgMZ0nwPpGPJ/N99KIUTcRq4s/v0E4o1H8OnSaATayLK60GHBOHkiVVE9BDuWBmN
cIXfZTRYSJfl3bsnvupg2acl+AFJ4GdboheX/40XoZCuhpyh4Bae/jcQwmlCip/A1tUAw9ZkW3lX
09kYpNQ4uRb3v8LmrKjw3SrnURwh0UcAJA/hmFsez+IrQuzbU3eYEHbudEgjd4L7iDK83ufVOFVZ
cpKOp7v5ldN6KQ2JbepS5/CPi7zLoL8a9zWCjHB/2gXa1le7963mExCN6hbS3opeuZd6NHz1IFbX
rwt04pNqS7ocqZcBR3ipTCQMdaPhq2OPXK7b+j2ny6wdsv/3pAb+RQHqPA1v6Tis0KYZR8cy/wgE
Ib2eGPUrh5FveMX0qeXkhR720EB7ieahJAO0MQIE/ZGOsJXjWZu6nQnZOnXEwyCpjes+zNMjB2wZ
P8q+xSEH16D00YgOPxD65Gg3PViz+ziWwYKq9OpgT8u4HsXvQlGxK6cN+cTYELO2QO6wDJup6Uvv
cJVW8P1Ggzg5IzeWGTn0QGjAb2+oN7rK5AM36f8FgZEA+DWzAq8yEwuKMjCJyrkI7/fE6LSobABk
0b4OIYd+hnFpkgm/Q01JIZ7+G55Vn0lQbQtqeBxw0eshPcYCw3Tdi4xKA87h+Q48BC8Xm3FYj7iN
G9r0ImqMp4pRV1Ojndq3cSOuY5n6vODQVh6WnGA3ETw+o0Zg7trjLJwEi04QWs0iaa/HNwl/xE6Z
SMcALIh8R5gTG5EuFrZs58Yl9M6WQrsAFoJW1lwKlqmmTs00I5pdYKcoBHwf1/RiHfroj2dd0sWs
Barx8gynMGk7vmlUFZlfA9LycEOFimqp2EjKAu/m0RFJs8eovyrsxqtXBTGRgv2j0rWNikf983KM
QCiEyc2HuuU66254XIGBzhIDLnHM3AF4W8LBy8R1XgCB1ETrcKHYMf+SH5IM9yytDttMvoI9Qh5K
83c6/V1hB+jqZ3ia1cIgl0Yer7EPv6ZcP1jVMEIdZo6J4nWoOBvQaFvQsly9i0s1PB0nh+HyHRri
c02i1CYH5q7L6bNurw4uJZb3D45KzZ1ZVZuFYQBo9Z2fA89/wvpvZ121dSyUeJRF83CSsGzSeR2h
CQbydz0TaX1oDGY6bDSiPGNYf5bx0Gf4nTIFxch1Z0FFAFyfWI7u0YIUFkJRo6D9MUh1nBcAbIlw
91Q3HHw83G8dVB8cnbsv6M4pzKtt1oUikiXl6bjrmxXlO6VyMMTiVrVj9PF84McfrLxwMkMYEiVa
EPDpICAEHe+18M0hQCZE7L4ma12gjlx8TuboZDkbsy3Uv02qoCp6fcHtTGAHCYNj2MZ3DXAOTT5i
YNAToN6G3onWyWURuPDi19XniIpR4I8kcY2cbGiTy6k2KU8AoVeo9/IkTrMVQaIZBvOY5CSlHuFz
mRSUoVE7yHdmGQOF+HIXYVI0NV6i/wEekRg3uXQEplUAyg5U+pPOEpBVGhN7MNLbg7bebchr2mLW
3I5SYc7w+hJ3uVW6ki4UW/n0plYv5MtpRcaXsrjBKMmEHevN62Yq1WJuvfmxiJV7GZKvUyoMvfH+
JJW+p4HxarOCoV2EG+3NBi21SSAMy5GJRIaFT01E4hrr/GasHh0TuuBMOPQa2KvSq9G1qyBvnwF6
KCG+SzzUXmvUBrc/xYd7utbVqxOaX/MjCpOMzstgPwZZNUG4K4qRxvia2tuDrXL102+cZHbuKWlC
9DS6oSwAGa3m5JeSfbeL+IN2TdJA5tY9zE0d5WU1VytFvhX6Wn4mOkZWi1dn2vsx0j0DbLC5HEPo
iGhsHHrPhGInfu8Ye2D8JhgoMg7WNDrOyHMvmnjJz81CzO0kmhe8KweIrVCDE/BXD45anSOjLXxB
GwrAC6Qij0fD8HGjIEfelYWBU4y9QQI6+O+DtFTF7GUd64W4RJUtYstdYo1JyhvxJqOWABRN+RKG
Th51Jv9Htnc7MJZZHFEI8NG7BtJDoGScZXOIDR5qLkod/sRQoGYx3OzeFzzUUkJDuMZPC1bKDynO
q9i2gc8ewH+fdkjx1HDwbT3zv+JRxKRJQqNLdSLgT/y0vD8aesaSYdNb2ljZICXC1VuZZf6Y6m1W
JPg+zUOYWoykPN3T6SMJRbwu5dK+EqmNvcAZNJd7b/gM4NFuysoDJQX0L9jSuOcqX/LEIDFGbRZl
lFiPWjEmM77YwIhTdG3B4SN3Rn5AU7AIdhawLrkZ8q1lGNXCbKBO+UxT+719GtB1AqlGeLARYHDr
TNOlQ4jDiKiEubDlszBiPK8/RHYS7avZuzFxNDAYXboTHnGUKkPrGR5srwfNpETKots2JbegAFn4
B1NGw378e04hTD2jXEgoRs39LUB+vSHxtHoZt4IsVEyb3EV9DnT1GaC5eZOPR6besB61ThkvMujx
f5zOG06V0qKoUOTcuGF9LCFZfHVTACL2owe+fcU6d+U1tDa41coklSchh+5782tyEIbL+QNc/ZPP
pmRy5/EjS6fjfAPIE+VteWKuCKZMHD/wX/Fn/n9xQWR5Z7tGk3ul3/3SzyUwKNR4dVUf8PFzeI4h
x4/n7s+EqdJFPyotSc+3Ld7lSVxRG5OFGX8z5eMIM1YBFAc/zkOORGMnNa/eLbWhtxA4pFJe1UIm
6M50O59serclsy6kFjW1p4M0yUT/N3AUW6CZiiQZJ3/M5uF/ohszRQLxAlCvpGlStjRZ1g9V5rkz
/3etYq5Qv6eshuLsHFV75SnnIPex0uFWEtOP3D+tbymGBfgcH2ZTPvHT4me2+yqEVMlYHp8fLHTq
x1anlVbYmNPnwtI3hz36egcYAz2vwXT3tYPlQlNgn1nJC48rW3jkuvj+rTBBPy482GTuuQ7wTMyL
yDBxntFXuNnBbElgPa6ZJpmfqwi8bhTyTuFeKKDC+/0fLljaxhEu+kHH1lww5p9iYnb7iUaNuTjs
WFkJsx3PgvXVII62aajQVNUUhrcJOjrc6Wu8p5wWSH+AiDi0mfcMZLBuWEqo1voxc+V4YvubIyQU
APYckGyxPp1B+d2JJN5431ez8wDPdUAeR6FQ8TvoLZxKwg18lJTbPjbsPV3zkXfLYOucLQUmWejE
bGMpl4i5Ip7pk+zFGfGIcHXujJ+tSANGvbdG9cy2Kh79PaD/L+J9bU2cuM/ccHx1TrqWe5T2agba
JLwzxFQGjIvohTy+X2tk2ZnbavbY7sr6byqj0r7t7KkLK9jKu08aq7qFPb5BwLI69mI0MXUx4pZ5
i+qztshcfd74+EcSCEy3YRbqvVaw4ptIn2KyjoN0VJHWRDCkhZ5pNGZjf/frmrqE0L7MDj2x8LrV
3ZDU1fq8XM5ENnaf+axZwrvXj+OAcwDQLx4BdmHY6yi/i9sscyHr+2uK5iAmoOvLhaGbZDb5CeeW
iyNCR5WVeoOJXOG/ZDjMnc61kQkEv+F5q4otYmFV2XYkZTZnG0APR0l+ES07NDVJNWozgmOGB/S8
UDcBm0F4QFrf1lSSrJ0DIsuztOVuz1uhsfNLqpB+OcXp9ESqpHSC/bAr0JnTro+BYNIwyNMKE8sx
DMtJnaK7vRQErpcefKmoR3VR1wVc4LkEQ/s/cJqfsUz1BETPN/WP/Jd5wPnLhtFAYdmUel81VsfZ
Ewd+4PkU0KYHz3PP4NhiSA4Qj4cRNn343s4/SvGNpl3iOCNF828m31bkjoTprFBET53ZdHjB0rNg
hHUX8fSprN0ORMwc+zYYnk44O3CEa8O4areXMwfdYtangarMJk10oneA98aWIua1RgKDmiNHFCZ7
Bejme7hvYal/OD9+Bbot9R98V3UmJjsMILf2jF8BIwT4s/ArdUvCaR+obkc/+PxcPT8ALzgAmDKo
c2cSgs2XShYkxmc5Osz1wGUmwppd/6uottWEMoBCXdJUt0Dv9mGsBQSxXaoUur09bIgTwiRMMMOK
MmwOzC5t2Djvp973nTLnuKP7sr6FXgeR1soRYpprWLBtR1gnL3srctRzKNbKASwie7Nv2oXqWjry
MukOCAENJLFqOtJpaM/veAGTKiqekHGsll7O+mklZDDVzCBganSfEoCCPygtO+aPlAd+ND9CnmoN
IWRx3ryTsXARyExwP2DLitJvhXq73JIkNQIpEAHx1ZvOABhYsERm56AskIjsi5X+Jkd2+ffQUIcE
9WQlAz/bJcGHWEIiA92KHsfIU7E/7toSyXFjD+p1o0ZJnNg+tsF/Ws1hq4qNR3ugJ51NCicvDRul
y+1AIYujJW416oDSfzPqiVUlyPSjnFVr8wXERjTAMaP6RV5GHtU42UcsPPq8f5xcFMvNum3x8Mfy
8qBOUL62Ljj/RBYjc7nNlV9arZvR7u0GliHK1OUhMVcJrjemprpE4CHbjyp1tsr1rFzLfqOfPUPb
xEchFlTQfC0lwL6VR84IxDRE7R1ikI9ZlzMyjmzIAEnKCeqoAkkWDEHR3rdR2fJC2ra+rH1axtKs
0LkT4f3Saga4adZAr+0drZMdaTQwcajilE6oIAZ5bVxW7yT57QjdYVrrHp6iBEZOY/LCu8P1kxJY
U6n6MF3kuyZH16S9MQsz5N76Cwe1XKgs2BfPz8LV60XoFxCYK3XUKy+1vn8niG1XT8DTXS7+xY3f
RA+g5fi/dpEv9MLn1KHv90XThhpE1cDhpF7DDpkoRDgMDAPJfJzgjNFwawTPFBVDOzkNlOHrVmFD
tsL6neXRzhTVzD8g4tARWNzIdh+n+1EReVwFhEF3yA9Pp0Flf/sLwKKqjKfmJQe7dTtBmrJQ0d6H
w0tpGNn422/g0Wdu7/Tfvj//BWZSCjernm6cbqXjQFBCyjaL2lugHPknypwsMyerHou0UZvt3emQ
LMNRGNN2OJTxnuYK+wHadLK1HGfrZCUakbH5mG3UePZI7Sd4b9FDT00Higvt7oh3S8S9dFVgb1Mw
jIXxcAoKqa/mCxiywdJZ8dmULwz2V0mhiKFHJVGTncr3DPdmtJ5SZ08ojsZauIWLhk8U8t5Bne/n
M0CHn6a/G7OhIFClduX3i8GSZlCMD9aYgVowT2aWOhNYF1UrkhjDN30wn5gijbwr4cIXg3eIZxj3
daypHsh5+lKvsUnUJGgl9auKDWZA1DuIRIwgWTDWH9FrBAYGqghSumc32+87g/EYTh9Jd/jCYaAh
Fgta9M5+3WEUDo0VF4ivawbgWEXkscr1vevoK5vnccMLKQPXoB+hkZJVW2U5AxP0RiyMnc2/Vk3z
d/OsJXu2Q/dTQP5W+w9ddeXsTNGpXU/B1fgKTJLKM3IqYvUp9PI+iZjxwzaYag5mxNBaoktt7mRs
xPvonOslwtc9eVaftZO6wPWe4uuctpHYQoZyIU5B4N9vUuMiHvQHWSpeo4nE5gn5zXWI+Jk1SWYY
OWjgD6YMbUM1OL6UAcfHH6f0+Gg1wpOZYPS5vh56ak+kvRudwL027Nz28yVVm+CJx0386gqZ1lpx
hKleWKsrLVNws35WrMvkiwQSI7JEB9prWcPFD6hdJPHsrWzXTfWOmvj6B8dDC4smtYFiNxJUnfB0
Qea21nX7BPmbCHTAMY50Vb9NkvKWz7ze2k5i52lU3MD1r4Sol97oi1zioYa9/voH7hNMrtdtd4sC
yarNCVccBARv408Q5mMEDl5pHyZGsWMvAnYxdbMA/1oZD504ufcCPC2FnazZAJwAZIb+4fY4V6Ga
9ISTyjfDpOUS+YwulxEIV0tCjQPG2PJREaDdTlmF5mt8r7KQHd0d9K5+BiT5KgdgbSMR6k7HvOJU
cZNrcGX3ItYGKAsqY/AmQyUpltp5lHaS4x1wwxfCSkIQLTEMb96x/1jNbUUCj0LjO4t4O3+vEDrg
W/RBXipNqmS5CuumTNmxGdxJjs4vbujNc5sSXuwfMqIUiCtAbDQ9gIN8rM3B0rvkmJxZmxd6FC5F
QbklNu4JWuW+f7XxIBmxtl6NiRCPsZzLYPPtQh6dBg5vXWyNg9krCV4DWTuWpgFk31xjtXNGbANs
JYeq0VjNk+H+R5BuwrBeOx83f9M4qLYA6dZ61uUiP6O3+JFx2znUJInh5UtCvSP4FWa7/2TYH+XN
yHB1A93hh3w4pbtcatTS92w9PX3rVyuy4k43wV+yD0c8hkW9cb3A8mmRGYH754v/giwDw1RGC62z
q5oBu3vmUsq0xOg85bbI+V6XXfJ6km0liwkdwrRfLIybICi3tZNPCM9F7BiEiUR8J9IXb55yo8nv
9mXRDOBYhm8AzgevM6sgRSex1I8jq0Vx0QaGrSAzIjn/LUeLnPMNHcf9I+r+ZqQxuJXApLYt+VbM
/Qewk4UaOI5RkGaIqAoOvTW5cdmLZ/cR8OUF8wjJKgYfHM73NYnH6raokftKHG3Qch1T+H6apCjm
Gs4jO0z0pMQo7Kem1zf5REjeLiz2bQCv0RPZqi8Xc5qBlbhbUnXKelT3lPtQdmzqpLoDcQ0TMtY2
WjGLCwsNvaLQty84e+/sjJS7QECxGFhEwcQoJxFxJyNpjn32ORr/TqfAWMjluK2Ud966gxA8ui+8
f2E9j+F/C6or2BWeVBCWNgBFCuzAGKWFbFz6G3HR1TGckF8vr1NXNGWKqpakhE42ZrnOXC7e11e1
xUaWvClP6P5VoOTwpNv05w8Lfuxecgi3Yb+ylcTboD2YgXskaYu2JocQ6D5WJlGVBx8XlixniMev
7lSde5UcCht1CNrN0RM9ZXsGhut+G4ws+ukifki3+399KO5BOCQzytR5gBXt2PUSRyYwC2ufWQTk
nbD5AObwcNDJ7ALi7oNL4vZLGmann64X+CiZFn5v4yZ1VEbjqKGMDPD+r94DnWXhx3W0rvaFoIzZ
OWr0+RW7+nS0kR3VU7ZGtHGLS7CPjHVtuoMvAs3jHSqPUkQ2myFInPy/u4xWeiOJ2RX+ZOO9YVOu
TqireJ3jwJnv3qo7OJREJY2ITdpqgM7Ud1UVMNXXmmb50SFaHeRz3zsY6+wTXR6BgUXCqyegLj0i
0wJzhi5MmquULCIpxMgU/vPZoUOwDRIlKzFPuvuwGyg2lBTRmWLxyCcxVkdkmQ5YbPiy8N3Mmp1+
xqfJRnCwx0v+FhYNzyOtyN70eKhhTnxgOJPAmEjSHkNvPfBI9zdAPYFAWzkPDdxKWNlgRU1geTNQ
cwrZy4vn8cieHowDOXGDCJkSFix+EgrJUJIT1EOSAuaRb4JjXvH/2sMcpeAw4qAyKAXemGnRYBgz
+nQQQF3QFvo94vFi0z1x+gOR9BdHg6UEGT3TYXLs9sbFrEhTh7yB0gIJJT5ATrRtJE2v/PDau8f8
/F9s+zbqtnB1ioaMiHXgf8Wn7oJzHg6BpyVxSa/ONvuCQ+uCx2K8al3fM3DSgjLnWI1unILz+V9r
lFPUQ37eLy/p3YJD7AD4sIBpyeuN6BXOAF0Otrob8SvVaaDzSObHIKHe9iKobE3nDmObla1IoJoX
mcOXMQ+WRPt5+RL6AfUyS00T8SFFO9lBo84yw9yIZHc5wyKdkU1UNVBSoY3UH720AC16TLf3S/Ps
eY0/H5A3EcwuBnlqnV4G3gAdrjbTyJI9AjE5xtjebWTH1SBO9nnOcw0RluF5/llu9gNEksQivk/z
7dH5PYVotk3ubw1psx3Gfzk9W7HfGDm3K8K7/S2RR1ARM80+AQMImJ3kYJfh6mSD0T7koxzAcEPu
rTNWkxWhoyDaWiIb3/iFuAVrpVhzcrWNe7oqpWbDjy+TRVeE0kypHxPB9cIzbivT0SZ5hwoJ1RTa
48rYFGch/HajBoZsXU1XYZN1ZsRoiY6ppg9KswRnVCo3Vce3GTTtFrX2QZjlNPIwIIhqSjmz+KVA
YTQHEAcvjPJe5KBwDM5pLoSCjWsunENNJ7F8+iPLvdfDni0W/bErgtHYGS3OSfYO28zyYgX+4DK6
eOZO+GcaTPYHHjFv91rfczS3WYuHzuYLdulhg55C98c8WaOPUY96UbKGcqcY5BiLD25AhGBpkN0G
9wJNPX6uESWJHIAKEhcTmNJUdC/x30r08Ij/jMpIDVcXsbI9tC+A6CFSkRZCJhsUTlmQzA3ej0IW
usHZ0K5YEzmeJasF0BprHfYxza6RSJRJMHw02aoWzs1ulsfgwwZB71oWKV5yontukENtVvpnS16z
dbRgnjCXsmM2w/6GDJK5lI/dTf7pTu/nvqkeuGYFjoHr0lyZbyvvgRydE2exywNMBpmeJHdsZlMX
CxepTxf2AoIC8kn+/8DNwGzkkNwXNc8WXMjetq4f5LGUHL5gH1f4t+kjLBHzcwUGahVcq2kJf9Yy
5FYDLqhmXRkDsZvFXxIjz3+mAvmyKhFRX0GdhB/TzE02H6VqNLdHE39eduEiQzqD0stib/g+QnrO
Qtx/tu9tbMPySWEGkRYzJAxTir2nXGxjCtyUb2n2jFvZ9fAfH9T0Nuk7Z1OVdYErC6oRn4UmdGwc
EyuYzabwLbt0VDFIdjWXyjurYt9iPPkJL57MItpEtTQEtoiDlDF5eOAMiXXDr6DHF4kCsdlFgG7+
ksOJm/PaEdp0LFQuSHoXYxYQIo3nlV/ITx4E8DpCiaZzbI7yG7GSYayS4d/8zQ1MKnah1yj92im/
oOiM9L/SmDFT3DYYglRj/Y1Grfx/ob9emJAaSiJEtUXY5F6W7xDxatVjurhP7ZRA8g8Y6gtuSj1K
nq+RpjjP+O26ZD8yYr+FoY9pdZIj320ezZ36fMeW0XVb/eYaQG9Mpp2GKqD0unkQEUsLvJtXbJi/
pQnNqUjkD9nqzlTu64+0MwCG7vaWnxaEpZrY2ZlY/FPdIHUEpr9xN2Pe3opPO869lQqUc7Q3pp3O
7SS0JGRgR9Xih9jZ89v0N4+jJ+ygwAWag84SWkFjgEzGOEcQEKJVR5ZGcCgZ4isH2BvZFsYhWUdR
pcmPoEThkqIgv/Et+3bcymKc070snhE59GpP13pdy0J2h4GmOfwiSwbH/lM2M7oLnnjaqignMHsT
/D89Mya1FMw+ceGcNxHOQLlJwte/IEZ6Iq6m324yl3rG1uFabc2oVpaSQylU1Dvd8PdoFVJmaILz
ZfhejrdiFCtA+m72TTGpHPLlFGsHJ5s+hCmEKLu+7fUOdZbh/7CkM8ZC3JxJJviMxy4bBl6ljm/A
UWunptL9B8P76wO41u1dwa5cWTTMB90QRloNL+Ghxot8x8XNFWbPlm0l5Kn1QDxPOTsSVmZc49nw
DVdceDUL/cqrWfOebzPIT8sZSErpDJOJBc3jBCouotPbo8Zir/frBv565zWVlmLpEDHWer/5pSeB
TyCQToUQbwODg2XSN7eYKw5C7p3/Hp4TbgsaE7KHMdfN+xEf/j41AvCARcTTdYto9s6Qj7v54ALu
BKwJE3xYL1xSZAyK3pYIJXw0qTsPfTayEFnf5Q5AyKF8hnLl6+iuKQPcQe42JT4IeNtBRKAlnW7A
DUEVU0ZgzFdoQgT6+ucjSYJnywMKsO/nE0yNj6d/J2uBNHfqWOj9x+ZmO5jfh8em8oeCzkyZM6g+
Ka+TGF6e+6bx9H8HtzqiNr32rl0p6MWW70VmgJFOYovp7FjIJieTlXBKczvSFPOweZURiDAD47g+
nwEvVgoGuOcP69r5TMlXWyEj2xEajaQd8Lh3d+zRT57vnzwTIoU+hujxLm2RzXccI4Rt+E0mG+dE
cFc2xFwgxWPfUO0sa380lifhS4BHFTGgfjuxrjAXD3xniFdWk1bToPIr4aGNM6X9BJP6aWFjY/ha
voTx8Rwmtd+uz93R8Bgt8YX3jRo+GrnuWtPB3lSnbFlTPcdSu2oiBqO9pw9tuwmPVTCA/k3PUMY1
y36pOIgEMklyW6nOn65RGXrtcCu+PGtDhwxZI/Cu/Mu3fXkd5aZOid9bzlZ17E/6MkNB1Mhbt/Z5
crd19K6LHYgTgAqBcQVqK2MPDRKSuMimBZ1YOw+6SU7D/d6lr57cHH+X0qbhvHnSJqW7+4Ho7nP0
Mz+IfLs3paNaBhfuZGEB/swi8roR0zQuN5uaq4kJKHs9JwtD33H+XM2RJp+Gmn/PZcP7v/cxEmka
FPq8PfoCXrL+fLlHuINGcAm+Z9ZVWBoC8Bul/m5E2M9M9nTUTvIhN2n4HDrHhBy0tjQFV2EJPwkJ
5jTLPk9aZc94TJdCXNRDAafSwW3fM+WjuNwPOrXBd1e1VmnNtayfz/5CygxfD2XAI43tLjnEe3PW
qD0qmWo8AG/eqcF3UYHxMw9Lj0Khnz3tGUTrVWMmhqUgvmS0nYl+il8sv2OgA2i7qPwKHAZD7qIB
FtJAxyXRKHxt2+il03j10Mq98/YlAHwNhxls1LdvZOq6x+ZaRQMDiVpFaW80e5q6WYBbLuWXxrqI
2BH3B6ehDdgaVAyOsz0FVMgeVE4J2kNyGsNu0OL8CRJJsbu7O+OOXQurpyljKVJt/6NGE5s6UVbX
EUfFbgdcmXn8/2XJarPj4s4/BK+WZFbwmvCS8wJDw0Q2dwQTbuPExhTW/lFHphgDDuaZdT4szJ1B
B0sLRa84uW1k/u1A+01mbLjTXNIvdpLSilI1RkTASoVJ+GZwfPyXRkhKnKe7lAe/un2mz2zvp5v9
6L+8uFc/ISAc2OvvuZqsv39NB1vbQ35vrAPrBKK+QHQGglLqsS1QhxAM2mgx4XSe9NZE2THSQSEA
7KTZui40FukfE++bm6ElK1WKwfKT5XqPTsMwrnqxOAvH9bXkKk5notGtTDnubwfSyQl+3bjstuw3
Ik1E4zoHVXVGumkayFRxjRLtcAtRPLA/hb1PnPuKQeWdWITcyKJfVGgU4SYzeWScx0d+0OPWB7EN
FmPcyFCbmg5gSxArfj2yhbCVqBqN3w8vRhgxJ0MFR9wlBvW5LwFHi8WV/4D22XAQlu5hZPZKMC7m
ihDPnjDB2TCQeIafznYs6u5jRXRi+q0E784DndWc3BVMB5C9yzAeAmuABwO4W0PFKJZ4Iwvkp0wC
2DPoicrQujJQwhLBVP00oqkccEgBtyFDJ/FXcCCirM8yVBtJzghNcFtVB73nR2ZddqMWkDD1ztCg
bT4aPQxHFo9QadlojkR/YKS/bHtsuRekmqQ76EdnGg+44hZFkTGL1kFAkHk40ccIsgwPKBQdldqf
VRxEW8MKS+e/sjnOQPcbk0nohDb42Du5JVHN/8sypMZldCBJuZ/7eaMuPRJ7vtvSeGykAvqFOcmf
cRiSQ5t9vP5vp6xsVrLiAwY6AkP4PzjJNk7vAmYFUO7nL7fcbdqCnxIzCIPgWo9N3NfDKTcWwvzv
FDIC4kk5cJrotlw/ABBrcGCu3cKhAI00vTavcHCNVYKgXUry1XKCG5dhMbxthglTTLyZ4OQjFeaD
EBs7SgKZWJV7tkrk+fwwHRTpg8Z1yhQ4KwVwnn9HqIT+D4Ycm00tJ9FKpAqgX+QVo8STNDCBm+cj
AofgH75fSSn809w+AIgYH7w5frX9hsyblP/CwFJwJnF1vm3it7ccehP/evMEZuEHBHzd0+OEBqou
l7oCCSTBDrhgw6GoyIJDQdVzgfViRcdoLt8Nqn/8Mt/ke0Fujfyn1Ce/kq1x/rgEHqLsqI2IgPNg
vDmkFdwyuKoli0zsOdXU8LIvApAgL4A4VyTTr3C25UYoiQ3uNBNfMJuy0vTslUSdFvWcugE9aC3W
y3U5TrHOKX16cng9rQQxSOE4Fb6Vn02jnMjYH1kFWRqgRMi8sQ/S9z+IzHnscyZKBV/AOzk3b8MS
AaPZrK9POlMxX+blGuT4bNjLY9EhXdpewzJkPaUiiug+DMOjRewq85rXNwJ8llzrqUVCO9fp3riT
P5jGOUDrlZWjM4E/9Q81P0KH15lh/O2Gigy0W+RfV9L5+rg81YmiDiEomzMUufnqEHzOHhtGlppI
7ZvXLHDqIsEaQa1KVA6ZNqaSm0l2v6GJDeZWxlnXwsV9tInESLRd0jy0N5mXdxD0bMgV8CYR3mka
sKqmITaWioaamVcBbdw4qgygkgtHC/tHgVI82ZRg+RloiSj+Az9NULfkyocygI0YLbNk/lRuYPsO
KLHMi/IR1+5c2saGAafO8AS105zO/nKLJoJ4A5MHnIqXnGM4oo+Ti0/yv/vzt5HMr4HaMcnaRFRZ
j1X15WwPoNDgfjFNrtceBYPlm7QwOzmk4QkIEkzKOSIyIvim1SdWIhtMJtaE2pqbfviyCS1m2YDG
E+SCFG8Ua3j+t5CjLiTa9p0/5Cjjc6mQC2iagu1udNwNY6RAPhEBHqm56ksCfZe45vHADbpub1JH
fCDoR314g5HI29WzisW8O99jmyCeiVZGbqibg9TW47Kd0XM6Pyz+vauOUJ9QF1Jm1CtnV+HOdSxA
A7rVRrNo2m/RZHeJxOMk4GJgEwAMRnLRmoc0xrHAxBVGx2jj06cVM2oyAihpM1QwXTp5+UYHNrS1
QUrLNroAoqSROspD+LGF2Z3zR+t6NqwRmRHSecUu0Daax3L4Y/evrI9BWd65TXxFjd3DFi+U4r4S
7LPjQPmeGUKzQAcx4DmASwR8dyGJ440sdjyWdvTSmeWcG4aEmtRx6p2vlw4j39z1XU4hjJvoEpZI
3DQd0GW2nNk/YtO9exEUW8NaIf8toCSDe1LUBQpspRU0NVnOD/YKshhIvKs7McE5Fks0z5FvOb3l
gLHXoeEL4dacK4zvuu1zZpb8NMqUQOucqtaSgZXuLyYW4h7YIvy4FanE7YrLqID65GjJNhH5sJhq
fWwUd9gnODWe9ur7S/84+/0X1zp0xWd4NUsdSLkzr1giU4VW5/Mg62t1rZ/BfxVjiPg3FNbB0oIX
6N29Zn0ngYAH+ag16vmQZKKZJooe2sroWaHTnsF8Oet8AvyqdLQiladkHQYq/IMSNULTmg26/nJr
6Il4QxXXwH/Hf91sro2Uecae9CPTmocYvnn9cLqQeQnN5/hgblCKZrFxVK/Yof4foSnd/2c6Bl0A
dmV1KGyI8NmTejrtD1tdobUUGanNXHNdG/jBonzmrUYspd74t8q3G6vS2MFkjFRBP3L6AKHsHyA4
RMhFdN7UqHYhRgC9XAoDp0YKiCCOv+6n9keYLh8Lfp1nnUgCiFFny+LD3dq71Z5CqcsFEddV6lwI
SFLVlwT03vUMfrNrkrBvRrsiwyKGJ6DH7QNEX5E7rJfP2gCtl1gEyFONfyOHBkesY2ckggAghUj8
VVT5jyKcc1jotuKn3etK2NNqtCSWMMAra6jNSZpjra4ADP6K0mezrHP/xNXQOBeRUIPciBMsipCt
IaOKRFDUcCEzaVSnpSAtppBJsQuFSWPox4ao3ep/xLOryW/P65FR+zRqyryyHjROm4nkPVCTwHse
z40DK3VQmqWKIC2RY9g3MyCD5QtCZtJt7Do6Giux1iqZpItRgNnOSc/LdSE2CicYGsofuSNZVr1v
XRQB226nWeg4sYQ/FIAWf3zIl6+aj95JdpyFwqUNmm9JOUp8NJZU6ADv7uhCOY68yujFsbtSJlUp
9RFUq238y7qPtDGYoVp6VR+SpoickaD8pxhup+aVMytMDXaTiJJst9Bd3MUm/Pg9aqSZNZfesopa
wBxIw/HVjqVwOTX/u6L3Su/KqttTB3DaUUZivO0NOzP2ARcdS/F4ayZeSPuvm0rgw9E3g7RZfOrS
Zz5lzKJ9P4ELBTE/Tw1e7KtI+FDtsufbm5CkwW/53Wahms/6Eo1Xz31P5vgbbKekCgSEo6aPMhp/
DbWAk/vnE3ua0/atJItrtgY6d9m0bS03M2HydiJ4TKnRMhHcym0T6vzd/l72Pqthnm8JzjJpoEOE
Iy4VdoYzue3zg3hMwAGmESVCMRqdsntmv/qg3q62BWoei3Yjn36ExTFr4pETeSmU6QXYqgScSoK8
h/6f1+G5XarDlBLG9KnfWBsJUeXBPNJNxb6MfX4zMO7hoMZpZrojn7d4BpsQx8gR6rdCdqqVvy9t
HjBUE+d5l4TXKHycJdd9+51OY0mw0vi13uIe+394kSLI+EoRHHnluDHyfPkbrYo2/nFwLaImlI6Z
V5nTmvIavUGvp9enbx0LXN3q6higW3zSQDoO1kBN6yJOFqxergtgo4lKxapdZrzeFEIcLRK2Q6xG
A6CoPeeL/fGEEPlQlZVl0ayrc58dn3h7WWCRl11hgi+qW4aUcRDq4cI2sc2oYB84ipJyRcPK5tTa
3HEfG34UsUZhD6+MhKZkg2FBtg5TJ05tiQauGMMAYOQhD/n41zJZrsr2bGCDe0a8VRSn/7EbsvHm
5ZB9REj8jeSKYrS7e1D0ao5yhjRjruu+alDVyGqC06yXn+ah0zLBs+Zh/AZ9+XguHhPGb8kQhpLK
kpNmWFSjh0mVEKfdM2dWo39vxim3dABfj+BCUtKsW3vb/mp84hx46eFvYiVe8x17U/vSnUxKuLLe
/jJeptQxi52wxJyZKgnFKEKtAOA8umttLNEOYDmY+IG1IeiMDKdxjqehR7C6+gk+husV1ynHljqv
a6S66Z8yRHIR+uCjrabZxX9b1d8kpO0XEsnzKpRTWS9hWwPsg7RuuyTPsihgkHpAnVPenVYoV6F0
fN4OeIVH/3v2ooHRGJ2M15BqHi7t2J3Ryjriz5df1f67NDl57bP4q4W3xqYIzL3e8xzt8RPRjGhM
T8BNJ2pv7ZBDdejU2HtrltefeS+ieHgdcEQ/Xt3G5PoKroUKvMf4eD7zqs1MI26aM2UFcMkYgdPJ
vF2Dzv5ag7F9vMn6Un6JXLJhhJZlUmjZ5XiOicNsV+7uB0g8zxTwvUz7uq8K1dgRpW3B+9BAJV1T
gFSjpb6H6T1OOJ/HATEifA+1z34tVOHF6J+T+tqRh0SJnFB0Bv7+r43s6IjBrJ9r5zKyPrSGRGwW
I4uygwqa0fHqbCrsZUwS65Mhx3wjOxmSNifnLwFGWOfaTXmkG0Fh44Ylc3QU7kSG4TZ79QOXsC2/
rK88jb1ZVKqXNfgF2KysWMDjzKYQ6tigxn6TWoguUAKfK59hrThpDOZmmHSsJfOH11QTbhc4YsbZ
6Bi70z3dnHsIRgMfGW7Jtakmzkc8PhWC5FUSSMD2iJ78go49ExUk5A77ogXCNeO5yTmeLm4KVZ/3
Ja6kbtWGTf8Pxp7J44UkwGkiQl9DoH5wAGGNroj9I2ov/OuQLjTC6aAn1yfhxt/dO/IyH3wcThbW
A+lkURgRbvjS/Nweq+0uglY0E5PxzrLM7iu5sJbAW8BDjz8IUbPM/etScWntAL6ACc5YlZGwTygM
TZDgsVN1gIdD/tvwMFz/MO0JCfAz+GEEVscsJPnhZCQTrUmuaknOMJz6sGW52WJQdC8CtdYaq+JD
qozz/qTwa9ywW8IZHe76tLes8iU2mi5CSiHsuWeqqxQ3N5tvv/tVIHOJLLmNvTtuYzqD2fRj/4H1
HxgotBVpVwLpNgWX6ZsMhujygMjZnbIMGF4hZY+Pq7cpKRaXS1EGDVoXQ2o2Nq8+buuvKymPTqnb
qhHkm1cWBukTWWipsJPcj9Zmgv3arWSct7vQpiBeH5Uy19WoILd4tKaOH1gQ7dlneMq3xEyyO/6E
gJ7a7bS4PuwbPkWoT+Ml5s5AtCrmvId83OIw9Z2btkcViJcZpWxQVWSoOokcZpNMKbsagwOWHO/P
b+XUDkaWnLTp1BPvdcFSccrYtMzc6VpRaVeX8JqpKjWNFEpApAH4TvdnWvbkFlf0iSLr7xUnsr/Q
0ebSaZ5VjODmL/DYPJd5rz9psyq3mqaAnBo8v+u+o3HauwqmhQPWUOLFwkMGLCy+LBZJg0FpDjFt
W/dWG9M3GSit+kaedYVniune5ULMCZkdYDWOHG7WKwMV2DEHyYyl8AJY58UeRSmgkV4PhswY1Bwk
qKjlcFa4uz5EsP9JqIJ9ACnNbKBRuYRa4GHHzA2MxpKkaB+MFCg43bvM9MQc9U403dJEtEY6X/L0
HKCMz9lStYNTxVzO6TejyePl3ENZvkwh2dXbqzBGbLajsACs0Jz5uLWJ+s0kmjxNvxljuIzKWRMl
fSllvhELORDT4YoKgdv1SLY5ZgrBUdko8L2bWan8A4MvpGKu6AgUkBk3fxxLsTvU91XVZtOhgge5
piBXdkb+TDgkCm1rDcyoiIwQfcTGCUGVaxdrbZ2kERmk2DhtMezhlRRMFtbf0AtXofUW3gdhMNsc
aox5miU+PLpdb1jLKu87cPSU7Iq4XPhN6kZvWZhVpbWDwTidUBqxMy5VCRJva6HK9fR+6SEtbNd5
wjObH0T/pb2WK/YDJYN096L54XqIuxekQ2ZDCOgNaBhhnAiMRDMFcJ70roKLKvojWU51bVL9yjb/
tTwq71NjG5iwz02Pq3cs+vesCCtLxrdfmQLuB9Psjr+AyeewC7r1MwHbjGqSY+TY1KW2YvK4rF8L
d+r7ZJTwhtI5WrfC+Nf325pzwVugRbGBArITVfVekANly8ZObeXH1ZPhrzNBZJZesD1cc1Fln7mT
9W1nW7wlHISdbuT5Wnx4Uxvadu6AhrPTtCHckyfKohyGwz3T5fIamdDTWTeGPMRFtBIpvF+kFCP6
0LsYwnGVNNFvPIV8fVglGjvIxNzlO8OZ7wHP2AtoiSePS26EbH2KCJzgnKLATsfrAYgVbu90p5g5
kcUBeur6TDFuyKERpY5KQV2ZV+qCAolWPJeczTTRAeOPLO/28b/x+vMlTmcybCf3C00k+NDYezmr
O/dmwoVX9q2bpw3/Mqg2Batmh9s5ADyZ+ObG2l8hfZFJC1NeUHLx2w7UnHW23FAJARkc2rUYMp9d
2lBJ9HofjwK3DzziMpzqSCaR32eqIdKfhAYFpVJNGAK34OIxRhRgc/HhVeFeyH0RzUy91rqwbiJZ
WsB3pbbtIapkKqRq9ukKzO+fXoVOueAJpi9z90HCwhWFb8cBnnc0mgLlNHoCLKdkVcVZ1oSpQs/3
MLzEQYaI7qwS4aT02FNtAqDGRferWq3Kz1944+8NxFSgYfMtsLyikb73o5pIZCyvP4JpbbIAAflP
+tKtTi/PTmGZH3Us8vb1WZHV3U+TKBgWgvlkX0gnN04E7FMJJAzqZ1zi0B0bi+ESUuJImdVqFh2h
RfHny8rXZqM/6fkUDnCIUul+F8TgWAhHW1wlPds27WD3chPvDgt31RP3WQDB3ZJhwqhmahx8mU2E
akri+Ck1HFSW2KOYFDzzdi1//0pPEWBSE1c46sfrEiMeP6OhbVDX/o7Wal5SS1EIfJC2ogfUpo56
IGwuVJ3xvhwvzXgQDoZubNz+DsdJdbNHIqbG8nCeLtdBSyO+RNqkQN+M5i1jR14EgEABm5sJsLG3
n6t3Q8MpXIzpLlS+obB5+nNS9N+7B/XBjLPEEWYWVruntWn7wt6u+MCQeg/Fv9rbSk32QSwKjIRI
5WwP07X1JsgcxPz2PuraaaScmaBVtXUfk6qfWdfzj6GoxAXqZ49FYo7ACFywQz7yeiWPfF0BmrNc
sCogFYBHk+AT8D01bR0xqfXYzNx9wl3Ht7mMBe3SmLf1bMuVzZxg+NV9ukyqXA4IbK7Xa8n32pJf
+c49CGn4qkU5aPn1R9zFDohpqnGl13Ckab+JG+EjWcqMmQBclqrKnR2lfphYExllVKBsvt2GfCrx
vSxrVoK44m2hR8xKgs1z87L3Ni2tS/U/V+arjE8a+v4ZO24sELv0JD5npX9SweTugJa7dop/ugfn
icB4g+5Rzh3RA6vQy3WMsSmJfJCatOA7fCJIMgrHgrVcrim5w2CtkbybKa0DvJAhwhjkp/o1d9Xn
GAmT8bRDpciLgpo/06BOTdTS4skuTTmTLrPRmWrNqM06sk4EmM65dpMCCYIbGFMgegsm0916eOwd
LmETe75OzcXr4JfJ98EnL4mxvZSZliVlgfFVulQlfcZX01NAVq1R2sA6Uha9cogOiKJ1023v812A
fxuSv1A06b+JPZlDj3uYMVwipOKEjGmvWh64Riz2Pb7sm1qX8UNgOooxVIV5sr245YD5NrmQpX0s
iZWZQpCOviH8hzKS3BV1MHlM0Hg7wozEGYFpbhbM1Ksf6enRFOYKXJy9tBLhIpOiqEFrZ2t3Y1Kd
NmZPrSYEJ72UuQp3ZxMUQqYACNHcbEkUlkK51E+1jtdih59Iq9T4nrSRs74tNVP0iRrLSCnQtL3Q
pqM/vJJrlpQRStD0hLn4MhkmBp4zi1PzSU6dwlfHJlJtA/naPNH+JHf/I94wTC5U+dNaTzQNOxde
3DIbKC8Zsr2RZT7qRPt5zTSzFPncB7ZBgR1dTpG4wkVSp8psSaqDS91xFykRrrhk+ZYG8oyzN4tz
7YHaImtAPjiCjcRltF7Ru4CwlurEkxZ9///phYEBdxJZl8z+mHuxVfM8bprxz8o0N5UhP8WEUdYf
HI3tWALkMzHYVQAlZ0WRvuMsGfIXTrC6sXLK0jVwMsoXrkUStv25N+NpLxGzqLf/ME2tzxdfBhWc
6vNTbfjJYDaPpGYObY97Ir1ChcfpJND/wHdSzA8HDR5TZDAS31lBrb7M1/aTlLQmvbV/L+WzIZig
AixtMY9nexSOvh+xju5ChuNFpFO2gDK5QV0U7tHP49QPZDRkoO3dEsNcFHwrHCBfAuCtBQdFdxnh
qVibAeSnCsKndyVrKo9vGgGBAnc2WwjTWWz3Wji3DVClC8PvJlNLO1/IgU3jGWboXByFVlml0wmE
L+Oq3W5YWqGK/KMkkvfpzr3NaeR3XdHSa87CMcv6DHT0xK02dGEE9daDM51+CiodoFx4gLn4hZLf
O2oq5RMaPMDtwUHtfsILWDXuBg0saF+Lf6M3KHoRoHHDyVqrgOsv0+hPlVi2yi0NS7pX7kjp9vEc
jrWSZrGNFez95tg+MXEIk2DRbgE+FTYEgO9AnM60KpZ5oi54wtc4+ZhoIhVglAIz1EVRsyPO+0hs
T/19L6eNlwbCevP6ylZ7jYRKQf6bGpJgvrQMOGdvopmOkH39CpSUvE1ao7IVPPot7dW7O/Dzya0K
PdqWLstCRIayz969JAMSDsbE3jsDVBrtvV85G8daQRbKMo7+wWohRZK6izuDAC9F14LWSQGZZ9F8
TsAU9nCZIHvaqwzxRFOR3fZRnSmYGL/dlB4I2KKj8OZAdHcuf/CG8iMaxmcQefLt2+gazBk3+yCx
g3C5bZ87p0APItLSq0i1WMFUBfNORUdgBf/sV/kJDBvsRwvkUZxiY2FFeS2XiQ30nuw6T2GkYrUh
vSXxDv5NG7Th9IatIPHfNg/EmpUXni8cTxn4WrUcZezG5jwLi7rBjMT17MQ2zFabT9x77B7AGGcY
dF1A1/lEr2sA+t1BQyX6HK3T+i9ylxdCQ3cfP99EqUPtsCE0zlK8GXHX1EaEoH5XF1XKd1nWjdwH
0hHcpMKXLVYsYBXmI0dBoESEwoQLoP5TCtoi7433gClUaAYQLEtSPHzPb46dcSMCzBhiB/Hjc+Gc
QUIUZ3XFdWtIJFsRS3v+3fE4uaSRdVa1tx4ejDZE6BEMQKUhV4qBrqmNTRa7UxfR9+ZgSCUJeODW
neYrSM4hyIj0ZqnlgpEkjROmIg8B/YSj41mGgm0ydcZ0yQynZvrEjslYEaaf0M53cxZjEONGXaui
fSHhB7kSqS9YV6VoyU75kITzhYVkIXQu2v/v5bHP94K9xuBVFT/J0SR5t7LP9g7e2E3naiHNxCbx
VU50kxWrN7b3zr6wFSPFucWIlg/pkfa14MUqm+SQkRkb4vMGeH/lKu+9erjJLmteJHarkHiN72wV
XxZc7LNNk2MxRTlxI8tXJH43oNLogWK5+L9XL4MMVYp+gdTOCNXnX2XLLUIefIcGBJJ6thJLitnR
4TxjTnTFQ3Vhte+WDC60pmD1Adf6Wdcv9fKoDq+8V29mO8pGw4Qg2fK1YkS7PIthfYXsRTwWaNj8
hqLJFRNWL1Jx1chWHy9kQpo27+Ol8L5p71e/dmw9FfOImsj8bxRJeuZdO25+O4SUJoNInPJs2D/t
O5styUzXmKPPEkxZjMO4cjV6JhfOfiG4/ED4VQqvJXZOzPY19rxE6Zl1KzJfhjwt9HPExrSct+9+
wrUJJz705Nc6ZNFyavZq6r5FQ26F1m31PTu2Twv+TChNeRNfd5g3hoRJGTgUdT5TwF1pjcrcP7eK
qyIfZq870E2ner2CyedyE4z7ZPZD3wEdji+Q4igOCXIJmIVW773d8LwR9WTvSTaMvWborYBXCHjJ
QF5DMa7rHPADzLvpg1iXnX053utDs68O/DcEODKN9i0WQ7iG0OrG0Fm7WPNRyaY+hh0akyzdnb2p
E2c4hgooBMJJ38OkeYCMogL4M6DRg0UYgYvFpShSkUj4m2Ss6pkm3bVDfEV6AMcIdo74a4LVakhD
qSWWuA1kS5+kb1HZtQRrmELjz7qrXd+wywtd+Fe0uVOXri+tDI0zMWaY4EAdndqp6M67qc3lujJj
m2/PZ4AJ5j1JlnFjVwn3Mpw/R2c06sbvQAGeJ58A67TLfFNdRZKS/BRa1KoEjUQdUo8XBEWtr6eL
/6Rk+GgtGN40PM2Soq0NRXCyzIJIzPS1ulrQD3/mpkxxMsrYJdfr66yuqCZDB5cyzyGroclYfLRS
dv8Ioy5SsfQDRMS4Ri3lxIz2jmrNzg9u0nq5JQIX/IbW1+rMnhSedfno0qNxoiw3jZlnEJYMREdp
CgTvtpGxZLhTzWMTgh2UR2U949tkAVJZ8NBl/AFUqYD/u5Yd/wTR1b5XOv8LyBrYru8FOP4pTTRI
/d0gqKn42+fB9EJh8vdImeX9o44ufmg4jtfp47AMJXGwX7SvCr6kAgyjmJV4NY5Oc82cy7v/QQAx
7tnJ3grX5rFw/3FBnmEJFFhPHhcHOuim9VZ3nj2m2SuZafwyp3J97Qf7osKP88VSqoc+vvBxVDcM
APICid84xZddR7RT3/ffOspHWXV2u7VpT5p6driT05KJ36kNIWf6Nprh40vxD5r5YB1todb/Fg1k
/KiGv+NLeW7yq8/WqbIHEGBkhK5UgmGbtb09jv/tIuZRBrIP36BjignZosKmfYSTaNAA0HE23Tq1
Vy6gxTj1AFwmkDm2rihDlZRbNxUfZ6imBSNNoH1YVCe1wmN2SG7i1jzlefA4r3O6/lrz4xtXQt0w
MFxOAOq4exsYLuXusLoarch9n7W77K7vM/il0Q+EyAbQGXHaG8vuNeQPJ8hsg9NY96AM9fLC43Kp
h2wRQ9HeCsxrPhgVAw0yRY+OUGxHuItN3HjITRamu+HB9oVjO3aoUzLNB6vmeBkXEXH0Db4KmNZo
TGTYrGNH0t6EzXoh1q6AAdwZhuJ1vTmRMiBQ+Dxa4/tQY/Vt/kQNUXhEUwbz41wHa6ipREowiUUU
RPWtubaTqIkAuWwvwGSdOBch6SNULYwMdOe4ai1k20pOzWi7hRas7SwJELvsN2LxKN3XnPh9WuJ1
iuaw4jlny7zVQVLHSLtReSrV0uAgDWWtZoNkr/XEWj0wHZq30UL7v6w0k6ykgxPQKVYspEAX/2Fm
6dglfmXiTAOGuy8jQH2++st8vHanAK9pICvkstmaRtwdSUjSoa6fhe5G+4eYQ4OMHbq14v99J/Rw
bP4YeLdLEuX//yaztnD3qBctRsUrp968/IVj69hXYd5cpf5ku3ewVM3kxVslwjOyQoaVx3g39D7U
CigT5l2MhsFFY44qGtMyzqMxIoRu8P0YAJq2hBZBCJU1GuHTBJ81dPD0rmRtetqrOA6qGHfVn2+X
tp/t7gSyclXm/Nz/B7MB8iN283CrIBXUHnTdCUfSeYqn8az9ybdWm8Nzp75qKAmVdtCEh84dZE9o
DvKyipXqmlLHmhFFV+TMDzeUb1nDbivYSqUiZ46Wyb1Qnq5Xo7wuzl8g8l0qsAZi3lU62xNwSQZK
aksUcA5WPPw0tLeApAvbeBZw1sZogL23EEDeI5945ja84bCYBOvBZnt4btB4P0TFx3EPITLn6AAv
6qDjGSlpqieoSZE3jNDfNtGsV59jJQROcUteRgNXbwDUa4jsB/mP/lHZWs11HW0SM8UGd8dQfrHr
VlUvHcy5CdhZJJjfC16B1W92UVCTUFZHVd4L78GU3AhNu/qDp2tpOHpqVQbAB/4rTNKjC2NhOO5P
fd4KtihZAzP/4QRXY+zRa7LDphq71EYGYJeb3HPwhDKj2mD9d9jiYG+U0xp3s4rOEDKgrBxOOh3H
3m8HD1WQRj5AH5vILfmJ8vcfzj7W9ZzDwgQ9LUj+yCLQTGZlKKhjVooj8eJMBwU5tpRH+Cvr6R0/
7DK7ili/E/k06p0En84yew3HLAhd7Bjga6FsOwcjQZWANmI1GrXZbZ1T0Ga2zCCDA24bz2B4rGX5
9ZRWRXCGil/gYygpKyckaiFag3Crv1DwMXQYdkTbfvOfzAjwYLWjefqiMmDcNobrJQzVPTKmTC9k
I/FBgvYvxJgLcAMakvIPpDvBwVEbh8XZD0JkRLxhC828ouJm5+xUgKHz5WvUktEensoL47mkcXaj
u/NwPISPuBn+vBk+/e0qKMtTcCC6O/D3tgqqE0ZslSFLFY9UgqLiylJJJaIsG5RlrZHlYHxJpx7b
FI9MHTka/8KZ9gwYdcr3Sxc2u8QHzNxJu6t8HSwSqtHxnVDfxCOYignuCp+PWzTt8N4YYuHl9NV5
KdOcwTbaGHSYG6pCWDThwceel3INg31lpkYZdsdGx9YhFLbtDFyt6hu/1tJ0dz0mjMYcaITnRps9
GFY7EKZsVGLDp3u/HkGGd6oV2I8qpdgKgcmFY5v3fe/hAyS3Gepv+0ByDDy/h2sGDDq+dZ3hKlUy
Rku9cFgB11m1N+VPefYvmTOe4Dhkfb859JHaIAI3X3gZH375hTUcDCGNyriJpu3pOZTCETH2N/W9
cIGrp+hr8HhW+RDuPP4qgSg3H6LDHFQM5uhnel/abSTIfakN04owT+cTIy8mMTOqycUvY/GH7JfO
KCq6OS/I0R96FP4CXdT8XpxQRPp/pQ0yjA4aDWO26mXyM3iOHWRYW57+KnqIh4MzOTmWWf5bseRt
7BFG+6iP7+qsG3U16snTw8c9t8YQUXlommZLqOk0H9JdHEAKFAyyHyINb/M9INR5tgmeqgNEdV6K
8uW5VTpXUbfCM7dEahJGnw3KRlB8zAqqYPDpfC0kwrN4gImf/aTwpqF61tXpvd2AOOvfk/EkTDbT
q1l3GK0Wa3S6JStNCg+vBJhxtoeFUl3hhEI783KOfusK/Noh885Zxoyw5VfyaNKlG8geHejp+0TZ
H8IWspIEc8FPNIN4AU9BZ8F/V11/TBAP3jUC25q1L+a4p2cO/hJBGMkxjQBBQevEH1oUGfhgstwb
0uDadYfGpuSE29ymAVWpxqOsiJxeKCd811keg10u7kpnvnqJeBvoNcSVf6cspiHhsub6Bqh5gMTm
dTn9RVND4UvN9E3TZFZLWI1r9qxDweCA5X1D9vQ/vDoiK77w3HxB85/JEiXGf2GKkxZV3jhZrfY5
D/kxyI3SRtkmafq16oTPYFOwcskcvFSOqrkusO3A1+6F/p2QuAQw26xIc+CHS+jGPU6YrwzoAIxj
CpA+6MKuPFpxCHgYISxLpgSzqyy4P4AFUnmiFjk/u+K8nMAdl3EnGBBY9QI7QJ2D8bfLjjx6X9W3
FXHUVXuXkmckLP9mOs8QC2GMOr2++kVKSNv0NbT8JT6nkzIfBwPSA0ECLm4wdUV11BzswJIFbyDX
R5MAgB19m8kMu4q7llSVJYpf7iiIDO+l50Bpq58M5KQhsIfLt4X8e+x7yivg/gpy0HxzMuVufNgM
oZFSBueXttb/U9ROU3HJACVZnxM9hXQI8CWKL55LyBWVVfSCVPbR+dfhuHas89kJgJp1Il5itLwe
zo/l2ybB4dmyC/7dLndehxmRqidIxeuDXW+kOeToGktEjRHkJH6lDko5cCebQU0D+WK5jeNJjwe9
EYzKS1LaDvb85W+ZRdioTWP0LU4qcvBMgNVHKTCprjfXtJVNPLMt9yiDZ26w1LPiqpA/pKqg2cEc
BdrNfGE8OBak1omcF7NhvWcn6a1Xt1Wu0YyqO+Jhf/cnEwb1tVMVuA0WIqcpEC1nZt/3vDwx+Ib+
TEi6MAhQ8G4yfXNAxj4wAOvlydreeZFU18b3rzrug8pJrFca5NOEelNWkVnS85EgbQUQEdlVxoIz
/y/hPLakPa6V9eqdcgWMhFUOTcEMl9O3/8mKlpWXKS+4TBAsL52KWqpi2cbxVZqUfipTweCv3nAf
s79cLK38Q1V/nknreJlKemBCUQVJNf4jwr31aBYHx+qXYIcTD/PscOB2MJeQWGceIY+ZF/5Rs9vD
IjZesbd38ekQ1D7/LQIeZlQGJmO+MADNrNafWo8tRcLmYr3RvU1iHsYak/H+Q2S6DSOs66HdCvs3
Ms+a/36PjQpxE5bavRoutnNYyZxRztMlqk0U/BZGCP5DJH5lB/6CUTCvoSPtrt+9/HE/179H8ZwL
tdaazPnDjX41nFYpkmUPVVALH+3GWU8kN5ArW0v6upho1yAN+TV9eThAlbHu8J3rjbNkXMMgd78g
s1W4XK8IBOGitq4zN7Wz1A16gygw1hD6CLBBgygnNz508PcT7NfYSTbGgCyuP+eGHBhCMeNJByeJ
hkTasDNwmmb5edVYeujTZiL/V8SBLz+kTs7WHt4I1oxhzNAQ0xDEp9ZRVqFD3rn4aWfpAtX+BfsN
VW+AwNA53/9shLyEzkya4z7fkPOSD5nSiIDiVFdiZU3pJGADLDe8N48aRuxppvR6PQrmhVFfJHuL
ItGudNA64rdx3As0is6Zju5RKMKHjSQhDFIBHp7Moo1cvbsXYPpvo+OuXfnlkkTvwR6UWbXxQi44
vKvfYFzICRqbv4Hn4+kVH6z+bUmZ55DdhvkpG9JtfN3tlaskApttA1T/OdtRJEvaUKTGnmPOdeSv
LNv4bAP9SoQWvPYDIsZ9MMHZezyILhZJk4E4NZA9ARsTyudgv1ulyh9xTT7u8ntkDXfLSfNZES7a
Ty/aVWle7gU9eKWSktyvVvZmkHhT7ngtbuDKGfwr8qwuh6bSPEsp9jyDSHy9eRqfkEJZh4Oi/m7q
/v+LhhbYKpuEDOjmivmj0H9ixdf9f/Xo8TqsaKUdmBk7QKUhL+Y6IHbTOU1eCLLjQib4Nt9TCHe+
YwGsNgKKf+okq9exx8HsAkVpQFvfDNgodOTzokuAHr4BwAZt8ZRgjvMn7l/dq+UAwVG75w31l4jG
9hk2EWON2Mw9jXT1z6Yd2C6xh19QqxaHB1/As2Y179j9vmWlwR/lCMgmK2ws7oZnkplS023c8/4q
2QimZ4kKLvk3VITUh6VRlOdmxSTFSUJrotNQf2TlV/0YCORTHujqhXihsa3UR5YyuJ9RhGb7YM6m
VmZA0Ln9jzPbWnJDGqnkdddKHINwCv5S+8mvRKQfy64AbRORIoP2WpnqCWQmHc5um5Vd3yTKC1uE
byFhBrngTwPF0TcLgtg9kBQP5DgzHUizB4+3O0tspIyw1gCfJa4CA+gSikOO58KviylFe5HPvyHp
ze/xJmw721gABQ021nedRQqVKWFvraURhmAzCWX/DnyqsLqD1q0YRkXVve4uzuB0z0e6j8UjsbSU
faONhZitA11K8SQK3wXyLoD2bvdXXSm34ywMgg3pzN0Gn9HRRvaHQwmPBQy9V869h+ykkUQNPqdW
6Eyxtpz9jGs+BjtXefHEXj2LUYtVhip5GotLcUwN0GtxHAzfAXV3Z+rngVxZUNw0K1vp0o8x7VTJ
zf+OPV7t61Lm7guweJWn0Wccv6A1b4YTtBJf8eY00Wyz82thrSTXh1RVpZFkUWz+iD5B2AeBabfY
b5/ahntq8ZhAZlev9AFw+71KAZql5gFZ6Dc7YoMcvfqU9pHz1a2UY+rQVaoOpcGkiCfQRRfALUM5
LtS8V5og5N0TJW0P2LDb6BDPesvWFtVMoY/P65NCKMj7PgzG1/yeaLWHYoZtEUJxjwAfalMB4AQ7
t6A4sI7V9UZQkfLQSFPzLgIyavnq8c+HIt/phS4dsPXggmZ0zj3ENHX6RILNxT7nb85i3efsb61m
rjIjLv5CSoroSC8HQB84mErxBJerTMzceeuQzF1a+jjP6T58Eu5xLQtWRoqqk3n/oPYOa6Lgpx57
Pqdwz11l/FRfM5q7q71gdqTcKivB+C9Kki4PUwwz7VVElnT77nNIuTr6EZj0QZ6xBo8ggn6PcEFj
UVz7hsJFd6TpxOFp3FmKnuBNXwwQz4uYg5T/NEDjpbR/EG9QJ71Jep7BUAN/QUHYMU3SgmJgi3I6
3F/UWIujNDGvA+ZijOK9hi03o3Tm0DOsi6zbKlkTFVQGdajTlB4kAziD2K2Xc92FG+Za0FSU2Cm9
kg7XyihjeFnuCYbOJteU/Exr5iIUgrqsSyzRmSEQ+1syRHrhmzOY9xuSvFw7bMtwnMV6REDC097a
uTaUvWW3zF2KzfUQwoZodZTro2N3qGi+I9RuZk3C9EhaLkIypBWl65392YQg5QE314WU7tcGJXXA
vm/kRLrpd04mC82u+dELndJ8tiYWlcMwRs+DpRbb8XLXLUul7jtZw72a1AQ5HPonRbB4Me2eOjbR
lFxnsjdaqdx8B3obzPNCuuju0WkwO6YT4efBbDTTBFk3+Vjw7zdCsKUIaLDrTUT04SFNbLkiuv0H
A2bxI9FNEMBFvBREAVUp4YRXZZPtqc2A/GEaT5b4stw5Ft2nP1BhkoTGxepk2qXfLjrh9Npxgygx
4fUBSeCv+gW+1dgLzUi5zbCfP+cqGYZLIQBKahLl7mD6tf9LYK6mdqLV+sltCKPErSNGfmfD1qdj
BhAeqaUwynBhwR4h4MyWWseHoeFPApU+M2SDqzfJ2pD8Nu7Z68yM81WKBLIE8OtLVTkejN7Hbfc/
fc7ffcTm5MXCB/tFWFwqOjPO04S7JGfmzo7nMKHYn0JU2YXfl1oI+jGN036DlVOMrvpAASRG08WL
Tb7kltLd2cV+hDtjaP/PmASyyEEDH8HmPuTcOvud7nVsnN5VVQZr6iHHgc1WdKbpxrpXcXsCOEaS
nTl9ZOu2JO7wrE34BvkVUPTrW9fNRrzEejlrqf9OtrhTHaWRDIFS5zDdmrOmisbx1WnnBv2klOND
ATfgwBB2BJM/TTF/KjC3fQTI2/hI1NDvbroyIWiUvA1WamRbrB9R/SZvjxlaLnfziLDt8zASHgW0
4UcXn8LsQSzNKcdUBaOUlwAgsWt2dHlUNdEoJmkkMv1XD1beMxwUvhIFvcT59LcJinGyHgUs20wa
GYHIuGughFYtzLMn3buGrb7T9iaZreCE9SAiWWWwZBTXtq4QkaiVtQX/Deqi6znHJz9GOYERqXqj
DEmCwqRqqw1WefjnhacZq/66i7NBrVwymYAAHYXsTEIpty3LF7qUmvqqt5VwKYxVCg7ZtgjWNGfU
2izt3J1IqWJU3vctcazWoGjRwfKBlXfwz4dC6xGQ0gREQxiPEGDMrsZsiIN8g8gdpOxEsaXQ7K2i
aqrooEzKlL76GwqS1mtE+ynHzddDNXQ8+Je/L0LANop0Ir59yji41F1BD3ZsarL7Zm8xYEKiqaRK
j2nyPUctectNwPzROTBytjrlX2OlKGolHMCgLXIaBiDWNURvTCmVqarDxucjbvMvpK0LaYJCI3gv
BmdqAOgb4zKTuPxL7YCdmaS2tQwY7/SvEsMh7f05tl/U6swMf2gE2fsI++kAL3AFb7LXp1vdARMx
y88UjfhFt/ckQKve3GoI2c+NJ6LlUEdtAlTuORKqkavERlV6507aPvpyGd6D9iqSwJ2ON+5WLxVo
Cs/0DkI34ViMdhWcjuMSm1s3fSQjKlNrBtqb9DLPzwwQ9WK3v7hThLereN3gZUzw2wR0ICIxgFEO
2kuJs8RQc/pvxP/BWN7sE7a9ktM+LLN+8wdheF37gFBcDN/FWnfEF8YJ2qiWTCQ0NaLtrfXYwfhr
sFsqqc25R8BLx5ZiQpP9UT1csCMFihS8cb2SoeZMPl7QHsvY6HXAozVk6XUN/k3KdJ40qfYK+GEw
1XsOaQV95x2fcacLPNTtZ4Vju7W/nfDSDcsJWhtQxrvIFgtp70EPtxs9V2O/rBv2Di14bD5Jl3sf
DKvNqehfRSo6xJwUJm3MgfHDiR48E7QcJfN9cB+awJMZFOC5QDvN/WVFvmYjp6qBenFcIFWSf7td
wst7EIwK8HtLg6Jc1nS4QxxLK8bUmUJrk9MC/hW35LI/d5Tr9Wa74vDSsxWzk/YzYxBoZkyKxTA6
RqscDWq5MdxAMdxI4+Rkb4C95RBR/Od6VXfEJzECPq4+hdpvDNmBH3AJVk78gD3sYcOLWm0hg6Lz
aq5awOAi7J95vLmqsiDbquwzUlMiZdlvNdU787Duj63JKQhmOgY431zF0PuIZtsjZnWmtf9wscv7
A7WtLexIEkqRMd4YgVn59GJ2UIReE8oykPRQBSXqnsHp1CgkedHxF89GWMVyK6Bo8wGcEIMB3PHO
/Ecp/CYLZjorJ9A+XrJ3k0C50I59P3NkuflUvZQLMXY/BwjycbNuwmA+1DDIn334Dr0Cv4tc6jDc
Z6lxY30ufjD2vgBGvdNx2UU8FSvayijyt/hJ8XUEPPvbcl4mIQWa0XFwK1WC98upb15N9Z+ki5Ei
dCt+UfOfANihW6HFYozPpnM9J+ws6ajpfOeiiQdePyTD7MmJWrWorI8uX14MboAlJFP318I38Vou
FRE1Fs0N0Q6wB3JFou001E7jYERIhZOv8d7C4gL9yU1WNNf+R6K9c+o0wOZXrX+xrIMMaQUrqiU8
liwNYQW34s+jsivOtT9jV7l5bRgPtoRUZFgBs6Hsl2285H+K71VZoduKKB1HWh1XXujaVAb+BHjz
mlz37Qxnwi1w8/u/SxdgHk2Izh+btv8Ngc2yfdNHVJv1nfLkvmzDMl0DQU+jED0huLAj4nSvXqim
fa3dofF5IMtAAf2RDMagEQcog7ITAwelwfiJkLlPJC8oXi/4bJzqpA2YORQbcYK+7QSq5ruPpNE9
txmW2qDJ+ORMCulhJ4wyQZ+VUWlVNUSJnaTU8nRpIItdxdPrtYBuUAB8xye3k90k+MwOj7CSwZ1y
6b/cWSnKNa2hlnVp+QqiP8HeKf6CL+4vX9vQmc/UXnmQS5O2tKI6qsC4VbgVCnnfonObGh7fcJCN
ush8FaZfdAsr9AAXjrttI8aOdFJf9CG2qjtkjtgV0Yt0RcjTFysYYEeLEYB2LLDRz1LNFuFr8joH
eodaZCU6FyShzV3786BnAvSkZ3apYtz/EQ1oPGv99oEtu40YjcT1afT3nPH1N0Nim8jTDm3iMJZX
O2y+En2TDpMenqUPBpennviC8b5/G1FUzH0fKCHFAUCNk8CInyWivM0GGgc0bFPS/1HIcuwRokL1
xUodhA0AFbbQVct2cfP6tzkqcJFD02NCp20+9LSQI0k5rzlbIiskVG4F3z7oSMPcJvs4QO2raWBm
iko+mhwlHy+MWXBTb9Oizcl8NvJ5hxn+4+VM9JbRFdZz5XOM1hRLsVwovOZ+if2bTOyp7nyk61Ea
e4bWQumfedxddouxVNtXpoBVGqimOJDbT/aQzIMUFwGQGNaOC9twtPhnYCi5o1aGbVR5qC/zIsyB
jtj9/m+SZbSrRhWSMAcqMRiB52pjTNpuywnHaTpuJarDaPmTbg/7MuTO1pMa+6UH9s8D8C1vADrp
XJ4tQe7OkMDeW4tMID8iG5evvb9a4TRnGAR18Ec7GSpQGB+ll2mxNYbAlGOeq/qNsjp0MQMRf2t2
YKqp4Y4G+Q/9bWnzHtQuh/G0lUeY53k0PdJfVzZCBlIj5vJhTc1R5X0BB8V7ngGri0NJz/TD0YDG
vAKGRZXzbGLy6fXOfkL2D+L7BKhzsbixPO0Hkf8JF3VU47aTPZdJWpZ8LifLrk61mNwiYvNSMFI5
WJ9RxwEo2zUOwcQ75K6ZJ4DX0ktVONUYvvo+u5FNP8JY1PYUnCPPSZXOAmEScGRh6XQj3h58H9dj
DJQ5jhGGiI4x3QJegFdu0It/opQXE2P3iPnmfD2pfObM/avLQnjkm+E7y+yNOP7NpzWZ9t8ZB85z
rs4aytSGTjuMON1pWth+tIeiOwYQvDZ99t+kRNMojVA26xQOWPUgaf1fTXPREip6AubFzrhjg9TG
gstHYtA4MrQs75Og5s+W8f+LYkBFRHYz+EI5kRB3lfzplptBc9EHoqngkGmfBxfg8GUMvpOKKryy
Rq5WWab1/80nRd5a/cCOfQJ7Mh+qZ+9vygKMe8KL9wJuxLK7OKIshZGlrqORcohZNDeCqsUTQD7x
wa73h08ysp/7wPST3NcWrFLlPy/kxe8BsAOtnf/ymiBYxVmwkSTyj/5OYPDefHA1pT04JUs6Ckdk
qG/uweniB4Byrvl7yPzkbQEhwGmXAAbRj7AWW1S2LYV1IMyquT+OnLo8WwUhJS95VAgkzw5wCHPj
UF2alwHVxPQi23OZkmLsQ56fNj1OPid+4BgWA9KUByUr8Dyg5sRMaDBbxfalr4/ZYc5Y08zDV294
DwzaQPyxcDCXasnzTO334d7yhDES8xUXiuxuF4NymzzjmYlA17VRw0vVWzG/4g5BrDfmahqsu/cc
1xjVgeeWLHuKDBGvxtdQKO69nI9UvaJc44DSguaalr3ygmK79Iiac6gWQSpwOZh96XogI1tmuTql
QgyNEl4ogwTsTrS2hnf3KD204Uc7MNRxbBibirl4ywVIiOB47hqLiWyS/fEqoU0M9ZO7CgwEz1gL
PvkX+ljcXLFIIKg+TYG1t2bin2ARldDLT2o3LNOVDdYmQAepk+5+phFbMApnDB6Ps4uUrDWVZmYw
eJf7pJD8I+dqxFwq4SmR3lmB0AjoyR9NxhJVG0D96F6tJ91qKRHNz2GUnNdiDu1GlJPYIxohzB13
ELVtDBJOMAbOpcOdQs5ACfNIWqfuLUd173pIDaP5JM40OsJDbfCnCWv3bWM9ZfT9BG/f8B+gutrl
/9YfW/6n0mBI1EmbbzbOnAC6vt3i36xFGXg/AfcL8kB66eeBGbz3BWUztf6b2QQDTEAqIrV0gp22
BCoHOzJXwoBxDmjn5d84W3SPF1Jo9+R3vsvcuRVC4vHXglwJJOMqlAXP+m0hzZ81EpWwzqaDXfH/
LhlN+B8pRY3gU/sBHCDGl3h1yr0jqgVDVzqjuxojZfZuYDbIg2EqEtoCKokT8120vzZXpydlC89e
1wlr6S1r6xd4HNQLoPFxwdebOQ6rmV2LqR8RZl2ccPZUS6ID1OOuM4dWcfMhG1eazEJ1Pr8VfAP1
bscmKlJuy5r+Q5xDOdABIEDCkXa48XJuBikZHO22Nz0f+joI77rdQAmup+O58DGkJIZPAsdaspyg
PuwcVvYF95hcK+OoHNuWsYX58GeU2rNsrzhY38XMXPy1hdrOA7ewrQi7QlYDSbDvagtN2FFfD+DN
ZnaKlSALe5fNcH06OPrMpSTG+xJce7rGS8QmUxErlu5bgYVFQtQfU7VxbYw8yHIQsnImUNEvqSOG
IqT61wT43npYgAC7hg2qEjlMCN/3MpW7EreDDPQrTEPe5yAktqGXPCKRD1w2DRwOfnwvtk8q+4PT
t1W8jQobVHIfEdqLESk40nUKz7pQ2IOIjmjZr3bLbmu5THVoC44XImtysIaTgvcW0KWi7X531Cj8
7alfLtJPiNM0luyoJgKmKNaUP5is+iXocGaoLxvKLkbo2qv1JEL9xLZksWT07sxgEPb7VfKU7CtW
SymS1LMtkquJSg98SewA+50NyLZjoNlBgby9oJi+fqa8PtUdVdz5x5g/StTEJOewxRjdf1kV79Hp
yTgzFbg0LMhYuzI9YmjZxOb2Dq7jh62VjtKsFF6mjneFFUvbsavIyCj4DDcL97F7gzm68FHH9CU/
PM8x8nBVLjWLgMdnWUADnHbX0wm6eTlhN7YhDRWXJApbNwhp2SXoIG94oMZ5KgorQ0TXowY0Qan9
YWiRGwEnudLmJP0UvNoV8CAlG3yBs7EXIxWacppd/NhHqOOSTM6/2f+ht+0ksliUaO6oIX403pQz
QswuRXNvQdAjaRE2dd4C0W+ImeXiqzH4Svv+ngfnZIdkGajffM56cLNpbZjPdl03qCw1mGkV5VB2
/olQvIpU2NfzQCJotXnR0LWyBRhKFb8mB/SvHbXEJFO+sfjcRL3rUW1z+ulyWpLSqSS0aymdKkBa
iNY15i+iztc7das8thAsOwdOTTsk96CfjAbE1pT/mEj8offvlpPyCC9c27zBSg7sDInJEn8HsqC8
pzbMdfZIQ3xe//o+Wj8Iu/CSwAk3bhknzolZA43vvefoBElBhb3YxOzVQ+n75tqRGAtH0q+Qm9LS
fZ08w5a7yGND2SmQQzFDx5CowqCdi9fhjIMlDmzP0uNLfpIzyghrhX1mfP5JpWoiBgKYoQch/1yT
+zd5CBb+dIVvbDyy/FcTIjsnYc4twQYNjqhbHlo/rpdNf8yzzsPnjFPyxkHsNQaoAobZbbeosvA/
uFfG8s6i8tlPmvjaOTFSWOVLVUCQuqXLDg7odEv3QVjQmM/FKTL7GS8ytKCwpnZBchR9krpJTzyp
7l9YlLb4qzXolBS7i3s6KEiZIBUyiElP+wbe1rsWrFViiOI+OUBrCpqTu1auQlPOSeteDZIi+Wdf
bMMsULh9+ysHodEMbI7XTIn+TUlxBeSZQ7MTAjsBMcgUb9+2yt5utfsVLFJCEeQt/2/HsX14v/d6
xT9v9on93pZFYSwMK1Yfrk2qub7r0xWM/b3ZpXCIYbPjwUMJjMN4kub38bAk6+NbnTbJgozYKZtq
fDI/GmDsEuda/kyQjiSJdc0QZZLNprQEMZB+oS3E2CTeLiEqzeAommBbh4/REa+IecjjY8H659UJ
Zg+sA2/TANVkhC0WNdnz/K0hqEWrhVDAYTacQm1N1fC4U4FxnL0eb5+3PUzlW4kZZFvuKmxwD8eb
mTN4S+HP1oQUCIXuAmrTK5Xb4eGsoZRA5mwSi+FytKZYOzvfxYYnas4TJGB0StxEeVm111Sa2x1Y
UbzpUwSNHYwP4PIXTXw+qpBtFRIK874Tqep+6e2fdvLqWK1qxifkO3GmR1SwxRkpgv2WtYhmQp6w
DuYQ+ZSaSU0pMnmrS7/DOJaOoveUi/J/wWfaatlmxdkfRAQSB24OnEKXFgSyb+nUjNAeYtKDjYjV
VT1D8A2vlvzAqZDgFav6s9cfP0+hZzJJYe5oFNr2AbV7v3FoY8zq7DTenpH4Zat4GOx+vZKYZgoh
nT4wHlLjpiBv1Rp4nagyt2avUEJlzRBz9hgN5h/yMLQm9yWIP2P9Wima0nhEoGVLoVqQ9gL+IIIX
HOA2vjl24/95GYkMpGmIjcHGtnIME1B7w9j4Vs4k4bZ9j1DUN63HHJ2c8fp3wwuRQ248fXsknm2E
UfVODmdO8AkqLeqHI55t+OvpWauHODOZ9mya4HFUiGJVXcIXTphCufUgtkb2QnWywQ+YVSi3yEPP
HAbgXTFMwWpYM8G4wMSQ+UgGlnps6O1WsR5E0Taa9ERjONpoW8dsCSwHu8emnl11n/VWNvim1/vS
NMteAy4I/EZBqhPmjs7swkhQ3Ew/gAC/nsPy+p1Fx+13jzutY/jqz06DfORZlLL11Hvx9kk9eF5F
J9Vi/0s/EBUK4aPMBx5tJmxkAatVs26Iam6491Y1dIv1J8HUsDFonDnjGZiQJ6Aymo89bjAQUgKq
Pnr/uq433tres6gWCRNdT9VyrhIjPAxhNgWh24K3dl0FRiKs+FM5BI8lO1nsknoNiESxyLcB0mbo
i9qwtvhVBDFhJOXEWYZxzbVTbcOC8jUBz++mEJWEaTILxoJWk/fyFwyrvDY1x9Ocle1mYaZG0+mh
TkM/0UNVlD/xUCbvpAcSLXemRwd0tV9t0lliO5k+NnO0nen0tdTPoFhMSoEpJZTeJ1rDk0RHdT4V
XGINajDXNJw78lr5aMzoYnJv3TNEIfhpPraOvXrO7YefDDy+THXA7oiYwG7GDRCjpZ2LO8Sy8ehr
8DXiMJDyvHt39sx83XuuX/yVVaD8XQbn/M91tjEzq0Ccg5iWC2geS98P+a6mLrLZ6HS0wpLt2AFU
fFogjllL5RYkfMd7+A2mg2Q1r6fPT8y3UklRmzaGJBPI+jvxadxzd5XJkvsiZ7NLtqrcwvgcuzkO
kgBob1Y8ogNJrUXCUqWCZ1o3wLJdBGNVJOPKdqcr1dd9Q0b1VR3R2RwQuSFN+OvtRzMyNvanovpM
vG1IDORRyz8uv+/Lzo/8Vol78NJ5jkz3k2h/gKqyFes7/QTsWC8o4gswKN1IhNGwqrlO4SZywWwp
VUPG1usQC9uq/EzvKB3gNu5DnzYyPY+ix2RwkMuJKo9+eHmS/4uYbrfCCOKQW0PjO9NfkTIkuiNG
LPBN/y0LngTUuhjVbY1D4XjK4KlvbczYToBnBOP/s3O1gDbZYqDJNFZT104yni7p1jGi9QEsKUBb
xU/HRfhappm32r5LAH6QxF9LaleiYOpsw0tcSBxhQASrn7scIT2fM6p6xRjTE48knXFCZZ2Dd/z3
hw8f/YOK2zVTajMr4ZHyfSpljUQf7IOVHWk4oNRfGDp6VGTERm4u69OOR00oK54hZaDVf36YKO8v
SsZG3jVZV2Gr/1pyJZpMtkWiM4IMXPkaZVyApaK4AcV7VPVkFQvYcv2pL1bl3ATBWttlm1NpB8UN
8Tak8RrSrWayI92aKRjeTcPL8qvuS7cAad9skd4e93wl+xNA2vqPpV+I3/igXuxMK7NOhvtsfdLm
YcKMtYJPzlygqiVWuQmVa46xVztbDRdVVkxqCMtYLsH2qx/bR38pBQv5Qik7g6Of4Cse2mvI43Am
aXo+LQwD590QFhdRwNZYjdRy5Su/9pcjE+ogt6Gw0FJF+E7Z6FhYUQSO93X2sL7vVDSIGMFC30pG
e6tt2BJUDG++dnkbRj1UDtwbTTbm/WGVPkO6BKTZEkt7VEdgrER+/dwfLoBh8FAq+gPzeUjPUddg
be6Z6ImSZVD1Brv4cm8FBp5fEIVPPRUR24jQiX4sJJaieh3qHNWbPGb/jl1F17kk53IEsJELHp3D
+hyn2+ZC+Iu36/6lfaIh7eLAbKHp7LV0f93iNaILhqeJM+qLpZ4VZbzUjFeVpxvH1dVMQadYgPbw
Tu/r0S6pPLYLjfZmtSPL7segNj78L4iMZlQK7kps9RPjWEd43oQ2mlbiUXjccEpm9g1BRWZ0PeMe
RlumMBcWPhSyN9RHCf3zmTwIIzKg8T+V+ERRAAK3mLvylY2Z4Bn7jcK+dMLP/qgrgrGL2MmZGGTH
u+/WRTAsWk7oajkjsUpDrw4g3fA3AkoQq8I3eW7ELEX8jZ1HEcb0S50SzSemg3gQ+Qp1iUAFgPy0
sLmrGBFvuvhzjkLynyuwCMu1ZFVCZUwL4CLCPQLSwVGSRnB9U9XgY1lLoRlm6ILdU5d//lC7tVrr
hQlnyiQgEPqn5S7uyqeIeByMq+W2yMJPkfPEfHUYsnsN+wPCfSdX2WlyAJ1yGZsCBbKfQ7291mPJ
18IDAHXgOq1TiCHeHLif6aowV4DDMhokxeBtF71S3fgqdwDUS8NEoPQuRxj86HCqWhy9PfTRkprB
iI+z/FkjEDrpm0CND6sTBXBcMCLgSXG+ZtCpgyzLWcAWZbKpfPJRDPrrj1kXjwGgo+UobztIcnoY
l3b7YSigHju2+MzavjMbmg6qovkC1ictY19h/HeYmj+9WPdhC4fLwk2DMnw2nhXge7pb8aii83kj
WStH1CLYkliFjlezg0EyKsPXAFLVQD2f3ZKQFawyIM69W5QVnM8j8KiCLNxdy5Yrw9oFj9GXpAF6
fgzjTWmSTG/2pLEkW2OLqyFiX8ZfHEiD6tUX3PI/oXUHRe0R3tuCZQuNkopKBYOcJfLhs1fxUbiF
YIAJIKNSqRDCh2U2yiIYC3rJHDu/3C4qyu4Xq9ixo9ATaK4AGgsPbAX/EzcRzsWOnBH2kJeyvKk6
ZJNPLDy/rjPbKL8yv7Yq462gQTw1U6K/o1DITog9IdUR0MYSVfcyu52j1g88V9YUcyjhqrF2ZJaU
TaXrzHZfpDW6ho0mrBsqFXq35zY6mPZIQLZ/0uXfms4nyxNNnaPT2SwbfUUA01KhCWN1SvvP68TX
quQShJBANeHfx+Qo419Sjs84scXnMolkdwCBe/3cEU3/upcgirjzK25Lw+UYr5oQl69DzldPYwyN
9Ls2MyyUogiBov4/feG5KvSYMKfpvSrJsTTQhcyASnGppX2KKwZJjC6JedKYXnvrJopU2qa543Fw
uhTMGdnyMawFO4kCh1owINgvmR0c4FWnSBQ1QGHycO6eTcgizzE8Dv7XmugOIkweilVVE5qCgPmG
MaYBYnY8oMsk5Y8pa3T2u0rtKRIaNmSjFVn/9dCozxtCVLvkmJvRDZGXPo1IIUy08QHnoG5FrEaX
GtDpYkCSrHe2ImXJlIs1N95ZVDNCgPvecBnG/qSuWrcH3vicIZPuirWrvq0ZOnpUkc96s4sjq1BI
7THoLhsyjvofcDGNwdNuF/ad0CIqea+HZruWdvQNzipdaUd+Lcz6fzPmF9Phh0y5bkZzfSrPLh0H
Y27xIU7F0rkWFQ0XcL/X8VhHUwbzCCeObqv3aIqbt6zVYfqPRBNzmt+0vNIzBmQBIhj7aEHhCJFt
hAE3+YIxmxAujka/vXyoSSYKC26Fyl4zESmtbIrryg4Q1UqDXT+azl2mMrw1251VSl6Jq9gPRHQR
n1TpFOpLsA8VL+5fM232Akpy0Stz5HuX+8zDU7j5BX3YeMqOXGWAMiox2x8267mHuWFZ2HmYqPeg
ljJdXyj1cu1ScNduzOiR/STF54BYxMDSLTzizQHL++5qxYapYfFbXEWYdMm+EANq4c9GF71CCRr7
u//DQpkAGIfe4m0Xqa210X5S7lvJDPbCqi6XHMO5hlK8Deeb/tOTmBTlQb0SckURMTcievoLT7Wq
I8DaaF3KSoIooSw4Z1iWFEtowra2xdYMDLn+UoD82dSige+C98bXSnKr+d4KYlt3wJsohvZ4Zd51
eXE6ZbcdXtHyYRKJ8RR8tfk+ODYBIDhyNHZMithyC7TjFMpWKgk65STkQXrz0qAT5yuU9cmWPa6Q
Hn0UaSwItD7CXVE/iqTGJEhpnPphZzrKUCjbOd9TFBJo1JzpEqDys4tT4dXPbEvA2f0pMQaCnZCA
XkWmKVkNflEe2IsZpxfbBhh7iyY6N5APN5U0MS6Nq48eyHK0M2FjEym8U1MDGqm5Mh8+SJytRYbT
fSKoNuvnvq1kDsLyvGEcIwOcIGDvtBADdY/7Gc9VtRxn+ksLaIkCgy5rgD0vnTNH0a1iaulOs9i3
CTPiI/1WhZgjHca2F0bg0gppzfa90o4oMMoSV0TQugAIIrr5k3S5nO8ysTpFqlBSg82lwJSPVs8o
j5qGEnuUrU8VQ+7fKnU3oXd/XAPPt1YjnqW4X02UDamGKY0THu8euMdu4d0ktIzhXAISDEHcJfpa
2WUPmbqahS1/HEPODTLbMaXIX2LhAaHFLr3PUbpCjB0qauprcNtYkHfCR23zNSEXoUpfy/ZyGTJ1
Bh/uQBXFFqnvPJqSXidM/gst1/Rh/RrhnCVnYER6G/tifKZuqhMJZx2Zk6RJoFiMlWo/l4OydS2X
12FRt7sT4B3qUGYrsngaaM2sWoZ/7wwplNzA7AzXsrXg5c/bxlM37tITqeif/PjWqz6P72CC+rri
Zzcifi2rOU2AFbLepcRv+FcTzj6d9ICKY+UqdgYmXehFxihud48/ONJxwSqOQp50fB99W2Ty+RDv
GNYKBILDBRfB+Lq78C0SB9ePMQ8A5aXs7wUaY9ff090riAxLudJSK1qkQsKuoBo+fH5xdFalhJXT
AdV9/+lL6l4oBLcfjWV478wUdiF7edq7d7az6Mxjfflm91Ow+Fh9GhSJ4EBXVsEvY3VBIHzgKGMH
mgy+oxIYTYVtsiDwbMbybl/fxYn0cdrPNyZ2EoJseIZI3qaXIav64Cpw+9HebihxRJfq8963jBRt
lhqwybTrwn4C/C2vE1N3p1ztLF/eZxZVkX898RUuE4QjqU2kICwSNBRMQzeDRAQpeBsw+thXU/LU
vQ2/01TctbO8F3b8f3mkCF506yHxRd5QEa//HKopFgUT8Bg+5vRbLnGPEDdfhaFSj4dnh5Nt3jVV
/2Rndt+UDdi6l2L03Z0V82IuvcO+14CpRVLRB810xzelIqFXssCdC2vlJefFct25lUZTBb+Fk8Pt
hCstI5qe9vkZW03HsUskRgIgFwHLuuR7lwyt1HdTXiqXObZLmizLJNeXzPPyR1tQe6wyz3gZqf7C
aDOzHZzu3VDX4hhgLZnpf20eAo8+fY8VdYvy7vEjCCuKwBK3fn3pl9LyLvltSjvk1kLRS2Y5pG5B
2TuyJCVI1uUxzN1/A87A0LzZH+XRg8SZD1q8dhx3sBLCHqfcAFiW01E9w/wrKFzWWArfm0SHbsat
LIGYnNlhBTKq+7OzpJtIaqyiQHizP2vsbGD2fUGadSU7zlU8f4lzcxPfHh9k8rc/OYmwDX59xjOr
OiwlAlWsBVhd7RyURUpjiK4P7YvZnj731S+xxcTp85vrWytnGbbuzJTAbzu9jkUCDPc8k0Sy19Ch
8gx5exY9nH0Wn1Ey2cia80MnGpCbsDfhM8WhhH/Vwl6QXQCj9CjpeVA8KbNFcFauK4uxIzb1Rb+G
0Zoxz8uQN7uGvuNFIUdgIfFq36mwiPLKktUb7f8q/PZLYNk8z3bNaHjLnjxQQ2fzSNJbw5Dt1qiY
Uymu1sO9HtZAFtIQtS1lz/d7sh0MitTKqWSTBeq5AIq7KN9GQM/uFNLhXiHWCcAFa10F995kmpAX
tcOCFMiGTYnQs96ACTbQE5sBCyNJBhi3Pthat4E/fYtgKfsJootI7Uwo0E8vsFKeRg2PRxf2twi/
3VWU/UbNeuQBUlvPfd0xO1cUCIQX6SKcgAJzsOJQapxpKFZCoyHedgTWsiMSrcIF1QqV8daGkNhE
RCIMkGJ+Dfx/10uwMyU6Vek6iGqz5RCgOMQFJQqdf/U4fS3z/eUTarslGj82PLHhW5ETyhY6fu2i
qk0Wzrcwi4z0w3GKDvdbhjyQEWjbC9YhUxYy9m1CWi+li8jn6J810aZC0yrLWpGS0ouLtPtYAY7L
xduIAL0B177v8J7BJys28atyelD39REtkPNIrR3GbnfcVUDCL7KGCkZlLXtfLgkx3S5YSBL1NuRs
jbdyPIUzQSN+2lcUVWkgUr8N/zC8D7ErehGEfdbLTnaYUBLJnIWwLU05qReLd4TEJTVS9iSDjIF8
EnUT2t2AlwtRKj/2TuGcqJg/E6ZImqDfv3Vv2ojGUBvATIlcFR8rU+eKWUZ7thfnK/KnTGRO3XPi
cqtQ6tU2m6XYXH2liWv/KdiuY0O5uU/t/vODH8U4w6SMFu9/9+D0IuKSer0nKxauuVRFu7rpTve2
CoYFbEi0dW6+z5Dj1DxQYTskBn3tG2WvMO29AAUbkAArp9q+a7VduMSgdSd2a4Y77v8iGq0kEtVL
Ivm/kPUl/6+fcVtK/6TYoxBTFaiss2rGHud07iawW8Sd7QvfcMTLJ3oeT22JuYcWenp06VnZ9Bmk
ZaqTT3DgMR9QidprG6kUL5j/qXFDYJwZBT3VQi1MV6mlUGtgswhXHjsMWG506qbGSb+Ykar9cl2G
QIW1k6gpDds9uP/+mdRTs92aROgv4MxlkKRzBsbe/FOxE18e6YlOcKthpbe4FAjgI1Tqrk9OR8Go
gRXKkhq5jxmkfDayfxk+L7eQlq0ozr2b8qIAVOmUEGLmrsIQ7A7YF/XH51HPWMeHt++CQbLi8s2n
NJMvw3yo1k6ncBfWEjjONRxYMRYMiPvcAICcxBOgCHpe3aoQsiyMw11TqYGF3xeggcma9nlxehnu
rGG80FMF2BeRRMOf6+qKG/fKszNFgNL566xWHEB5h5zbSX1I+Wx7MPdCerfFgfS0YDmEThPvs8yo
7ExMhNzSU0DjuIkkYHHtc1FFhrtWFMN0d/ECAm+Ns91hXZMCAOF5z1mzDMEvE9erIh4/4QDahYm9
Ybqi4GLvN/+l+R/iTWWoaaiVn0xixUg2Ex7EmPQTbNNkyy9EV3/JfvwD6JGZvR1y6Z+8hCPLP7hL
TlmTQA986oMJ7xOEKO2ONiZHsTTf+h1SW6RYePaGGsfNh6bJ2a7uDBTTGozqsOwYp4I/R1Vdi53n
3I1Mk3/Jm/BtPlGk6FpHAPA8BRs/RbqhrgmafJoyVrXouVjHjU2EBUiXAjP4haN1uj3HFWiyW2hH
dZ4YDEOhADK1dTMUYqsBEUu/sq56Q5elFx2VKW19ztPlaRkhy8uOdY5EFLiHTJJOjvRge/LJyrAN
A7Ti5OwqbMi4U8oJ0k3bMcmhR8Ulxz4U45o8QcxynjYkymz15/dj8YuU85pQvZ6H5mUNqHgiojZF
VwNlKryM+ea+58UFYG2GWIHewbCWLhn3BYBi0urQseh6xIxI2CPeJ0xOIJIzxZdTXeYzNMyd/hVT
TmKqm8orO0OTjDuiHrm7eNBu5qdtUSSQAYi10h0B4SPdkeZPo7FZ2FdvXvHvATQO/4IEmJaRw7Jh
I0kCnd7wPH9V8dHWpBkMJUARqB2Psh69evGWxnG/C2d5325+j1gMTle7L8akm53sACBK17SThKTI
hQUT8csTPpU9A8H28A4Unlfa0QEHgFtUmFk3k76igJRZ+wzZ2MX82ii/V0tjc7J067jRZX7Hb+F4
uR+P5kNVthdbE64cKfNz3vkQLubmFFe+7z1rXGpjOVBBibcz0LZqVpLbp3t/K4omsDVT7+JnAvrM
6hXKsE57Nr7IcoGcQXryvgB+qS9OxV5iFOH3C3YkBQpUyFvS30M3+B8Pb+NxwXwHLldV5xNW+JSL
xuqpgL5PyhF2V58tQxWBG089wRfDQ7owRFiWbjiZ7Kbm0PpBxlEbaHHnH0ip11ekoKZv6ak8Ozi+
p800jD4mU/LKCnZU7CkFtORpT/YXbWgUKsBCM3g5V6trZV2nEtesSvDJAJLYEyk+Ng/OLExk866J
CiqncObjpaUvFIrbQBcTt8MySRDIW1xyFeqUdnByRzL5sAxHg4mrL8wcdg+IpN/7QkwRIxwo3FDd
yfDNG96lf2HjvjJTpDC9ZQWcVmyQ6nr9SaEs499wG/P3LUJ3uTyWoryH8hIsSZ97ehp3AhMK6CL/
iwLs4MqYA/zuhAVlhc1+mLpMwahAbNuX8xBTKo3CGl8P0Od2SD35/cb/V7IBduRz3+fWjRnmDomi
NvHx44AU1BwdeiHMf525BvA3Z1JmUD6RNsXexYaHmZK0hzX/S51Vzl00HW3iiU/cxpxaLS+IubCN
CQQQ7UlOHJROIZk6cW/f0XBcjTrTNBnZE0J59nYmXNE1ip529mHQOCMrNMbEXDRY5GOOq1ywW85/
kFiagSsrmupT/sVxiZRV0eysroztKw2vZC/s3VRlhhIqZx3a/XObpPg8GCJCB0rDwqQ8t+TU7GSK
kzogzehC4vROxKrnSpQeOy/1hD75hKIB9DUBVcPf8VfNwnYuMDaeqTQlOl2XGVQhACIfh003Wnrw
PuYUTXuPjzLanntp8yxGduOIStDUiz1vJUy7uJ83HwhZCYecpPelPwVNmqD3bie1olLmm8aEIpz3
kvjlXjfNegBCniqf6wrBkF+5mot1KGQZi3eZTaUOTvZ5E726cWU12oFzZlE/pfHPQoiZsnsUPeeq
Wp4KGORLsX/4WVEroi+p9uvfj/6AsgIPad+Y0Dl8VpIW3UYIJtNkpXasSAv+kh0cT4KJRWEDx5UF
Jhkp6Qo0S1VnyNUOtpe9V+a9m/5u+D5fxQmbxmEmgpBsvTfzGXFB/iEQnZB7Zk4AacVmIBWcVgOn
5OPNjz/gbdrXFDe+fU/HF/i2rnidwGciibtu7pyaGfbjrJfNTJE5BNxLDZWp/klRbNTSK0sA+4+n
iBGto3lkytgaDAFeMYPtUEab1PgbzEcFii7fnyymhuRSZTEct3G4hMepvL490Qex6w6jyfqRvY4+
qO2VCv6i+o+jmZ4YPGL4ebALcqi52R7miALXUgqZ6oPb8BD6DBdkcBeP4uoUzGXBqn7QsfWBzADL
ceApVX5oaj5FAwJ+iyXHQ1WTM1BUON1PhLQwXsGjfGyBFQnYIoS9Caxn7bO/wSmaYNnPgtiNi+ZE
tgNksAxwJ0cB8p+CR1ujHgWPtA6YmY01EYK5ts/+268yxAR+IZpLC9gPzxPGRMqj+fI81t0C5M8D
CRpBu2dPiWgV6u3Zq2uZmXMGs5bGigYnCPme9P6uqTGcprj9J0z5WAIpFt3jihj54J00TVWxE42I
l6+tABvS8xoERoOOhH335ho/ojqnKdLUupkYfapXYKhhcqHi+aHtRolJOU7aVKfgCPW9z/BuIPCv
HaxlfPg1tdF5qF6pqUl1MtV5ysRHl3j2Ts2oYYbH46rKRXhQPITc/E2Mv05p/oAsraWb95LCoJZ9
u4DYKgxwL11hKSdw2rF8A7Un2df9jvxZRPGFGYl3J1GLIYeaN8y1yjzmr/L6nDOXXK9thr4/o89B
iHv5qIfgHVVLvi+XwmlTsspEHMehRzbdWRNJL366ZZY/pVoyIMdj/EwGeh7tynZJGc6JlPi2kxeq
3foVL7wlAOcR0BxI+BHF9opFBrE5tcNuynS4MB5WeZflQnqyqj5RVaz55gxxpzUlQ6CTiFEjhpM0
HRmn8+d99UKT9ehfP3+0Nw76DKdyrt681scu3s8AABC5X+0yQFBazoYKzf/PmqW3nIDbhJkf9+5j
LTdkT2IwQwnwlRgG7BKDmK+Exf6V5fGGM0EdQ6jaZJLVJDcJytHYC5KR3Kj9XOCRmHCe3kUK+1xn
VG2HEZPK9Tg7fRgVk1OFLMsgsF69H/Qt0qfptGY+Bhvo/b7OpWjlsW1aCtEqoZsTOrXxkmSOYaC0
NcdzvFRza5YLBN7I1k9eZXsYmyd8QgC2UUacuaGsRAvZ397U2Mm4EsAB2tKdKQe2S05n7FH5iQ4G
E3QfRIqHoEMXb4mt7Zuy+meph9BXIN2DK5aQVYkWw7Oss73sQVdr21VTXx6gR9oPOYnsD6+17YqO
wVvHOWNKoO6HwMrsxncQqcIshOdIrlhGaY+QltfRvF8jAWCG3K3DMRYdJEUTr0zQSWTM0Kj9CVra
pl7ibn5E/NHYrwCCZRaSYIV60sKN9Gfy67EneEvYzf3iIFV1C9ZG9+JoPcoNyNp/qjRgsDz47Hb7
LidK4BQqVj8u9rqQy17fziwYTWVgcMuBb22bVyHrKMTqO4wTlRKEGeWP3zMt3uUeJEbwPBo1XBSz
QA4hx2xNP6WqZo10HLqBsd2LKsHoKDFWGXtNoioNPsgllXoID0KDP8VGWnK3OxrCbz9JdE6/poTA
Hghu/vYzMLwaV5gHHFjFd8TSZCky+PIHg3kWhpqyyrIeDVZRIgLlGqpjYl5E5WbEXD+K3ZziJzZO
m5E8lib0sHFURLomhnysgXI/5J9Y9+20somjVOn5TrO3U9OjdfLaiaB9gw29x6YOqcMZdmgNFC9h
CE0p8/3u4FDX49GOFAgeKjjULVUNUtLC8+qs6sMKP7k+hM40nVWvzyqRdAoAPB7Naw5Nl8Nxgprj
6WY62x0Jy2bckqpyeT2yKsrhCdaOylf8izXt9fCZoNKTOZQYQAzZxIpJsXZtr819dotRuZe1xu5Z
faJsV0fHtn51ls6PPHfrzCk8/ZLk63p7Ql6CFyVFiGieKxKUhGHCovKk/eH0HjgMrBBtfyDTXB1T
B+A/uFTV5AoufFXS8+xoGpkLWnAQZulYJF8g4O24PKhgTVpM9bGBNSwoUOfpcFHQspwnzbJvezMu
5ubOApNbmTYIaawhvuPixLW7hr3twemQYJPy06L1gVxWvUOx4iJKpeb2204VXNqsI6a+UbI5WV7L
hwhoeHX/Yj4xQSmHV8gvp4Y4AiguGq8NoJaT3kleQc15+RNLpl9ABbDevAGCB7U4r252QRTiVOj2
MwaqzNmR3aJnqkd8uaRHNLWM+By7eHd5mZXgh7AzJYRINwIydpO2OrSpuuhN+ZbvcMHZlpsYBJEF
W55103D0hql77QILSPQiQb13TLs573yx02QL5D9d+/obxlTRNXu4h8jW6B+YSQJOs6ZxsCSX0XHn
RdsyljGG4dp5r3PU4xYNiPlMFEV79YZ6so1sUW8AJgf44/EAga4IDez9TalKruDSepv15o4mtt6z
e3R3uufUKkhyjQRv91UwWv2fgBaMTa3Dec+8kfR9poxX1hxFfgMxVXKdJQwpp/loTZOB0r7ppblw
wOhMxnobTtM7kKHHWW6OXM8bkRNaZGtBZg2/LL16ltyvr7mtHptSjuzH5u5lHle9LqEf9xJZfqky
GoTibN+lOifkjdNE2As/0sE6hjohZQfHKQn9Vljf7hOUI3UYKk7YVMagTiHP+qnZq2ivKT4KA5rN
kSGfWCMcODbSOsXc5eVmASJ6TEhidNRQb0YIoze1rWKRiUNAz364nLmPcJ3jOWgjtTswmbzj9nAK
XqYFKekmTrwgvHdW9AgitM+iDtXTE2WIV35G+T6qcI93Q1RSpDtUqYN2szK5MiMipq0Ow9U7W0tJ
/49w4bh9S0I2DFXmm2nWtQa2+K9Sv7XzNKx1uHYWHpDdUz3w35XMgGY4ujas6f+DdQzQ7yW2r8Ge
OOfaIno8Eq3RtfI8RBDPNAhjnJbGzzJmECUGD2mgHtCMetpjXUrj/mWFaeGx8+JCY/1IIgHCfX6w
HH6X/6sJA1jfd8vgVkul1PSwfTVHDqYfZ4FsUSGxM2ERZMGY1dW+zIbR7QQfGILIsllVI2M8O8fi
XCqoE+E2D9JTNN736C5l98Z0S67mTRwFexOIC9bvBBm8v+NDhMgT0Np3MUs+fyT2OwNEgg+PMb9a
8zIwnIbn6ZpVUebhThjPTSwby2ZxHGLhx9Mv5jQye5KhNBLj26tikfdojmF/5U5pnjvnwl2IpZkR
1NT5YSbpw9lPMf6O9X5vJOgx8jGCpIOUJVauXh8WjGdQC2Dc47IoIUtyI+EA1jErNoVl947/CsjZ
iAGeMCIndgy+511y9bOjTe33066LghNpssCdhyJNKq5NUOe/attsVgHCF0cqzj2THoICxdd1QuNU
VrFETiXN9f1/6ka+pkoi6gbneoc6tOjQTS/8R0Wj/W+vEXgq5qv6lnFb1j5PmBYkuHwexodleXmY
AiBMqzcC2RzqHfLliDMl7z2m3IiJwTBpsHlUUiy80hp9iPjqd+ubBgTV8WMYYcrr1YhTewnHZY+M
tJCjw9g/J68gL5j3ZnpPMntXsBrW5tJVq8TiYuH3K3rIvY4dEtHSye6k1foZ4djHBwwCY5+0a8IA
H8Xl+bLJ76RQblikO8/H4hpAUkzGKg/ja+Wd5e4A/FEPLerHmGIBLiBqw/QQ51qDs7pQkcRjV/7n
Ip7qlEWp6y474J0QGvW8ZjGO6y2rt8/0QcWPFfqNcG+L64FmJm5fFZ+ct7djoLXf/PNdL4y//5NF
c+XJU7Q26sVG3mkh6rD358O7QY+UObnbzRRPRWXy0m+9OT1qFKdT1WCV30GB0vk8uHPIW5rA971u
LkLTCBkiLAunp1P2lFPIGEUMSVNYYinniTc2FMhzSpDjKmFs4f9wdE6GGgyWKebEBNo3lIDiov+V
lHssvirTCRZK+WS5nqzRz+AibCLkzCQfgG7xvxSt73JrXssyEcgK1dDcmmHh8Rczx1zsvSrzGsdB
RYXhaBxYk2oGU1fjGtPlsv/uLYQ3OEo6P0ao8/xmCy6FT9XHcryoSqj/rBpv1s1HaF/vE9fY/Xxc
Tu3KEXDdVaxX82SwgDeG2f3cJTd+k6Fxd5n5xH/fwO+bhs9Jm0bcbdihjgwpJgSvd0fv0SIKs2TV
lqoKwDvOzZ3Gmq4kRb4f1aogkb2V4GgNsD9Pch9WwjAbC+tuX9/+V9tTFI8HvFj4C0ZVNFjjSKj7
Jc6sa0E+mCDkZQD3CeZ19PgEmP5XsNlvRQ1IkjR58dLdutkymcQ4Lmn9N3H121qqN1mg5Qfge1PI
NiIAnlNgB2h3hxvg/Uln0VjI5mbKuc/gpqiNSukiEzkhM9NuCNSlA9sHZGRF4MPPJIE9tnJOicxZ
hcSVwgbFO837xnVocKHxbKYjQvTjmIa+Bx10pKYrZE+jkmWPeK/4fjHZL6VvGDUPoBaWKnrVY8c7
xFlDGasqyaW76Out/xOAIIBqiUBVDaPjOPcXD0T6vy766SPig6Uswe3ZoJ3oMWfYaz211jbR5lLs
gslBWxmcR4ulleSgnPsE34JI+17FFMjhZL0s3srVt0wEreVCMWzxEqZfyQ60tIVidSPMTYJasGqA
cM+lLUe1KakR+jL1Mx6Lh1/O8HGMajpFtLOy+8ocvqHxIeZL1wxto+1xDKZik6+nSJHxQbb9N0Yr
4DqzuhmfMKZYxv6SFJhXosHsCTKTLyH7WyzTKs/EP1Ny/yA0qsre8965mtRLIuJSCIyHTdNQtqI8
V1NxluYkhKrj7i2dXHEy9JRAuVE/7iAsPd4oVH1UK91Pv+pl3xBTVF9BFbp/Z8+vfmZqTUqRH2x6
3eYgiSZ0EmzmyVIXXVLPk4bOTq53UKTb1n50eV+QEPK6E1ZfqgNfzCdtUdpfBhfAnRmsnDfqLp8b
N9jKPX96+/QflJ2PrNOsSaI9xkq3OQwefMnmCT1rugGFEWIokmmmdatyDcA/KAyDUbX9h16OMEul
7Zcav2BL53LxymcZ/gHXEl2ARF925RhZjRcy1ojU+s16rAC+c9HXt8ZyJ4w1wlIA4lJtGDbL+w64
5jWU0L7fHuSbTCwHcvlN1UzSwbdVT2bUEyojP81H3r5H2MofPmSwTDcVelB8kWJm6KnXcPQ53oER
LNrnqI8uB6I3qONYgdRWqXkesQOrJKs4LiZEMvOYznYQUyoytvwZkhtbTag+Gws4pfTkJajRCNqk
VZ2mzxk4nZ/sVLoTV5Rn8n8kc2Sx7rk06ELu7dNEHSiUeDgHvUFEAIwWu4kB4X1htXIdq43INAjm
yJA99ALGoCOu5UVP7hIXdoi/due2WbsVT2iZiB21Rj8kHLOPMdy3O9JvVWJYEXWnlnyKjHw2r5qG
npV/3Y3oBMSZR2jMR2xICK2d6FgzRKguXaxO6YAFSsoTy7u+W/AwgI7CVJ8y8dw3v5ZbORmPXqI1
zGvGBh92RVnSTbZo0v15oNkRpEk2qw6nuvXl/+eClM2+3CX9ciyW0QyakDEIwA5JwxcWak+JvEcf
0ee7qqasApq0z840LMYnyohC4HFpuqmJsSgm76Ju/nXVojPQfHOKV0Nnp1+sRhTch70TdiiEnBoV
7xjjo0nOLgyuRTxVQ8s6cl7l1yFgdUZT1jA5g/oLH2j5R3Q3yAPM/yLjg9S9OahUfY9RiO6M/G0W
iqpTwwXQvrsgkyKYlsbx5Z+E/2t91mLZe4McoUXspsgi7P5sOh8ccBaSwEpl04O7sWWJsspN/pP4
psqCkxuQc+itlSOPXSn9gDLgoEoe05ZhOcE28H+GtauL3LXsWsawl0KtpeOY3tkL0hwo5KXDuYPG
3ZYUqbD+ep+KPVmjZLuTSOIJSnXbQemwCIemGPXbZqDew5vnbUyd/VLD0miqknAwMaVBfhEjF4Sh
e/aDDAViaX9E83RYQauXTzRKBxyX8fn/S2UmWRhBwLbR+WLVLqZ3Ij6+D9WV9VNFKrr6NQme/i1A
kSRpmjwHKryGFMk2xZr6Vb4IPi0FOmfnivdQrnjA7kESs8IA/3IFHrujbTlFxpn2SFIHN6mBkBCC
22Wp9NSsY6yf1se+FPot62HsA/HRJZYUcL6QK6bLSIuAukQiDBwMe78oc4hRQlXKL/MBej833uW7
IWrkg3l7snflZeIhoiFB49NhW2vA4rsb6IROJBNU46Ux5gdVvQOdr72G1WYHj06rVWKJxrhnh+Qr
QTc4vluv4vgQfVV1NtBc1an+b6XLgoOJ/AlOnZyS4aimAJdFW4i5WRRs2d3EBu/N3ObeLmpt1lJ/
0dl6Aj1uCGM30CJ8UVurYcDbFRF3OZ9I5y9lz4hQHst/HOsjihVFmii9aUsI2W4UldXz1u9ETEog
AXVVcsgq5LyndTJ9X+ZpLVQPC3sOThqIk07bcjYXPcKWss2STp6g3JNOTrepSDkvLP2JMhPDTVnB
/ePa8wYQiW78qYiBb1PsIeOGU3BWgqxFzffBnjC5BtL48jO+kC/bzFjAMxTlmRJzqcSoDNAdtG5/
mEEz+TKm7VQN7wrVybg/am9nKux9X+ES8CLZHCiB9Vo7+xrDhonWo9FgO8kOLNY4EJRgocfWJiGa
XYI7mEgZDYw1FIDm8vs+kMJpW5/3EeRVtqcW4q/E/pnPSBYj6H+lmqHQzCnLhF510Q56ZTnGWTis
F7gwkkUUhNiOPt9H8Pd7P82yfiOpZQtqRszv9QUSL7QkefJREhY7eZj7GoI7bE1D4A7U189t494N
li7P6F25Zcdm5Duy0STtvRZXNI2R+L6CkSDP6v29ijmiQ2Nr5H3Ov1ncoJni7HJog8R72ZWx6r+a
ef651aNJhlHhobjKad0nJ25+KurxEXpXow9Jy3euhcTA1rlNFlgfqrHAPq7hUxB77w+g354dv3cQ
1j7LsMDI7Isb9XwpzhUH5HStsbpwQDTdRyJLgzVM+HQYrC6Q0dOY1GimwwVB2Wy2Gg1VUIkn5F9R
jbGH3tWBPugLe0Ec//F+oY/IIpGQH+drp/1ZfPzbaXViOrOHfsM9P2H3YpLeaiheAmnvixeeaVdv
LoRZEl91/caWNoU96zgydkymR1uaFkNGtUl9BNEzCUk+8AkWKckZavJpVoDs2/BBJGPL3qMqX8G1
Bvdrj/PA9J8b767k9no9yx2XzCrOwMUWOC6HSOZZRtO7wVsWXUeZXcZwApK24KhWzi6Y3AtfITSR
40MaGd4rgkX8PFS7PPPsjPvroXlnvtInr7ljW5xpOAwwJo9mwrIs3PRfr1CeP1ExVsXBkhPzezso
rwQ1qqPTupr3v66cAgRCMrQdUtnztgvXcepsbAVqD9Oi2GoAxF5bw8pAUG2eB9D0sWPv1GNhe6Oz
cQ2S3rEpb41f8tMVmGiZ5Gy3BzCWPk+70q/+uj8E2t1/PjE4k+x011KNApsWvaRy/U5D2ZDdDGCJ
p/BeL42YWXh7+FrR2+78AtEawT9Z0ieZC0JCs9yhL09qz9FowY3ebN/NTej+k2/jWKIAYDJH9KVD
SwQF60DD/F0XSXZgP/oZ5phtk6ZUhzDURPKw53JAU08EHbHjKmMBSZTfV6Et+vXYCQ3Z2e4rQCn/
iFnLDo1B+EdnwWWeJhzuS/H07YuixZHqhyN7arbBxr6bmfJQWiUW+yD11eRyDWfNMVpULUv9Dnzd
M2WssmBUAbdYWD5A6/hK80brgFz38Gvooi4pweCP6kleph9MULP2NOlE4d+8yqKufwIf96RddCN8
1Lyfq0NlAyA0ru5BahQynBv7XQra4UnO3CyR+rA1PKIz0sU3QcvqJMnxCWscNKFVFO7EgvkjjK4K
5cvN6sSfQDRhtsHrR9Kkulq8b+7XzZoDtHOXJTWfOJo8kbpmSjOaNoLNitd1owBp/iIq1sqJ435L
QV42UydfIhR5hG38erjyx5tdT86b1ald0vG5m5IVrdrzI5cYmR/asgl5LnotJom6SGSEKVZyvcgR
m9L2hhVEUI+fKrMadzrRheq4kntwhq8gapBundz52NyqKy8e6myzyNwgq0jvOlHI67j0LEWDnMva
W8tzrZEGCCytcfKibgZIWBOEFGVU9SdiX3/MyZpguwUqMjcm16pw4DqTLNmJTOKoDdoYkPqnoM5X
7OrG1eYF28jy39yRQ+K/Nc2XjdEXcp/y2kFXjARYHB9esIvCezzsrh8rdNLPEseCSih66Yboh6f4
khtm3G6hptjHjBy1qRr9ijj5Xi+YFWyhlZn6Tpv1zqBbvo69wzE4lTruBp3RHb6EaLlJhxCVhS/+
Un+IVAAytj77w5tCeZgWNz8a3P1MTFsJD5TklduHydu/NOYSj8DYGRhboc2V6+kPdvHX3ItAG5dy
Wa3v4e5zzfB3PqB5NR2QAehsV7zJTlghJogbDgHQxvSCQ7ggnOB9gwbAcmpl+RugviYXk1vdGA98
Fwju62tMwtrxJQV48JKVb6JOfOjRAdeu96UQqXLl+Ow0CVv4KcewOPaM7IlJsejP3hCQx8IaLm7E
1ZDbcT29rdUzpLz6NZmST1kgtI6jf7pa9sPVAEapYTz1maDxbDyMBdPwRadV1qIkdGwkNXleDrgA
kbGWlohhIBDppcyYVwBAwzQZ2it8ioaGtcScESJJcm6ab/iiUqE4FfimI34y7Aw0UUPv+j86X49r
oMa6gbmrzi0SK2h5asO4FY2bPdy/m6MSLeu0xnteSvp+ENSbTXn8Ozqk4/RSZmBP8/0dTtWF5yze
OMP48wzepNwejNmlzYjD9WICiIr/eWDTRWK76cBK6XqTJY6JqQhSMlVPWQA4gTrNDOCF+bReJQgN
A0z1AoOLMCNTD9E/7ERdbSWrV5I2zNP5C1K2m0/Xz3ZPuIfcFdcG+rIJSQjCz7Q8bVspDWHcURHJ
E95UA0oIeMGAXfwZi3+645VlSMuZA/rqnDtPUPb6+dxkhYHr//V0bG9eqz7X772c/yDqcmDPuCPc
juvesfTKqWduX0kGFi6eS4/zJKzDBbhcgI+LQTsrye9UMfeHkhvgpX5ik3toAbiBahuooWEekrUZ
SyYASd0u+UpwwQXi0dp76z2S6gkpw/a7/u8ivEX3eQmer/YzTeG+w3ypfL23vPD+reAkdfMyqwT3
r78uqjSclWSuBA4DeLreh7Uo1WPZgwiFiC0vgnigCnZ666341YGTbaSc/EP+9PZmyJ2TIQGAtSZg
71B++A3zfWNCIv527VKHs+8CUJfoTtdSokXgTEAqFKO3Th1YqExQ9/5HY70i40IzaNi5yZAdP3QE
EGuieBZEH1Agztm2Nb+X5U4K5gBnqDK6Z0vQ160MHenKP/MXmysIVhPHObYFbHD1Ud7MMt65LdQQ
obiWNbK2Psyppza+tEdlrLX0bj4sKLGADV2GGKni7QkE4BdqJYWsw/YK6pK0PfHsfsZZzVP0hxp1
SQP3WirTb7+FQZOwjGL8uZMEtk/pHF82N3PLqodlKPaquqALiFn78EWahQq3kYEUKg2MgUn6P0Sg
yCGqhlDq+02mINTEZinzB9DmARrzx3zMDcoVAcN7JED/DnbztnBEW3vPyoFzONrOXfWsYESxkMZ8
g2uOGiIWcIMSMZ6xmRDNjidzsYnN43CLU4qFwBAAYsrRtboPB/GVYNN7ZmXbHxzwiCkna8hADPG2
kNzydiZbZ5BqOPyg3dxCWTjjx3W9l94q2tX/kAuvCokSjBxHYI19nPG5F/vspaObCArcxk48uqeX
Ba/tUXzLsHJaUvPc94AhzYhcG6fW8fM/lossmnPzIvmbKa5Cd9JWbHXv7DCQzAb5RTbPH3Wq6HyT
OmuBRrQZwaxeB1qevOCLdGIE7zp0R0irOBBwKBf5HpZXeFO+u33a1P+2jT9mapZU/rX6jgx8Kb1F
7/g48LVjpzqhec04mDjwLq0oxCTZkcierDJ11NUv07bdME80aTSYiYfimZDzEQg/9NcEWdRwTj64
aDIBlUvGaLqH3nx9UBVv5+F5eVVqX5E1l3ICS7PohPDcwjg1a6zvjB/hUOeNHD6KqmkRktbRUa/1
w+kQzlrA6GufMy95eWnZfOCyJxCIcw60lPkQNjGgezBBERIPyN8D+qEsuQto7DFhqw9QODZpOEK+
gEiBMLswoZP1VB2KLXIOwd3m296mzm/BqOeQujgU5uf6Qt0rb1hZzIiXDlYFNnOYVxOoUrGGyLcD
yV2jpeUfd7JndOya+k7/ITh+AaocTII0DV66+d2c//56RwNstMa/yrJ9T8AFJyv0gjJ7MK+Ukb+P
4he3dSzviQzMc80m9ZLSRR13D9XpEzuMp/fEMlYiIXiP0C8uayhC/lRvpqc2mcJBaZ2eWtvLY5/3
b7ALVUe+9uerMyQnejVXmAoJFtHMleBnsnoX5MXE9qWDFa88skzi88YDO2P90tMhpYg8R+ARx0NT
UoClF0hIvfEBiHrpOhvihkvbZLeh7DgGkS732Xw5o2ZL58K/ZhAEFFwFZahQnwglMxNo6IQX03Tb
XFpNTo5GgpvCVX67u1XCiPKS+Zc+1LWuLNFlqf/W+hcg71iVA3P5eHqcNHXAnIkTLVDVMprY0PcR
TWr182UUcltpdoUsLzSds3YWVlVRlrx3i8KyMj5J0Ii+6K2wf8UzaTuCobXGp73o1pcOig1zcTvw
gbggZzTtUPQXBh53iPoLwi91ruK6msspVE3AsD4jtNj3wyws+gGX3TC7YOE7dfg2I1zboEFOpZCb
cj5YrdMigtsCfKZCVSv5ZLeDskoI6MYMvzWHWXRJ9sKo4YInc7voUa1KGK0oYXy4LXaY0ekHotyZ
nJgz7QPIUfYOnlDil5HqL/dNMLCk3vefB0rwKZEO6q8ZCOMOkubedhhhx7/nYLQPqXj857bGPYMv
e6HK1BRgJRw64lePu+MG5ap+hcYAoFzncRuw1cofdSv6kPCEVcDC+DKNPtagVU+lFBX2HCWeIRrA
j/+9R1LxPD4/3tIxfVcYN40vVhWXJubETjAN5x2SdlMQcbSjvvK6XEcs/+k91l3oRAARbXY1D19U
+EJajEjWoZfdbsoBAye8OEGNQdu0Vgw+iqMopYMtY2MwHac4N5n5d52qOCJbtygHyApIvobyW1/X
affKivz3nvYXcmlI0INwUu5Mgy5I9Ddx5JbfgiMBF+ltxZqNhWxGMbyWXCpVOfCx4iuv6D7Gr/oZ
7/EA6zmDu7pQ1RJfkFAHswklKq8AjlgEB4rASE2ygaOWj8wXWgvziqWJRg2kxei2fel5FY+FIQFq
/LAE1d8JE7hjntXUG6tx7yb4IRCV6woz9xSnh9x898iZsUsmCznp5Ou7UVuyRjHweHuJhS2Oz2Zp
14V3Q4YJJCwKpYdKeF5wDFBtKQ5cJGklZ7fflRrVLKi2BdCT6kwb9vJr36kuqjZtzjn4JTmxrfiF
MQbGGkCb4fAyC4W7oC00YJjeQ90fLzfVq+5jCFz9cN9geQ7P7ig7KFkLwoj2OcoQ9g4PbxfGkgS/
NwiBjnnn+0jzMjPyYuneYlZ/wt0WG8tVReY19M8vRU38osBJyzAtMPuWneZtLkMI9BPe9QEjXMy4
IHvMKV931qx+GUhAjy64o1PJ7ckqycNsXYV0xS/q63M+nHw0IeSB6fuXC2vQq7zYRchjm++efKmY
Y1y0zoegB73/eGcZmTpyCGCT/0j4TkyPZ5QXNg77DA+NypDh/eSdPoFiFGV+1i0sahLSOp9P1iDK
3gj42iEjOvOIzvKILWAXbd2uhEPDu25FL5STC8tGptv7o5rKhXWZlwigAbLtt0/Wd+jOlzgRP3gT
qDHC5bgxZ4bqM8fgeCbPGdqklEeJ27YQQ7c0NJN6/yYzm3/J0HTETarBwBy2IuDvnCAHPrhwaenc
r5ZRrSrASF35Slt1qHWENWZo1qO0Fw2hQ8TSbzfVwRQi36Z1M2tYajX256a3pcR5H5JygyETeISd
Pnqq0IFXNMCekWqAmIm6XPT9Tc+pzVJALcvFsWt8ZEq9zSEvNAaFknXRnWky6JZn7TEe91/Qvqfn
37pa5L8n4IlBiK0YULfjEp+PDVQ4UecDkhCrs6/DuantLGa2ohDDucPuPPJYRi3qF/oWlcNAd9Wq
konGS6ShvDOu3m8Rms8jTiUQUnLzUf5OSaMxSOk3a/zgEzFCbuVOm2kCQmqkA4IKyPOFfHBWJY4n
R0gvQoXy1LUrSmuGyhabLNdq8ZgoYo5EjrdQHvdQZkeE7Bo9eUPVGW1zUbaBC9/9D/S5r6BbmlxN
j9kKmXhkvLhORty3iQdPc1HYeegL6VC3vLynUPgR1r+A4QGiurpeaks/nCwQif+ia4h+LyQdK7qn
1HuzA6rr7jzpiyxOuH9MArq8jydz/0vXVKyW96gVb1wCZW98A5vFa/ZDuLcYoe2y4G3pFZfPSolE
Wqe5qCC3wiKupECNfYH/Ud/SpGvMXmghha79roQD9rrJLwld7Sgn0cVwYyjcTd4LhWrO0eouWy1Z
xjpUdqolgDCU0+hBTvGtwbXe7gX+vWOVL2sNea6yy5HcBDO+fOou3sNFNVLzpsHgGMR7VywWG/pE
FYf3156TDC69QOTuZ2n6IWVcrCWZWlOkRqQ1WnX5QphL3oWru9drebZJxSgMoOWQUtsghTNTLrao
M4zE5r2UR2PxKWH3UmoKx30CqgNFEzOuFXiCZfRSHE0Vn3mrQnIorrER7RKBSKdup3mMuqzxIdas
mGYF5+JD8Pd/Kua6/7sa4+ctA6yAVNqz/0RdlcHVsKSzFKNiLBB6fxQN9vTZr9FKrF0dpq9hLdfP
aum2mqNAyHj35t4IsUSVVgYdVSdP98h/rmWiGloBETAOIA6acH7Td6+zzQThSzJBBZJNWJ7WiHOV
lXiTYaTE+y7QqbsmJPLLXot5A1EUh6VMw63xBCNrW3QnnjbdnhM1q7TsVTAvDbYqAzHjQ0XVtJBQ
esJ/xuClIUG7KZdkNjEI0K31LTq8JSQbBzOAt0ariEEOfbjRhNTiPoQ9vCUKTu9zlxp1H/FFDKN6
6SchAOBmVlgpLJ9986DJLXdgZrhfaITNx0IvUXBIEATSRU5wu+BshelvRjI3r5vQ5sG+6CIZ8+05
8gWDEIhP8V2H0Qb4rV3RYQCGL0Ca226SSvpmvBbwmJFIbrWUThtmJQf1WFpzd5MBOaeD/foW4B9i
BzT+2P6E7Pwb9wOnhv4vmNATgqikkUNgweMyQdFHVhcL0QyCwIPRl2HxX4O4oHm7GUFpIzSHU72x
a70dDvv7kAk5iI4l1EWcRlDoJQy8RuQDH24riuycZT0cytWYf8E1SsaUTbpZFhRPeP2xhkCj6HMs
zwkdq6/UG7we05rVN19UY3Z1i6nI8kR4LdbdWBXXjRznYLSfUrys8fs7RWlzimqL4bSBKMM7UbyQ
d0TcdxXerPrjZHR3XqJpt/ZUoLUbEYzhbvQhbvz05xfzRFur00GWUg/CLmIsSCgbWtAMIwmbB34q
h/VRCjqYh6PWKckKIVcwd7Ya5PIkxSWhQBOZ5cVf4m7rFQ8Pq2xLTWU7Ru9WqU9PDo+3x4/tw+h/
KacGMy60zKBYx+DwlBossVcD50UB6Ca29NopvrxKx1VsVcmedmKac+HdRuyVF8L+LTyNVPHJ0Z7r
om0SxTiHzSAy9ck0NKdYmdcofehJEgqazHogHNI2D9N7ga+JnNTth+UryoPPGCLfZGOptyShox4F
X2F2iSFgLmDBX+TWS6HicaQ6pmvMoXpVbpYY2lujLQQYvKGA48NDvJVWfagarXgZ/kZCFZ0uSHvE
GLH5thd3bQAtkiVe5AEBmBSBMstllaMz71GoddFpyQGj4PSqzUyQw8cbV4FtCjXxuocWM9Z4RMYB
mGutbYqLzy9kHQkO5nFWwehjNH4SGbHM6vRnV3aGHToEVKk+xtX2nCtK1bKlutTk9jMz+1uiFXfX
jFGnQ7JhkUHAr/n3YZz5LgDCzVNbwCVvbSSiVAKcm9hI6cwC7lPljx6raGW+ZdJGW1HQyAQGfQle
rpeoVblA3F0vanHxAIOOjHA7ckFsniUN4ZDQujLi04nQDvcjy2mdjHmKI7CL6FtpArsxuuktO5B/
vghNjOgex61qU2ZMkF46P3yV7L30DrfyMizHwLi9AbOG2UA6uZn8fs1UG6ZWekXetmhX5jbOtxR7
1xb2ZW9tutTuiXp1m/VHUEHTsHlKGSKVzFDh5v421uBq4K0tHDGBetyNEIUeIV/Qi743G6sHHP0O
DFyAJeUjqGIDy1ljTAz4ApYyUvw99rDhIjNikwfQUEOTOy1zgU6K65n3MO63yQCY6YS1IiPjNhSp
kRzLVoAncsVfLu6Z+ChXZKvsNW9Pkv76T4yTiFZYwsgF3hgwSwEv/Nep6ljwNS+wNhhV3jIzn20o
u0fqt0v1QAm1aP9y/6cKIb78wqGVBPVDpVg0+uqxby8/e+FbBWYYQKUsSG83RmqAWqi+ToLUBgLj
b92Sv3W30S8OyPlK41dHP3uTOwl+hDiGU55ISHwxdAwHff2fmcZgd8DDN5cihIq70Sg79iK/ZL1t
Ed8VMG1XkVFPYlQA+TXWX3gpTA3fn8KmBSS5a74Wx6ZLRUAPridpKBRB6HSVVeY2d5+GmxjPQESZ
KJEZ7xOAsBojWKGVfopv/4tgctnM6mSY9O1qRsLAHe4OX/VNExpHv1N/AZh4xretag6akSa8pI6s
J4pdHBEpwJrNptkrl/SxmPUJksIxwTH6s4Xaecg6Gf+EuerAgrBMf0gC31QCjBQuPqgDDy3hvzxh
28dVudsZGkgg/SxaXxX2hl4OK4XHlQfjXppmPFfaqVLStv7lkXcbfxY6WQ+CQIRQk3XagFjI0g/F
Fo7fJ7M91zsoqSsMX4nBJjXlN2x2ItcnO5CjZJCJJPO5uMug8hc5Q70mSxcT7OX47NADOEHV8H3u
2Zfn647xHecEpYF38qGF88oyOjgQH+Ipdar9ikj92oQFPmGY2sJgfL5h1QFQDS4GtNTaQnYTcNkt
O7JDEySeu+goFIfRxElmAPbSGg1bKy0dfKZ54CEmibY90wyNYVPW4sPsYuc/uOV29fN2W2/vmx0Z
0j3er8BF2DQoI68k5ddtOz8xp7tsylNMMwjw9GBN1dkcfUSge1+SWdxUIYwVdwKNF5cdJvnGS61P
ghTls7nZsVPGkDdcqRcwMd882cg3XWp9cC0r+M/uF2CZDYN9hHTuyDOcy1DOi/7jKhs2wiGvG9su
c3EAUTR0JQaE0WZBh2uQIJ5sFNxVFNQJcYMre3mMKWEL3m/5HcBLzcm4MKoIlMGZxEvF96j3NLPO
MXUZDZ+GnZGy9p5RECYcNBj7Z+TAbT17xPebNkOIRYQb7kLEQL1Po+Vc1KzNJlgGLpnmAkt33rN4
UHoGp6ENRyp9hCGjq4TLG5l3e12J4HaFNdxmC5qUjIfnUsUTWdtyBiX5Sri/ONMEzKXUyvQb3kkx
8/Ty5w7nLqUX79gw3zt+/DqHSMAPrvt0NqVxdCAx7kr/cA1JzeM8S/qYlczD+EW2cJGgBJ8hk3zT
zu3i/lqIRN0/BD/Vaex4TVk3vbZiO8mY0fS0sb7Oc640aVJwPOqoBRPafcMn7i6vOS33l39uE0gx
7IQ0zSBgJva6JtJmmexI2mhS+VJu2w8+0ELj3FLcUHraSYLsmP3GXrbKagLrgGiF0zRwKuvUt/yu
VPxjVmxZAovVVdpcc82QQOiPgln1DYtHhVjWHuU+sWzR9JEEUKShGW3UZm2ifOdz/32U82GEYmuF
q5t80UthopVW0OFR3oTMVcJG8cGj6JQfhmk1HxxFOB5Tep/wsiTaS/7Lvc9oDnVHkfI4I07MuxGB
ADRQQEvhm88CKb8T9N9KkY4JkAJUTDdUvivNYrAZwvbgtFcTaVG+lbgYZL4xOgagVeSwvwRxnjTD
XULmYOmYuuKf04uOlH7DFEElS1Vk1n0tU7h+v/OLfcOJyrlcxzXbFboRhuY9LoN3q5HMrtyyjMoK
fytW3FpUhzUiF2z25EQpCAUwOGtSx9tiKRsruTCWIvVCVn+mAVr/So7vLmtsEqGrjd65IicgRvCQ
nV5xDKvE8LIrawimkCrsqnm7oBYYY3nq5t+VgXdY7DJQ2JPOI+eIVW+wwJOnSliwXmFaV4dgcRtx
22mdmTgCbC7cwkqFpEbQypM1W/wfYFvRK3hdF+XOLCOR2oaBj12nIo8JtCHnfdRyR/Buk6AmloqP
kYGBRRnoZKRxc/by7LWZY/lDTz4/duof7h+vkWVAlyUwB41VDPskqI2VJaznrgRPYJGftyypMcDs
brZ7MUjhDRF/lYZ8QAADDJOfjukIjDQJNEnkw79eglD+BX+jdndR5IvyqRp1bf2dipMG9toCckE0
0+prV12so4pnWYWGFsvfYgtybQ3CIQ/wyIdvxJueWzrSd5E8mzF2AeMOhlrVB5Mwf8BuTL+JuA8X
Y4fDQbUxdGKIXf6xB4mkUQsHPCWxUTwRve1mjziZnRpPLQ4F8TQpAEHK2C+TJ5LW1+Tenk6w7nff
arZzD2nys+eLg3xNWIFXu6Oc3rgKJv0eSp7xrzJEd+7BJLRSzotZ+6XahGiHYuZo8MxSjs/OjyWx
tqqxA0oKQUSLDT/2bI8o9sNUi96D8ge/0rtUN3vMfc/OXLM0+Xfqc4TFLBdEd3GwaWf/Bj7txX3s
rx+DvaM6KoH/ZUAqsGfP5CvmFROELFIWmdros9Dm8XlOy8btXvEHrg3iLIzwRoISsFrgpmNWuzT1
hXmfFFTE1gcmRIfHJJ6Phy94g3KUoEVNXQrOmHQjdofyZNlUNXaYX8HkUNHVCu4IFfBR7UFElJhh
/PFaBxAJVFhtIeFZBJkhIKD+XQxhxnLOvHmm4aqH2C70tuwEh2er108POGWhX5mHt8JSJBjVPjFo
NEkUuLXA6X8EdPOJS8ogZDV8MehD0XRPN47ACqjlGQEvJD10nueECqHu8U90N3DMpaYQkmDm+1Zh
2/1JYADEyR77UnzQwqk4RjPcyiE+f6AVappO3DBxIRdLrNw7MZM4kklxd3tKMnqewXJ0lzSPw4yR
UL8Dpy6OAJQ3VXt9HPosymO/v9pbe0E2KBslf4PncADL192ZTg0znfazxkXHR/RNOzj0mhPOrZyg
7Dr0q17DRphO/FaYWA7+3/9WAcoDG48yt7ev8GBQ81k9xs1IHH+3Wkg1ft73EjwORvVTjrooATc5
xKgp8ypgpUmedHMI1iAp7VCvJ7PRryl+KxLTDzbn9RnhyWaYmDzcsBpaaTPuXEsqzV+jYYLRtVfS
1csYsBCroShrD/fvJAuZEo2l4uDVCFswqO39V8tBRoYaKmLk0au9cCilz6Ifatet9mZiES7HyooQ
gt8+4R1VtnQ4Xl2+qiPsnqTYDd5gtM3Fo4ntt5gkA3YgL7+Hmx7sXO2cfRDgRynMxXsFZa6nTf/G
XxuESwEGyBLMCiZCBSxxsIQsxvT44ZyKPuXaWp9BKKTDFyipsV4i4mVe7AMPjAxK443/bHYAUlAJ
Rmd2KyIayPNr4cTJICPwslaZzSbsVtyOBUzsmRiME6/wieFXk1cq40JR9Zc2SC288FYlO94YrpV/
V6n7nur/ojBnKf/8C9fjZgKQAZTn4JsJf3qmOvxqICNp8ox7aBXCqQojSgJi9jtqgUtc9xGWU5pg
Ut4nRGQkWKUNNcD+6rL+WLenB5KjhLkFVEEemL/kDOeAc2ZwDPJzv9yUEuX6x8dy4nmgLaahRUe/
lBk2vKyBqKGJgnIVm9hfvwLBd7fEInppFrzYGNcNkDUpuMGI50+hGcz0GXlmw5hizy7cohsWZyQQ
e4Fj3jum2h2FvKw8dThTZzAhYCV0arXczpi0c6kOXKQg99da22kbuudSCsbh6YUg80cIhyqhZ4To
aCY+aHNZYCzYRoW3motFdbtLjP0fe4jNwlsQAgL2fXycoe0HhCGBq8IDCOy4082ZIy302yoNSVz5
GCjEv4vpRrLLEfMM8I77wXAfYCcXapYnktjuq7ah6UolthgcTduECAgUvAWerhgyyLs5UI949W4I
cP9THPP0M9w+wrE7qBjQjQvchMz6rhduCLT3WbmG5eKo7rJ/c4bkaiSe7GKrtY3rQMI/kmfXHpkB
vIraYFwnnoRnBZRYiogTIr2icf9CYsb3NvLLf9en2pUuHwdsdBxXA5AtkEdgbpkwDKuIbYT8yHXq
8fmN5yqLyd9dXU3tjyf9m0QApFeLiID8v8AFfrGQbDCw9R4970SFKTRTN5yLaxWw+ukI96f2Na6X
tTkosk4O5DMJBX+E6JmbRtsP+/eah1/dSHgHitcVaaBh2Ygk74YEQzz6jJzfm3e2IylDNi9O45+3
311BbJH5IWamh/M2Y7H/wQzQucxybFdDWLfbp/xzpjUoeTA5dGxCEzr/IsdwFdl5G4nhReSmy3UO
2BWWF+1IQnfeeuykFeBHRB9hHy3eQwHqEhfxtAFAUpopBe+ORexEQsTDJkopa0PNSwt3RWpAw3J0
wHeA/Lz5AewXrPQ0hhIZMWlkW8wW/ICZUJb5JgGOjLbLdDfXoGG/BcTJNnoJj2xs2m9XedXPzEBI
GP+nc2yGXp9Xfo4O8qms5GZNgqxcxnstgQK18luFDgQ3+0CQUsDnJo8bf/6IOjLoWvSfqf1HOv2P
9yW5uoIk0sRcsP2X32mCWczkWfRp/0aWWawtQCxkEYT6blNpDAER2VJzfJGLSVWtULhU+a/evoSP
mNSVBw+86XKYJgRHkeEiZmkZFCF+e9TlP/XRNydRQ2jsc+4u8K04kFWn8Y+op+UdTXymcyM4ojPy
WI3ZSQLXlDlbmE80oUZHgCH74+RoEozXWW4FUQ4QWNxR04UlfF8re8LdpjxtVTpv3ykdV5Kw18Uf
OlRiQmiLHxNa9FLtglIiWuFQzM443ph/wWqTF8VorHo4tRvIDpCpNqjteWZ71Ikx6FZGAwJF3yJa
6NLibSbrli1dJ9Gy+9zylfy1vjgFQs900WJmytq29DpKXPk3REDJr7dmH+7PsScmBGlUAIe6i1y5
aD3iZ/7+awSx8FuYAyEpoughuweCYj+m56vcvr3wZb/40j6nqHaaY9XZHfUNgJWHR5ctT9Nrtksg
rN3hU5O6AVZaVapvwuoZj/HWrqcuw4C7WRJCr5+5S6r8KmVZ94sEPWihTWyMxzhA2LBiRJwf4VkN
BCcHJwd8OLvlVo6kVe025Hu2wLev76jCA0C5zWMpCRfxtt1AcsVwKWaoNRfdKyaZOr5j0ycXFeS4
sWBy9+gfgzaaq8ePlbscISi61eYdKJ1K8n6HR3Wxy54KUzd/NzgDxOceyC6UAOUaxuGK865rDCv9
n8RseQFuez+jGVkhXWYAaF6AdDXRGb0yp+9nCHc4XCh/jrwxCdg1DolCOjsFYM2kJUGc2OZ5QbD/
V/o8H2R5Z+Tct190BKIeicoEiMuGsfwKIsFttdqOsHPX+NYa25CYNK56dzhdorUBGS/qw3ID37YA
DSkLLnV92C+C6IFcswCwWtiYE7wPtMlq1PplGDO2oX1H1HF2nwDpa2+iJa8vjQIqND5ykQ/SJNFt
CMUCfGjDRs/PWmJdbN0nzyuMftIdjWNDoDYqYroUO/fKjQiYsm6/H2R1LdjDEtJCKotZxenfLbVZ
Bhn7rV45CpSLvX45wPmqcjNFrvif7jdijJLZ1n6bLKwJwdYH2WdXbmkIyYqV48BXJfejjFYvMgDT
XIrMh/AC4F0gDRC9rHDiukhUnkMTtMyTbTTINBhORQbR/eMOsU9h0o9no/jYLVbJm3nOWRLXEEyl
upVX4u8Q20rs+OuEyQM/NVff9eWFRtj8Oa9XoF88hFrRP0AtvP7kgBZuHg6THUBdnPn74BS+y6pE
aE4Z3wo3Y5ASfi/1UqWDH9zJlYt2Tg9FXRdPqUJHdpomc3Ttf0Mfmcyl0K1fBpf/oAapbFJ0nAe3
7/ZhjN07DWpm2oR1uAhD6kcmstVI7+Z6xvp72i4vRltggWBU3G0zZX7EoGSU8Ou3nbf98ZaEZwyj
2kQ/fGYdlViCB48GPrGDPzruEPYqrLmshkd1hs3XcEE3YGXwS68n+bZoeabtRr7wzVaUpN+tZrlp
wFdGAkIUf4i2hMVWKEr7ztNP5zFA1UtR7SZVbPDs/NZM3j3pBiS2fGEj3++2BYLsOfK5wEMI98Qo
ap5EUMK/47U7CP25XfiGYHZ+7kZgtSNQvV1SRAjzYBzWSve9bdBZMh13vUf6ygGpTClzpqSM/N2f
wKy97L4f14PjJqTA0D9KPxBKF4zR9JvBoPkJklcWGcwXevR1hZIO9xZBjwXFhj4eCW2sd6/Eb6l8
CfPoVSr0mDmaNvgCC9HPnzBNN8BDQ1BkDlYt69qbzelW/79gUMpV/8AX2kgaiYXqlM3beuLU2+u+
+s/iPGKwjUDBW0VDPkH5eaIpCLdHFlMCxE1tGhHf74WndnXdqrEHI++mCOb73YDHwsAu58UH0wFS
PzhdB2pIh9xesMPh6LbDGhPHzDrO/r5Bh8l0mCTLwQtTQULzoHINE35+bXSWmUM9/syoDYpjtjo9
M1ymTqxSVmfHtbQWBwoKH5OL+nrO4/4L9U2tVO8Z8YVJ8WQnPzNmiV9vfjiIUfCIO1kTtO75+Z70
L/QX+8FmBJN81nghP0kUGpveiFrYl4YISmOoRhUmTC7X3eKHzg1Ivsv9xDGTjEggM5KXkAmk5a4J
CBZV1b8ZNm6OSPqMKhqLKf0jNX0xRto//PZ/CQPvI5RXzSEaqdzDhG0uaMVKa92+OoQEyrEyzoOQ
4OOEjJAqHp4z56TzkKkvV3bt4tovnWmsiXuqaUUqhqIYE/AoCGOQDpe2Dcmt8YMplDRNohHB3xdb
orFbZtrMMFKXWUdbRvAqh8NWaAH58FPJ8O5bEvVoT3QzpuFae+9ccytNx9r4babOiDskHwt31Hmr
CCBMvHJ2xoAG2MkU+MQL02ELWYME0Q8EWiy1ekoT/bXotymDuktIFmnUrqkxVZPqgSayNZqURPng
EamB8tTywYDPDqP9WTgf3pVpbB7420rJxEUqSAFnDAdb47fF3+xBhzoZJza6wzlvYk9LUrqR32mo
BmlEA3i2h2VGsniIZarchBmUT0CvjUe9dzN/MgvStfLhprGtNWL25nH5AzopBjtOUKAOvPeM8QuI
8wyhoW5kcSowcivzDHMJA6wJxe9V8uxUlnJ/PV5qwgH2uqFRSCUIEGorzLZ7YW/aM/t8KU0Xd0Wr
zpzBl5oi6Yy2YBBcf88mL4IpAs/kTY4mL3WzKgiPsM9vv5EVwCT/A28WgWXkminO2gejOTCtUoZp
Pzu/Y88qm85956Le96yz8n2mk4F/NW2PkiLeCBL2eWqF5gThBWNTbkqI+5Ym0OYzeIoexSgcMku2
rVUoXo/CO+uGfmmLmXbVuCo6GNn17tnMIAp9tsrRnB6GYB+HNlCmCu0Iskxz5I0CGPMfShpWuEXm
VsxwOTvY81kRFeIiJEcgl9PZzKvseR/Jb8dTpy3bdqJ71k0Zi+esTGIwnzg9OOMkfaw/40UZoZ0A
0YMK7TZZ0M49ESjhUVbvD/hsmtwa2rKj7ETe9XgWJ1RRuu/JPH7FYgOq2On0QoHJid7IGPznTfEv
xd+GL8U2V0Xn7noDAwmRwOUXpnMTfkWVkNBh+fAhtLLvQ6bx9GtqQbNmcBJke409+xbHvmOfitJo
yziwSX6HXeOB/lEwYI+xDnPc7VRcP6XmAIHWRDNaxJxrK0S0JuLpr6i7cGQCNBSMCNfWfC+cjjxZ
9z/lYhMgtMBArFrnTlDB+inATS6JHRVEo7/LeXhTIyOepwFZaNmOep6mxUnIp1U0yUK4lksjLrIr
L394ekUXI8BdoBLofvwOF3MD21H7el7s7c0aLTF465zkBW9wFhA9nNqY7dJcap453lubGXi7A0ch
Azs22KTC4EqdcKJIrpYWqowD5asWFTGKa6hPaXFOd4i3UaLIhb4obCrp8mf7X/e19THeLZNFrb+2
X21cnbxb6cNVRKlss9Lhg9wAO57Y7TT1tr6cUSyV9uF5UYeAPwIHmRJ/dThp+rjE6e2Gu+cLeD9d
YERuYs4IMpGwPzeJIuM64I8uX2B/skW4vvnFO69EganByKKqZG6Nc465U2uUA4lWOHehw0asFzny
RWNmR5+REVo8c4W09vLzWRJ6oqovh/w/4hd/eklKo0rj6D/I7M1whfPhVzxnK4wk8XSZYveAhe35
8482FZlg0KJEpayrMYuULf3Wih6jGoN4tOqJZzmJAtNLKGXQ1rO1Gr8GkQfh0hNk6lBByvqjcgR6
LqehIWEL1N67f1bl0hAClRnlQ5FKBOod7sPJVjv9p+w9mRojdBbxe4GKtc6CcGtL99txI6D+GxFz
jJeJ/Gx99mKygfHfDdk5KkOM2r2+6ylcWgUFPNsfnl2UCUv89AmpFoBTQQP76y1tOuYoB8OookFY
xzKVl+4fvbeH7h19kjfJuRlANS6o76ELc3GF7uS+oozt7qRQarpPaUp8MJdpCnVqc6BB9hU1HPMT
hdcV94/dhw90iH79A7XhCpruQ31hyVCwDNTbNDDOugT1OJ16Hdd0fgC/2XxQXxO4qo8Prxtw4vVO
BigJmCmGjpVbd7DbNmSR+E+EMCk4K21l8MefeNypHqdrzllLCPlA71pTNT78fEZ3vbnJDKZGNcyg
R4KnqjSMHSk7s+ijWe0wIM/+fUGFp44Yp/YCoo9FTdBFkAcnckZk0SoQaEzyx7veAzGgbvSEFoq5
nY4OZAScULM7ME66yQr1P1Kziyk44pvjCDfZP0Ez77h2B7GimcyE2R40Ad5KmfQkOZauJZmcbM5j
+cahI6mLtwTEwinDu4dMLBaKtZvYUNJ43ONexFFnBzmd00KBNFnD5EEj39ojJMjsVa3IJDq6GMNV
qkoYQbaCkg6QIk0Uz9I00yRl0bSNeVstr+vLXhnmw5Mu8/zLXRBvDjnNAELwpUUnRMYoQHBSFwvK
z9WW7L526uEvI0/G1CtnnzjaSscJzDJr9kkbMcMm9ieRt2FmZ/ixJmmcYhN2zYJkn90oHUCy0+vY
ZeXGhirk5rKQh2L0cgldfaeqQuLt+u3DWRf8jxjRby0wbh6/QgEmL9yL/Q/uF/omm+ecbN8bJwem
HPFPtKEhpafbiok6QyJOE971YOfTD2bxUVIlUkTgWG7UGJbpvKvNn54ehZ46ftZW8ZFEUnlkfF3t
OFmMX/UsRLrhwa5zYLhFfDBGKyNDScFPW5EF4eeZMHL4CxLlLBB+OxRYRFJm+UmCxEZRMp6elMiP
jYRVH2t0qdFYXHDbjCHcVrv46zzj2LxL/sEhCfekNMuzcjkMqumpIW02nisweyGFeHE4GyrbdLdx
TsW0wg1SfIFY55zQolrkxT0Sq1Y4H9Db87a7vDFjCIbxiSiTqYpEihl7SR4hFTc2CCTTWjMGul/B
DeCa9Yq+WbFddAGi6JlFUOrlgy6bJkYxFEHHjnVEh109FC9YlGftzJnuAqEQy/mUii+2gsLuNo00
GJW1AlC7SEjmUskPjVGUUXlJKHfuXyRkpfGo9MmZ8sHuUaLR6umv7GugMCptDfBch3acHqTp2i1s
T0k99JTRHbG7ycQzbn4HqoH7/7TtTlI2OC3fMScrUQcekSyAm8tSSK4l2dnQmD18x5Id+0qaI96l
N+OHZ2LHIIlrQR4RV86LABmf1MNy6w6VaQQQXimL2YBk1IW7YAP4KtuKSVBEAprNF4Nz/lUWBpR8
4qrEtXaNkouG51JBuVhfDCPI9OBFm/2pG47tXRyReYg0nyPUnIUj6Y0YGAzS0gGtiopxoGzlJ4CA
mFLqCxU6ww8lUwhTkJMM8KFXxFNivTObvJ3sKAMd5FROEU2Zz06Jaoq1qzljTZA9HoafEiPvFUMg
kzZr5kf3m6FCrf4FFNz/9aPbcIMmUK5RE2IugbsehadCrUbWAatdRRDxsodvKIfBuynSR6lgns3x
MSMqkjXFJG6NLcX+WSQCaDSY6SFdhl20ktMl0ezpyxmtPdCcffEIlymfwMkAFgtDa4/tukv9tCL5
zZveZiPRXI5qGSSKcPfNFOJ6rpE0atFbo9GnF4I5F+KKQ12koPDFt99CTr82DVHpPfwtaR71wLxK
JoAJzzl1Q2fNZ9R28dsr0ZHpYSvWCFzMLm2G2xEAoezsVBPY4uNz/mgZd6ym49e6Zg+66neyUD0p
kMzI/h38tR3RaHrEz/ULOdyaYgqB38/9Sop2PVOYebUSDoqHTZWR6Z7PMIDq2Of7VhUXu4hyc44H
xxpjwNRfwxLoh2LCKnXK7rM7fkxzchzsHViGeh0TaYemERgAuVnQfl9FsCdWtuGV45TFz7Jwdft/
CyrZoIe57Uos6vrmxjPXSulZN8OG6JhyFk2749BETSzN9CO8nRPgQa1meogP3i0ZSvaCh6C6NHk9
nxcF4an+wkAjC3bSi0TnBoMQMo330pZGbsP8Z1Y6wNWhzE7OqzV6uFVZbQl+bLixmTEky5J9a03J
IFSASWqIvFVUJH7URa5QcSsUbbX35qnUveWG4a1ULHs7PrygEEDwDv154lNVKWp6IGM7JN85r997
oW5JeeV1A1EvZzKgqkg8DOyYVSuWFiC7y++a7+oeFJBpGpWAoA2JhrRxls+NoQrQyZEPSfJCHghT
25UW9SSRN2aDRZd5Y3wRAIMOUFZ0TUA4yM3GrBF0jle9IujB37bB/Cx6QHRW7BB0e3hY17z6zIk5
E+Gh0irm0lJdr0w3PBep5Q04Ol/tAYI7T8zVf7oB/f0MjQaaAIQaP2IVduRBKoT6ox8H2fRUICo2
KIoVDN02epM0D4SAgzd01cn4vx4YmLgZeBWhyJOq6+O6teD0E67D+8NBR2K9G5f6aqTxb3329UDf
1XbsaL/Q8CRyKl29FsJS7RvsFL58ZzkZ7PgaXRXftPbuZLCxW2JYQcGRkJheWGgUekPFPgw3RxXu
2giD3CHBrGZYRcdimlXlyv9FvPfXuq+c4A8oYod0+iM0lvS6VoQZnTRI0uVQK6t1yY4yjRdSAkSJ
c9AONtdQxYMojG6z8UFH5y/FkS+CE/y0Tbkc8K1RMYiaQFfVsZjiJ58On/SFJWpi+WpfHrihck6o
zj8vg6sNkNnNPdRLoDscEs+PtY5XHICH7u6NU6nuzMeM0iVG7AXWElYBF7+KgbPlUsNg6B4LHjHM
3SgQ9uaM54A3cA6QoNMHAlFYSCrYkBggMbj1TKYTm83SIrQ3+SxfJLa1U8+Myic/kxLKDc8whSiq
ym23yoHrIFuQQU2PvlOvDbm6nXNVugYJYoFEowR7DNbJEhvFit8QyyMcWgawGNripO6YSlIn5FmI
6c1RaTI/my+O/Gxx1AJIPhW3VsWiC+erY3y4/pLD9cQdBD6ZQgDz5AAkURgLBJCOgZT/A42yGfqD
+rtX8KdOaQeadNwtr/Ak0xixP0lOtLBNhyA7bHa7K+mBGF4GHj0KsCu0ZWDazlL4+pt8QGvLHM8b
NdoI48F6pWabROjJWa4g51RgkDuAKpom3KU0JOM2dG7mmnw97zRSaW/cMSL/CIrg3P4tXCxWCXtu
2+8zDES8o+KF2xKggI2HbHdT+dgCzlz54JnGE0fxK+4sW+ykkKp7st7m2PkO3fZ+KO88RYr80VBf
YdjZ4W2xQ+rQ9x/o5JIOmp4Wqhhg/wJUN0WjpXuvD+Hvn+OO/rZV2/HCQGk/DZjLrmjZo17Kn9sm
2Kf5N7aHb4VkQGAgJGmeB9WqFrZXKjDZzNp4Y3cMcBKDvCRjHiljqJr65mnTcSoMc7Fd5xro+xDF
30blUuGTuyMqHjfle0323+RcbcwCokF9XkcZSKaq9bsMARaKoYIaMOQpI8DE1j9NPGZW6DeEaImJ
2n4NROqxK9CUerXRL2mFz6jsOVdOm8L2TwKP6P2AG/ZrRFP1RITV4lACmWGkKcdF4eIer4HpVXWP
oUQPv3PBZqVD3ql+3lG59AXWoNqIiYKV5Adu+ZWSBXdr36KRNegrcVAJkHUFOqCmfjnnZRj1qerj
Ugq7fMy7zSmJrt7DkXhlLYIMwBefW9Y/7w9F+IiyLPptQYM+UFEFhpKWVw7qfaadSp+ikswP7018
Mz1aVRu0and51M2g8okGSapeSTZDVgDEb84GDjjv2sRr7QkY8gYFp60XA5+rE+D7tPmGIYzeCgtV
iB34SWRpYJuXx5aI/G6uli0vHya0D2HewtQn0czsgpvQflPI48uL2M/N88dozmk/2Pj50UAN4jEk
9en+kjAj+VvRt+7HinTYQgMifQTw2uWuYp0+jYsCTHhrR0KKlv//NKWgMKNiIxtpJXFSC3duUwqj
/EEx+EubrY+/zkwz4aPhE/2pSIPdyMTpsRzQBuCQvKJIxgaokNrSXHiohXLWj/eLb01mAhX84mNz
fszFuSwyb8QQAN4ynZl8g2u6ulnDvcveanLy0H8z4nwvWLrdUr1OvWLfy7lksibD88wfAiSYH5yu
XkV2XAIikNEE5EO35pWzOUAgBcUCozaHave4eWg2nLiZNJ+xorHSiqmo1ypJZNUxBII+6u8KZBWB
FKv+OurHsPNwv2sugf4VZHO7bdARLHEoCHFOvxs/zUdvzPyyA5PpZeTuvpBcy4Biy3QafPLQiC6R
9tmWlAyGIM+WJbgCDTFmyKb6seu92s1/64J7l7HJo8d0JvoCHXhD8Rf0KsGmqfOL5FcwlBcw+OVQ
FvTBPmCiFY7Xsbs0T6KjWmcbE3FN4eEts9y6tTbQRrUV9L961DjYoswmPJ5G+wC1i9pnARh9/umL
XIqSRFNf4Lhq3xulS3ZqKOB8CAErAEwWk40DCJFVhJemsy+n1c5HdGyWOl5GPJm7d+Wj0XDsT8PN
VqaUhYn+g5U3hnKt7yXp2F+2WbRvRyPkmlk6RwhpZLSvwHS7D0ZnB7C8o+6pNYNq5vTi6gmywR4f
bIfsfv0HSU/DSZSZPDRieWHu1lAv/1PPxDdqRSrKkRPHRsSoHg/HS/Szd7+2PovuyLsOfD4c1wxk
xIeoYnq71SfvD9iZVazmux5o/3eJ0ZUxXjqX5yHf6AhvTFiyHH+8NQFUqcyN018qynl9w/my31hG
qu44NsTr1QB+WzujuGC+886KcON6XmmXElimrv/9Acfwbv7cNSETc5e7TU/nC1pWCPZYyiw/zsBv
l3KSpCXWR3LpjGO7shZeR8pOMDWW4+bfLLFCAVpydiFiBGRSlayl+roI66q6CkI8oRoSOdU7mHcj
Qx7PuCVXaHCkzKrLn8/0Bov0+l6If6+Gr9jXWH3KNW46GrYdyVI2QbJ1UpVsPYzrhw0tx26WxyK7
7pPdlFIb26qmo6PPIh2BHg027N4+ntKp6woQAKwu/nYeqe0sNgvrOeEMmsG9gWMFdt+CPO3k3mx6
7EQvzPwDNII+EbuLq2/Bc5t3z8wi14/VIqiK/JCTFsZJA7An6Yu/zgldXY7G1TsvOmNiaKk7v8Ej
FnbIG8KNsRkW1PwF7qYzKtRa8rdrCBm1UCF4LBVOnHpf7sOX73wpJJy8Rwb5l9NdE+ALCjvIaVJb
YM5QGrAnMJv7XA3BbzHdvstV7qkKdqAgZlzfV5JSGV+N1mFXk/YG1e/yJn1dHSdWQjsPqcP/kSgv
zWABGKypYapvXPWU7hnqN9CkmoZKHvT5qwFP3vrP164ribseTverp++KDY95YmuzcTSw4eAooidG
slF+sKpCXJ3tigZeN0fEz2MV7eAoRQbWeEEjpSd48BcMvTF08G6dDT4eZ7Nq5HUBSCUM42fxI98+
megIebcRg/gx6KkAD+ZBSzygC2owBperhkS0FEoZfFJ0X5Z4laSwbxFAQdUJct134O+VYvN0vuWI
/Xy/w8Id++7gO/2pqFPpr8NnikQUkfhM4ieT6JzK+S2Flr3PRldmtUsWjCK7pvZ4QbbW53u5I6ja
Ro8GBOFI7cRgWHix1p1USsSUWl/qGRqpElWZikwHsIBgUKq/VsHNXMcD1SUn9nigYJP6OXazX5+o
jnrY/8DcwMGu38asA8PIXcoZceDMMcp1yKe+N7BWtSQFvE38/YDYC4Qjf4Py5KfsdGTYrrw+2/0h
Oo74FqNFSxoTSC5J021OfXogNdqag5SGocSWfBDGDiCTWzzZ/0oqFSEnarH7hqfhy5CwITHVseAs
BU5s8O7t83ME5tAWP/h341OnUwXPDTaGnOek323AdQeQKydEiBKzPqdNMnPAI+jvR/XQvCMf3B4K
mcNTvuGyc1oYsF8NgpZVWLR7k27t6btjrHjsVSe1lkY7omF//DcrGXai94iqg6QnFxLM0L+Gcxu2
AZ239o9Wti6U2+CUVVgC9UdRjo6WmnSRv4NV8Kh+VZyoIiPmtxJfQ9VQvUBLyNLyRl0ITMPy//HP
E6ZXzviBA28SCOSZDyU1J5JXFWeStNVqaHunO7+gIBv1cat/aez7+NQR4CDjwpSlJmQZ1vueV+4w
YYuOS3inNp1LC8Bf7bhANfbdmiCNKMCzdbCu/zJ6xB7KpkP0llWM2JZJ1m1zRf18L0x1A5JQMqlV
TJx/9HOv+QFA3Zy/n8sEelhLoFqAXD8wLmZTnZ/BFd1oIHeDU2kHfvtNZVw04TKMVl5YmXQkYfDv
KEGyeai1WZDmi/RLTsBjb0K/toX2N/MFWuCASruKkncWbI4gJzdvVX9cQcMjUzeopdz5hI26dC14
C17dPome22ooCEFGd3n9+YjOo193Bvu7Q2MODnAFb9beqIwKioAg9Q0fbodtCgiSiWoTd7qaGpYj
NwZ093mHhEQaYO3iStDCE2Obh7Zrs1OT3gxT+0Bq2BzYN7B/amR+DZNQZv+7cc/I3R5GO4MpTpEt
iAPMBDFPCwQQ1pLLNwN9qf8sEo1gVddgadFsYEjRq4PNAhuSoHsByphX0DwCHGJQ6Z164ul/pehS
AuP0iztZ+qfRKve0X2+pha5O5AGVOMKj1j+dzGbLU1W4cTNN+WwSl2J6fzqhL5VKR47l+6WLv0OQ
1ywqlTgM+5ir07tkQXzvi3IggXi5Q8b0t/YDOleuLdRIK7ZSxlmkRwG7O1A2XtpBCarPsHCGZlTL
wFF5Grmr9REgMypfko3kF0HKdCCTNVHxqWmTk/O42VvZkeQzyVgwKR0Y7BCwaCahY64pQiaI35bj
VTaBcXiHvZNEFecchoN4ZwlxvJdL4IFXU+40voVOWiOrkfhufSwOKwHi63kTh3ShVRR4Umi40SrV
rHfTetfS2lTMAHd38Z+4xG4Qv5XpkaETy3uerfLUfhE8AqU9D0xu//muKUP5A9SlyZRzW1NHlAFc
zS/5OumOvcRv51rSfp84U8w2ZsZzODyJipBAbBanUG2QGx5+c65GWX9vWADURx3+RICVrXeQgMBr
u8WxhBoswBQClbnmVXHzrj39MGpiqvP4S1kI3jqYJ+7NAKX2+hfHaoaiq8/aQacz6OWh6xnIwBk4
08M0OQ4ollLjHb/ymVoJvrE+niajdDD0hXB7Smgd0iU2FR4sV4ySuAz9uJfbySb5wsZ6vys7B18A
pjGkEaRIDP9VL4haS7Ed0/WsdEsoZv/2dilxac9dUEPanFndhgx/RjYz2B/ItvIhxnpoEL2oLZ0S
rSm9PiuH0ln14q6Cu6gQnSsnOjJ4K0nrIRtfz+X7FqoTZ7Vd8dpCAq2H5gHS9xjBXaE9YenWihd9
/nAlfErJgP+vIMgUuMf0SPIEnnT/9SLlZdseNso9zOIhUYf4mMGlhvRDHVsPTqIkauHeeyD0AthQ
TPz/p4TkqATyMhhsG5xZ2rP7Pk4QPC4VnMXfyUwq0YYVkxX6080gugIOoLYP33R6km15vXXfV5XC
O0xt5OvIgu0mpJZJsi+JaFzmBE5vxAZ2Vt8Iv1yp01zUXYbtKXh8BFdDqlVUTI+UiXnmClfLt+Pl
Ng56a+/E0jp7HAVBxd5TXOXexEelC5jBfd4r9B8AqqMpaAESm1lrGWKqRT+6VgRP0+ZKNxEPw73V
YTDb8wPXT09tF/oqG9m5P54i7Nvyeyk/1ds8W5VBgNzK57kM/jfdr4r/7Y5NrU9ShyygDaUcvhgg
7qHsYH1IICKOMLdNs1OkoGZ3C19Thl4zQ5WtTdCgLBA2S+8bSMcj+fTSGwCtSQ8DzuTpBXubIfv+
GNFOQ6M7QOka7my3S4MYE+SCDnq1LyoIclVbLwlMI+afIUBhS3fh4mGqHrwR5alQZoJXfAR3Ab+H
OTLAdRehoQQjiZIL8HHt/M+LNpc7zyMyVN3TEeif24P5vxbeBpdNOBgmcwVgObDlo4a3jex9DLqB
Qs9yk6Ld/13/0sUgQpEr5yW61lJspDFxg8KsgIiKTaQqEOQtYOL1DFnMHwW3cIhQDZsE+cN1HAiP
9S9xB2cW49JFEkymLA1SCJKPFeYCLjme51T5r/KSQb4dqCF67LlAPhsMhozv/ZeloLWYfzjJuFM0
18RfaLD78NsjrnVFJ7k0+zqNF2q9xad9P+WzhMY3xvIrmTcCVPNS6+1QXo/VHFzyGQpyb7IHPKI6
ZXM+UOYNPy8urwaQkdCJhqPONhAFHyGFAdKMw4Ol42jsZzipZUlGuPnXHA5KajfxaftFzNzTnmkM
JndYS0/cVG0ihZ3/RUEFNQF2Cvw+53CshkuFhdBqhfO9ES5mWSruN32qYq+etHphJe8OJmxXZBFa
XVwuENSE34LQBS5R9BUck6MCBm0z02ZKcM2CXFtaHa7NUsLp63YP8am1mL/WoLAw+apDFLv2zs3F
wE7Ahg0Tpq3N6eSOmy8ODML7L1P9+Z8B/uX8gYfN76crlkgZ8bNT01of+wr4VILZYP4mLiZUGJdd
gARGG4haH13VilC1EfEp+u8p3lOZIKufHHm9+bepps7XC28mDt5wBtOxb5i4679rWLymO/uBYcKQ
bhvg9xvSr5br/hohhJwX4DfxvNPc7cW0jDoNn/5eJ3SaIbC0jjoVsE6rKXmilbv44CqjFijRkGVk
Z78vGtXGeWs+8aQqUcPa0HTmxOmxGnq+XarOwtikCQJxP1W3UY8SEZddJ5RU/VYGHAMG9/dXygTa
Z78mlIzxUUTLClZEptM6T/9hK69oYmqp+t3DhSsEeoGkr7BkuSgdJq9OwaDNafTIS2gSaUDPNJeo
EQYYWFewKmBXyNfnwlhg2dsOrMzKKIDz/nMP2xnv6tznO+A/RjTTiEb/galAHx4BTfLCEErUdpre
lLWd88TqYKooW68WKZdtEuQ+ieAqXWSPhkyJJRvT/v5IlQy5NfLDAj12hHhDatvG1iuDXFJ4bDOd
aJ7b0NOVip5+gpdaGQjnNRmUc3/yyMhnV5UfuWAtG4ylNwsvhSaOAHDtXiOAE9HN6D4YMTy0doFW
qoFax2H/XyU34Aa+nNh9ub4cHYayqoF2UWi+eb6CnjQGl1i+90umjZzMQXm2d0C67QHbkGXJFM3R
NziV3Qy4B5w6TfLpQJUOcxdFyIOUFwdp9XdLntSNa0omnkZgt8oMf2uP4XN5ZrpGppjXyvqqPlUj
rgxh7SI+81xWei6KA4Eo8MUyPsDbeWjKCNMbosHkU1nsYrtMV8IXvwYlNXt6Kd9j3gjj0+bpsgor
BCMVlVAYkgoZnCUrjJIm9GRxxbNhwaBfE9+5Ws4bbmyC5JjJ+YY4YsaJYWc2mgCWHiMUhs9NaA35
vCosQbFgKSY/1wRS9A/5kcSwN3ODMgRjzQFz5glrdNSfM1yZ+5Dmxab0r5aYpyVjn9oGRfeCeemt
V/Ju8pt875hxjWKiTTpLCOy3CfdWRkx50Ud1/Lixz0hPqMebCfs8iBMzpdTyFaD7KQWbYbJWxLgR
lC6xC3FiKFROMIjRh1QGkqjcFom89d1qLjnlgYPkCvZ9gVOdQFE2v9OG+OR0h/aaWKdPlXA+qlaR
SkoGWPJTUmQOM0M2Bto0H0G9mVqfOxhd+XPtDNljT9RxsZS9aT8Aht9YePmDbY9mt1ysGyhMV4H+
Cdr6WJqHgbRIyyTTuB3rKxYGB5cue7EHB5C96Lm2Y8aq9DGflScjo/9Cp2E4SD+pGCCtgwCyd5mD
RCrqjBT0ooGaqwbViHFroAnO+mGb1YsRxiXgyr5y8SJYulmfDIpUzmTwOxf0WT1jw+x++95nt/p6
1Q13ETKQNrQidS5933jRG3FHuiUZJ9emfVEnIvSX6lQACf9SOo4DEsD2/tzDcQCvf+brv+wp2kpp
jNuEHZsz2cNgaYk0uQECIY68fEjyFylOKdIg1mBldS4BCuyCqp4mUdaIoSKVd/nddCvYUsEYoZjv
7HNQ8sIF5aN/j9y0cJhErHL5mjgm4fX5P1hmD59WrnV4V0Aa/Ij7FVQUvi2G/puahuzc8bDV4yTZ
ogU5L1uw3q+Eiggd9Yu/MoA0VFZBAb1Sk+Nk50/SJ67H5r/Rz68yGLD1Q9lqq67/wwVwTwqfftqD
Y183Npo2zCcvHXMYjFQMyAXo99AEVkEwHHGegvBiJCp5oPQyCUr+4scKHupC7Vt4/IA3kmVAwjpB
Tizuc8wAfsBxCLIZt+QxhoAiDGqLh2R21NDvBr73Y5QL1ewZe7/mpEalzW8ZhJwWIYq6VC/Pb335
rUjOnSEwcV9nD/JVxxX9qbRyDtV/UD+E6hn2AZqINnbElHAFROYjDJnMq6F++acQ9SEY1RYOk7ah
t9LI2GFqTB6RzJ+dwpis4NP581bbH6LEJWTndMpTX2g5JiL8nVmWt3GUjvhs8XmEqhDwDTRDTYlp
bjedjWF8oBzfVxI8HY5+HXgtDNI0zAu15y1Eqf+0YgpngAmLTfYGH8kY7zvWCNWzmHY0NY0xAmqT
MH9Rqw/GhqiSzjmee+yUI9UYb6cySu6NAbLc5w5XOWnFEU+qLoXlSF8za6PAPRWJ83qRr6duruy4
IDtCe1rY9cDGWbbtGd5DXNwEF/q0Z12BHNgnhyefqlJHmS6shIUS+JWj3J94XnAt3NWX05z7Y13O
osG189zX/MC8ilYjnOpsSL1HpNXZU7ubaI/AAIrU6VOhZ3a6sfoGhe2zq9dw9WAToC8ccYuvsh3S
jE0Y5NtJC4TfKnTP2eZSN+cDP+AdVY/g1s89+r4uwN6jISBxaLs+Jf3s5pelYHS62IL8Cvh/GKHs
2ErujqYKNm0zbwjYxY+Yuv8cz6+ThgjDeSgQBMrm5RIpc3kl03TRC+4tmrf0Mf9rQhWByuR9Cikh
/Zy+yW7PS+I/soIvq8CHnVAfSx9XLeq0Km+4mr43165lGwgC6PI67dJ8x5fxbKNh1ZkIgvs2lGHn
vQrZbfvIlOyheHc1zUN931Z43RVZk5IF50pOBv4fWEi2871KvGACI/sUBhnX/oEebDDeSikmXZDv
aHj3eAOdEI5Ynp+OJfRSCNumIszRmrCNSMCQvUvWeWCbolwC016PfUHoMVy2WQXFgRuq9sFmFDhf
wLn8AS9lEmvVk7QeCEOALiriNWIYb7loFOtHqGp+QM1VR3B8S6TIsv/ozBzY6w/wvNhVJ0F3Q+tM
4ywZUXsGbaD/17/VGNzebM8K4HiU536n9UA/5iekO/zomTfHUXE1vLih1NqPiT55HYvp0qZVJSDe
5+T2sEfBOaXvwjRa36KojGOgJbCWJMWbLhWkS2Q/Ip4pDk+2VZq0BXTAnCF74/WlhfsVScOJzBVE
LSQvt3TGyNL7u4KdNSydPGaY0cGzC7KbGrEtaQ2X2JqxvM3xZ7pbiNh0/YWK13MaJ/2cBHa8PKJa
nvsiulxBOe8XCPMwVt+akJ7ajlBNcGIRSo9V922m+88G+EyXcg5lN/jIfM5Co58jfxdA2Kd/2qsr
zDL7EX85IG2AT0hzjUY02r2H1FCsm4JWOQP5Qpzt0mj5lrdd11CTjJ8ag6TIyCKwWamwIWN6KVJx
xfXn2JU5FfqWFcUGLU620dgHcqVjdytG935C2NuYOOVA6MFaEFoMK0GwWBPn+zA2wAhBEwYyqVIj
d7qKEBL5Ojdzo5VkT4zbinchExqrjNJdwxnPT+W03G6iwVpeHB6cMiTidqhRTR4hgGAEI7Oti1Ga
1TAA92aEhe1GVJdRUJixD8WYrxXiM1+zDSvJO7sfFCWjSS7I+plJyRa7TSNB0WQyLsT5qQRilkzf
9trIPnBj1gJufDNTTLzYElNmrBc/lIZenX6nP+qvmvstypAH2vpAIBkUybnIpwzEL4N4xrbSFRiC
nue02iWUdPa3NdTWtRf03CbKHvXPss+UN0v4qdpkawrS1hfW1A/IKpjE98kiA9uL3TJNFQ2E3wr+
Ca+jTjGv8IKDyluRUM5PLf2anWiW3l0VILEBCHg9nIDiIkBR1NdgrC7BVh2YHIet5T921rZUs42B
qlKANCKgvw68nbGdyXyd+Q5cz6VOjAqcrqjAyDtbF0fgD/pNU4xYuow0MlpkZG58h2mJrVjBgdh8
ONb1Ne3lGjO/YQOBVglGsAp99BQgG1zL4B0NZW0Z7VVeAWhZTJOQfrMGay8y+xctvl6f1wY1yYxu
I0piYBcbhY/eQovIPTgmbhIfRaPQVpLjhqO3pHZ1E5T1a5UVShkaHdRl+RrUDgKvrvtIwyv/75sJ
Z50pHysjAfhTxINoXfua6vJ8Na0/WNNEOh4EPA1lkrsN5dIDOvc7R6PvnxaYrKu4VhKB/F32rgGJ
zHzB1QxjUmQ7IoBW2SpbKj7m3Ea1WvStCt7H3cxhunVrmljrGQEZN659IyIm4P3qJdtON66IZkIi
sPyNmLJeb0Yw8S9xw3nZ+nVJMeKbMCv/IpamQtmLsYXX86vBKQ4DiIc8cd9+zHltNe9KklRHKHOr
QDB1Y9K+0vq+NE6AQ9ku0pMoP7hdCL7cATTWatputLA10LtEGNLiHPNNwLS4U9Eurxx4GveaKWHQ
xwXoQa1pp84YKsj6sTTqXdRdxeMggKlC4uTvaBbSSkj+PdqUDNTsAkFvPCcpYHLVo9cEgjYDhKnc
Ng2Yc2wh72nv3dJaoFA/8GQyKM0S7v51TqRoz1mT7BQ2exqJT8QR8q4ZxmiTl6lRL278pMDaLCiC
eKsUDflKY1Wajw32c2kg9QwBATMFM5cVg5a0glZZlROl84zsBQK3/KUUZW2w4YtwDX1Nlz5FQmUs
qkWFQ4WnGwj4A8D0HAn10ST9Lb2kCYS4+xii/uOKzJ0ZAAoN6MvCxcJTjbkNAMb71HEDV6DoOhVo
OEUYFWAyJ/Is+YAkJPRBW9III3Oqa/yS0sX9TH6byyT7PBgyTpeg+ZcLWasUcqVNTKvg7Ba5dhjD
omnolOOSbIvromCNEEqCPEewNRJDoE5sZ6hQIAhGWvuKQgrW3zOnMZ7Y+FZkndUKsEXf/TZ6v8Lw
Wbea3VfpjqI73z7qkuEiZHpDOsVAwZNpTmFTPPfmjUahFTrc9f1qipib1hYQABQwtE51eMK8g4g/
SZMkBdBzOY62t7nnl3WM6Bh36hmoglC4F+46Tj5poURzZYdKTRXj4iAy8+UKZRW7o9jnsQvcf5pR
cUFcsj2yPNHFVMuJcrastiwYpIDnz5Zi8TM6l0yhxEYE6TF4vu1UAhNRWGqlt/COw/nRK5lrvdTE
Ia0okdvGvOhajE/LnN9Co3zMIfegA/9jTl1hfMtOGAAkkk6rcC0g39i/IM2Yfr2NDaRIW98OGriQ
AP8O6v+CH+8CawChtOlqcK7x8Kod+EHAC12IvL3hlLWuanFOdnsfu0wATK40UnCEXq4nF3YUUZ2W
sNiS4wp/MhH+ReZ+onibCB77ypATx0qyXpLZlnw4MMm4T7puIaENlxP8h7i35Gf2YfV7Z6Cgs0ro
NJsbCrdqW+fJteBSU2Vh7uhlMnc5V59KlPti9lQA2OEexAz29ge71SptROAgxaNk+DM5FEz61+J9
VF7WycePZ4yhM2+nBu1IvySlx1xF2+DJxYBNRZImmX5neJ6vXY5+WrgufuDbfMHamKAODH8CdDeD
BKeEgow9k5x51JDCYrEFozQw4zjUZ1vTUVlkTk9FciuTdOLP30LR0ONhT10/DO5JqjvUK/N1VBzq
5ZI60Oia5n16DX2FLDsD7frde2ONEFBx25vahbF+Dg9dPqwwP9Ip3wh5DjZdhfzkL+qQtfTvEMRj
DivQTGMq19qe3MpgutmWXYUJJcTtbKdOaP6/XvZBOq1BdorvIf51U0/TyxnjOFvXtqzc+PwqH7kH
6EBUym9v5RFl/m/xr4VmDWcnbeo87nb1rp3a1n9FerJcLnuYBls6RUVDq96hAd43iH+E1cCQHGsm
lG0iTl/V47geStAMFhZzGiYU+Uh1KKPOcH2nEl84/yUOR0VZ9Slycvn3rUg2ad4LHOWuXEw/KXhh
6GVZE/nd+4PlKpPZo8IxEBw1VEtN9/mQA96t3a37DDnrZZbfuk/vKegfiG2auF5Y/+5vq9Ft7/1a
VcKnNRZpYRpeBMjzoOHvPXzJAxFx28jgrHW7R1DZFNZFboEfe1WFiR6iay7McPAHGhie6MRMOGEB
srfHb6ALwhjMF1Dh9ALhSK/q9KWwJDCvFRLZ8pKVjyWbIft6w9o/hHVfNsOWivkCgqn6HwvpKJM1
WGM0vh22uSYNGYGr974GEjqIhBlg4L6UqlxFP/aa5Xdh0ln4/z4cjpYQ/eZwcT8sknd0v0fo5pr6
drkXANkED+fmHN7VPTKAEJ0G7abFRtYNStCxlM6SO/g5zHoT8gJisofdr9DqwV1OVsvM//jaHAT1
blKbv+F+/YyhWqqtcHfdjq5RpO856e2Tvp8r3g4qIqOCjK4vnJYRT5ijRnq/wrPhtnjS7cstZ9PL
EwGuZLPLM4jC4n75FNCjp1KrXtBbOI0azE9Rc5OD8k1dp68UEvwYRY0TEXgbKqif9QFcpnfG56f8
BdC84i+gt6nbtvefOMmRqNU5MtqxiznTsyB5RAxLAjrmjInnYigpUhK46Mxx1/fx+mJxirjy0m01
747+FXGJQ67ayHctC94xWSKsz8tdn8xBYgY7KMgc5sB3/sm5V8w6FzNmPfLuQhErn+Rfdtr2Jsw/
kRZBiUTfewoeiEnW8yDf+qeC7ekJFkgER0eqaP5aUq/DbD11NZQzsmJZ3/5qfeIJuKMZXmUUltlB
Llw8S920wen+ue4cr0T0rlwGJosP00JFADO1PID7o533amkbwqXzv0CM685ud/jp4qGx8k0zDadf
audseKrKjJXG+RXoKpBDBc7Nbx/vMLydJ8oDWfdhR4kCp4kOSfXTBn8MkMIKvzLRLU4c842MFqvJ
a+LvOfGVrC4twGiBtVO0ITbd9/o57z9OnR9xboGUHuT/b8GMPb0fK7DsWvGX5XH3/PGRAssiH3xS
P9QQKNAVO245NH589tOVDSTCUtY5xQwxA74Pucum2+t/vSOi4acGZ5B6U+VCNtOOMHYG9PCaup/l
SO28Ik9z2x2tuU1nYDqrXlCdYQFwR5NHms7yZPUt3I0Wh1SLJG3B3F4vMJ9hnFypKMUWylfvSNFB
oBkcwU/2YqxxEEaD636n5HeuhYsyuF4T88UyxG1Qp7b1eyCMTIUrv0ajHO7UfAmribH/vL7vnT7Z
gAoFcOAzZTKMlBi5APqP29sFm7p+v4z6Wmay9vPqj11ZXbwbhrseBmjvMPgM+UkQkyHZB81qkPHb
fjo5tg7wSvn6f9k1HeWCTjZJEL0eBeVAH1hGcRY43JphsgHFVyieVZ+0q4oVEB+SqTseIvl/UywL
lRgs/C3l63luLEp32vKZryHFK+d4FrRyaojqWT+BklvfwKcuXsLjhmLR4cBRzjlK90jKM5EWVMvn
SjUkDk8W339Ju0MXDz8TRu/AILqfxms9jqvHcaqlA8pgum6Mp7xgXblvRtlE1qp1oGvX+9CWj93u
kcR0v2vM4VtM7D9JMvKZDpm7J1MCIKsJnyXKslXynAVTYd9A6P0C939OE5xReGQpbQN0kwFQBycx
j91Xm/kjh4q/AKeL7SEgep9b8T9W/w9oCqGJXAmvydPwruvLp3PZyNaUu66ienYgjflbbSk3huEv
mEvl/gXRls/XvtKV/zDt0rMmyEJOY5DIX/cb1J1+PclvBmZetRnvFPuvmncK4Q3fHo++MqYaI1Qh
8lKW9nHf4HuKdGXzkU3a3vHr0zoSBZS1OC1ouVG5vRWoSGYyR0gg4k2CbzUovr8vUJypMaHkQnPl
0o9UYujPP4iOeoNecYiC7pzqd8FvUGO1dKRi66JP0WZwXg4qIcRvfQH6zQUXh7UZzbMecuOPOZcM
dBPKAyM9p6EpkVOBcy817Oh/WK+Tri+NCDwN1HJ7GxWdMuV8cIqfLqM8TsAUgcg27+GHD+s+kN7V
pCHe80EfOLjO4eJpoXzP0P84DPduXncp4E3RdOslwHuQmVE6Y1qNUCd5HWeSy0ErYgL3TyOGUEXe
ddfwyjNhzgWe6j+/14n3NBaBhfMtDinIHoy8ZQjLuK5C+pKDT9S82a7lwnN9WdWlaJzFczCrVG/o
ExgcMr/3uW/8I5mURkPnup6InXQttrYBp1gIA8Rnbp28VBaTlZk58oKx045X1ESmPEt34xSYtMfJ
obDJ88xGrrIb8eej+bmNFFbeCicbdVdCnSxLv9ELjWu0HK1FrL+XUwrY19GwJ4OHFE3Sj7tgRTrN
0T5gf527DVK7z9/MK4clOruNfR19Q/Z68U8Va7/WPQFFW/NlP1DGtipDY0VLeyb3N089xTo7QRTP
CGgbufgHDg1OivW45D1HK1n0TtQosH265DTlg++4cZrZWOim2W6z9Hy8dJNzsim7ofSFIbsab7eO
8irz9ZmwQOh1vYurGGqGT2mQ27zZI8F8dx89Bbch5dk2uOl9xcGO70r1exObLFU8neGQNgsp7sfC
ToFojRCTM4S8RhaX+wObNWxobz2agopA9Um1gsCY1JYR0XKb8YANrij4aT7zoR5QmDGPlpm7rlg8
42UcfrvncGiP/WwPNX/hi/HFnVRxWYulFXsM6LnSuNciKA7k+au4pyzWYQA8wS9qgc8s127qGaqz
t9y4Cyj7WvUWTu8v/BQ4He1jojGSBD6Nl3U7qlbE1VdVDlYuDBiWMdJcvXDFgxh0pz5O8a3eOkGi
YRxFahYAqhmworDKlOl4Dv5p9QG6iNjOOXQL1bwpDCfH9qNWoO2oEZ+YLDrXky4JMWzAdIo2tmMv
89tpejs8zmLtmc9WgLwgih/9RAwHwORj5w+IsVyAyyd/zwA5sS2I+CTzjvqRpVphaI0tc4k0AKAQ
yxgljG1zgwzhdxidxPLBUf0hfFAUDJXUrshrDaAnygOIbBjF477mc5A0vO+PbdJYh6v9F99m94wu
qf+Adc9lsnoWLsDrjHiZSoE4AxDkSUTMYP0bMpFBAqW00ls1QWVDkzmK0+Gi5LEfNtkqUEXMdnyv
cFGNINxesm1HXtNTtg/hI5vMnu5BJ1gdd4rqbGK0cWqrlLGL4bMFkROMtIO9+A5U3LUnTMnVVK7M
eigIo9PTIgZnCXOpH3tIjmXLRGMftiN6lz14LC+YMaoAWvYuczVjMipK3TLT9ZNrUA2DI6E70tgj
VjQdU0+HEEBBknFq2yL3vTS+3N/Fmmv9oxmcHugWyXbnmYInxOknVG0Pbxv+DGbTINF/7rUuhKn4
hPFd/qBBwkTi4ehUZbC0a6mrZ6WVgJUupE9cQjIc4nVcyH4RgPVSsqKpt+8bCFiCcfGFMC887R9H
EnBta8ZCmXFUbiRk9FyKDS9fh3H6yvHvZ/3+Ll67V7ut7Mp6ViZeTS4NHy4vHOWzCd+Q9SOCuKbT
/rqhfZacorbzSXoy0nEi5AekMsnyo5MJukZ6Zyhb3u75uTBbUexvhmOzFVFESw5obVsUeEBbRy9a
2cMrn1TSDMWzTSkSnssJNgmPEz3y347dJm53LwlWkE+n64y8yfHzwVeOpSPLDOsD+o56SA/qpFYl
ddzoiAw+ganaXNXMIcGaCJ/KDsQXQqFj+aNypPznxSr7id9IWtAJr9UU1vnGuxUF7ljTS4FM+H2m
3mZUBNIZ+qokivnUCgoIsv+FlV5uX74kmFzKD5d9lGJUh8UJpY1+paD/415CVR8T5bowmv9wOhvS
YCmlAC9UwZrpuiND2xx9WniqmGMMK+NzwTyEg8lorEC0N1g0rKNGv+awl9zcq+0FdHImVlVbyuAt
IliV9sKkg7cASu0yGEoYe1+fkXeo6gzquaR2jt0vY3qwA/Myxk8rVlBB70DJWHJdtYxKaf04mdGj
/hfbbJ1ac+NVxp8bBCc+KRWbz83SiK1ZL5mel0DDiThIfHOsveLIukgDsS0pDk0Qb8tV7HC/Jj+V
e56FL/NEwxahw0xcUgr5QiNYJEdCmU/oSk7uDJIQz5NYIReMpHY+FiqcoC4K883w2/tTCmRQY3dt
Z5vW+QHgQ0UL/x2WTU5g99me3YECgkZ8Pwx/K5sse9fi9m64ZZP361l9OFcO9OJ+LwvCVOW/pUkO
PXHCDrCKk5LULmAEDH7ST8C7r9Y9wVTHrwxvjVWeGngTc7dRAe4qVQDQty6WFtxZyiGfVeZ7F8T+
qUdiOSNVhmQ2FxegPyNC9sy05EZVA5SjPb0xUUMfk2CyK4CXDvv1p/ywEFDmm9jONurbVsSmh7Ym
/fQzqFW8Z+0lRDbWl601NNP/Ly0iayswD9WgHgjEHzRi1P5Mt/M+e+FIB9U0+LyZ8bjXW5gv+88j
eb7QfGalcItTwRIRRM42oZASmJeEneMFeGVbP0wOS76TTnntD/ZwSCBDb3yoUHrX8ZLHq4eFhnwk
Ictw8mYMb+WmbmvjzHZ4yCW0N9l9ds7Xj1yK9ktP1FMvlQS5LPOt6VMlU9Q0QsGigcECQisE/NmX
NroOnWjKdtIzJPOSJLEDOwScScXYd+hVz2U3uemS/3M7+1LQcZwXrfORtMmfRVaEq3thqsY5MuOR
opSln/D+9tsl+iwIawuK3CqYZH/Zc6bSYLrrB6eKk65yepagTaHrX2FnCj9Q2LdHDE3p0fZ+Orwn
YUBcJD2GLbzwXsSB4HFNcCDPud/s9aqsj/A4OzRv/0JKUitsZ0shfUnxq/Q9IJXJuadalGkWW1d8
gcB3mslzBGvkB+DBH0/eAv1bPtuLecSMA4KWb4BS2krxzm7aVt/JFfUGWeFxuI2fz+Mfy7jcuj4n
4H1dbDdX0dcEceD5kSUVH6YdoJdyfr3TNRkPvkF/oHtwL56FiLHL6XTsJxsbmsOVe1owRm7wxUT4
YcCFXFihOazmWjd3qLGUUQQVycXvUlhv9XsL2N16ysefDukRd9nAJ34+jfmeE4AnjYnTQg6ypbEM
cvn7esVtfep7wEFQSi+v37N/urh8lQmlFLFF01Oqye8EZAke+/5KhsbrmbVodlh9rEQTeqJkh56U
JAHK1r6qGNkhF0lffGNPGtkqMK16cveY3QUOAH7L//T6eiux8d2TkXOdRTkgdD5syGzzWsUyJroE
vPufDBLgez+pIFB4HTTuUVjbTqhaIdjPtKH9jztJLzqtdikjua4nVyU9dlybl5NrRgppAX4yS+G4
SvlgoF5DcjMpDIV7W+l/+SFun9g/ylQ0w1QUZJnlie/aDxdvnRvUkK2LeiS3w9qOnk6nUwpXu5eI
XJ3p0lKS/fI5KyirQiJJCEJvRc8c+jsF5RF1f4MlxrBBdQ9f0B35U9BNq5QhwUPjoZW9wu4C6NT0
dtaiL6V8sJve4LEh9mhFw7Xg6El0lSYh6RlMPNlOSgNYcM0HkbHqt8f0EzT+lJ++Wwk8r1oR51SA
rJ36gLYitZbthKW9klNzAreufH/bz4u4UEVX0OutwDt5msNUef2UM5Wd35uhgyv65dCERuJUnGz/
Lmx7f1vqjfgMTsj/QyIY3/AnAxvuKb0GfNyUGp8OFpJApNdDs5Ytm5bqtQ8KEzoRYgM/9tepiQI2
aL8hVrfmHl71yAYCFJIEi8nlY7e/AZC5JMfQE11OZbJmZEsoOQmlG+Q3BITUwSCHV66/4+uGVZp3
nRQGrH88dlk5rlCAUiokx+L1+Z8iiE3rHI/6WIJyGZVVqKDX3SMzDa2+g7ywmfMO8PYndBhbm9RI
ZBhZj7NJ0CiFdBNgUtSqHXUNmAZC+X7YIpWq/j2waKhnZfBhrq/qxr6kaTLuBYiSPeFnTIRtpUlI
k70zlXwGWx1VA1djJh95XGk2dfl5sSTZquaH+QiOnlUw3DHCKLFaoqA3bu5CXfT+sUtC6+IXtk/w
4WUXkFHyUZf1vjQasXLsf46Xtep82MWbhsAigbuesJgv27663HBOFbLr4AYYF2SSWctf3SZahbBX
LXFga4G1fw2Ec+UMUA1jCfMZZnDMq5DwaDMxCkZerwsi+WQwD7ENDq5dZ6E4TIXHMz44/59dLcmQ
Ic4Z7LvGoZ8Nyu/T4adMaO9iGAvUgShdeQnFZjxvrcSgFyvb/KRQuRwuOc5ZatZ9Z/ziTRU2Zi99
S6PcKLYtLXVziQdkycVeOQA0cZA+SbLBiSRU/S2raGZ2hCSLeTxpmTW7yrRudvDH21Fj0YvT86vI
FhBqN5Gy+GtSP579SYmomDafbjFQ0lBHHVBpeESinDiPd0BLkb1zIdUYuY8WLxHpjlZgEpn8cDSJ
1WkOMB/yF0b2c0X12dZRR32JtkPOWFsbo22jN9nqjTzVSqirWVwNxptmEfw52dcTcfmTvcOrS5I9
Ipo+m+ykff1ACx2yQxmgK4h1iXsttTagfdNX/O1/wOC6hZJrz5b1QqbOa6wFAoiCftWUWJkDEM7E
OPmrhbW+JitMzypsFe9Zh0ejl2K8Rg8FIrkofg/eGz7pMqE/wMdWnTJ4a3cPuzD0l/lr0o0qrbu0
GmJ2HjP/5r7mpUVb7CxeWAQG3N3hhc7WGBtBNfZhiTAGzbPQHOjIASW5B9cTA9YTZWJD0Yltobme
dAOi9NMw53twRfA2iqXbxWRXLjb58jxoYBMEragtP8oIpON3LXSepLs2VA5FkDuJHM3qwGBz/XNW
+8EFHlbhR53cnOvf3ZiO80CY3d/K7bxx5oIAShO8zOn7E8pJ5rMLqPqwfRDN4w1+BTTAo2UQJF7J
rQGGGsudIzG5dfjb7f+h0aS2mym0GNAnM461n0nXM+wrMsGP+nuHJjAlNrsVifZT7XgxksVYPrPW
cQRqf1zhTbOWRY/dPHrmsc+Cc50PuPH5Wb4o0cyEXvTxlnxm0uhf0GqaAdRtnPtPS8/fzL05+VpL
AcLKfCUy4M3cd16J6SysNaW7eEjGB6vyNTeFH2mvDiqC8V1V3+7DCFCoXd+FZvx7LTcMM4HOf9Gp
6FjZL+4RyyyA2/KC4dFSCe+2PpsR21uU2khFwz7pv9io54bBbwToJeRmOYBLiIbdiBn3gvVmTxeO
HshG1YvaynDmhwFq8Mw0jIphiTg9gSaKiURfQKHV8brrM/Rl6ByxEaT3rmmDPjqMgAY3bBV5+cUw
e37vU9dk6AfcBYb2j3byaCLc2GDsk6geY3Ew+FxN1b+8vcSI8Pf4aYiMg2CQTikwLcsk2i1QD/+U
NP2DjHUmtAuPjwDjDGTHc2I2Sm/JUG/nTRFQt/0dXw6ApJnT0SugjtMMlqe1cv5NIYdtGrSVOuo+
oCDenjYpzXlMkhjCNxV6F7+Z/dMezINWHPCy1haY6AFGJYTEZ2/yls4GURGRwXqsaZX7s8k6R4l3
bjwtngXDLzMKl0ZRrcTLbli/1rpSaMBMFSewaHxsnA4Xaa0xWbTff8Gk8O3RfdbA86O8ogJNVJtR
CzlJoEIJlWfoadjjlD3Jw1HRyf05uj39KjeomMNn9fOFikJQlncELZKHqxTttkIjQ+ZkpY8l+2ub
C6vmuoYlkr4dv4WlHfc6X2z4xctakSEaujR/MHUD4nSW2sWeCxUnlipheG5uXM9lpUKzmmsIAgaU
PcvvclQZZB+2SlKM1c52uHVInQXZ5c+ZSWPzI5/mFHsDSZnyHmtEz6XDgR1Lf2JWDnl1vhs8Apcw
LIOgSGMUrQMDyJe7R23QP7Cu+Olz3EyTWPfYsJYd9nJacVHaOVB2o7bzp9A3CGu7Ajf+XDNtxztl
zYtRIXk6FVIGrutUZR/q4Rxk5Pr9WzzWZeApJqIUwRugFKTbFe7Eed13tZXRcGQX3GtsU///i11C
KPPml1XfjhRR1s6ap1/1hAIkbg4gXwBGlS+TNhKGrkowxYrADtsCFNzeFiAOtWakCDYFqEcR9jrv
+X64C4UIvys0FhQpdKMVRleyE3lKBUSojSFZqSS+BKAenCKPkPetqPvjkND3VbYPZiov7+McMfK8
HGiXraeyXrsTq9WCrlHzSSUaqkqfskrDZB1ep9F14jB02XWieQUP+gCc0qlTuMNgoJ/geNMkTX/6
XM7kwfKBO3jWpk9sIQgMtCsV9pRprGj/ZYfJjhOQGSvSddPH3U9bO4CNznn5mleGHZBcNvqXtJRu
SiU45n1VLxmQlns93JTNRUBM2WSdvQG1VzhwZWZg42/LrJUztMYuJAQe+VX+jUrsmzcyviYXcuFX
BydXQkWuPmKMIjSmWySnO5nEf0SwaE/DPARqruT73uuhPbLxy67ZYFSJGMU9IKH9YLfMJnAseD7v
JYcoSE4igM0HQDoTnSmUlmjEhE4W4nQf66CRCS6MsNgdFxWAz5oAN/898ltr1lSf4DbuGBRwDG82
rEWrO6p6gmyHTfBGp8bkdbtpFJXEOEBjG91uR69z9qKiI/5cmsZv3ttgQZ4RI48w5o6qeCZhx/88
Oaqqe8zZF52TQH+iUNHUTcCyfWTF1c3w7h56K7LZTsPn95KkhiEHzEIindgDirR3ZMSVzJi6PTdj
O/VdFgFjeK0oeVSh/oyGG+10A2WznFZFBCUiBH8N9KH1kgYLbc1RbxF/csoKCvUqVY3pQmhKj2gq
ijXUmJu3AmYOUSrMhxVUl8G0wcG8Lo96eyHUqSsxZb5TQwsiXtmqVpQNPAFOvW3SkagUK3ApufbM
fwlI4vCC3pyiMTVewySZg2A0Bn9D9e9y0HSl8jJggXWvrFVz1ZMpvk3+yu4RUGgQOElnk4eUtYUa
6DpD0+8e0/TxqHxsTi6IXSg62S02nd3GACxYLhZjf1nsxmTL6rG6MrWMQmUMTNz7hqaEAw8YSniA
hfCwnrvRKpCrQLP84sNPBgcZ0IREnmPzq7aHuQVDRpwEHwqUVlbsC0VIpQLX3ONt0eoYm/Z0+yuF
PF+8YHmzzjus86dpZv2x+gN/d2w3zY/RYbv+gG8ELJv/i62qFgXu4HtRkSYTlSzLy6eYCYzFy79T
T2hjABUObO5gdca3r3KgXrPUA1JR4FeXn0FfZgAGufU7J/4/gwHfjBy1yv/NQfMPTux0dG6uJwYw
zQH+V2yO2TXkd2ZhcfC29o2eF2mxdhMOJq+i3yUrUTS7HXEgPhXP7naQtAWhAdLHVAoTV9ObGb2X
H6pkcaDY4hQ/2238CKUyCBQG7BKT53kL9t499UzFN/jato3pa+7ddNnLjgtRO0bQV9WnlqffFj+I
jjuR/+0NubSjkQ9zIRx7h8x+3i5lQw53o6jWu2Cm1WaXWOyzr2RC5l17BeakBLiyHBA1tRY8ZhqO
C7cLOLKspReFj0xBGiGOXAk/zJS4x8HjuxKL72iFMMdUAbJDJ3JIbWireHshDboBi+esgTSU3kmZ
Wfha3lP+MT1sf5SUvSK4vzxzGSKsqEsDdjLJrL45LH99dyODbs7Drn0KlkZLM62/jK/OkqFX4/XN
BakDOVbU7phwlTyLB7NNfN151gORxZKwYervBCeKIWrGM2F1kcA9unJys3OWfZ1cP3KPqw9UPG7O
ka0aa93xdafPlA5CjKuPTF0VMRClQPkCXYa6qrz1FdwmC3CtIZb42xPEAVfw7oRERUt38Sa5wegc
/Uj165mVsJ6FSVlpQmkp86esApw8xW1qVp+AmVNZWu6O5c15x/My8MSKYYd8RpB3Mjx6KoBgW9/D
lI99jE4cpT+UWEdD1BRWBpx5ZhIOJYxT4W902jXBhqnZlFAOE3KT6BoBrNnSChMjT3/jTdjhVcZY
0sXkrY6yM6LH1dsxmiHMuIsyVzAbNjshxQaoJLXyq6n4po4Gqt8h37jvDQ7iwWATF183AOn7eeHr
dqBygKJrNTT5+W6urpfFK025uX5ESwfWf9BAB7QfUMRbrC0kQjfX7AY6ISt+Fm1vrq61NrWm4Bcf
uA35R4uz95g9oUVXkwGwdkUxq/DmlHqTYkpyaJryrHskbr2Z5RbiKDxF1bQq6xtU4lYd6TD4pDN5
CQopiFiqFLr/yUOLLVPl7sABfC36oiAa9dJQeigNJgJjbQEG4KG8zMduF+zoexhJn4CsdQnwN/jV
XR5E2OEHYVESMfOxYsNoA8TRoZ4sL0IA9JQRdCw8tOTEp+BkOMqlE/IyxPcFP43VS3vNHsYE15Jb
1ZiFbYN+XQ5uQ/66iRARC0NwkhdstzPOetX51s01OvHufKdWiiNrZV3yzDaP2Jtw5iOF/JNQ7Nnm
agYIA0ZPr7RVZhglpJSrxbl+z7/kgs1ClVgE2F9yJ1Na50B9hdYm3ovztEID8Cs89DaFRS9uCel5
zOTl1vKhvA8myuarHV/MqFh3IPsx+9lus/b9aoFkPcjhlyT+gSG2Dvjy84yjapxMxrixlnd1RkNh
g1cLMnqvxST3XNOQLxlvEuzWDHVr+cpiATZIiMl4uoCnCJbn2hk5jPWUSB0sUEvjZw2U7zE7VHOU
gZsJ6/vliPANISnuXdoqI7uu3bQmnycB8x6IYFKXan7eSIFbe1Kgkaosz0QYBmfoAMZU7VH+jcQt
1AlP6MHkWbdgn0Hd98D87w6kd9SC7moKRkvyBbUx6ubEVEBCJMb47beBj75sYvjQU31+F1eo4uH9
07n7XeY7TQaX+//uwIAYGHLXiVXOSyBIA0I8mZkdndnhO1p6y9OlfoxHOFHYoIB4RqTYcSBVOMUX
HUlRwx0D12b9PzuyKxkVuCfYG+snmx2+mqf5GdtXZZaoPRbrKWX9xaH1noE3r7Y1NPiG7w6EGI6j
1+CiFN5Swjzyog3RyD3tzW4fGxl+63ZFYNMiNAZG5x98cb7+kiRDI41Ix7eKMi3ITppkQ0aZdlLV
FQshGDKP5IR7kObb3yZNmx0fVs9T6WtS/+7qxDA2FiLTRG6q1ooLxSRddxuGVZftsAvJ1+rLvebA
uW3uTlkbrbQP8RyMBfLYIlpTcXfs06VPeN8oBNcpB7eJLtRtcTdk3Qx9C8kjMAcNW+WBEhEVEZ2j
++m3e1OG6DuYzRF9h1XdKYaTAyO12LmL9ylXurVpb4zLTX8Co/nx2oj6EQiiLKNej/ufds9ClGu0
X0H1NNuEt31lCdOQGjQK8zl2Unuv9YUGev8ExIN5JXknVw2XpPaIoOw3rN2zpbunWH1DjMwAfzNK
GTzEagB0T7MPsn+R1QnWqglTNogM2G0cEk/ycs7YiDrlxbSQMnhQljjzSV2Ni8intT3ryGBTmewc
RT+9SbWNKMLXZFFVxWShQqiAeqoFgSKIHhE2bZ/WXeyPiJGKQ5qQZjd4MwQMCWmgdhFNScU/p4im
JqhJd+BQwk3AeWVHjWhTWPTtns0IE8WM9JTPprx9rozfInlOsAUth6uS0itc8i7PcHRWTD5MzHqD
MG7g9NWn+FitaPobHTkAeh1+zXmeCDgNnZRRSZ51S5xfyvbnCeJAU1sPiXVj5Ck62E7W+mrkQEam
NiTkRO4kWKVpTA7Ki9eU82TivGuUvT5HBG6ZHR8GYmJ1H4CnBTf8yqb3NCyKEzEKurP4mIxTu+Ca
fcBT7O/YGyT6BVewUf1cJMdw4uCLm4aDbEuQkhzqx/orSYlnAhKWMMd/Q7gDvlJbyqq0Ig0t8PYj
g3lbmzCO3tY9AEWqkqRN5e/Z5N4QPF2H+IwYklPlCb3FalHeKU/lKpnX7t2d+mWKyax88UV5OuCO
EM5hlQ818hZ8cgaT5AyYKC6QRLXZn+4/FuLyjiI9OLEfiy4+SzxicwiYovwCQHIp53L4MbKitwFT
ciTiqS3F1mq5m2PCq1HufNoDtK9kviANtC8yWjvbxEKSTG+86qKJ4EZ6/33M1UxoU4RWQoTh88aN
4tdRQ44HxrXP1e6jeZuX5V/Z5S9vQm4CPDXnjAQXD0iBUfbBqdK7BGmAG68pXTlWtr6r5VEccIlm
SMG1+gFfnvtiEHzUB5GripW7UyhnPTvZLwd9+9zyMHeFdsOfWOJAi3mOspnzdxgBOw50v+F8j3l2
D7E7aA6LsfOaZn2Upq18vx14UdKmVZYLKViWL1TGdeQrwUv99lzCPTtx6MLQ6yY4GlQ/nDaDfBw3
aa1Zc7AA1ehHSZE/ZAcTikMzRS9phSKeUX7fgwzwY6CBKOghfDrOf6VArh0kOEC9A50f4ENwqV7V
KMry3qFNuxliod91xtE0UdeHHu8vl1aeYvuANT6Sw7AJYkkJlHq/V+F1LTjJMkRYKOQeErGY9Uuw
OHo3nr11uNYMy7Ce24fn6thxR5ACSkRZQSW88XFBwQcd8i0rVCwmjXFwXVsGhXnguZxa5OOrSllv
vBA4CiSl11J7Unn8w9FxLYAT3XYp0hf1LtkWjI5+JYm33fujDQLg/iJw9m8TwGG8uZ7xQknTseCK
fuwv8IFYzgT//5v18fTExkSLzlDXgdJRHIy17gUTFziHZKF+aOhtEBwQE6xfSMri5P22gcDTjB4G
dE0hrkbIzdnSg6zsDTmbA26Jgkqfsv1Z0DgS1x1dQFI924o3CMdYVP6P+S69XkDPIf3pGvc7zFTw
ZMh2Hq/+myxs4pQLEgYF1wnchPoWCoHEKs7sQPJnORt7h+yUnKR/GjblmOA1U6wu0mdHeUhoxWpT
hzzKMLYVnBVkVldeI+p0UMux0IUkG+Ftvm5gqZBfklJo7GAgdKROmBVagfuMGRNG1JezrN8R5+nY
fKkmMPaZPDFtO/ZwP7KHZeO7ab0sMyzOW3LwyVqxxZ8xZvXMqdG7XMGK9kSs2PFgWS9o3XqJmwOM
eECLi3gEDR7nPh3iiFPZOf4uIzixZ/KTB/tP0lID0PhGoA7KEHG5N8ndcu65xNaoQnC4Tmdljsnr
0veNo62g6IU9AyzVoRVzmg9hTT7vFPEstD+RPPRdykadLImfckMlnx24R2I1Ngh4OqoMxHOlZ42b
ENScoA76h7ydUF1Ta/FBN9m847+biFVP1Cy/7jtHuzB5r3T9RoloZEADnr3I4UeTihXNOZSTHHqy
EsNfK6+AqHcp3ygSx6bNWA4D6opJ2gWP+h3qev/Px2JvI/KQ2U7pQ4m611MiVNa8xOUC+HOmBkEn
K4PAuR/3iAMOhF3XmjE6V7rrlHJ1lbdTjSvSjlzIJbfgpZlG0/j5/g7H+aHwkGJkVDWDH7yVTyIx
tBhQ7Q88avlekzSxFu2JXt6EzIk7woSEYbqvYDiDRrWoNUVTBdn09Y+14n2X43IJOyZfihkLr7QT
0fz6koVD7BGElfs3AQh73rt/CJbZOASQzpsDmyK/xOjIkk3wWEWFdxl0StkDgEZblQUIwDB3tssj
0e5+ECOQsmil4qI7BPrvbO43vqqX4XM9Wu3//VdbP8afx2mv9W1fH43KxqF6pEFsgIYEgZm15Jmf
90IZeK5tGhxddzZTwGIQcfOARyfnEtEbqZ78X78vNBF2nK7LG/D5J/xK2rxTt1my8Zj3H2bSLtNK
xoMe4nXRRqEbxGTgncoto3Pn8uZrR+7ahlc4lz9/c+BcHILGWBfJMuNogkXbrsP/BUsbWRcFCbl/
O/nbiNj/V626puop0O4GF27Yr/RMfW6VVtA4E12maRXN0EVQxaolL0cqLczFH3FZj/cyd8THRHiB
mXQrREU+yFi6ZIc79APnlWeg6Vy06I7HexR3OHhViRMpkQUULOdGz7vnMIxttEW6lCbaTlfQsHxX
GqZu/M+7iL1pHR7AeZcumDf6+hN0KRF+64V2+1Uoz2qrcwog3aeJ8Oky+/D2VUslHN4L2pPVaqtc
JygfLUTI3KH83Utq34jlvoKtiGxKc7ix55sI2/0uoaUX6h4cgGvROVycIQuwZ5Vx02NhMNbGbZ27
hU9GFT5TQwA3TWgeQ4ickiQB+oZBfGuRZ7E4mjIasAS/xEN2WuMmXb5blYupbU1B2lBU6+5LPU3y
DzKEoNAe5ZLkRfiArI6jj1EZBk9mhepwMd8a09P09P7FIjiv+YbjMB+x7vM2UyNbEzTq2Hnvof5Q
dh0fYfLGP4c8UBgx8NEZNS1Nk7yxvFc6TjDPdFfSDxxcp+q3PDc+LETjTq0rVj3jagN8XUEb+aJw
vQSqBms/jZ3KhI7d+3jn29RmJVXUoLmmLyfSzU02YYYGJO769ism8R6TLkqYnC61Cd3m5XNbEFxc
oRcIj03mS67eNGn/QNO9lP9YENW1xQo2Soeg7rUV3qTkKmWGSgGHuPVk3B1xPyvkMiOuuJrP6MXD
KzmZ/Ojzqu17asQku3gsCggXy6mBHV8Mf4mC4uSHGuqQqgryMstleXwdFhgz+iIvl5HFoiZbGO8w
SfPmduF4CxlSe2bcObZ8a7BxJODkxxSh3W+9tALKAQgd3Xd3nZxd592QQPLAexCQX7l6SMpmYrYr
JzH8qu0wJeQG3lh792cQt5qIoL45DM1JzX+oQPv0XSkFmJfGEasSFb01VeavOcvpO12ZpVQcpfxX
h8KSlMZ7wx8XkcN4jfGBNLmZEOXI20kB1OS7eivgf84HMea4LgMiiTzUstEcx874o31mqsxeL3sx
NW7wcTE/JM8agrNJ8G/N/FPlIDnzRsjyWRdBb8oCy1ab4liDPJf5Mcee4ARfS7xBc937Ep5tSTiT
cfq91v6UmDJNpUswYI3BU44Ww9m4pLYYMA+vT2zeaY0pEH+lePokPxW4tUOsLQ9TX9YaCi9EM+3v
TkjIqe4LwCPFFpYgJbtSXlWoei2wk3sH3Nhk1Jcf5XdmBQdYEVWMbj5nR3LnkC3qoyPY5z4syuJ7
RoyveJZxyCI9vH7lRrx3eM5Zx3Tcmar073hz+t9Iu79AbK4wDuwnhJMy6kFXv3ZNAnzSynMEaUOp
40CTxK+VyT7VgARw8tpLJTTOLYjHEEvNnyIQG46k4JQjeLpif3rhWMrhqbkrgct/l9aM5bssxAFZ
pjkMKJeNViPhPyo8PKcuXP1FeduvTMD2i/vaDwUFVPPjH23zfinxFYEwE8Ei7XKdDFKrvgqt6ufq
+9EaLJb9wypMKHN3o5ny/cwbw3YydMMMe7vi0nHrlQBmgvV+LPQaKM7tCHavK0XE9CitdPaytO3y
0hb6pOB5M1SceorW5Jv72bFDTfNjD+x4S8ZXVQF9Xk0YExUdEB6UXXzDyIPvyZPyDuHlGfcJ+AXG
x7m4CVXtKI5KnMWYSUEtSnJUqCg26VAskyVBBifQq3HqoFILhvV6djvTtwTnsgQmV04Ri5ki0DnH
Ieg4mzXoWNH3nfyJPEcYJwltBBr3/nUGJcfOIAuTsCiKV1MdKJ6eYFOOy8eDeN7jEu+V5Jj4q1kt
72zzgW+LK0cBry+B593mnU2PhpF2SHNskGuCFO6Hz57816lhgvtd2EUj3aaMp5HCRtTg43JEkeCA
XD5DMgPSrKYPMCSDcpXJJZsGDlFe5X19Nvps/Aq2kcTqf+cuGXhVKNuwl8QAjFbeHj6AIvuSGMT/
tkSk9LjHF6PJ4173SWZrgbHLX5A+E4yyLpIv+roBJRYjNwHRwPsD8U0ZjRWNl3c7e3KvMEFxUBK6
Wpztokju9TrV47UT3Uyh6SE5v20PYOd1m6HrbhVaVekg91pLDF/olpEBOgZ9Xl3CB15kyKzpVcQH
0BtxtXRsn4DeEkJHu7gdjhBQUZGjUI6qgEpWRKy/N9LMUkDZDhroXsCUK9+Kz2gdWD9CgpqwMADU
UrRXkW1MFXW0W39ZaR5tkogYuu5E9NF40SvIt8y1uy8MEI4kpQ71mM1Xi/Fm1y0Yxa2mr3aqfMQC
oKbC8kKeQbYsL4NUFYvqK2kNGYu5Btq2shBX0NU1KmCEoZyYNFN1nP+/LanAXVeLGxh1gXY2kIEp
SS1cX9BalW/thQm6j7/4lTY4m3wJ8D9vvKomIX0CpivG2fjIMhOOO4VFwe/aZGa6EZe+0IlgTQtA
nfDHt2hMd7Xnv8Kk3zZtDT3urhR45tb9G9lfcBopAqKthH4qKxXi0n3viBPrq7anI7VMViop21vp
5yL0uI1ePX+4hQsRkzuqAwTL2j5yK4d9O51FpKzEZSFKA+80FIRNW4y0WbXSGm1gh8BnWilxv7u2
SJ0Qx8qg3gGa/Ns9Z3RP31NyhY+qHvTFXeOY2FXYFKmcz9jy9xaczj3ksdNlexDVfn5wln3ZqyFf
Esol1y+ctFkpCKWPWSide0645kmMvnW4ypt+QCXoFqiwJclHL0gMozrZZjqFGMtwXHP/7Zq3Hgm6
r7tw82NqtvilqWxEsZemg3dACgq/5BIZ7wFAeUgf46RQI6j5fZ9Gk6Mz2Y2/xjlfAh0/NU1+l1D5
9ysFQaSEUNkEoMtWjzJve1emjKpxcx7kxsNm8CIuntv5DP6z20vo+BqjES0lBbw+aAP+BnSxnKnP
HwDdbtO0pBUWPG4V656mzbi3IbW0AEWk7uSbn3HOu6cLyc+dTSRrrRrA0qh2xmFa/6SkikwGwe1f
gcOI1w6a3RWAkTA3QEhtrPxfrqtv4i9tv7TaTv3Q520GlVdQH4k1JS+BhRAlBcu6aumpxK57YLZA
6i6dxg73ecVrJ7XNL950EgsUAS3stubhp4k25EK9jPq2gjo3srqu+b8qD2j85ZhNf0EdVGvpUjgS
P8OBpomoVEigSFk71aj2LeWw3rY2jLcq8TWSz+OZ1v1UXF9/vrzSqO3PJQO7L+dryAvhtHeDxWKI
LB+ixTPP3djzD/4UZ7nhgzleKq1ua0YEwVvxgLtqx4pcW5/VJQO9E40QmtR7ICOSkuW9g/6OvRER
V2hd6CdzCJrYJLTT7hXyJ6DyCp0zqSD4OhLOtNoIJTqJgiv0UQNc9dnZZB/ycOky4iHhy+h1YVKr
yZgwo3PRRgPKGUPD7TtlZno3ceUfFGoSVtP5W5gTMRLMFfryejPHeAJsqucEeQN0V/BNP7zpuk7q
fe6cKucTHRYd6lSy+5CkXj3gBzsJrp94lmMG68vh+ZrSOGBdeIV9bKS9Da8sJ0loUIQTOyseQxbI
skWW/aSL6EpOXKl6thpMRj8yFJn0FR5KgQmTPdQ3svkONDiMFc6El6fB0wBSK5QaoVBzxCEQ+TF/
OkMzGlQ4Lp0k+S54OpjL38Y9XswiaAYpMzksZKgQmc3b0VTdjyby0aUgJ7oZfpqPWxgROmnAP3CN
Acb5owe6typI6AZLtS/r6Ue8qjlNvedDq3VflJFfpdACyJTuPqbkQTI1kT7eR2mN/Q4x0zSk03Nl
YX/m9bNJ8CCbuyjyRBsgPM7IDEfZ4+uJtsUC3gK3vvN+ZaCjGn3/+dkdqsB4BNerrudXsEEaYAMz
iSrNhYm2WdGgUBCy+AMULZVGsFnDKUHi8HIt0xdWcpqM9ijLL/3WrVHaqDlLqstGH1HjnueVd/OO
kh7vB6Bu5AkY+q58pDJJaDNPucf3kdUb+Pl4xbIl41u3KC5NOKkbRIQzXy5HlNFf0YY+wsDGzobz
qloDjsIq905XZ45q10JUcp00XKjDEmHnzM2t2oTpTZoDaxUx4VZ/+YPVt4pQMB+sn3ftiAwL9ag6
JFDnt7waeaop7Gj3OFA+FDhU/EebhwoixAaqJjTpIUFKDo7C7sibwUP7iMBf02pawaEt4VJzOboO
pY/Gm6ECFAU+RCV8SQN1uopd5cWf6lCoN2vP6QOY8bZSVYOu3Qeb86s/zxhZVFgUtnVZj55IMSgi
EgqJfJA8JI0ck8I2zkgncQRhmGMt302DzxyIuOYx2bzOrUdVPtQCiixHo5f5JKwsaY16XtflAR83
+Eet/D4BaOOm5LX9FqrFc6LNYnv6dJ4kMPghnqyp+UguhLDVjA0wwEteTiHMZrENdKjT3VD2urwO
/ocb+oXP0DY8SZtY+uJmZ84WbVal9qJg3lcJlYVTbF3NhFL8pmEllSqNzv5HxMMjGimMbpqvt06s
LnMH7piT6YBpoNgJyntGwMTQHDFZjyn5MlJdzRs3S7JbZRtFnxDkw965qlPqGdHx4VrZNXrHEx1w
aH3vNQUxwHZ4zg3y/rudjjyUO6f0cxbAAPprb+TbRSCLVhOWes++QqNdxShOatM4Q1mSWcruT+if
vv8NwTFFD3DEIQDXxnDvhLl5XzFZZysFGyJdhRg0oQ/3tBRBc1oJV9ji9O9jAlTaJu1fUiu1dy82
SiOkM7zPtL/DomNlEwfT0z90/PYUO7O9rJe71y+s9GeT9E7ape6ftGE8YLPIge1A18ZAka4V4Lhf
sPGIGTVQDKOCvN1kCrSt0ihX17AYD9EsdkQjfonXFASoG6rDQ+wLYE762jrX3UrpXbgMjmOU/5TG
tWykmyIP52mzqVexDgMvoKPz26v9pcMaRqwRGxXnepC16FvzIZhV7vk0e1vvUHXXgpFqrea8oTXT
mPD4v73JiYS1P7MC8lklj7IM+6UecnclIcivVWY39693kR2KRRvNk653b+G41NdiS1tZy8Za7vhV
Kuy4nrdmmy5PcCAALVkpr7gawLtzA0FiVaCfSUrLk17nAVtuSdT441cCI13zaMhPZcAAJ5PO7xXW
YS6ir5RKQGKNTbBrC19p/9nyCNRHCNOreOqZHuFs+fd6X+T1Re0ZPoGg06keAx02fkpBNtyfw82j
dByF1acXTqQMCFHmPAd5pP9zmMYGeE9DwnnkE9C08kzVD7sINTSySMzivO6i/wRFV2Slp0i8geZF
zbttYL9k05l1FINmXxuQklem6dstxE11U5Qol1Mk4k0URgBgobrhe/BSoeqW6xELXL1xyB5UvJwU
nbBmWSmk0tbamgA/vRk6bg5RMNt9GTioOwEFCuwafoG1z34ZiFO3Hf0pr2VaQwJCGuxFjQGlVGU4
AvOgJT1vpRin+r+KXzH1dh6kkubQj99bItGZx1dZ7lxxz3ZiYVfnV2LTkSR8lZnrQNb5cogAKqJv
VtxQFSN/64xtPP2IoWV1vHz4tt0M5i1p85MSJ/k0BSZuj5rBSig2lRYF+loShJeUE0kqpVHjtgdZ
xINjiPgwwglL0b+hV9lJDj3NKotEWEH3ry6HsscLmSJk8rB8KrEmo5Fone9v7Eamr9VEu2jHuOEx
k7ODbY63LOvNKg6G6TBw+WtyD9YzkKahr4SENN2jef0VTdMtsnMJ7AQRCIxK2LzGtD6hsN6XoGwM
hvKtLaB+8oaWrbgvrTzSxCsqPl7LSn5/lt3LQpYEALpp6CaLOrbIzuOE0mWFDGOZJCiNbyTL9Gzm
zu3IzX81GwTM5EiLu2IQFEbl4bE92u+I5QUo7VA0G9R/3XCwRGfydWyQPi3zpKhrugK2gHbZDSJI
vj8/OaS8PECybCecrb5TUqy6UM7ZZZPEXM+49uWaLyAqGHfREgQMH+VYrF5+n1w6lTB2L6kvR5Tn
REuhTEIv3G72wTpqBKfaYZpVXmePUpDhq835tf5ot7XRFRvdLAfPnV72gm/GUUI0168F2EJZ7Gwq
InubXX6hJ81loWHkOVLi1ugVH87mv5DfhonjXGJ4LSUiZ+KTq6Jyn+8VoBo9z2RdPnb9ld6hNnsf
Cj7GHko+zzZ8b9OHsgxoTYbBvFz9z9zaua7HoMqxgwffx6CVpwbhoR+FJJJi5+0o5zwyCL5M0n91
wWEi4EbrgmxAACAXAFjClmLHt3XkTKqXRe7232C2ItrxngTYn233b1sa1eNWcvX1V8evGTqMkbOy
EQiFyvjDa9wtdDFOYOoZXGDvci9vHmhBLhN6dL0qS20CRxLspIt1sJVZcwRf2yR8dBbKSTn4P063
vGMuyScEblFHAjQ/vkESRvG3PE8mDmBgnemUXpqBj/bddmUe2kVTGYoTjeJiDpn8vwACYPvGBzGg
QqXzSXPYblakUs7dp46PBf1XLMTXu92fYX4UwgB1gJF/iEcu7L2lwI3hazMEgSWw8wqQTl7+uavF
CAHn2KdY2rR4snX2mVAdrT5gy8+E4/p6rzklFel59HYQbNu/ltPfmb/dCmBXjEGLA2w+JZZlz5yv
3IGGywNglbiTs5zxvIAIYvZ6tdVhgm3XQauPRn+n9SFLTPZ9+gGoX6gLv+bkUrst+uKRxG/SxWo7
wS7muojvGLm2DGR8CjKeJFWIFRS8wT16mvDxdXX3dvYHMU2JcNP/6YEfQW7zll/hkNyq4wm64D6f
LMX80X6MgD47f/hq5j38bqeIWjjnOrjOiUsENtYFxGxcfpQssIroedIdtzyrIRmnZnLDGZKhZZuO
TpcknRxFyzSwOO2k0hJ9lwzzCUkAXFA+S/Qlb/yJKe1zfQXaR08B6a0HW2PWIWGBBBxGJkd1G/dI
yELd+F/9ZJ2/jCg6HHSp7BF/hNSisco+eKg8x+/HI2Rr48R/K+Lo2zNG3r8+h9szwx4HKnFlcvQA
36KMLv7dOeAc31anG78vk+L68auak1rzq2WKwW2au1LQD9RdEP/5S4BuURcQhlboJXmu44CYY0NW
4JCc3ud6lytsaSxk7g0gfN3Jm5pwfDc0o4bcG5ebwPnslmbqROfOzOXEvTJ09yB0W2g1Yrjyfn/+
TZuOUTd3fQ3FBAqgfoKQh5CY6B4ocfwl7nx+7VMjGR5F9x47QYeLcEcDV4baOBEaXHb8Rdwec+6e
oVRqYUCMuCmA3rrsljoOgi0al3ezVxUFpbIcYYnC7cMXQuuyvql7J2vmNbnFNBQGFJY0yTHh6Q+Q
xnoALzy031VovmTN6YDGNNadG6z107uSop+xa5PzRmC3QVpxJzx6tPWEFkbEjxRGQC4XfcYSoYQu
air5mev5YpqroEr2L8kRks+zHXcAs3la/Y0chDKXUtEdjsU+nkuOZzbAQVFyq6ULJMbtuWaRtSKK
YgQZeceFB2xt1sGvqIB6vGdmjo6ZJ0KKFL84ihstjDgQ4fDjqtddkoI38DRO6iDgZHqLuu1d7/mj
zPznBYN+rzsMEUPBg/hf89TCYAPSQ+aJXQsrbaHX4V9dqZDuXKemllR1PNQwjVji4Gai6V5Rw9b8
IEkJ/wXkb2UCvvrlCSR30nlOeI3KLhptW417Ty7pv0N9GV/gxqGA7tUzInNE2ia+1y/+5S+9UOcd
S6bmiubhkK3TaeGCiMASzCJkvqmXaYxf3E/SoznYSzc7JAE83CiYnDk+GPZFS4LlvrJfqq35y6Un
ncFrJaY8gVjxZ3bUzsyWB9YhwSVgzpwH6ZUeh+pGTbCHvfPz6mpkPd+NDmXaHSY/Q5Jaf+/QzL4k
Aht2u0hpu+Zy5zqqkE1R1K7aM4k8JTUgkUJ2cQj2cRB7KtjjtvTU84W6zINfmmAo4UIM3bdiEPNH
xJM3kNdI721LhzYfpjovBhJh1+E8cWnRRIWZA98dcwracFNWTutH6/V8EuXFGLg31B//5rLpfh6M
77o2HccpHRBSC3VzUKTiMZgVSqDpakGrUV/cuLqMOuIR78r6n/UZgq4rd0SOu91xFEGywMDPwEOd
Z3Lv02+kJM870qrSHpH1tEF0c57LiiD+EXb9mGff344RwduMBgXhaD/S0Rqtjyzdz1L2BeH+MMor
KziEiDZRmLAnAZII30V3yRWMZzTzGWANbCGelfs8UXRZVyBzjRpi+zVhaMoENdsjmazPGzuBQLE4
K330vqmt6AvT0cX7gPTpEt7HsU+3EKkZ0Vb1Unv8OT39gxOxTrLjnspLLDdWsIr2QgIL953iEaKm
Z3GsUW5O/J7Vwdzk04oEHhXy2l2QTKoDJtuOpm6Yu6DZUSHFEw072dVtUdAoPxxNgAd8QCNz38lD
6s91x0LI0W/IOj4eSRBdKYie0lhe1d/mQwEvR0h2Ua/lqCOsrnGqT3oNqHcfd+t0bZtnTk1CUhZS
PJa60Tm/IE+4qLtbIxW3Ib+3ESpktY33Ck+aSXBdfswXuIT9/25qxi7Mx7TtN/xp48rOTIZrU1eb
x+PLiCAvDZb8sRh8ozRUv8lE4wtY/MeG36v9UI2Hqin0+aTm/EXt8jZNGwkUeGsgqzSUbYIIo2mD
Tn+4oP2OIQ+9rx3M4d8kRzBK2Zlvij7UYwzZvI0Pzzqq+TMyEBk08MdW6Dq3l3eJyvGe4Zbolxu6
QjXt3vORvrMwsyU1d0fQoOio0xAqTXfJRreSJBIRSmps7yTrB9o814b+erqIj8udLhgRtOHOMCjo
qwKrnKnZ503dcMhQPBIiPIngSNyCyKUDckiOpHhe1oN988XgwhQFuQiAu13EvWhHZR774wLANyg4
IHWYymWwGwRQrbkG/WtuNs16Sdwtl7mLMevtQ5UXnYC6lKlwlVwOj5vWNd6NrcCiz1PPEuk99dnG
mjP27F8afS5/U6GYXkmqgGVwENuRvUdE6N8DFsdNcG3f1X5R5GYHu2JUmpo3cSV77EBLtZXiLh4W
ueE5DxpWpvpK0y/JLZ6wx592xd/oR7yhTt+jzYf5UR+L32DeCCBc+T0bMs7kwJVTfITqgGwI0R/B
2KZLJ1+oe0CCxltB8NwetHZgLl0scTcTdAD/A4J2+9Fuc+S7NoLGc7cSM0DBHZJYt0DQ4j7+TaQl
8CqdCX93J/6JjRRWXavtQyBqPGSNFfjig4pSEt+PuQvfz8F+r+LF6q/vT+yzzZ6uU/dGwudKqUfJ
vM3ptit7TkCYNwIMvO77slrXsjUn1SuKock1bnaJ2HErV9yyOcbpbtc74AyFaOA+S2pUx694lcRZ
uMrrHws9zFR52Jo4g9hmZ4wja32vUXOnLptY7cnZxTFDZjztEYCDqjcLifPo6di+3A/NVPJDuKaS
OUJQUErLAHPLdFlquevHORUoXC5No3o+rIzCe4cuw/6Ut21ajpXTqCeHK/vohojYNnfgFXjMdHtq
3FbWbUs151VBg+A73oYbouFErzxu0PvnjoSZxGoINWfsW1GyVXWGFce1rXKE0++k6axwSdsckzTZ
jE3eH7XQKNfUQwuJYyev1+fymw1AgFfyW6oTZWONghKaQRYjuEBNoxfGwLQSWX/9EtRw/jBvBqgm
h8QusbldPSCEhOTpFJD3ouEMUd7pBauCUa5YVdbSyrx1Ii7fTMPs3BuVlNYqVpPqHuE6Vy15Twvl
hw4VBg0Zk+9Q4ciFbNosqNubuUD9U1KrhE/tJVbEBN7u/F3ATLlYIFo+1ovOfGRjUFMOCRbBvS2G
I+5/FCSisOPsQ/rss/FBCYq0rblwJNNpTIr7DwqeT/dhAr/yWBdHd5qXmiqltLCMtSzf3j/GM8lX
svvg6SRamUafg1ua4Ufr78B37sqWKx+Iw+PMei//Q03+ghXoEwun2lYXF7sFnKf2VRcd6lF48mZg
9bKty/G3msx4rAwj8E/49co9nJ5xU/1ZJzz9xOsLG2blcoe0nk3gUGxvVvj+kw4ikmJ3iE+9tOET
5iH+SluMsSBM+a+Cgegc3qlF09z71Oh+5rYowyiKPYLhquHthpZJIzlSpGGzMGKMmeKpJN+wlq99
UApm3LyZGqyc9tgx8nOYRzY492cl1xbO7LzRGNeuvCaXEcS2+poO8cfL2hSNT9FjY+76BijQlujN
Zc2r/Vs9V/XJi9bE7136Jp+N0HtwWTQBupkQ9fS3L+LeR/wueeOrXd7JU+oPO95a4uIKtK8xOqOA
FEYImpUUM4NuPKvqvYTZz4ej4DEDageO5TSVA7zci+izTTVAkyvw7+jv3HluAQp5rS7DTXWj2QTF
fpYYAfZPfu0ntQmsK5awijVEWotdvzozzwSYHBBxpbe0UwNJEPYJ7EtSX+O2ZZ378elSJDoQ5ApK
nr6dwdQgObVNvhJRsx+wO3YgD4oaJ2/daH1nWsDPQZxRNStQmb5Z6l4sk+5q7mMKUWgF7e1nu9jY
f5g/Y0m2T4RBfswqYkyONWyDYM1+imWkyPIwaSMoc25OtIWP+/VV7YwI5sCOh4yA8USP44S2HCkx
/7kosttN76OTKXHrLABNm/rNOg5dZSUlr66qjSQhZKSd/KB3n13DuEodbMhSTGtONZa7QMiR9hHA
YU32J+/b20hluTCFxK0L0jRMzsBgHr8zQByOJvHsvpJM72T+mf6wRBIwNzDSWpA3VPtnifPcR3QW
QJ1CrLSLDwc6CPbjYUT/kh1CIvwavvOEl6+Fels5LoNoU9nELI5dgW1JMkV9LDqI0kbkneg7yG/X
RwqrQi0T419cBq/fdIwebzTVI9hTsUtLPrkppBsIJTMkB8XCUXKFinTYs/cA5P/AVKI7cDFDWiIi
tHYj6Bh611cixIh4m4lkvu8H219Q52+/U5JuE9F1ZL8a5eb+02GOmux95jh8p21HCa0xEa7mnjs+
dtLDYNyepTcfP3c2qhti/epDS42ZtFy+BFErJyT6lYtFwhIMqtbe5mD0ACK3nsITdzW82TWe35kL
AHerCYCQlnF80tjwG8gKFPWbiBY+5PJSrxReSQlkQMPLTAMpypqLc/Y364Hn/3oKsgAex+4xsstM
9fd5UZKUrwB03NCq28DpF+WuvTaR20hEEfRG6OoBT+vrLFTKuzbDpWk7gGYLpev4bdtx7ljdp+MN
Rt8BeIccZe9Zo/OTYAUXZOLS+/Yo9CPEaZdp09xutKTeeWRTZqBSTgTj0GWLg8P5pK5HGefCe9VM
VRajbHMpkHavDvdk0uEIxUmKCZPnmj0dHYNAfFPtG7h5dRsqMykklJ0TaGvdlcT3N542Bf7KeG/G
xQMW5//QPfJ30Eg+At0q8bP6wx6Om7ibmQd5DMdiNsCbkoskhe3sPuMMILIqwv68ECd+AfMI6BHN
5yezTh2vPS14+wTW6uOlk79h80TNywD4MuhZL07FGfQm7+BHYZFX7vVZf1zUeRX/Mn9NoG+mGHA7
/5ANtW1Ts0xjcgrtrW7SVhq46RSIjxLF+RRFgdt10EiDwzlYnlch/jXqZJPg59495A86xEc5Yl48
6RcFnBcPo+j1HiDpJAC5R/FV3xvdxBSm2e5yGW1ORM+o1UoHucBvd05SdCc0OpUlJZL/5hkb1iaB
Irm0c32teWTAupjFvWTWR+RPSY0Prl42MG7tKXhAorje4IzjZ6IhhVDRX/S9oIVEyQOP3LOfd8OX
lq6ZH0Ay/0h/TcQE9tvSjFsuC2pc4K/tkHaIK3U/AXppvznmceN8LUHpQbkhx/8cvixzd2i7WHDY
xJD5WsbZl+0M8t1af9FPSKVZiOKKO6WiqTBVQZaB42NQLVd/fU9toQmLRN1HsHhuPFyNSob6qy7e
s+a6cScYi165WHeZ5Vy4n5o2w2R6qpSKxCRkqh2pR3lbia1xAJz2IOu0wY5MZKcLtci/Z0LMaVh6
wtIipPsG6uTTGedgICwaT6B/qrSDGLa+hEazr8ii65mtG322W+2CB4igLr7NgTP+ztZ6YLXaut+q
MKC70ibLr4W4j7vY2gg9ox8tyqy17KWQ/LBXdgVuu8gKN9Fdqqc2pI07k5R4ImGVLKmiOojrPvXT
QDsOP+w0Lfu98p3h6hG3E6pU2XCdyNRrpRW0/yZZkfz5/OxCMOChrr5JnmvfOtWM/ZWovTxuLPxi
XqCVVdYUmRoJ3IifSB5p0QpevY00Wf1F+eh85xmawCQYoVC2Jr9WiD5trKAAYaCAOouAMyoqlOSx
fpf2Az2XmngEI3c4oSj6LlEE6zOZ6JTa/0y7XSsGTvibIflDjlMs4ILgzXcKwlt79yTUTwTo0bgV
ZtjS9//CTT4KItquZyj3jl3fzq0O4ykF9LHCaVFwWp3y3RJrlamlCYt90OStX3/YHf6IQl/d0CHW
xRxH6KSgtZL2VodZ+lyXWk17olv8QJj80jS5LiHcl2eDCBQ4t0yC0QeuDC2gSybaNEuDfUIwEh47
/DcO2jSeClIM8K3+ZmudErUIxcNdOWsE8OxM83P+ZKMKxHcwCy2G/fBHl+9Xb9iMC7FkR6o399E+
tG3voW/3cGxSGiSYgmoU9ON162kjNCKZ15bxdQyhRUn6qck6AhBRVCQ9foHeLLcSPZDtH9b7WIO/
IVl/mJnFl6tv8F/XQOfZpQUVHRb/l30x3tXlF0PW+Xvsubqx4HjkeVqB+/Q/1ynx8pmm/wiudZu8
3XWSuuJmzCUlPm6yr8RdXfkh0B8LicJyIh0et95Bla37xRDQYx2B1N0nxHHl15VIVVUCr6+h6NA9
pYMM3nnISGCBzmzpJpko7un7Xdr9c2KCoIKfw0c/qPzyH0KhJdmvzEoD5Tf1HgGIKJ8338U6sA4o
vMofiP9+oSkuSQ3yP7Ma1GxecJ3VJRc0z/wCKrdU4POTxd07wf50q7wJ2fWYwsVrcLLXvetlqTYv
ZzOLytv05qu8no9mBc4Tdy6zD6GC1UvaPueMZul14JRLcS9/wADFJeWSg5eQHOQ3FIGP4X4Yr8F3
JeK99QngzVOtfBUzoZ6zzlaDEPgmMOM49chxN2yv3tjea0NV9bb82bjBuxFChCsNDM+jsp4yqUaP
ec4YSfsncFlmyWw+mAnkGj5SacAmoiDFdK203UeRXeHw63GvYBFl010TfqzINFqwmue1pYBrCYn+
nkzsc3qD1UdEUaXUmcuz/MpPSuzPXpNzKl/tbX/8u4yM3kdo05NTzTSGMVcma5/PfZVsNgjgWC5C
7RyTd1UvMGqVWoWLwfhCqoTCgJN8n41I3pxFjvsNefGVHaRKJys1rO7q06NeEvR216DcyD2Xzz/V
55wYqCk030JwyGqdQkQyTMNO3xuGrxo6cX/Z74h2EFl0UAWai57B+SOrmfGB2lQPIOCiWEUDasx2
pVx5TUSPuyrDCWGmj5zdijROXGZXppLe3nphE2S6bTiCDrO/bkxfAXKjHw0mDmJ4zgwHOFjLSf9I
xA+loGX/uTvibGcsEGaS6bHVxLtXyKF36cDUkHk3jUUwbd+4svKYX+jGJkGuviMHCHeMzaTt5sTg
KmiHYxL0KGP34eCm3PhElAF08SHx0msJ4+Uhk+cbaykq9qE566xdreSylUupqV6+VU4Xwge+FJ81
amavfI7UWUMVjKUO4sw4i2TEINvoJePK0WE9XFJkoJFpOmnzz5wqRDcK9Xdl8IfZVpe0oEDCKz73
AoQwo4qtw6ufalL/WNw6UN/uzsKJvSCaet/e3XE5zIK9x2tS0SItQmyRt4mNwbIyK8iDD+LUe7n5
jKGHrsCTKaWqimK3KvbZvxXLp8H1VMdj7z4gaKxO+VkrNcAeiFZyI1X+Ikztxq89V5MHFPX0itmV
F68ktPYOlfEDPdtl3H/ynsL93poSvW71sSg1me7rHpNNfdP4sA+nv7k0Dt0typr5+w5YieTt5IC7
tYGLz0DiTFrBSHGc0H0I3pd7TCI3JwUTz3dZyrqiuYfa4Frrp42ahaGxBZ9jOC+w2rJKBASBPsU+
Ayqwq3MoLm5blb7o/ENa8DLaj6Luh5UwBZ+JO3HeE14+JzlsZBn91l48y6uJ8tdKh/EZP+ItGcSj
rCkOxSjSJ8qjguGcU2k/EKzi/HDhtI5Vkc374egI94G9FR2NlgNmUrFmNVSOFNLXFLk7OHc8gVRc
Npw2IX9Uaa7V/IqPU2Z0PU/mrg2+rTPtAzibFVwKfXZVubeJiEYih2XTY+i2cqYPI3ZLyY/EYiwk
Oex/9Ra+BbrUGx+pPsQgyWNq0xARnsASitHiIaTApYaC24ZZ1S6zHAmjb9Ss39SxnM1wSjoxFm6z
CyBv3nVM4OFpYuuFvzl9eSjeq0pjT9svHPco/txoUXTIJTQn0clSsyLVFr/CtEIpM2fYy+r6lzMW
UIqrjbFCmqDAavMVerC5BCFLpbwi2AM1T5wZHTwM/roif4fUPZ5pOoG/yrrMFHpJoF5RB1iN4o6q
qCHoVdux+N18qaCzeKWKjnR0wNkc3IOzp3eR5vglYov+dgqOfCnvARMeVxcz+eTAmU1F3UghrdVA
uihGutyGslDiDoc+BaT/3i7XNInk6RC0wHDi/5VPNr/nFXWBQ9/4Lm3ckqxLa9z+lhScEzFXk3gf
eRSzQYvs9Bxlx6yoh4DMJRuW8FMALe2gBgWe35Q8syJAnqoum2CcN3aTYSpmGle4K3KXphg/VJZU
sYzNhJD/EaRb/J4zntaDd0gO68jnlHmMtQ2XPW3YSzz0JNQKHQuCFbHhwUS4JOkN0KgAR4JiGkRU
/6YOOFl2EdJnvYW+gPnw+xmY1TJAbXVJsY8q2j1PDT7bJ1g++mncnM2/25YYAN3Vba22NsoPnCAK
p4UJp6VIqJN4oaHxVFmZhvuUiXd7KQtlNI5Ytp4f6fXXtVac2FRdalVKYR6Xo/kbQHsxiaAgjq1d
Az4v2NDgTKN1qL/dejDQnti4rOPJqEVfC6LR1hR4qN1k2OmdSkqhoOvc8d8CfrnRB8HETai8OXQP
mVBjNkolDw23JdcWkqTgNh//9ZvXoP7ge1qaNf0YDBjqULXawIc7GZGICfbVh7XlnD/XF52ek+/N
ebtDXrtWcPqxrkw3NJG9VobmCqKg7dR4733rt5SJhk7EY9H0E+8fxNEWTNk4ZEnnMGj1aGIdNfF8
iRKLe7Y5AepZONgOdTuJaSPUmVsk91CQMqKlqkmLWsZlLgY6a54FiJy7IVJIW/ZwuLsygWPJgJFm
O2lrq8afJBwiw4ro7DmO729Xpk+86H7HMl/BlbkFJDnsvFunQMtWZaaY7yGEKNKgwG7h+727CZPR
sYmzw09gqWJRA0fcQ2nFoq8Ma1TRAOO4bY1GSLt2/VRFbs4muxLJNEYwoTgM6ccVbsDiq87cEYMo
xYF1n6n5T998WmE0H2GMpcjNUTOuR+7TXrW1Im5q8zWAhBN9GemVRWEClZlE5z8uMmIN5uPsOj1n
AKvV/ke10PZel7EmQF+hLec7CXd6w9HQnGlSDkeBFuTimcBpqLDVIEi5twBikixK7dbDM1g30Lvh
jlMQcGxg8hIqqowHZX1JyxDS4pj/UJyddB++4Sts2Rc0MI66H1tzJP/PNFSvALIhhoTTJ1nqZm1w
3PkG6+CC90L7TsQbHOahF+2O+DHc4qPlyPDLyn/KWQpHXfw3ZrCKcpyLWwPLkAP9zmcmm3DgYpTE
waSTD/F78+OmKtDIspU89udle5DKWHHo+bsIV3xvF+1cXsGsTphnvFElyK5f0m6Ko6g8XF0Q20Ow
6OECVSCWTXZNGdbFc9dUt/zjk2gbE4PGdmN6ntN3tMTg0w+vz+puJFj2+UucCZtunBfR6BSm9Ypo
n+s4OUOpZq/q2/ldWBJ3Mbsh8rdda6KS+x+w2LSJmHuiHPAcrrIUS4rVCzq7k6Imr0GJ6GhBQtnz
njO8k/j2DZv8TYGAgoKUrhUcRavVlX3NTNOwwrcBkjei52WTW7EIOU+sddq94bhH4vez3Efg8kSG
2vNCqO7bZMpMX0peujrklsy3zJyRkDiVhIxb8qysUqQct4Lc9EOJ6QS9aGuivtDghOTTZuntYVHi
bMYIC3Y3MfBBjvBwDLZcQ8FbqZSzDiQ/YFlxNhi2RQQinBF57N879yR6E3JB0rfrvnwmOPMnfZYD
jNyn/4sPzw3G816FCnB+LuppUdUmvWkFykdWTXd7w9YIiT3Yx7nDxkUeWMJSDTaqGgJguAxozaQB
/hx/a9x9qZL5eAzmUYhTNXVRESNmKBH041aqquMH4Ebi3ltegKt8SVIsL2xQiSN7sz9hFrOeMRbZ
zA06DmxHIC8tDSqiRFgawkvwTnMYlBWSRtKZRu6uhE7lEEO4BtsSpv5C82puDUTuFOnk1cSoy0r/
Qvvs4yXaQNLwu6nn2bq/g/+XAqyzEQo1xgqctqprErjaAGJCFlSIhc5z+h6iZFS+nFaFX426K4pj
yil28s5qzz/M2x6HqA1HI2aQ9OPsUtLYKtOKetPwtxyNaFDiosnjuLqWjb89mlUpmqNJYwTagSRa
bu96Cn3HxQeZZh11fJmOAjpxkbh+nBkBh9CHs6HxBPme4CxPZebwrJBYj3MGV6Un8oaqBatRTg0n
h/IPb5IYEY76+0sCu+wZENtZf2vjzvbcARSSTKDzdEX0b6sG/4aytFBW6vB4M8mbmX2bSfo2C31/
yO+ngJa/RhfYRA77+cYJDbI9RzyT6cfg6NV+vIknnd5LX86dDVxyqfi6ovurR+1OJxf0efQooijE
sceDl1GgnZLPxXv9XCG9oxqm4IscmVTYD98ZjEiIWSIN3iBPMYj+B4NVmrValfslvfDe8x8Zj1e1
r/feRGMLuwQmGKu/jhqM258Ou7xueOtH2u3eqg50bC8fQqwkeujUTUOzH6YncLl7oJWkZH+nCnuw
GncHKSR36Pimk7sUjIO1730Qj6vKabwzTHmGgdE8/d0RTYG7N1186FavykgtC7NNdrY3JDIKaN9C
3bwY663atHMpNnv5IpdvUTyxNmyA8MDEfLEJwZfrEsHFQ0Cs8HPfDmbDD601iJKIqvV7sjiK2/n1
auecq49TdSqK0gwYaAaOtmSgvfhuAM3PUJ+ED1fcuDpAbn7wXuyNRWS5pDt1JdJqvhW5KvYVwbCA
P+Tyw9rC9AP1p+JKUhknsjg7NhKvBWgic6h/0NmzkLG4zAjjbsCCibNCoqjS4Q/Wtg7U+IZFmbvO
6StuSI+NYYChGFWKX0LEBdLMYPYCj1E4S0iTePk4AV/RSJxp1oxRbBY8YZT7jjDVY1AGCvwK4FWF
gQD0hwjekLSNVjOfahyg/czeJboNCGh5lRkVbeX3ecGYiNvIxrYTZCCvv8DPHl5rJtDtUE7ngUBz
pCIrfIx4eiAHHHtbL2bOyR1KWbL11elFCBY6KBP3YjVfDskj/xI8UiiWE3ZLZbR4oAEUdSRFhiMp
SbR6DIkLHTAOZwtXMOo6gAT7yMR8HfQiIXrFJbTY0Flrg0ZuJbUj3HZNcIF7ElDNhZ492Y27HPXe
XOc1giB+fuNo086JjIHv5DthFmrdDVtHNJeC2B5tXMDRB/ZXzWAXNhC3TrT6aWlLeJQIzjTWMpXz
dRnwQbYbhZ8P0XL+c92aGeIRhM1pV/qAWS20iuFm/yGSY2smwXD7Jj7o2KG+te6MFDgL/7NYKzq5
qAQ8xgyDVuOE95gQboc1LPlqkxkBBY8NnEJN73zV84hEWddUPpXwE3N0rD3/fA/AokYqfLSC+FFj
V6fbEHlXpqE0JXSDMDhbJ4bjE7FvuaHqiGZHwQ2/P9IFQQJO5bGATaQGoDf+M4OTv0Ke3D9z2SYQ
5EL0B68keyHmehC8aqFSdlqnnDbJWgDNWEO+XCm+Kk2dqvpt8mVGmvZB8TnbJYM8FScedjRI9gDs
ttKN8P4gXZEKlWjXcR8AQrnana1T7GXVIPCz/bYKdrdg8FEE3dRQTUr5UOPu6pwJzqK2VGNhS+kN
zHuaTx4nTpChcgCsmOTWUstl/avo4iaTB94wCCyi3pp7wS9CF2uIPvvfUAPggFlpNMvak1uI3+Np
+YFrphJ8kJiNC3n+sVLdqYlX9fwSF5SUhyYiEr6FcWEoxlzdY8NeJTc5nxAMfYODfHJof2LNtxa8
Q9a0HrhoB2vKM4X68ROc3+s1/QJtEl3fJYk70ascgC/3e/p2cH3A5wVTZHkXiyCQZ0c4QWnVGsYZ
FAomrLzJeohiZ2LBSyTduxfgg4APfB+Mi20AfZjzwCquAjyoEZx80dLlxWYaQjJAHgTfQDTmoBvk
Eu5hLInZ2lxnHcnd3MtUHcwndFWYZgJtKAYQDoJ2E4qg8FxT1md8tv5W+mY6gRxZ1EET19n4G2Vl
sloCX7/UXoBsxSJzYnmNyFGL2Nv6ZlfqezIf3iCBc0kHh5DPKoSnIad1yJi3QxqpgVv4EoJ171m3
0K5dQgKcUkF1CSxKRUX+Qx5N70AJitDkTAqJGosTooJIk7lIymlNXZNrSYti43lEvwp4iZbneDkU
cQnjTyt9EKybtZJg1+yg7GP8RWhJWkBkD5uFBisfNa1dTSTexzhqgXXg0Wp1yv7lrO2fJ4J+WxW3
Xon8bmC9b/XMoYEUTR3E6FhKWlzX1Dx2tb7JlKaVdjRsfPRMiY1uvCunikzTyaLe9aRvFk8tKqP1
qItG8XUixKVJmAIAOLU5seKt1prVe8LDaZVWoIwcadpO4DS6Qrq9lSrFzC7288T5TZgkJwOvOvXh
M7e6yLGDn6IdGFktNCXyMq4rfn59Yo4aiyFCF51ogPrdzirIgwxzj9LiMS4kxAk9WBbBd7yLNdHM
XOm9sKdUYSbXzhxGtf1thPVIQWUqZj+gjWfutTApQU6Zg2miFEpO0FEOHh/MeRqdYfrEUMyTCQ6C
4nt7IiNRtVcJbV0AI09de3OwjiSchFAzh/uCPDgIxeKWQ3ZRUxl0YKVAgbm3DLxkU6UU9Gn2C6+T
3AOMBg7rZo7ECUnySSMW88dNYX0rrZAu9a+5GJVUo/hrK+Ak0UPiGZWjGgGaLqt946zJJzB4Rv+o
rpuNoP/haBYuwxblc09QEMcya4XRrNX+DqH01n5USrgUaYdJG7C66ciZldGCncItzIjCrhPtjNmQ
4bJv+uLGyG2Tr8B6vGXtxxc1SBlfCycBDpGGhE6ssU2gbXE19ESAhD1R9O54KLaGeySaWARYckII
fBr4PcNrJ3wzILlNxea5+53lqm8YF2luYAGF/MZhw0AHb0jKpqA7YXEaZ0bNt3SKzM1R2xSlzAgo
ZfF6kPrSa/p8LRelju3+a6oMWbCaAQnt9Id24ptqFq/cKQWNQ7VujpZ+IE921cwvYMMa8QzNSw8T
mvgjpE04MmDgWR4gSuGIyMn2E8d41MpVYeingAfLIwFEJz3JjqGxxQKUQ1ydUMae4UzZBnTiBuAd
Eeqye+KYo5Ubu0IrMbNPeLwQLkO9tWp5oLZ1ZUdABzQNh8bm9E5364XCLpaPsg9qQDBqqHAqYf2A
POUWqw6ixFqt10B1YhLwpOpE1/I9FdEcjO0mP4iCmbNdnK5HIYFrIz50UVTdv79oSDGELAFTYci0
xBnx6LwDbwd/EwhZL6jwjMcEqZe46MXEL1O8/RbWSBtPVFILSUmg8K4S9qK6pRU6qySlYynlC0mM
rVG8caQtTPkfcDFIwber0kchGuPayI4Pg9V6sXzlJefpsBlL96kT+T+GWysFbbtusOZSyZxqJKie
wdPT8d9AVl79zB2j1vnubToXnELLpNJgChjIZMAh/mcgZM3Bkx0ngOjswzeiLKWLWBTzb38G7g+u
TCr9dOULgrgyO0+BTX+6b4te4W17zEYf+huKeuitULOcb+KnB8vpo8N+uxrRTc6F96Js/wiFiftX
wiIECiXrTXjHoMqz1LLmBvKKVeqMdleOTq2fBiFIO6SLPkD7/CYJkAydaT93LZ5HefMPdcEchAIM
IZ+lVYojkUg5IuyoT+JaJjSw/0lBpi2mLpl4x+2wzj+XjfKstyDIXMz8ooxEZYPNcbScZ/y+/4HC
A8PBw9h5wONCzfSt40cGZ/a55B/gj6RSuCqU+df6u+Gt4SVLBmk7UEGH/EIcOcuRtdxF70+uVlQv
zyWz6xN19Z7syuClkizaMh474uZVOo8eyJGAzgV6k4u51p8OEXlUI7YCjfvn06VpgV7pKf76okXC
Lg2qK+TlLsTKhpQQoSJLuPk7v9wDJUch7XPK8uPl+aQz1Ue1vfPp1ptdt/nq4MdstQxRoJEJ+xEc
c5KQMjf7c3yi3Wvv3xfza4GDQAATR23YyUl91inWT7Suw3v7355bqUUHsNSqV9XpuuAdmv1/4kBB
zFIdPkE3zefvtVgBKGyruZn9BfNmw8bZd5vJHoXgXy4lQ8JyngK6ouoafyl8z1vnfkPC/wPFaFOO
EACgQxy9auBMxgRU1/bBV51iDj2CRtbk3X86+OHVeZDFnUtyqnbijj3URycU44tHCaoQ3yoVRP+z
t/F+3E0Re9vEQehD5SMUxLObeKpbg7f3vWAwAogrWOCOfKhk8utWF38+Dpf4zutCW+P8jhEdjure
tmtjwuxh6zi3II71I0LlUepfrQ3Mv4L3VeVHc7sVcUT5hyAQ/wRZ8BhMXAs+mTO6kTSWYe05k2NI
4+Rp8tId32yOUECUXq3XUvmWmLaEhKe/GOJCXKmFNVWutOlRiqkfaqJJpCOTsEBeiPgS7wSrcEQt
HVNB3MicZsq+AIL8Xr1LCEIJK0NSjFM9L+JIZ4cgJg6BEXLXd2L33FdZneTGW3SvuH1PowiJN2sW
VobqJbz5WtR2pKTNz5JriIDigUKx/Qey0x/Ei/apgOgj4EIEYTxJUGrnhA7rzp8NyQmg04P1dR/B
V5pFtw2gEj2x3K4Jdx8yUw7b5ULMFYVwdknPgHJe9LQ/sbkj8/vybMEj6+8jmtOJMLojD6dT1KwQ
KUOYaVKFMKtn4oYwyx27J9M4Fe+WtnbG5TyJ6IvLryd1kY90A5PdoLyncmerFytR/NkBJLjj1IK6
zFpxFJmKoeNRkmI6bDzL+qNY1D0SopkMI5Yw3K+TVOvhxYbIe5bxr0YgyhrPMe92j3qmZFAB443N
z/QiQ2L1Pwm9KBd4kds56KiTzwtJFIMJ0Aajsi19StPC8NcyXTGWpCj7xZEjKMSs4zQg4WZTzTLy
8NtKcXfpGF3fXVB/2m9uDZ1+w2oQDokjOIJBj4wU6jpnf35YHJyYEokbScnAUUNjWdzIVoCfpUYZ
5SnTBT21ZqyQlDmWJB7jAR1pGO/BuadDSTCL/tAAxNPJLa/r43M/+Jr167BmViWnMyVgzsB01Xv+
6A6SIoJtWYmCXx/korJsd8MkCipeJYjcSHQNyaA1Iv2xxeYQ3Y5GNjbW1nqVGqX87DOcWEYcGtnH
CCorT9MyEtbRc8K+7d3YtFYgTJdltxn7NI6JFd6I+Ue3j4uivuevdE2m8aBk8s8In1qq7f1B5HVF
nipkGm34eYZv33ngmK2Mt9kFoRuQZPR15JjL2hNOL8t18/z56nnjyqNfeQw2Gm0kgW4BeXKPZ4CS
7Q7gecVW4GhQb1pavncaD8MUvZ1IIumrupz6xxJoFHxAHuXDNavFKML9SJleQuOR5yLXo4j3ayc9
4rX0jD2Ua+DF+Faz0FEClX8s8mz5O6x3Lx7xZOMAx6eeypBPPH91/bJ6Y0bw+JzavvrNStZ2oslP
B8rZvSsf3GHAZn7w3b5C9uFTdHkxu35sy5E+4BLYAAMkYcZCcUwNp1CfLa93X5YwpN4Y/b1ZeSKt
OwPMExDWUdu65mhDKc3Nm7xXUBRxg27CVtUtAptIOPxk9MW+C68r/ROQ6+bwLa9OcvPLxmVtF3BL
Um8CmcWiUeSRAJbKrASvVsvjrDqDq3xBB9gAyIccsbCGbx6KbGKJC8QyyXpFbyfCivB9pllvGr02
+GQsyGP6D93yP0XtBYu5ZLdmYLwoyng1dJhgBON470YenTjfqFmf56TOPrSB/TKvJpWYlrE5ff36
TfLsmmpeXqwJ7CdeYKBZVIpXscuVSUMWGmx4ofb4vfym0+G6E751xSROiprC/PTZpZ/1nKjKGV2m
P0xMrI6yWwCDdx3irZh7DafZPzUVUQHvw/BQxXZ/X8m15/uwBJBpHeFtAVzG+iEjIxMXquRqLnkU
6HwYwj1Pn+x+JYoONz1ZljnWYafDUjGa/J7SmZx1Ssb4sC3ieKq4hD7rSHIzYvajOqOqoV2ga0bS
eeHXAsNSS7+iAfsbFM6izqkn/ucXcyh05FqYP77I/T3fXPU0wHJIWjufgNKDG8s3xqjJcFqcrTdS
COzUVeHbrTW9W4V5NX/3zdPNFeaW6rPtdgrAKHV1Er+ONYrdTcqL0VPuUyXJ5P06drQHQOoPqqQ+
0Bk5V31ylYgWPHLbKKLYBYOgI9CM3m3rcZ3Fmx9qg9HJcs7ofnMJOeU4SeHh0+Gtw7D5O8C7Br59
0wVmw4SI2pHqlgHEm4qCypJmOKhC60eyqX3fN/0ZqF2pYmwp4iFu2/IHjX2ZGKpSK0R5kaer27i9
982ambhCgFRcEJ+DuhHQk2xkB8SRDPWmH63chi4V/lvj0axebCMOlWiKY2TeadvRIpk9XYtebq2c
BUGKt5eQpKj7VHSPdt/T0T/hdQGdGlY1nTKXGZodKhp3sEmxRnbSdJpyXJGE9OtLRshTxUdKg+w7
8N4KHToTrPVeIBOUojfPq4aPprGGnjVWASggZ/BPc5gwMhZ94aV7G+ncNDyW9rrsLcj+h2CzAJwR
3jsIfoyC3pXrqapzWTp/1e853Ud+ykABowdXG7FOBiP84racpg843jKShtBWLWpLOsUTnKrac1rD
YDazlwuP3ywh0o7uJcBXzYRGyx+uU6/B9aVH6pec2HWBbTavZ9hbR41mx+R990+vaCE/3Cra6bYC
1945tCTIVMN+8qbclfq85MJA5l4adZPZ2PNToRqYOFH1gfhbuC0K1cak9maEANODHOHVsbfA0RaC
TWKtZBURfZvPGg+J4iP6+gQ7nCGuYrvPsMWeoPu/lPkO3a96XOQH4KWwVpsXLuR/5ZJjUSne5Inz
x80ya4RzT7Vdl9f7EHFiQOVCVOF2Gd+RwgBNfA1VNY32ebhFtNJjo9bNjzsrJEhgwMCiur9gaaiF
aQJwyRvCe6HNLECHE1pGqXYrcHNmzIS3gQtprXX/TjOh48cV02JUwst3hBpZ4DLdhaZNzxC474Wz
G5L1nf1uIb7mtcZhFV/Wt7k4FVUd6GS6u9GFn+OTW4Nbsqij0kmFT2V56kHapvdOTOxW2xCZii+X
5TPoLpKzlrg9IZCBtR9LXuD1rKF+axLw+vau1PA9CQY3lWNSxQQWvDqU2QCroD1g3QzIQ0K9CJnd
h/2R3PfsHBLWQ+3NjJwmIz/xugPQcQ+Ikyyi1gZzX0uyM9J1VTUIybpSKx0sVyrbxvtrsDHAS5F8
yIH58IESQ9U2R6VgkJj/gP6JFyUqT5kxgJ/ItPe4Kk7cvPL5bvbHnAjurApWQ00/dRg/2o+17rgh
CnOjGYWa4P5gWI/3CaAT0r9rxIL4+8KnCmCf/fV2dUEGGjHIpoOCEB453BXdUIXT5JN2TKxGLagC
vqVvPjH8Q6fQW/F4ttN2Z6cXFhV3+cxhiGqdfQ8KaLfuRZ5fxKaQU7ZjtlgG4g4JiDTqGbifgB+D
ikUcZyZ5UNy55yzgvc2W5LOF1kstXxoGImU1Tm2p0L/Y5WrEFkNy4m1EawTx2bmzqFxfBCfGOWYG
X2vFLVi21F8J4B+U3m584n9iLt5XjTFMyu8SRh7MImsJo79af71Z2jIxCZTQdBAtRWEFEtvbkdSX
yv3WhaRVsj1vldkfQm5ebOKK1ASs9Syq4UewORmp+lHS/ItJ5c8WB4xAeC7QrWTb73IiAwOMIDpg
i6FMYj8/2TDfAuMWMWcHa2pcByqu2//VIsFFYZtOj9sn6sy0EaE77Y2uBbUqUTSJH6sQxwgayf3t
t1J00tINdQzfIC6Fmpdjx0mP9yQgHp278FkqEwG8HLnmo5wl4T5XvgqS4FE88Hsh/rP4P/jwNdbQ
hMm0ie/dV17ucJqSu2j7e9wQL9RlormjvAzCVWWwmtX92xD7udrM82+/huOztP05hCXB14KLlA50
1dCCg5yiPsa7XfNkjtIVN2SIf8LNg8TnM1hLRP2ZlVcAHvIuv9UsxV/us90GdHPp11uiz49vRh3/
stwaJu5smGTgwJWrotQPiqM6ZG1KX8GE8zNFoY/Tvbz1qhFo/CcUSzt3CcDga36cFSlS9uzvL79h
yZSSJVLGZn3uOEVaQeBI/Dj7zSU/K1rvAlwepsRI39ExbgpThdhcUHMnZA8gb0SQ3edx8XsRMKDv
OelW44b1vl9i6kp+zgxxsE+fKQO6fPerlFRnNXTIBtB9h0lshFC97fdHCAHNmui+c6SORvE4NHJy
B/lXqM/pRn5iStw8YiNV9pTHNEFSMigW06WsJacnd0flCY2MDGTekzd6PgwCvhZq35OipepcI2Ni
fZ0z/a/jrWEPibBNQYLqaE4iXmNQm9gL/oreSGGRmdXHPGqSglz2L8bDeGgpdOCGIxUik0wYiKKF
B5v1G96ZLlKz0ioccXMuPCzlUNOc0U9fNpYmXJddSIkr2rv0VX5thgEMios0PNaax2by9rj7q/ic
a6klRWYoC79ko6NQEcyqia9WgRJk4oEiVZCuNxblbFrJeaq3SLxcXxnq1a44QmRvUAMssZ+NJvcO
GmI1/IW2zHcSnDkRzyICMkQoq5Vpa+khz6e2DB66FqKVhp+EEkdsZ6oMgggAAfj0WEvb/szcjWj1
HgCNIXiGOSYnXi00SuMtxIOlS1AQPhhpT+reoVEUtEY3XJNGtxiGlpjthAgNrJwdo1FxNfnqsIPZ
1ix9CGURS2IG7QHMp0mXmrRpph1e7HOCuR6WXWbrpSXJyT63jR6IjV9ZuEq20Dcewh/2qnhcB7CM
3dZn/GScHvYYTw6QXgxQjfOVRWXE8jjfStuh23pBbcodId4lhhWsTNp7ayF+CltXmm5Qy/LEbYyv
sFgggi0xO43TRc62kX9c3SmGQiNxNvXjMUsvnsSRsW8XILLahJmkWb2jz0tbiWI51HB2GBMVncfl
TvgKAgl/WsGqZxNNn1r4xWWYQa+OUKeWB/qr0zAsfijYLj/NpJBDzCFAMlZIUahg9aCdErs3qttb
Ib/ykgh/XHE5JOS935u/rfR2xPq8qrLK0Mpx19q1t9mUJuFR4Z9nV7WlJu8NbMCXioJcFkrC66sd
SLXfwnNWnwK16h4pMbCT3NHmucTiicwbDSQx53j8aijUqMfghSb0GqiXMkxJwbR1t9DjB0Bv3lfw
jyzjcrGfKsEEv2AsRLKFJMW2rd+R9UUTxi0VZ/1FlMHd1TpY+1vJveseLxlQoOwnhYVLpby3pnRI
+v3Ltp9XQLV8CtM4QgUtq9XDEgMjcT/NXdDaevMCk5QPR3/5pu66g3kViZrBN4clEVICQZJW2XnE
u7YzeevXZdczAryqdayF1l9YSqd/0/2lDxu4i1MrjFmRl9jGQHLk1i+/QudV+wpiIIV2K17yt3tP
mCo65RsDMxcIjhWBFpz2tG4Z9O10MH+iszcLePhamwtRZHNVHUZs5zT/oVtNAz7S7kAXK9BJStR2
Jcl7I36gm83DhIbVifhOV38blBvQh63Adm011GovCnoMDEO3qCLIE2XAQFUWVzivAaLElpbkQVRV
FChX1KaVsDjKFi3QJmhu9fy61msa6Vmy7VMM3MYDTkteYTeDBlTxGMvyIYvX/PYSQbuifh5sgRUl
M9rrGWAESwfzQqhDPyrt7LidIKKiKy6I0YIB7iNBldOh6h/QcMuwhlaQg8yt7kEwjm3fuSYsoCpA
BRCmpy+mQW2PAJlkVpLgr1wN8tZ/p66lFre0zzeBYjcC0tGDu3P564ztASw7fsVZYmRPJRMkk8by
QlJ1UQ69pqjmAfmKVsuXvcCeBErEYFxOT28wHCPEqd2NfkyMP+K0IyTmntoMIY8voHgxetgseOOc
Ewzg9rNI1p8n8oesi9HiSw1tlrjtMqWDeHTYBE1yVkxCEap6oC6uB89ZN1Oz+GdD8vSPMXGSH/n0
JcvP/CDiu8F9ThhFfc+LQda7OWsgguzauCW9Wm1APCg/I3vx/d0w6mJDZ2AYraBapm6LVU/4bfWN
bnRMFIt8eu7Ihi/mWiFvIeOTTRV1l4eQYJlex106GwBjMnR7X2nGtF8OAfGgLnPEGPAxnr0FdlSx
mDigoqu7FTrLIa8ZdjxRqJb9PzK1FAUhR7AEFIT7j2Cxh2+dMvyiABQeTl9SQvgYrDRV+pe4vloO
TKS+VUeny4k79cVX2s1FgQxqgyv/FQXZ3D/89n/+pXHuAwcxbJiN0Id/BKejVUsPGs9Zed7xrvX2
nBaGwR2rTPI+SPoU8zRZStuXNuBW4aJ2BtMY4BjWzb3xCpBGqQlu26q+uUAy8ad3vO/8WDskUT4g
Eyo/iVF+TRiJjC6kfWYxcqZEGsnTvNepMBCL1kmlFNali5YBmfWQxJbQy/VJr6saKz8jMB9IvA+y
hcXJ5UvrdtzY0PhPzWuOViiJalJqC+S5UD4l/kxCWVCKHY0UUpa+gMrSECMjqgEV5t0vcKSNYUux
k4Bi3xCv4V4bgtlJZp3iudKeCfhOSrjBIuWlvZobL3yUq6tUVRT7k63rwqzjF1WnHdAbpUvIMD3T
Jd8hoK50NbMtQ0D8kk+XSKUVAgtYE8C8bSzOsrlFtGYGm8W3lTQpWkTNaK7IeastyFQx2ZD0tNeC
hb+0B8vHe6lyik75f3nSFyRWFXR8qSreDztgnotEi5IDcOGXOGXQmafVrX8QGZyubuqoTUz7byFw
EGk2rpiNxFc+hqAe10AfL5i5DYvvIBmnf+Xjt+XLscx8+zZf+eqcB2R8Hr1oUzSFlzraDIF+F5CS
aGkBm35S/h6bFkggPeZ7g3TA0zTnQ55Pgw7luPL9mN1N0j3UJRyYh/jMD8SQ18oi2F9qKLcWL7xv
mOnMGKJtgQKB5p1ZrJn08vIN9do8+ZCUUHPVPn3b+y3O98bgOCqbAJ5XOWSiJpJGbTKbf9ynQUAe
BK0cZn/9uLtzPhnSUbGvfVwcQ3c0gKwxQl7PR84181PUyXlD6JqrI+MrCCWvmCEWISNG8WwIaCPs
joFTJHKXCBqjYSd849MAP6tl6vtM9WkFFx0FvF0ywX0lgLd3z/jHjqe0x2iSK86OxHMGc59wWPcL
FOHrlBY+h1TDw8E9HzEAhu3bJFmk1Y5e4nTKwsV2SqZ5HbAwod0pRsJPfw3d0CYpOHFDg/CdRy3d
gqZsJSksKoCNHQyVgl8GIEUun36boaTCYwtt5n3wkJMErp11ZOVNoLjIHT6D1HIjB9uiH5tohgSf
9ik7Unp2EeOJX62YV01Bh1v04SC8xMzp5smfAn/UAOGBRPlZG8RV1ip4jqb9aB94/Yp73RYgBAd6
Jf6euZranvgARcraEe+l7sh3BVLVwbEM4iC3XumsFdtAfiuwAfDtbhuD8KTeAH1OR+uTxXs5jCyH
77Hs8cj6TmSyf92azywrBwp7shooUkY3a0Asjqwo6GRZyfljV+D16UtP7SnS+ROE22pLZ/53CBA8
j1YmXo2+SAghZViskyJaEUVXdmM0t4rtmcLiHPpRhTzx8j0u291AMHUhfy65Y49GtOYHjDSMmMyl
WLs6gFmp/w7z4ukrj4VhQO02Eak0EbRh2v62dqmMpZcP5oL+s1iSvjwgSAgNOKq+AQ4mxleA4kYF
0Zg0HQEKU9FQVBX8KRCXYFCTJzCoD4fKhvLzL8kSMvvF2wg4a2Nd80IuFtCsY7Y8oojZJGe6y8PU
/FEUstvz104l+C8Qnxjq53+CnjZOhkmyHgoGS4ONz+gk4ncISFuHBbcp9KhWXWNcJSyvGqdxfg5+
ivUYuaaImjYgW2vuOE9+c28wGZY4xl74cssFnmmjedsKoSkfUKUdjAirsApC3+pgOvhOjmMGZdjN
WE995yLGpEx3HxV/7F4PBzjKsx4Tztx7vtLTxChEFf4exl6QTa2jWC2ewERp1nsis5he/Ec7tIiS
1mpiJaA4CFAhvwh12+mv333zHGU72bJSau/JgYXxwFAHeXnnDK8KXQo/YPsb+nNcpLKPBtmjJVZc
uXWEOTJ8YUNBur3HE2Xt7vmDlbZD6zaH9HveWR0k+3DbZhJ0NbKCJj/HMIw2oG/iAiHZrrgO8pOF
8oaCypvMZhNwU6SKx2hUnhE2AoOIQzY2jVIiff4Xu/5YVONb6qe9WWxNzbQWeK0OdIN/UvFHo4DE
z1fesmPWVVhe77fm4SdYO5p8bNvPiYSl0tAzHAhRpZxsK6AC2i/JM298LiZ4vXIgcW0MlgidmyHv
EuAboanJuNneW/4bqdpLfJ84lx5rDMLUCFKmZguLA9LWwh/rQ7MyWqIYIQeg+TQZFP1ryv7fYxUw
4Wmqz3PZpR/NRdG3XtvIf7a0mTuJfeRCxzhrxqagBB8ITSQWvVJpSuzusP4O3wrDolX0mEPmCXdQ
TWBo0/J+DsEfp+hKBMGb619+9LZhEnXmjNnDQRbqTqzV1SY7xrvCnct8Qa6sO1YFb8MgQCFhy8Dv
nmZzvgHsuOTQIfhgkslwBLa4hXc70EmLtmUdcqh8Pn01/wvealKRPa+R2pBGIxlehZ+csKXA4V1h
VFGzfDXZh7KKs2N17JvXPu5IwABXSeFxGyUQCKhz69aaO8UBNCI0ls4sR/qXB6oYkjRrMzwPZ1os
ReqBbeGhQO0dJmo1HZ2doXSJlSH4d6IGe7nKyKPfGmQKAwDVpe/AC+tZpCOj8MMjTqceESaV4Njo
k1iXKosMjnpNLR9dY2Hu/oAq9Nx8xp9EQtLiVRWbHTI+unVXscoQq2oiAQa+8QCp2/R7nOb+ipmF
Ms5ITYePi+oyA8LJcB2sfk2xSRwm8YBiLnd6iA6ZP7Fk3Xl/ipKBWCAnbNaGk/9ahtWVX3Kw5LaY
6zd0PRkAI2Le/jLwWSMM99+TG8H/vku+ZEtj2rh3QzhO7VZRlH/vq69Knvi3giVP1XSKtO+/FFE8
2jlP1QVRZwuTwiVxhFTvbLC35kjAzyviCpHdVEiVFfZHmy8iAcWmp9YEPbIILd4E+MH/JYlsx5OK
CqioGA4CdLsnRwueVYQac4TIxcPPKOjQ0KJfIAYvpohMUN0lzNUrugw6SvS7aYEEAa9P3ZBvk74F
KBZQ9uWefp6VI/FTK/YLgPuUNjkD11OMtel4QLxdgO4PBQcYCI73rKbmNLar58An2BXP/lukJAUF
1SEVUW9kPQBUd8YkrktaQZIfx7I1bHzLyqYwHjGribmRItoBMzNSWLFNDw+JvriCIXCZUWiKZS9b
bQ64pZ0EHRSHLNvdOPHrXv3rTC0Q1Yk0AeX8WsJlWdG3lQnw/l2sIB2NZb6g3tVLs0Le78g7AZjW
2Wx76jvkATmbgBw7hvYLmY425BR7FvNIbo0jtQa+6PHG+lFSxN9PQoYKrnvEKX4pW0QXWZl2H5Mk
SNZgAoeNlDenxS2hxjCZ/h3C2R4GjG+/4Gs7WzK17/Zx104Bqe8YSb2Gd1CZuSmRCmFq7bAxdego
bHnB3dZWVFoYTKGu2gKsEvEkczEj/YmqOz3N7oVnHZHXpwCSum5ryUcu/PeLClbkQaNto04yBdaE
EqOLoWZZWuCJAvHx8wPoYGrul4mdHQFKo3H6cSgGDPDtwWDNzDDLyuIjuQ+oCH2gSLZqK1IEB1W2
wQMbI+5fiYkn8qutrjqSGULCCgvax96jjUhc8Q+LAf7Tdqi/I+AhN7jGrXkLYwyexef6pzmq4y59
2CWpS1GRyueaCg5dUEOb/NVYg/Opi3z+JAMgbmmhG0BLnQ4yDNAxtXPUgskGumjPt35DDEgN+H74
tcf9vN7GlUJ4YvcJt+/OziljcXeFxPtpqQzOLIsMl3jM0r976giQk1CVQpSIA7vrgauZRu2fw09+
9TkKQmh5/bJBsL/slrf6qu7y5Cj40ECTJdPCG/bSb3It1uvpLGkmgQCa8HY3JS1rvE7xboNdL06a
gXDSZcC6bqEkLZE149zL/qxoMt3DfuQrrJKSzHv4py+UeHm1uZYzi/QN7QfwuTGcfgm0C1V8xzoC
6LFEvvdThOHjt46PcYIqb6vvfP8bSEBDxRjcHbliXLiH7RnC7cS6mC+kN80F+4KuQWdW2wkvsROK
UQ5bmYwmyjaqsUFp6Uamxe/YYGcGhwBpGgDmLyWtGeOE1Zx64NTmsYTzVgByy5asORH5oLHz7V8C
NWZUuLeX8CoNpLor29ApAnCsRn9Xx1eiQJrYYIMLthBiwRjesRzS6S+intauTVnVDEv/NiJV5ifD
YKR76fiDGQpWgscurUPXrJN+QCf6CmkP+M80B3YKDYwFrHxW/kKr9ak0sWkIYC7Y6Xsys2rqFlx+
A9982DlgTvFa68BuWfnpJH4YYtqAPdvNtqIpZAxau0WE8SY+NdIklw0h6+FxLwHpbsA4qJKHQGZn
0MCCspL9ZVFJeFNrnqPI/lbz5GQXEczY3TkNw66lbT78iFiB09dC8+zjjCkBI+F13PezMQ3aommC
MUcIeoGABZxUzUZzka34O4j6luaBmwekcBgCJp7uh7lqh8m8yzK539y+8mQI+7glnq42aLKKCjY/
Aznd1BqlgRl51LXDD68NfF0RHc6QgK05jFBDTZ0pAOAEu8PgBm89jqhXwCnZQWjMMp58DVHcq9my
x2OPOU9h3UaiCO9hSl5t2xYtHd/X10z1ZX8hcdPp/sfwNWCuxqdMd26yhu+RmS27E3aSV/uWMZGK
SLno/QlkTUNsYVMlY/26mMm2JJemC6J+m9YGFkl6+tyS4UUc7mXQyS4ZB7RwnIm2Sm6FNZqLYU06
PFdR1KfAr6TrhUEJBXRCPokbkYp8YF0rAjennWKlP4KHMsM+E91760GzNLNRR8wQ6ABEy8s/91IH
xz52wHwocc4Li+lOSO0TGbXMRjfoocKmogw/E4gqXqKCKHOQE+7n8a6rBgWk5HJCUf8VocVN/8YD
/4dw9yMtYhoCutTE1wYSWV/3K2XSroxCBQi7Je7uHBl0TU7KBR0p4ypvrj7KHMlnxI9Q8Z8BsFbn
nD6AWCpWTh29PaMnjvaORhhjK8G5Z2GfzH9AOsDkrnawdI5s7OmWa3348mwU5GFFJVy4PHGBoVho
ptfZgngLoKKK+aAmzgnVikVzLEDqhU5FqrB4Fzgwlz+PWgkL74lNclPDFNjevH50MOBtFsmIiPS2
VoFvRa0BZoIVjNNU9zYwHMApORzc6dS+04cJov3IJuSz4FFIlcU+wU2jvjRqsvFrW0fKFX1x31LD
Aa06fl/TwSxHpWHtNsz3brhJC2KeFZ6jZJqxrl0EfIfqT2Z+r+pzm5TqZheB/4zNw/sQ0agbvUP0
2xv3vgbD72B74MSGZ5PgduaPATRTdFlVVp6nuap6+oe2kEEdqv3W0JJeqUbyJuWUS390OqX2z6FO
h9haHxvATQs20BrfD0vt+yuAPPrCzIefEU/dMxtF0+1O8h/uz7nRWtGI91EBXxoGNprke/WHQ6CO
OHzH3m61hsSHKReO0Wfsr5tAk4qrOENhzy5qbeugSP0jXpQTkWbnfzFJRaGvliO4nfPYiinJarXi
et5dZ6cNcVxnR/wXD3XrEBB27gWp/XSYfF3DbsOuB5cWdRBPEmrcpARZOSVqNtA6TR9lG0lYqL9d
2m/ZA3v93v/YxsPjrjTxhndPxAiT+6DtwLz9HsJqZl0cqHG0jPW3XW4mnisBv+GgAFyCSZt/ntCF
1lm1XL1jcNJsHTObti7dnyXL5eVMM/0VPIZJLT0VSVY6di3mAt07AYrkBUIY9nedzC6IY1q99IXK
Ekyg0g2UnsW8S3Wl0SW8mSfkt4y9bvdW0bSoSr02kJJ/N1SO/L1AOZrhN2VOPwIuHqsGkpfI9CPs
V67YfyEYGeNNQsF2QWVsVdTwxhTciqCeAe6xqOQZLAnAEJbQxXLrvUNViDFSM2VLgfdPmIW4pEIE
Udkw1T26kv9WqKhEDctw3GrTHui93nHWN7+6SxmgC1Lgz7ONHQVNFnARX18df8MJ2UXMeAWrKVZP
cwn8YnrXm1mqfNCvODao1Mz+l2T8bMaf62TOX5B5HHrwR8auZUyfQTLGyzl0wZM9Of+r0ABUElqL
JPJpmS2aW5trg0RFgabRWUdyJSKaoIZzYtN0sErdfdQkM+x8zetCqhpM8BdjTnmfyZ/7NJIRJnUJ
4INyjAQ3zlMA7jyD6YIaNYGGipxTx7+ZNQiVC/1QMIZB7Ev+v9GpgOMhcttIGnZjPIV4N9qLl4Db
lW/X+1RzpNLMVqpjdT9R1Eue3yZQoADfrSkjbvUTbB36o7O840JFBAdNty9QH1C/JRyvrLpkhy08
pBgyfpD8Sq1oP0jrmp7jAHaB15oTyn6XwBK6kW17VO8//3muirgThhm9Pzy7h8GNRhSnvWE93LA1
knskb2FM4w/2hspFHQZc9PiJifNI7cJ5Y1ukYYsx1Vp9aPwnfqna5zQmMFDEKhBk42MyKABWWFpK
4U/ERT3Cv/xZv+XtTcO/hqoloD/exwVCybFI0zwJxS4bKgK/eCPwbcENgl9SghuZsxoh+V8e1ZhI
gPlN2PhGJvZmQudz0BnUNpcn6pGQ/aoDqpsXxeHyU/GOfCd79RnkoC7WqxMUPNANPMFM04N1V26a
4kjMaGriA9LKORh1cmPEOlUpLKscWh8tl2hZtoIOwI+10JibkUCLLKRl0YxC6w1LPVV0PE5y8uc2
WuLdUkhIIBjnUsswS7hV4tMws2FYbdaYjtYjePGfrP6VfPa6EjTRYwPHu71IrPYP9qJj2oU8gHZn
+40nPzeVyXSDQhVWqZPUQKN+UcgbtA6FEFLZgSjCP37ZJXaXduKIrRZxJjFTV1LwBkotp5uamwxV
lJZABI5XXp9aoA8KXN6U9IPyOgwp+OnZ7fHUAIlhq5lwHPokC8D50UYtkq+WOrqFxxhUyClNpp5A
2hIU1JzYzvw8abZJRxlY4lbehhj7d1sI6hFPO/ppd+vwod7+OJu5kd45+C34RD6gxoHDyWhKOAIt
Of7BxsFafcUvlL5M12437MA1d25BM3Mrx7GyXOuo+Ax0eCzqj/LDfO3yqhUWMdc60iJMIvrbDItt
KDlpzODZsfa4B5OOUiNfyHHoLNDZvXLL6bOGLDGVpfL6mDVOygjTQbMtiaTLY5yYyBJIg+b5SM20
N5A24bQRUv8JFfzGUpow1a7ugBhjyRNGZrrQXwDCs0kennl7LpdSnOnPxmC5ompR/lCXmmHo/uqj
YD6DTKWX3Mh2rl9iVbstw0NXqmdsZ/U40C20t+nj3pU0fS1lRM0l1EpLS5PU0y6S8yJOn/XtPuZU
XyGG2ruALEuL6iwmlQuk+/BjWaIqlLPoWe4U2xL9Q30SowqjUIOotfuxLHjxRXKuiTQlOjNRD+v6
EMwfeAdVE7DTeme0/mnXdH4KtAqrq0d9FQyoP2crosrBG4izVKO07p1dpiv4JhUS1PzJF7vJyCA8
pLb9iwhcW3gGrkGs+JUAipI7Uy80ix94OQFB1PjE3GanHHzcF+LlY8RUhWlWY/wvWlwdP8+7VFzv
EUVDFXkScndlK0mqJZm9/ehBXUbyDTaMDVXrzPio/bTjCMFeLUpnKCCEyU7K1TDBJaexZ2JfDrz+
Br8MbUzdv6Ha1gz5QNQ0Dd/r7VmtE9gZig9PrF81mU0SVIHN5diEQvKUiZn8ZGrfCN3x9yofIp53
0LKH5qu22G82j1lGoH/mTX0NHjArSUf4vo5cotXPxa3dBUBA72W7hFgeAJufmCmBwTjmhikJ+hld
xHUW+/WIbnrQD/Uyjtv5QOtlxu5xL6ewfp6TMl2zmnZ5C4kF6prO8M2HFunVobU4Q7AM6MfToxtT
JUmJVU5kPg4dF5RMpnrRjr9sOFbx2yX5hgtewFQ6zE+bqPXbh1KFDcFXDVaLriqXOiJQetNfK/hp
SX339Bh/Vui3HQjudSeeKfH3YIcqovr7vLH4j8q+L3ZNHExcyNMQev1911t59bcF42GawUxgKUl3
miHZcvcMTSmJ4NuXm8blRnsYN0iCOTxlA+woBIPnHasXPPyViYLwF1MK2xTXjbw4v0iWNyvBE/Cj
iSHqt2rt0/z1fO6hXL7QmG6LsjrJdX8bgRpXOBjstglT1Hh8dJ9lsw+te2hgkSoTGTH5SnNmj/NW
lDDdOst00ETfQxSgsbCeAK/+2NgnPiMFOejwD7M1WJBuq9oeokJPl//FXKTHmlfJ1Fmam8isqJBO
eblJ9n57HZ8rINEm6vPB1ydn0O5xGJRnGNiELnh9hUUNarHTs/MJJx9CrpTxihiw7ogTv3SuqTRE
ZPpqtlKryV0TDq6iQHz4XpOMNQOb07UsRV2+dF46KuDNpVdfL7iZuVkpLfw+FEI4EGzn7RE7jrAl
7YzcQ7jnW2/Hdwwn3z/AexEFEpD0dlQbDeETiLJCmI9pnGFjqHkdOw1zEJYu5WbIyi2zfgkAB7tD
oYrhkm9Cjv8mX5ye6a+HqNWP/3RYbq6T352NrttMcUKojkaCZr8W6mNCUcryL6z3w420WxQzfSvx
PkO9++Y2SzkugaPv6Y/n74zTkfRWcTtEQaHc8v9WvMVMgnC5574/ccYYP6wCFvJxQ1YLWtKt50c9
vt564zaZ99wEuRYL/FKa5aEnDXrCaw9IQP3bL8n0oNOrj5yPRcoI0uSqIghwZXrlRCRGzpuWrIZg
zZ0bGH3d2TCzpgyplVLsneHop/yalaf4K1YzSSRczFrKs26G2DMwRDC6u0iO53egS/D4D/pnPJzV
cXx9urnWrUiyY+CBQGuhxxSBIdhFYIFP1VWQhVRSfVKdhxuChDWNSevPTsc+hY7KVH7dTfZ5GkxF
cZ3SoJnwsG/njlC2pkAQC9YuwmftO1zrw/4BlMJeTRDOKGKUj6WfihKm5yz9GPG18BzdNoFplsIc
I8y+eGqDFBhOvpHdQCCZ+ZvsfyVP6QdMSln7XWi7GFKVW4eVsoD7hLqeYXanU94M5BGLYTgjWGk1
w7OE9HfKFETY7HkYptwPCp8LXrqtUeKM4pJMJmyVCJc10Z/9Y60c37q6q/+bm5CfdK2yTdiEMODW
7pIaNZRw3nYW4thueco/DxKLVDBW8hcrUwIXn5iToqDcVYJKmYSz/HupsHjf8xZSG/+zknupbSKQ
8SpyG31oHDRkHPm4Wlp5ZVvEamfzG1twgRWLxUEanNCZktXC+aeRVKfwiF1AOrE4RhQhNpZQc0e3
5FwOoar0CaYgtONcX9LbIwQqm29le5v2IrkFlnKa7exRZe+sncX8MmfPwFdEhp9PCG3zdsN6styT
lXDgWgM+bQ92TtwmSG5lkG3Xei5JTdpL//MuqdxkYmn1kFODK3SZjPxTELSpcTcRA9Vzgfkcaggj
1gJ3faLV4AI3DmDH8YREH1Nmyr/DTdiVmbV+OWaxRRIYI9ScLDPcdS7fSfvpXcgp4Gb9NW8mtk6e
wJCcSyEDl8sdE3SAltrvF/C01F668jsxXY5xjRTAtCMkls/8Jj4T5WWQGSMVSJx3+jSQ0z4qRqGn
eEBzDNPCb0XVns6hRWIffg14qE0lWuqW1mwsNcaLYKsuFfZWot10OK6ViZV5NLMmnM733/0dvOrQ
MHC9Anb4APeS1o/mDQn3YO+gXLsCa0yeK84oCQ/V2QcT3feVhHyCTdsxcji7oBFoTAkPR5BlA+me
OH1y9+5wMPE/3wQ0mY5TI1yh9EHCM3uYteyy9m1YPFoj9PvHkagqNNN4xIKyxaQL3i0Q1gDccBXh
dJ4yp0ax/S/m2EpS+/7GPTCx9hYV7KPKU2Y0hNY/a9XLjkkdUjDW2Jgf23aNcb0UHAxdc1iyO960
peo7PbgPJMOGYGF1Gxli14kgJahNydk+SHMWpDqmT/XaSLR2j3V6jet8tX+X00T6yY8ywXWaG0+9
K7JR0XraIrXeEAyzEld6/IT2m12tR9Z0VHsTClHdkvC2ac9qbZrOAejH/us+FMsnFfcLyocHIaBZ
hjzjlNpFOKGOTdb0BKcaBdZFIP4NJ035bfQ8HwW7GySzuS1Imsj0Bdh1rbk4esUa/GzYqPclm6TV
NrIk4Jx2tkCFM+q+n0d9SJd4vrWFfuSQnEIIe5zKqvsoQ2aRyY39T4J94VxP8mo2xy6jKojqq5iJ
OszBFUZrqihGYOMQjRIZvLk+wQ0YByOtIqmjjaWfmCBRAX0nnuvtEMHiJ3z3Kj0WSwYAS7JTwZZH
DQtXXI/gVTBn6Y6kr8+YUXrCEoB96MdFdaxxaFMPzVzegJqYHGwnhYUDJwRcps+weHDmCuHiFeeQ
IiMClxJVqCK9UdrDzycznqJwFROL21N2mn3BcZm5RAMRr8jlcEZCA21gSfefuN1aow1pb77jC+n2
AI1t++h0vOOGws4rmkC37IoD1ioRFVOFru+7atMd7aCXjct4ry39wKmXZJvFyTmnWfd5/kfTzjIb
0JZlJssfON8Vh9K+N6o68wAM51TIu78PhZ3RvpVqqw5twu2w5amydopf2XuQQG9V/dq9ib99H+Sv
wX6YJ2/pc/JrBQqB7hOMiRTy3NPrMcOIDNvGJtpCoYDjhbO/ko7IErHoki2qDVIgtgcN2vSD7zgG
eW/fwG5WPa6AYV/XN5wOAQ6apVcM9B85hU+4m9ueXZqF8iwKgwLKCL8SlSZ2+2Wf47qzBSK829SC
yo8Kv4VDGiuNnXx8kbdHz7LJoLOTEFnLTDtsp3tGxSm94jg5ZBWYDQwFGMiEA8PKbCY6sBcttc1q
0AhLHPXQ/sbhuu6Dvq9LZeSjexDnRrDZjmAYBR0a27qIu20FQ8WHGiDUaXhkpO7QeFnZmXC2tugI
9X2MoG36d0dVi7Hmd3x5K7bBCSBH6FDwLduZ2m325QOIjnhgMVbY2pmTGEj4ZVPn80uYhzHBEtdo
BYgLJlR165L4Xw3ao01hN9ryu+Y5Oqju0JOU/tME1ddVD73VYjAn6vAO0C05Npp5IhBYREDv+hsx
EhDKhMhGweWB6UaHutcP1ng99G/BxFoX9IMrT+oUm4gUjlhAaKwv/9aK8lDuQUjFLJw4nhtbEo28
XCEp/XupZTKbxvH2+1qnrIVxovklwFdTCr0ty2Tdh8az1jtqkW9H6mfgz3qAHGUJSElEtWwyKDyM
nJIKMm2Nd0Eg4ndlLmsDUK+RsgxEiM6lAjpfhCCz5UOi/ULmD4+FWZ+82tykcJRcPJ7wHEYJSk+U
du1bxlSWIDx7AwutUkx8LRPMxm/00kN8m1gc0+kguWTHUmk2s0YabeQLhpM2Ocp5vHE7ZXOuQot7
oFgXFYUDOIS0CoNgNCE68Iex2WpcLI+As3iR6g43Hb+cBy0aYvl0KtXxvbIgqqU3sdQLh5ry9I9b
4iPCyMKC3m4zdkH6XxjluxB0fGlDtFIy4NKM29ixmv5s2YHtVXQGRe4MUMsHFKHsPnIlvSBAfExE
0Pi3QDW/9T9XPeaoBek6vVdq8Aaj2jJ4SXX/evhHSWfN4N3/IrnblbQg86kLxTgHliy5cqRiRRc4
ooBZt94HxMSQMfh8ZuHhCrcfCofh/dkcYzcaBWJlaWr6KDzWjQWM0RFu5ENYvHCObU2shpgzRBSn
j+5kCFuZOJYK7RPYjpm3C0mlVO2rH8NW1jKVBiGv4LF1Eo5wgRIxc5F4d3t8abKoOBLd51SbxhhE
9kXbpldiHNacprgmo6h++WzSoccJDIapY3Iw/KEgjifod5LluKGoC9E//m1q+ihqVuXWkscURNwd
12U2cE1lzBM/ryty/aVQMW89a+LE0KfxGVyjNgaEBmZYmfucmjcGk1hsjWEB25dpHV+W64eiO8Ix
G1PIORDjv+HBskC/kbzPKDAfze48OUlwvYjIRdcZDmS6IagJoTIp9BJ9Z4olD86m7YiRu5sW9wCW
rzvwYSLkYQGxmYBcxopQDLyD4O7fhS3lOCEIoVNmnNWZBMKwUfrP4oVn4uu889CRmHFkfa9DRhup
AVde4VdWULTjeLv6yypBU1eAJpG/iUy/V5TLVlGrq9uhm1xpum9aEC+ABpsbj/46k6WI4NNFzsbJ
SrXQ6f9GigHm+v8u9I+YeSSYN/TUg7csO0jGDzhp3Vf+O+kITWMumv2YsAuHH92gyGlYu/yu3Z5X
7GPI4S/SCISWov2n/tti5+Py2KD/59HUENaDoC9qQLSLrciqRumB6Z6lhoOtqNG58ZQIVZQjV4H6
TN/MoGpgT12AH3Svz6LFJqlw0HbWO13Ejaj1+/IORuMV547FcaDOfuqb7TD56pygeIX708TPKhRo
qVZ95HhoN/AHHVWz1Zkw2UD/y+piTNC7YeGcN48Ue+ZrjhifCmFbWDpuzsBKsM3TzkIGDntZx/K/
qTZbIsyzx9rmon0tiGkFRyMKLI5CtU/ZMygaeORYuT5rlb/Yc9S2Q66Y03mIaqCrFGj8LNNVBE3n
BBMaIFxRx0HRNHM53kvPn/ukU/6MQLBd+V8wAIXI0DlDv52PFr8WKpPnC8Zne+QtKq6KWl0JKwKF
tvWiE6gjvSz//C5XgwU6Y6+EplVv+w3eytdk4YbsW7VKfTSqxNdZfk5igfyJHKfS6yOQ+M4j1IAn
5zT6HCTRoKb8jLVSSEGDfF20jqDakBa0Cg5p0+rM18Uu8XJQHCgxnGuL/sSbs5UfBSVVXZZZ2DHv
T0fr+5eMy4HsTzbWBgQBnWE5LXNnC0PqHFfBc8MK+QjlaLAeZb5cnyAnfraz7eT4yJ+01xwOvQCz
dcaOgqw/WxAAq0ZtMDeeruDQCbUs/U6uSEix77y9mCz2kQwn3P7KbaIzuIVp4W+BVwWQuWm+uK40
pbiu0RCOhT9QxnBY+HgYHyo8ijw1CcWxWd6E454Ipkh5prwify3ek/JbnaPPs7BhU8QeAd9OIVk0
/QEy8xl2DGWD8ZbF3KeUHjRJlEQs0suo5jwqex8LyEPpDH20tlR+9GMU1V/O+0mXwJez+N182yoW
w6u/4iemZ2u/dv/fuaJjbedjDkpOQmmJNQvoHeRspGV2LAgjxHD9C1YfKTvHIDR4pD5q3QGLzj1n
7bRqYeeYjFsQrS1hrkAI2qTsbWve08w6HBUgOM8K+Da+sH9ijNqzp+spSZl9ZnI0wPKPCcKSIlUQ
u63KiCXrbQ3vgbv1OJmHp9Yt4G8N1nDLk5pI326tPRns79bTl5ofnN+AhKwY01JFrBsPLnWuv1Wz
fSPpOFBPEoUz8g2iFuh7rqfPaykNF8+HigOAZAWo7HoRJlSX0oOuDqZgsEcbmDJvm1XjgXaA/xKb
2o7knosTUefo2C5GDMbrKhZwdrgpU98vWbUcjOZwacbkK61eUfpiELhzG4LdV1y1KQFRUvGNOatC
sVtpVfmOWkkstT6f4VsnSz43jfDGssEhEgE1jcJRoGM37mVfK8bfrhK7GiCguta1nstQIb/muMgY
vzZYuq2jAA7LzmGomIf45ZXAiBQljdmoQBhp4+KzEz0z8Mt9S4FXHpTHZWTQCJxg0LMbx/gDuyW5
u6oQM4jXt7AQjNSto6bdc9pqT3Hd2exel7VkKonzz4Qzoy2uvy6kmnszYVUsYtKPUvsHqJMdyFGG
r9KGn55E0V+vkNZczZWFkuG6mDGBn1w9rDaHLu6DlBh0ft3CgqHe8PzA2oU1KQMXCbcCck8HPTtR
/zyqOGTz8D3QwobxPA1xOL8DwrKibBocnj1t7oeAPC62MOmzA+y9uHg5fitSYw1uezzkWrhq076R
+JlE/3o6BkCmaWcxNQnKeYVj3X8sm4nbBvbhPS52CjGrpYl448nnqhMclTr4VlKoJdFVXAOBr688
QnPP3aegsZnZaoSBx5BO4m7FMDTnW0F/0sHo0WT5fvV81XxeyMH1N6tsECivsxa6Uo+mBfhGi5kg
bmGH2ZmUTfghf9iWRjKkHRqLGPg/nsamru+VP/ydBzSJ2VE19HhgVOKdGZClC/QaaUgm78TFA/6g
slqR9ZDbe7/oa6beQLVDyk43MQUIT3omb0wO1jYZHEBMkc0myvyWW0Cj+yrZozNDK83GDPCCCMyI
4vvocdpDfE2Pt2jP6BGA4S2pgqSeeE84klURmsUJJV2tYX31x37N5VzAFiTefqY0dUH/S3yPlUxn
/AIIANXAu0PKdLxCscG7/H/BQTCBA/nl4yCotVf1ZeO7pQPg/DY21m8oDJ2SIlyC763GRrKpjKop
h2FSseFHC5WxzKZhMhW/RwArIJ26iUHQ1+TtGxOgRHkzmG4bSNZR7q6E3/xhOd1/7HSU2wzlFA+j
mskWFdnJVKsRGyKX0P36Y5vQMx1NhGajBo/c6mW59249xOXYn+n/G0211DfW+j8MeaJlzvr5IvhH
6JtQ8GSvoHY5mDCmDjEFdLk5X+Bp1QofU5Tycz4GGVrp4IXMBUF1mLn1DE7fBMHijmUdJ6hHNH1i
f8JmmDNP/sUdZD3da8J85YA1PMLXOKh90q4YRh/SAkuT5/LLlFfenohLBFor9u5y+yAApdYoJ9bP
nzuYn3/ojL45VdE2bFOEprfyBJszMDLPUscRARteunVJvGUecGZjuQ6wELMomPTOjCKXsFKF0Eqd
lx9gzYeMIiuTHgjkjEtlXygFIzAFfGHVOqQjeXJfCoe/970ZsVCTdw9EHklbwAFxXDKgMD/n4z9y
kMlOx2TSen3YZO6kG2gCPlWQCl8Wn3twVVyTNcQjFrzftutF0Wpj9m5+Gu8YdT6KO9qPWFfddhee
C7Pa5bLCmMI2NS7OTLs6Yux/7p9KeI9cUSdS0SdQ5CmUnm2NfWaHcgN5cG/RJLae5RsIZ6lU7vK3
y081jjQ0depn+/UOsQTboNjk8MzrphIgEfohZFdo90/e5tRqA256qMfc+VF/nUrEUj0BacXCeABK
r4PfjNxhrPsfJgBecIaaxYKm8TCOUXhP4XpsiSo5kmHyQ0l1GNDAHo7qrgPUXX4kjtZQGCbc8PZm
FF/F9FjQGnh6JvJf5FViA00ZSFrIgsovjoM9ZFnzBVAD0UXnURSCyVCVc8s+PM7xC0ytxQ4M3qRs
XZgbC7VaX5E5KGckdNk6+oBFKCiCfcYfZzMibJNRfaUlVJkng4R1LH9hYGKF1/y6YrqjhWLoHswI
6A/BkyORzub9aB0oJ/vzr91s7QAmi4i5rkosvl/L4RDalBeVfcOMzthk6S09IPS1bGpht+idSbwD
aMP4qG89v/gA1SZfnyBkKpJ31tjA2XXTkBjlZkS/H3PKVxHw8NxeqYUwU3HTHzYysdWJU3mYqNuj
wVcVkMlmAN7dCeH/NqqNB0Ldj3EngeGajzRSKdrPkdIbl97UVWLUkI0I8UlHogO0r04ReCdHmbA6
+FMioE2fAl7fu0/nLBYB5m0mSqQWpNiqvlnCzn89RJbAOpWlMqE1wJRZsaIiNHOL1pv0JxAg8u6X
4Kqf85B+Hnq5yiv9QxCb+zWflN0z4Uv0xL3ruj0xxz8hykrsNwLgMAyWN+zouB0aA2YxK1t9grHY
BsmpNwUl7++n0HJiQSfYcwtcyklWxENOJcKoo7TeIpH8xkVLpqT54AZhcMxis+rSD1U7oV4Y6/tv
BmyKRjKRYWg/nhNm9c2yDDINfvLRjLRls/gzKCNlup5tEff6iQqiGLtJBllrHqwTidOJGXZBCeLv
+iLibEXUZFGkEX/SCaW0YQT3sDvIyMnbmOatI5Xu8oDE5heh9lRlWlq3zHf61h0UdvtfVkBWct+I
dTJPcyD0S/hiiqXC75t+TnpPwoF3g1CfUfcfAcS9UGXbV33GQooAcblPfEHzYv6+98ZO97ig7tFD
P3Nm3ZCm0OoOJC6x1Xc+KM0huToQ6YbUjEt5NmmWOyLt+9vVy83Kzmmd0t1LeBg/RKeDJDDInzZH
ohMZCYkQFiqGK+xSmux7qfvKQTfNVlu+6ERfmKLb/f1D48bV24tzc0vYsEkaLo9kUlYq0u+2zufX
iEy6XeqYD/lG5MAidW0XuimLJRsZE0/P0UdQ4taWjtaX/lFBeWpsbymmHqvuiieOM3DtYyV1zvH0
s8muTQJ3aBzIY9VzhsZSHednowbs3yGraFq6TMu1AdBGKZGNVzKTnGGWqD1zsu9TSowZ8UXefhWD
lz5gZfmIXXzoFQCZH7FNmxDVEqOXY2WXXP166x9QCtbFaNf8lgni8r2jtb6b12meAvEH/F+ljFv4
qeHCap0ekFtjWyzkMEwnKrF43UnLC2IziJKgSQwtrphRlmxutb2Nvzxxhi0Oesun2hzK2qhvu44t
Iy2aI/0By+QJ9hvgSRCDk8SDw/tWJv5Hvd4lmg4g5Je9lUdvk0YETGC/p0onleFFpWwrEJ27EVqt
/s0eo7CLr9JtMyoDTsPj2cZ0yCtBAH/2fsFUIoIImROGO6JcuG/4x5b6Jk+mOWo4UyDCMwkPfuFY
T+vHtef2BSDHkgxPCzlvrNHLDDAPbLsb4WGHxvA48LOacRjG0G7f1cS+ksEW7YmaA5rTF4Pxrr2i
SVMs4n0Vz172NifR/3UCU4Pjsfzn026wGlFmb+XB9+4GoZJZAQxxa2ZM6ARszZ80m/GscN7oMYAb
yiXIRJRfGRjNulhLK5TAHPD9yo10yhxXLCI2A1XTWOcDJgPnt48HX4dK//HMfqsLpfd1MlEMPLqg
1vxas1izZP3+0CV6UNmIoLEWG52981RvXwG7Ho0KsfexzTKS8CVxLJtkFh3iY57QM/weBf68j/K7
8e6Fw9l61P1E/RNliLcBQPvEOzSNu7S7D2UVPthRezbscEWIxjmTXrNh3qUjOyiaQM2TklOtrTNv
bGrbKcnV35V+FfrWeFC3bIxnLeeOio5CeAvgUNvTAgMJ0YYGtMq4m/Ic0fCSH0zLp2JoAkS69p/+
uZQ7iVysYfME5tPadeKrAad2OX098uccpDwfDaYp671XhPuUpg+/ah4PqwnyHqQYjm532pFu5svd
e5cD16k+re3Sfd/SKxw3Q16ZGxd4jNSMYHu3FG63FFnAC3YoGhey6zYcQFvFZsJHXnrpqpLe5PgC
KGTARtvsugJpjA9s1CyD+G+K7+QToG5H+QazzwOoqttRJFrvmH+4X8NavWmrl8nMwkSGqoIRyOkY
8i7x8CSsCaRvrrC2WMxe10aRorak+zyHneGDiniHSV/l7N0IXFCio/ikqA/LD5/1ZsDLVMdLR68Y
+HGnu5n33Mc1raySJiOgazt9jmGJ1+VomUx7I1ZxhIFKG2MPS4OCZSmhjxFnvuMwM71l+0YzgR55
kyMjnp0uxwu+h1WwfkrdGRki1uplkgwiEgZ9Q3qOFub9anKtsXi6CErQ8EfH0YvX1axJm3Z/eW8w
eUtAvb70M+UD+z5Z9Z1u9zbQbhJycYigNiE4xYYti9twib7z/QV64thAcIK3HHzRxw9fmJnUT1NY
lPwuyT6P0lohBOhxHk6whFG/aCBWQoWps/HI19TQxkVWX2nac8dMRYPl41eLcmRDmB3/nQl9wf1H
HuA3zw5guHg65B4rPFtdA8gREpXm5OUJ8lD5WjSoV1FhlPNZzsVTz3I2L8tD8bKr8rWUJvDtXNlP
5CedpPkHFxtCWb7ZXPNPhXnRqYuMaq3wsTka4KAHNOfKAA1fscBxL6IW590FXj2KlSRRZ4gTzxGO
5dn5pRlL1T31KTxySLSJCZ0IOpJnAdGNVZ5sJYnvFRwK2o1Q/eOBMyvM4mOU6upt5LtAa7AOzkxL
9CMd5ojtY1lWgEMcAqsmcxZ2eVBVbU6fFf28E9kaRw2S1huPCu9DjYSdraGvQs98D45NPb7CkCHM
t+Al+pvDw/adaOC+T/lvUxAgpgR7fXIdXDdTFzTvcnONX9bO40fRQxAOR9WRu7SMjMAvCHZ7P2gM
MUdvVWdQCfEdkU5tKEvrqN+kRKNa0g1nxDmW1L1kvp4YgJy4WNreh7sNp6poBrp4WtNzoN5gvzOC
7C5gghcDX6LSh2EcWTmazu27kj7ie0VB0epzJYaJzxBnejo7+qi1A4TGvh/UTcH8lgGf33YxI9DH
3kcneat7/m5bP6N7kV9+Gk0CgNt3eTkVRNfdOdNVVx0FD+fOHsqN6EWntloM4bE+XuEx7pdErXMn
27AYbEzM0FCzgMj2a90AQZTozr0UFe/8hZAlMbKaLAnorn+uvs9yhbS8m8IPqNYUVnbIRN21xThB
JI58auCRPHMqp42YlKrOmCZDCn7dTKt/D6ZyGvykTCBUp5h6742mTUDcRYd6zYMrLHZqbj01Pxbq
ZXHWfBs7xpiEYeQMgp57OL6zXgdqu9ZLtWxFaQCpWKm5IQXSC2dDPES3s46U9eNX/s6Sj6L+IbLr
UtP9/ZRCXy/p0z0QFJpupjmHEPa60RVRqK1Gh/c8NosLRVXX9wJ7my0igH+erTewjlVqSlDYXIkJ
z56OSKEQF+fQbyDu4gdnjupWa/iYQrkwqjPrr2hPIFxQnH58tSJ95Lh9x4bC3uFgreUN5jcaJERZ
SLMa8mCnCprZbBKxmXxnK1euGT8lfn9e0mfs+rgC9e6piVkqRiCV3GmS9YVtkkGuZyMZqCghm29h
PSYTWPwFvP3Unm7epcxjYNMeS6yFadv1ZJTUZ5ZWwGDVelqClZCbBP6G5YnpXwg+xGtCUPcXg1iE
sBRntu783b3QJYT4Wlxk5/OhzdtWI4howJRFlvX8cXdU7f2Shwciz3K2zVUcdvmzaWxQ7u3uFvvI
8xE6eg2gXmcOD/XXXM8G6WwF508GrIGwRU6owV1tUC+f6qcYIDe4bU0IQSYOjZw1tAV6Inis/Lrx
XW0IonlKJIuiFe93XRaOuTdzyoXi5eup+B/yFUOJRoz/C3jHstAYhf7dcxfSXfVD0O7bMug4o8Gq
zTUU3kmefCBRNgeFjWN+a+388+/sJ5KNTWzVcAnTXj8g2C5+RxoOSf8mFqWMPNWgzyygpeKOAZbZ
I1YYVAK6g/qFs4po1bF/bO5hL9OivPdliNqFK5naKMgz7ih99JOLQ96qyZSKkeUtSExyDyz9toIl
Gn5Eat2XeknTjYa8ThCeBokhRSDW0E19MMRYqShfSzgJkbqYgKUnj66+l3H6YzuS3YRJzA9RH5mA
ptDQtkAQheebIQ+MJR4Xhv2Aeb4NeR5mckTQodiWw8C6gSWpEogzYNoTFz5XjIhz1v6lLPGNPzLN
4F2J3pM21qirhEYET29NyguE7ovCNMX903ixU8QcurQJVYVtuhHQf9e+1E9iG7IwLvzKEI4CLzaR
zxOEyRbQ/FpfQnk/dckIFiKb/OPyQ8kqgeeR2T1gllx/mOZpOnaM/VXeBIPHhfdhlTqScJo/Nf/b
rHWsan6pFsm/3HnKimuC0UXjTPRNtGW8gqRHlcCW5B/YH85ERRpvSZMrK9uNE+9baU7zZGTLhKUr
JE+d4eCZ8fqHD2dOo1+Y4OkaqJSAUA8BuIflsDYkEGq8yuSuOvUr8jrqi4KtGJV7kSbgdN2BuLn7
I2FquZKyjzUP2mGS6CtpGY1qdWvJw0SC4iTcnB42wN/Oj6gz8kUdidpMw1/GiAuztYcAn7R+jWlb
Up83McK9Znpsdgubb4A7HUkFbbAvrPP+VwX9CXzEk1hjaCjjut2ThuUSlSZ23X+16KN27Oc/HYf/
e5FmezKstKQ+Pix6IKWBv30HNWc9PRk2oxGcHkx8HcW1sjtTEO+J/4VKU2Brl2sUY0qpF5wV4LEh
n6lP6LnmpuVTZTBE6+h1Ya8KzJnRoBmYrKKC942CeoAxNSKDgLNj92ictSRLnuf6crwL5Ju/gImD
a1heiPTkQAG/JBHNn3yJBnh1ZEb4Ora++sO0wePnz8AYfP5ByK91dhYTHz/xoDrAFg4MC9TdbvsW
Wtv6H/hxAKH3WtNAZCOzKJcMoQQlpIhy6dQJMzycHm4Htm5UUvxAJZmQCUJ7JNH9NPJYNIY8Aq8S
vmJG8KYyk7+N0AFaAMrQG/uI1mu4yBm9lBCjjW/U7WFjV18kO8SGhzVNBvXxFVkCyqHsj7qmUq5a
feu05OBvYakACbNIwMJNMbx+FV8VAN34mHXMcydfcEPk03mlGtCdFcyTfrw3KgqJ1Zdq7ncd6rRr
bGC6HLL9qx70AcABFE+qz0z4cVICYf2/GBwxijWVEHbdBzCic0U1qouFvy6Qy2SzgHGpyDmwmOde
nB4qfKzoF4FVD04+kBVOgKHUILwJHF4b64eIsYDxE5aXtz6Upo/8z1yYB+tei+UKlHsBOAFsMLXl
qsxOpC4r9N5FBenD1nn2hMBwemCNDdffltho0Ool0MP/rNlfmdN8VM50/NvfrYtSBWiNlsgxR9iA
vUs9Gb2zMEzXsG9crzGH6WE1WtJbBEIeLxMqSUjdKNWfD0k0G+7LEyTOD6KW/CTU6Ny+A4d8bff5
jPy5AeJgD+QEnhTRq+w8avzuU63NUwCD0Lu632rWiAzaZ/trJUMTOVYbEC0C39BYX1/bn5KdJSaX
yWC6rBJftG+i8f4xEhQN3ryOuh4TE00mvZIsE/wvf+3WmgK62nSAnskXCovwDaAn4UegMrmm9Sal
uN+VOuF0De815cr4ix/f14g8TuSxuoQPtemyZj2sS69kI1Is0eiPLkpXUBY1SG5u3DC2uu1Azxui
BFhb8V0M4k3Fbil9WSS/lArXMMGHh3Rwq5WyChvUfPWNzujAfK/309RL5jkUS8Udq8te3jt+NOW1
sHAgX7YpAx7D/HEH2K2j4Mt20LX5wpcdx/WQT/AOCg+/6X0tCW2GFQZXLGuMijSbGN7N3zwYeJxT
+9yz0UZMkyyLIzofE4e1uBWTMVxS54ZiLf7QPJReYH4hXn3H5zMTrdTok+7OFwCgd943jC+Mapnm
sf2xhlzxeBXjXlsnkYOtFU8OSxY32LRZbIpWqDR8xvuDfNAb+WCD0U9MsDV2dflbC/zLVK+Nr91Z
tVeOMSMQXRhwRw+cIlieHTGXy09UYvQP33Wt9FeeGqCBQHg5zAz1I8p3YUjgcWDUaaXKjK/4UxKb
KQW1oP3QQi8zDi6nYASpD5Fcvg7UdAEITSQ19pg11vfmW7WyMx9iI5xfRZifNPByWje5mICfGSK6
dkCwkO+97gAhFTtekFs0AhATRkWGk5VrxUAz7GFB5bixjcZ/6y/T24XGJgkY5SYfN1OD0K8MAnh1
ulri51BXV4JK9wbEJPBtF7ehjlT8h7fUcej4lSqxqQkrXml2+8dzq/i1CRamW1+nX3+KMBq8jEu0
4oJGq3ACJU9wJ1twM9ziNMMAAfk4YXwXbMATXclgrnF2mHXPolt8wR2qq5sesWrudnmBtXgx9dFl
LgJz/E6y2R6ms1O87NgMVIQbOf7P3pIqtMKdA77atBbMltNXewm1itxRptU1UfTrvE4l6nz0O14a
X3osKUgtUQts8Aw3nhCs3FeLJGUdFGz9i03UvFz4KZhglGXhgmk0Z4DIVWrYdDb9fgs3Mh4GkSIj
FbjlaN25ADwyUYvF6utZ0LhP9gOHDRzR656f1JL9mIVIuszGBkwiCmwh7XjTbyPnI+DzbvtneYRi
97mUjEOH0oFLbQ+/YAfUsxNJb+qZD9to/EfOFwtOrtpDPtr4Ba8oUb2OBOcdjeE7VpyxgXGTqNem
zLynKJPG5DG9COXe+iW9nQMdbzzzroYi9DVFdD9BEgyLwJ0A1M4c8qGNCtN2/2tSBg8yevRcjs+U
f0UJ3UNtcE9UDireS/I3Vk+P6BhHny20TOMdpKHYOQqsaYIXW2w4742BMXzz2ZsTx/w+mhhL5O7R
Rh/JRzM0ELiPwyX8Bo7s0ZQhhUqHnOoKgqHTuIK47PQizE0ply66AOQaNZY2LkJD5kwcPjtOSJdW
Nz6/azolzreQrO2Enxsm4yQIAGZ4e/rhwh+364zXM/2VME6OBbhQCLhwY/QaJay59dJtOMMIdgYd
b9Wz8hOYdqLusQP8qH97r6nlo2jr03tLnyjYbY0gP6NV1bzLEgcOkKbRPEQg3UipnMlk+cGUBIcg
oWDLNmsa+5kK1GrE+a2mMz2MYBockkoOXcaow26kJV5AqptUSUYW7hh411q+/WIZN3tlFUKzKoOI
FGldZ3zOxHD/XhpogZbRNJYk5cXdD1SsLCLcht4AV44arpO1IlzYVrM7VRKx4i3c7Y7dvv6MlcAW
cJJzhbs2V7dujf9SBTZv7+e4L/IZd0lCD6YQUhATxNzQlDTpy3BRFGLe09/s43QO5pBiriMyDi5X
cUU6p4NI3ht5cVvWP84dU2ALnxAMLZy0mu75FhvpiMTWERpuunHVcm8QLwbWdg6ge7wdWFURcwv2
XBX808BCQxPQp8wQsfHropIf69ErayFxck0F2x8hEVI9hyXGJBqkKsYpuVCwqfsHqLIZQTlJ7oD9
0nJJLeM1pxgWeUg+B7dGWnJUnN9phDQMqzyg88rBnHdt/mktkgyPh0qaF+A+KZTUTV/F3HtxFTpr
wVkPT6z3oWTaxWsSdUokkfYHsv8W5rxc6EplWhct20sQdSxaqplGWPd5ZYmNOj79Z1OGQcFEpOtA
TBSAM4QMmJy3P8ZzNsK2DogLzRjvYTvoYm6r25erhxkN0C3CHJR3nJ7NCF3mFpiUebblyZAOJJ4G
V9b1J5xuLkQl0eTuU01JdJ47tITqvb0H8Y953lGYcgy/wzAyV3ksxnK4jSajUPnHFYzyvoRYiO4z
yLXBYU/1S5h/7wNgvc2D3S+JqNR5KASyzCURQHs0oPKy489fHBN/TON7YGE67qHFIjb0/odMUIcH
DzjOKCprdYkoRegVpq/BvIaHSVyfPsMjBiSO4/bEL5uCjq5DGfzeEhGhPp5Wt7YvV6kUGE7EprdE
d3dOMx3pkdc39RzhD9lLrA5kAek8HOQBovmbToeht/2ohAWO1X9++Xbt6T5NAlXaXa/NdyNmXYav
T5ZfBUf7HenaJFLHeQ+3wlQFKybXS96pSDvQFXe9rR9COVgG5VgV+DdwPoj0vIG2TOy7wEl9k4Xg
wWP2htZ3xqQUwNM/AHlikRfoi+RIZvrvUxofyv8bKBZFjz3IjJN82EHoMau7lf7hmljZ7blSzOvM
VUp4GsppJU85+M1iW4/ze7DzD2pBfEvoJIWvrd2rwfrhgB0vMbM3BEYspLtt3IlPrPjoT3TH8tbe
VsMvg5HtCvC6d8b6wpyDB9wumrwy2SyhzrWTdlR829597fXmGcFSXIZwXNF4MCSxKanoKHC5jC1l
eVgwoYw2FDEW6FDtR9RKNHQ5LZCEKJ63wvvIDVnxQa44DidKSPbJSzNiJgqc0BzqVoNWbhym5iyi
LCZSb3/K/pR41Uyu+6ti9mJRziVENZIBwoy4RoYSUE3Jd14c5/HBLumQJMWeZSjeVFdJww0yIVqv
1bktQc0QA1Q8g5f2CVkIbE5RwO7OpfPEktZgv0uY5OIi3LEhnDxgyBY86el2WPxJXvjSkd3ScWit
8GPpc5PzK0gO/PEhG+0c/NpzFF0X+8aGU2Zot4+D30DE911JiOjiHYT8XBBsC1fDH3wn8tBlE3W/
flsj4lEZmvt1Y2zO3ECub7RZRacDc5vqrqwykuirr4F5YCIqiFvwZrVsQIBIhTULYk3kinFi/Nd2
526MPO2nSmvHAeqhmbywXGacnVJgOJXz2Ca/fAoB2TCt/kUsNoJo6JerUyebvRoqT9G5Q/gluyrB
faKGAD5E9Aar4/RRmxcu6GqESB9F/qPOhXCHRg/oOQW3U83oEvr2fhdWCONtKHoQlUuxPyys4EiO
zRw4gn+zR8C4sZ2lpFz2eqPOPzXwL6lSHx9/Gxtv2Xd277+n1DIRUSlzlsLjakwafXL9FedfL7xb
IqOIvrjWI/40/RCrZqXgdwrSPZVvWKSaVJ+4QFUy2FdIye0CftiUVjZTawnuBXLnErPsORK7uRq0
Ghd6bMJr4r+GLQkS6+Nhwqe/vpowlCvj41hcIrIV7+SYae6RKEoSaW+diZ+nj346W9Fhkli2LgHe
mJ044qZ38pbua2FepIvadw5yXPj+/VCJdoPvNtg/jFqCHuLGWsKg7fyKvskFoEngaWhXBySJgG7y
QZ9SVNFhsKtYbf35O2JywnEK6od3rOJ+du8HsWc8UuWHyjdjkyD+NevL2Ef/xQM9s6bsxUClCVt/
ld+kPRAHirUS5lMWM1z45UC5YhA0is1UEe5PONkQDFhd1Rz0kkrO12gifACKqYhUiVPLKSxStxrp
SkXyjWp0zwuXcc8P/3x4jKytPWwLHtZQP127Ubh1sctcXI8MhQJHmc3EeWcWMIXlM59m0FowNuSe
Wo3fpZscgITXhjEEdEhiIrziOizgFnfrQL222AOGSrLKPd2AuGEpWiTuOzmOD8h5UYFKg03VQTcn
rHQHeHl41N2PasS8a3NdzdI8K15fI/H+Gu3Y3pD/3hcEIUAmq9F1upD1PxQBbmQ5RHdSWFflce5g
QHHOWnVByWP12UmPHme5G2WvhlfTmArJDihZ3B5rdXbpgTSXC+wBTcXI1ACn0zaKbbOPT+Xp2Jry
FvOc+pKm4eBEC8dzVFrMo+CFVcKEZLXK9KHnOHoWya98GGhBTPUGqwyEJ5/IcAxt+szwYT0lNFi/
LiSnw7mYLX062SDfBj+vK5zMj+LjcmPDDWOi4xtPO00nD6OxzFK3heufxegk/eZWRuMAwd5u6tJE
6Dy07za35JhZGXqJZl3CeXlE7ti19URHwNBAchhD+fxKGw8Qt8bWIlIzJLdw+F825HeWOIddFya3
kFTfBMrj9KMdOJrjgeJ35qYGcUF++Zl9Q+R52sp/EVZ/3ZCJozecJmVry+3n772rKZhhPkSx6WMs
mhlfl6ekacmvr8mnlUetvPfwikXjxAyMYi2wZjF7BWpogf1qIoW6ir9KMJ6jaAe9pI725VDDwJ2R
BD0tIr/7NO0BgW3yfYO/xfLgnPH1Au45AFtn40N0P0DSiSrquz7u6bi+1u/5nri3p1Ch2nxUTLvU
w+nx9FcVhauu+qpN3mxSwZD3QaKdDTJAL/PfbFlEatsu/BjuQ3ZMsi3cWcFtxGKW+CVKrVy+XPgJ
Ie5KXsJbikC6oOnWV6HsH6p7NgTBsYMt22PlX1qK4/rcFvPtXRxZB25w+m1wKmjAD/iDqisOzMVH
JhizcnNoo2RjpfSRvwmBPed4goFUKHFO1j52aJkDwh3ho5qpkD6rzAwzdB0QxaGHTpXFwEqjmp3n
eDZcau3K5FsTm6T8iWKO7DfxN28nyxASeKqYA1v52pFkriAI6zRyiWmgTsD/25LJnaXlp+K/Udmv
hHMpD8FqowxAgtk5CHDfoX9RYB5XUeqcvMgn3m9CjPT12XC4kZ8ajO1wHvBCEH0FwXUrfgpDMS55
J08Hd7j0ET8b1MJHYna3trRMZzirGHVE9uNV4iPOmxH1z/mv5GbyaqUicEGBwRrXPdaXEyzK2U3e
7h/UTdP2LTv2Vg6RNyqf7avpBYKBwz5QOisfNd4bj6kpU1ZxcvZF0iunJNL7tzPQvEw2tIiUK/dL
AeVNa+Izc+/1KMrvdmP4MpmHG51XBbWhlQlpSTb6NN6MroF0R+YoEw3NpmJ3cu8attKT2b+7DJeS
OG7L7xTCY5g+bxr4NR10pgsixCiyGVFH7SbkyGvV5hrXwq032RldDY+scvMsmhonaSbwtQCp0Il3
dQo4CAARieIwtHc48WAUu+lvSb4MxTAcipf1UkBesVGtaa/VZzS0vheqSn2swG2LADFS7OGaH1xc
sR5REaZfmFaNsA68xuORJxJWQipf1zILBq5w6lh3CKsJHPda5KBHC5yZTR67kXHDoTRqIM4ixZPc
P3jbvaodvH/T4BeNwHvFbv3GzVRg3YM4XGCwb5/NkSYu4/iui+mgaM5Z002AwfiGnl6G5at6PkOX
bK5q86aTISDHUs1RP9AnnbDGOECjQ2FHUOVUvmUUK1bY11A2/5V7XTbJ2nImDYYHdwOB9ZKSkJIY
Of3mC8083RQZRBGWG4eknXJ7p2PmPFP4Vv/wHwW8OphYO5rX9F1++fJpY8mwhzzAm/NpCSh0olrn
4ntfy2YJprJ9PBKBtwOdKnJeWHZA2/Wbd7vEOah6di2Eo1eZzzw3lCDPcqLSSj5wAC4vk3xu+htf
LwBVRlf0zBy7AvKnpOBQqdAiCXVTBefbGH5ck2UUYK/SiY0L+uOQyPNGrvP7o4oB7hfgWH/vVPjM
QO5exicG4wnf73XC4Ne08h+GPfAF3KZ7w8vPT1lw6Ep0MLMtrgzZhFF7gIIq0/evOAzGBdpROj8W
PgiWQRA0U3c6iYbVSkBhhkfwSGDaDuM2F6jIlrddO7aetqSdt9f+4jyWqBzTf4fa9HUqj2+QvLPQ
HEekBM6Bs3LsZR+fWvJYm5WO15m8HT4H29TH10TrbX0yrfHwxUTvgwl9CNIaW3HBm1xhjV37r3KK
xiBMU7hzAeTnRwPvvEXuQPXc7ydJkPQAYpUwgsckZhMvRM71DnG1PMyVCWVhJyExsbseLqS6MQvU
BFn2oQRr7AUedrfDrHrtUnD0vK1Xq7kfXAYJTOxIRxc/a9TDBjvwaqj4WckHb7DarwlQVnkyLFtu
BeGbiijjvchFLrIZlF9+wF33Vchk7w9LbhVHqfxDPJ7WCWVfwD88HRpelmtfVpg/3HVHK9432V3F
N4BsqsfEBvAepaTIWyHe8RjyCzk3egLQ/K8ikO07lsRW3eQ5836t1ve4TkMXXvvSSomuKKmiUB2g
xLou/kM4oPTZHaqqPgRqIR5QL2AP01kciH+wFgzMtU0R8XsiNp6nnW2bGRPdUrxcMEqRm2dXzZ4l
dCRhY4HEDoWcoOA+fB3W9sJinmrlT+qRVqa+mdbiqs/ScMxnbbJIzfIAlbAgFs1aDz+dl124GwVs
zhx0icBAXCPb0oFGdeiuRvJXOe/Yb0VU8ZwEizmqgFKfyfMyqBsCLiGKApbh25I/3AwLG2QODMSu
qhSP1eNdMvVObHBcUz+qXIslpYy4a+uDaP7D17TUJKRH2I1C6YO8ffQkoVfXZIwYZ7dSy8+nhbuc
9jOjDSsAzqygMaCeNNIf4xpRrNRyd/NmGACWdRmbgKzw/CC0ZG6IeydsUlL61QgOdB1Jqz4DoLr0
NCFKHpnZ9WM8K9uH0nUlXRRqqRr9H3CCdAF8YMkMcJpKpSFdEP6tfXnHq1ItyZ1Kvwe+zupyCrkr
sr6HwpBhyqSI4vV3iP9OOjy3XtRR/Bn/as5GXxZjChI2f9zVZh1fku3QelryZYGzpGZy9UJR57dt
8q7eqEkE6uDKMQRofphq9gjB9hz7U9SrUBn0Lx0vhUsTxcIb0WNBWnT4aGmtN16QePRaHcLsyzrn
mNgY6o0ACcb/tuN3UphlLAmjFKhBJeJPnDA9ozYPqOrlC2gTUaMneakxU2fAclzMEtqqoGkULmWV
+y4PqtytbEgAEKwyi/sGxnqXs08dyGq2dYd8zgTbG3CMRfB1ZsXvOAZU1oMWcwiVbzCHM+Vy3tyx
sRNdHkr3ruNsqo2SRL4BOg5v8LCae7BqMHST9cuzIO7izZLfTwtsWEemzGPmWks5GNNC5PS+3ll8
Rk2bUAtZ6I8rahqJEXF+Iw20xiS/VJOP7XIGI3qnMA/JaE0USVChWzfXHLq5r37WQadLGlxwBwZ9
J0LhGtexVX5fYMmJppYaSRov9NC4z4BLjD+mDy+1uj3uUQpRziCqpKgFDyVELrldDYB6ukJFsmr8
8z/Yt7+RP1U+j/22hRhzbZxkilQiVrNeNBChX5XakihREhvqPOf7ZghZfh29ON0wMvML3YTWFgir
hf8Fo86qYtIMaAwcqPWPrJ4Xxn7m5KEX6HulKwsZeHicm4FkCXrx25h7rTQYQPDNHY1kTcy0hPr8
dPiTRqV2qvTcPlFZOnxYFQhbjloKl5iC4gSN4Ox1K1eycoFqUP9+NfyanyKYFtqHxNq5sXd/shYd
lfdR+epEtSTJvc5Kg2SFa5bxEFWGBPgDxkPziP6RHUDq6vjCvQXMYwq5rKw9bx0iyafEA/FBhfXN
lVKK225635trb/z9U0drusfplXJxst7T8hXP+yeWqD0Qac9aQEgv2xTxLaBfzl6Z9DSBCQthxQxT
rEVeEf+jkc5wyRDsM+I+WIjOGtiQOXK9J2fDmrMmKwMmHUXEaoFbCW3F9tZLlUe3OMwD0i1ZZjrg
Xc3uv6kFYfDRpwcUJyzPZz6zVY26xBqgkzAARE8jUzYvpKexbwW/dN3WS8ZnGYdAge4p79qsxmB8
OlEOJHnDLn/tAt2+Ey4JB7W8dtQkvh+xjSXijC6FcmhRU/KoY/NuSpWAqxUav+2O8eLLFvkEfa4s
IIsoxR+3pkII78fOzYvb5uezvDOLB0xshR8ZaFZB1ld9UT7pXhio6OJvpfxOwmgbYyT9CUmIVHkP
EiHzutUsbBhUyEh1ee7ze+Iwb+esaRsCxGy1XkGTn/H14dv4hsdwSbPO9tcGBdBncNgCWT/XQPEH
f5voQh76Avj1+TYT418QdKfaiH//d5KyzUAMAplCQyct2pbVWFu4ReW3ruc7ydHekZVWSIVBNKbN
Yb0Lrb4cFZSqNuaSsCj6MeYMUGtq10smv9u6D50R8eX4seZWT0cPgEe7zl5XYQxc9m5geMKMYRhB
wCa2yhKOv0WCAynMRfjIGmMV6DTlUjeIYrPTmi0V1xqZG2X9bT6WvidnraesAwGJ2TOAPmkbnu6o
sO/C1xDstbVxBFqwVPVX2Sh/tfBCxNjo4gQK8qEvRDxut07W4ioVBK7CWLOSw+sEU8VjWdFAtaQe
/Rbw9R/kuVad5PoLJGDAnEmMRWzRuZMNU/fdxJfpUpzjXbrxLMqAK/gnpWBwN7upo5ezjP5Dj1CS
72cNI7aKTazRx39TZWiun3vUY6UQXCXpZpAOZRnm42MolbqWMCJohY0r3pc87z5/8Brtnrud08Il
D6Cqw7/NrF2vth96tMIGlCK3esUZ6+5OEGmEEtKaFoCy/TQr5GD3uSmJwC0MeyzUeLT6KviFBcNK
0K041f6BHhPDGouXQtYMAIr0hG8l+uzXdHu5zDN2FDPTy44VbiYZWNNE23Qt42MKX6CvPQvYJteG
0IP2oFpeuZyt/IPJHEScK1UbGf1Mupn/sm4K9xt7yoIVSA4VNlvzkqtNgbtNYLFfuOUVb/sBGyNM
u9udOSHuUvJUCaQSNJN1E7bkM361dU8mDPYVY769aEm0EB9pmTF8YEteeGzXPn/EWVWyEi365VLc
Hq1ThbiDMUR2CnZAO6n5v6P5E3AIWU8/aokOD7qcXUjmS1hyDveTUQSKe4PF1VYFp3NB3IufBvgM
6g3M7ILNzE0kSm9xoMaREcW5VW6yezOBzixUzZA+H8Z2TpcNUWXWRf1vEpzs9MT63wxjijSVGMIM
QPDMIvtMaizVjHYdH6mC0c/0hAPrFDoCpXeJS6dYjWcDOq/wjxgjzdTvD/J28e5C7+eBj5AJp24B
1EMmSBZnGrkACnfgnnK7Dz6pJy+MVGKYAEWm9I9B08lGvmJ2esZF0bySi1O2orB/IseZnG35xwjS
r9jlbRIiBSHjbYz8CcugRY2MFBuzoH9dUdz68KxvZuRqDItU2jLjTMyk0/f6U3GbSQsPiHKkSGTJ
OC1kL458hha+3zzXgkIRXuBUxdSMTq3L2iPZcl16wmYXpUE8tTQ+igxCVLXKc32W11ZuJFF8lYKD
GqRF/Fm8b/hB3/omPKJeL4rZh3eZcbTmh7BPeymSlVvYb4txOlk82eoAwK6eTMsSbIlfG0+998Mk
/DhQ1ahA53NHFcm5yrm9AbT5pGqi7JBr1Crb14/0y2vLoPmlu7MiLoXWUHgsxkf2rS9duypIx7ZP
VlkR+nppsQvuXA9JuR1omfayyUdKU49gpJaoNWMEesQ5xcKVqh81qa8mbtG/RlkWsuncnmWlALIu
DNrAdtw1WP90TVhReOWRdln1zRqeh3LnFHjRB/JinBxo8nQmrZsUm5TNtRHxKK6IyGKpXXZBlKwn
qT7N7NhjUTwcLVjYdML8hhAzk88obF4yz5TSUtZRtSMuK3zRpGCJwzNHWJysEcCT5m2gW0Ii/68W
MDjZVVCs6eOt046PF48rB5nNLTNSlizkDumvJsYABlklwgk+DGN8IzYWenLh3zGDMTfc0zo6GxzK
/Nww/KqwLAhHRWPQA4NnFVp+Ku/i8kDr3USU8s8uJf/paqUHVMH9rf/eVSu4y4UfnBxZJL+dt9B4
Aom3Bm0CVMEfIldsMaHpSpGbbeiXDQVbHlX1PcMraamyBOPBJgqvKyiieKut470S83ePxKSo3nCl
LVY+j6OogCl1lEVHK/NV+/WBz+Wt5dGSqrYrfzjZVUqTE894igWVbOp0RlR4kO16W/qogQ5XobD8
ajX160V7VflNDNnMWQIq4b25CBDGs9u2Qo+ZwvCk77+ElpnI7XfV7vG0ivgFGRS2YSnYXIP1xE4U
UerIkrtxOtB50r24B2Ve6qu0o0wrdt4mLnrxW5r/3UOjcRzYnAvt0kD7FZ6MRWVs34fotAtf9XeO
uefrtdbNkecC3xcNQvdEQRW0Kl3zk3aYIlSQ2xp5f7NoOVuB0UrYbgi1xu4Vw2iOUUnXExv7MNdE
T1Zdw+hTrH/c3+QrTfGxKfT7wCNEslr0knvr1LVIdv76a1blwbQ1DEMtIxpszSZkVTFpgtAmefIc
bnVxDXJBb3MD/1zHTSs5ewKuRLBr+5p9kNAHngI62V4fXHhc+ozAgZa0cGXVY6XtLWusyiXzDgEE
ofb1eVh/bvABlSU9a4D0Z4xAUhCtBk9V1rDspgfgeSBKouoYxiDhbvzPgtA3B3JWlMIk7GJx8x12
UJUlUDHFetOA0ebFm8qcS1xmneLqMC5yP1pYCc9yVIYmCjIAgAhzJV+rfF4wnAzETfX5UZFaBPsi
y5OgFMd5ldm5yGrPg/IIiWggTlrklJcc3Tn7sSuKztciZBBqZUAQ7ML9PqkHoseE4MTSUuxHop2u
M09ir3ynqh11FOOkQlm0M8U2M2GYzncuw/Qy7J1AD16i3PbveTOCPSFv72vNrBAgmAv2cgcV4J9O
JcRbAlw7yIeOhV/PIRv9ihd3A9QlvO1F1W54/usk8l8v9uCHU3z7O6yIQDGlXOCYXV2FyECvMJr8
SYvhtbWCHcG7ZM3Xy/wC5seTKAJQJ+GWpN+R61ZFmxBeAQTaX5ewZxbcojC81HTy+acVJUwdCo/w
QX2Eozbp1casvrpHy9tAgBq9f3rcsUpu063ooMpdyKdtuJb58pfgpTnqvCkYLO6Vo9f0RyNXLnNT
Zip++wdYzbzcXN+YHVn+Mk+vwfN50sv1md7WqP3U+WmzwbUyX1Zq+eYTcOzG5KeEf3B50q/dQDQe
xX63A/duYDbxk7AGiUQNviB0EqDXpfFp6sKYUruqVDMRZSD7zY0eZ5jcxUFfl58tsqWL8kGKkGQI
aB9/NOJXtoTVL2pDc0O/xZMtHLMwFm8NwWOvJocUR2tZcKEshlqBag3Es6LPyp98NHoOmG4FJUh9
w+kcj1qNwkA0AxDsWl32ovqihnQ7OjuXIN+HjtHfjf2sbeCQpXod/Ujr9UzjKedvQDlM5w5sThxP
r89bhu3ZUJXgAeK7dTBManA8rHzlIm/C9z/pd9ddX3zAsE6XD7mryK0e/hcqW2AuPwvHcJwE/W2T
GGCZ5P+i5vhpKZ0X+vChKmvWrynS6TZhPdXdLS23+jkXXJ1fa+ahCbH9+CTGNv+qpJaTE5lugP4e
wyKJM1F1DunfHmssAoTw2q6+/A2nA5EXYQ7v9O2Yc/Kef6kIOAH7vb8HjJjxn4fflpvxuj8mMh3U
Mxlm51WGZH8FA2m+I+tlkyzcdDYPdd73mhQgQtHkNiE/lIa+Y3LvTuy3KZVtRaxMWWyxNg8Iwtz8
1r/BOEJgJu/MJ7ES+d5IPYcZAnpX2IIZCb0Lb49ObUuKkJToGG/tD1kdy9QdparDQw7M6lFBjqKD
flElTguHwk/OLZxxBH2IYPqJUWxLpUnHe2OYBF14F9r0xz0wjNlX8vCPiqp40+3Jn5UaYjPIFoVl
6FkTrT1xWPdAW+yaeLrwXN4PL5OgQ7j5HmxnBGfxYcvVjZVPkXaeZZwsIbbSr8/adu37hPdOMf9a
9ypbqm9t8MOnwbV+j0+i/lEwuDByVKkLUZy33axzdHggc0kLiLLdhZAFBd2KjLvJVAB9tB7grdIO
rhaHg9tdLvLwo86DcD9pjxPECHE7ZDf0DCKHp5pKoPHOhYanOBWpesIxrmywfYwe8UkoHyZlol8u
6plrWK1Jxhr5mrDt7J6jE/3uEk+3S4bUE/BvQJiUEPqmDBBwIpSBz3yYVILhplxu2lpLi7m7pIPL
F5ryMMz4nNPsvfS2Vz4Q0h1HC2FQHzIKXEOSJV7nEfGpkvEgTsxdb/oK5DsF1c7AdrGSXLuThlSE
jbS2DSjHhEMhvvLKFoKvMo/Bt1D247yfBBgI2A75mJiBXWqqOSzksfMqxTwF2900csnbT4KTu337
VwHQLtAs/8jzei/+0jg+bzvw1s88XyeZy1GHlJMI7n/xwzdTqnag/ypriZzft5pZRKqAVq6H5hgg
HQGkdEoyQA2vQK84TllZ4ajdhXmCzHF3AqyDuZoNieFOEnjrye1cl2j+kKoohUhbQ+CH1wekzuqJ
A+GJv6EiGawrZx+VugQzUh6rUrMpZoGRuJYgwnBnzU1GiFLvHLadhsQlS6VYL3k5v96QDqx0bDSX
SaTfllgWVe9JxluZfLp0Ztj+VzIcvx0NB3hnz+EY7/Efxs93s1xSowj68SrzmYXayKCasE/XuwSv
CVFw6JYAAsd95fzttzN7i20tSFPgyWqret/ow1pE0wKTb4koaWjPUlK7Nvz1TCcvBW6F6dhqiyXZ
K7++S4I9/QSnj7C5xZ4B8jmhzMtLQg1qI3RBLEVCuulcJJwLGDG6JxRdUifpKp0NMGNImVhpndDo
NYgPrnyRT1bn++0UOjcy36oR+4hlv3dhvq6D4tX+yLyQMtxkIx9Sw54FmY61Kd4Cy+821MhOMq3e
+W5tYpz3Wbmzb5v1vUGde8KBjeHl45n7oGUw66onZgjJoxs6wpCgzveBAiBarzjciCFBLF2Ro2QD
VlzXFG3MxI5FPbSwPC/31JQRhjgymMBd9xNuCtf75IgrtergWvLjLC5YlA04knvn0S3BjiIUSX8F
Cl/qupZ8G+7q8Qp8Q9c/7RN48OYYT9w5Hmw/0oWS3qJipGnSyYEc0WCeoM0ZRAMOtMmTsqtFsA+D
3n0p7EFig/5SBYXlbBQFH5pbbK1E+DJAKnqScC/F/rSLnqUmqeXao/HRtOcWyu6BTIU1dEzxZOsY
97n9rnaQSkarKNYWoUUwIE2YH6oSLM/KZV/i4M+elWcFbsWp7Vhbj5scN7M4ANYcNZ+Ruf1hfRcB
6Qy077ChHEWoLusXsgN4D6lSWBQtG3r/ulT96+BzVoWWyJWGCansmE3F0G7K7SpEH2e+YEipo61q
jou7T3ftNcMWfjnscyIVo/604PWoW3E91+mFUl8sEXo5IylOsfcFG9OiFMmhd7V7uUKLeicJD1xn
hkneOdTwmTXLOrs9WNAhJ1quUe4VTfxdIz1PRPOPj0d93dsfA4hjYEShrFz430miyxWPO3LqMp82
l3WcejsIXvFHjUHWxW/tjUUS271TiugLBnNLVy6gmbQkfpuq3dkq2hfkkzE0kJdfzyDKR1z8r9Is
/VgrUT9a9qM6E6SRRA8A+5LN+Rap5tTTZAY6Ss7bUSE1kxlb3vGDUHqb3pxIzMJe+D8uwOkT7QkC
fsBmOHj4qRSi4AcRIqeKqmJjUO0b5iy1PWOW8XucLpK69PVPefkZwb3Wma2Bn2FWgpsk706QIQQd
SDYG6dRNvKPxyjQkLDVJEuS6rMOslL+KW/pG5CYI3e4vxdI2s75nHayDugtB6XN2FnSb2gj4Jc1h
u3qwXzbGpiWDcTcmmhdEsH7qgwu4b8jYCJaAX/LZk3Ie36caJSY1rcDt0zR4YsfHttcwmdpYh8cx
F/HGOU9Qz9F1wtPZqn3rr67oau8tcOluqIp1nBmamMS/MjKNerN5M2hrmVXF/38Fw+ChKAj4OFpo
ifpve2GFWfPjkIfquPG5NkcFgjmt7q8AAlJ7KXmucJ5taICsQWf/49mdU/eV6FCV1598g61B0bgG
mvxi3PF6WSNm3Jq9JWr2uVN0OwWGkpQwy1hOo45NuybUcAd6Iae0zm6w+LI39vo+zcomwiul4ZP5
b+R8MaZGMk5N6YqX9KusFiTR9sLMkL998GsXOFFr0hu6SkPhHe24W7P5t8oav13V3EvnpY5BU73v
ImWPsjTEWl+fIPhTQFKFxx89MbjZqH6PshApGusQo5HlOkqQO62UDCwnMoU14cud7lUen5uAwGhC
PbIBFM6fpVs8DvLGRwvbTqh5qV0x5dHcpqKfOH2/6eTCURJC0kuzUQXsxVNtrLtBvrAYB5TprYXK
BWD5PQbkBQq3BFxEePZV0qTcwfG8ALtw3B557bo2zPm19RPH6Yz1kq/qWHty5k0CP419HrzOdidg
RQiCSnt93utFx3z38oe8rxmwXsgGmNQo+gC4lNMcQ2qqu0PeqsHVr7jIQPsa4lRxppdLZoNzGRO0
izQK2MucNhjt/1r7rRF41O7f/g/GPA3CkBgFPr3xcGvEjX0wUdfT2eyMfCfJKw3W/qqubWTs/y4J
3O3OecF3PFmtqPMpzv1LkcF+zISyKpIeQmHpRh4KuP22sCke/z8yR49IgewUYOvtN4akwFYGEFMF
+tMompYW27H7VdH7YUH8leQC52oWCN3346IfUBCk7GWngxhjV1nR9Lmy3h97zJdgkEGnzJA8BHzY
duq/VQ/wgGiST4l8oya1BfixuCb4vMp/isVAqc+5GmoDDvMX/INM95qwwEqpW2VKKFFn+Pwangym
lgPv+3OQ8p8IZFuwEZ6Kze8T9asSusBBmOpDalRFXzGD6qn67urSHkLtQXSScJ+LWxnpW+rzeNtp
uGMHkNCTpoYGIttZufodkgz5FZF0vVhuZwMMHI8NP+ZIsebzXd/y72iBhGZw4THj3z8s1nza8Hmf
ARJzbOpxJvk5tDlai3VSa1IHKHtmV3fhNJjXm4Erxh0ignU6lnnXQa4I++GbP6ERXnpZx/d2TlkX
XmrJmbTKIZlpOG/iLnM0uXN+Ps8zDht2lV9I68uvJnNEng9HMr57z7YIupDGMPR5LLyIdHr8raBE
4lrxKpShy3Xwe9qdLM9dvakzXrdq+MMYqTjoHpDyGeO2bcL7Sbdgnhz/fpH1lpOHc8zU4/Wd9V67
xR/wBXDP/dY4pAsnT/hyPoVkgIaqWxjvDD6V6EqWKadEpNS5mN6gR9yB7n4B+aa5x1zswdcBakH5
1bPGrFvsuo52A8/QiVtjC1CM6oyRP2owMngfYWBGiKNwkmmqBqq4tahs402SmceVLaneAhBL+QLr
J7JCLzmeWz1lUNu8HxhMNnd+WOj0Tsh0VsI4q1vePidsVOWzcgRueJxBOejoKPTKeiwZiQTUc/hi
kiwWAQzysr+z0MC8vNUhoTibz1hR9RclKmE+UAx5kkjEXhVv9Zj7t/l6hgmpBDuVoVpmUGHlJXcU
Omhw0nhUCmkqI6c8OulFU9lZNAOL8Dj1XBiLje976MSvhaaSK8MYccFSV5C0VLkZMRaLPRyTSG5e
zX38LKGDA8kejkru6rqRhLmSP46vQ9lrJmBfTFzCJpbat2upslFlceMyWKN6LORzmOnUQUa3BCfy
ueGRSm9XoGtWBrH4++VfdaKGmtl1XsI4YlWJsfD50Ns3ILFbaOrNN4175SN5JMFiq+2kl+rJMFMv
nzpPE0XAnK2TSfrzHB59iDrgM7GycyDIt5kG29RG7e2RUxddS5QsjnczD5OL8h+GtHzSYraZvYfG
6Boz2QdXh7AaRPkSdjfSNlxEmfTkY1gCrDoUbIuJLRQQ+7J7/6gCOxAGXNbGbd0QDkZiMzfcWDlW
WP0kL19C6g9xupqW+dLqTLfCIKXubN2cGIcsWm7BxWlCg+8mia7VAx/Hegqy6F6K5ruNHlaZNEu+
z1ykDuo7AsAxEYQMaC3HDQFVcmVlMDi46iapF8AUNJKqVIdkpcPzL+hNH0tJ3C+DzuoPxpQOk1eM
2VuWAS+O6jfKHCBgv+dQOpUly/BQX9H1t4M9Kvj4T4/EvOgaVlZsppjNjRW0cTwbsMcvU1dOLEjs
neXbjg3E59xsyLH6MaOoyJN9AMhXdy5qsaX6rZWFYgzKwGn3CtxyVpSthdVWvEiySeaGDaj5EEDB
n2XIlc3mFKgl5631FCQyA/9gLGfVEzzfl29a8K/vvyZ9EeuXYNHTq/UN2cqaFDAiQKCXEBsTwn9I
2I9pvofIwBQWcUPEh+bWREEHV/3OOXr1TaPzm3JjiUvHyFl+Iajqm2/XOTJquLK8ye11IblZsYK2
Y1P+kBawpCtSY3SpfUVyXeswIVie9Aj2n7s6ep4o68chXppLX2LTvknnE2JpBYPnO4xg/57OqwIn
Cdexv6B4qyxBcHhLhWVXrxsdDTC4+Sx3ALXaVPKM6uIQJXfft0tOBIqHk1NPf2eBn+/qTaC6FcUN
dCHkZPOj//TJQ9axLRdYE3nNtmKq0SNy8GSlAFaokSImPTKmzm+Tu/4KkVVsrI+s303kwzTbjCCD
06AWADeHfXcxPU3z/j2Fdykp2LPln0v2mqL3UkGIBreFjI0qQCMAEDSuzUFN7Dd/WxM/9XiszUF4
ofpGJioepx+W7BpkP4G4FabLqzgDTQrDyoMjQxWEiuQhTkOVnfU16+6aMFDUT2wd6+c0SKsdLyQJ
nirWz6vIQSRuKbwP5J0IEnSxB8YIv7OpzKDqSAwu/lL1vloOn2KmPzwePa15ak030lNLbLIowh47
W12BhGRtKV+0KYr4Sp9/GYl7p62RyTwG65pe4NuC/1N8CASTz9Zr+gfhdJWRPBCCOHoCSDb9bYea
KG6haj1HwaJQ+a2JvuOLLNtPZM4cfv6JAE70z4oDdTpMm1qIT9KPn3m5eT6AJkdeXvfHkZGKA46Q
dmFOpGHNKCrNs5X26QBKS5LROhvv5a4Qv81QJUZXQMG5dX8NkIbU3TEsmivX0iP5H+odIkxnwTVd
A3KTUrM0Hp8nlHR5BEf5O42O2HG/bSwQbjqX0EqVT/LKl9vCL2DXzH/ikVxi2bPAv5F8yx5LG+hc
G++hyVOJvM3W+H+u9irBjarnZKNGPgvgznonhPSoCG95TaZKrxifpxypIlrJ7kjvEcPtcN5aqaHX
UrQYW3NO3vEBf/NCG/W4jeRAB60cg/NiDltZs4+N/y0ET5wcvA1qxibYGjBM96Rw84cprx5LM3+8
KTXh0Opy/dT8P/9ZeHI2JE3NUYzesqom7zvEQTknjzyUKEG0JkN2qyCBJRXOW6IwcW2+7CRsVq3X
gtx38Bhlhg/cJzlubgR8xvAvIbvPR0Yf1e+dKbkTrBqnCC6M3vqUwv5JqAW/97tfzcI1gFIMt7RY
Y9PBL6vxrW71MxcRB/W/qNj/gxk3erILm72UkYSLy1y8WX0+9gkpsC9kREn1ekVW4GE0n3kTwu1b
L5OFAZh4WOo6Ik134c/28S2xGJqnG0qIk8iZamYF4L7LzPi4EJZWCieetXK2c6/BRVsPZI7ZZU68
ypbIqq991kAH2k1IOvW3Ig5VUYlDQxlNWcXH5CNNDjtazyoR5DcYKCGFKGG2nskj5kSLubCtPv2p
ZBcjHigXoB5YLGHTQ3/xgg3bLVsO6XyXWIQXd9nImzPKiwi3Hq9kuQY5gdlw5kdW7Wr7y4oRkvMz
KwP8AYUyootB5ZbS2kyJpggdIA5nbux3Nawn/maHUgSTpOyTbhXUCwKTlx11fdkdotFH0M6II/W6
3IDV9Bi1vHsCA+QP6iBkJ8nc/Thgi0NsNgzgYfjTcbDxSLhViqh6FePccTkdWkLKgkpHXH5YdebM
p9H98tLOTTbet6F30Vq2H0drskGS6zNByIU/vhxJduFzmo4VBKfPVaPWWbEZ160QSRNolbTW/vHH
a96GwymNT3IjptOqfpAkIyHic6QpFDCjWAxsphBH/a9qjHLMNAIHUD49ou+NhI4QXHF4YXnMjYxR
WA/cyhkOjPwg8KOqr4ipKSi/ZmVTcTbq0WQct+XCUcL/rUjcS+XNEznAXrw+vgHK8yCs6ROc1B4z
Laldth1NpDzT5FFpvvIvXQjsXFbHrRCTBCeUnuLujejmnGKcFYp0QFODGabi5NcE2MvuW/ssF1he
NFmmTh7WFhJHxo87Kni6l2LI0C17MZ+pNPS9fKMwx/RT2WBXTT6Mxv8FIitK20QIcWgsl+KdreWn
mYru7gt3e27lV0tOzPnTSkP+c3x1p0rxCqJtajzNKVHa04vFWqDqBEjF9uyuvjuWSJanNfVFE0mG
ACY0c9uF4Fqih/K2WWbOi5lr+fm+4c5MhoE7bEkMm4NqOhyBi18eYS8Y8MC6rWD9s5XkEy0aqc4A
ZDtV2aZYLwdmiz89lA3GC5fD7tJ/qKChtffXYyEhOhfOK38AabJSoQC3MVDCgo3gLXY3NqHEzOQH
ptzF1B/9luQStaYYgv/u3ujYHre4NkN36xKlYQImZjELF1flUyFmYGKbii/y2OQbVCt1lrwLEGOm
L70EBxbcgdww+6YlLDFOhSeOBaslEVAFnz4EKdiNtmFRvJXlUdzgANgeZCMHFf6mCQnwQMHgmT6e
wPbPq/5PgYY0+2/l7/NEl1HRVTS3XT50WU9jnlSjePSfzjty5gQkNqUBmj8Sjr9KBXmg/mVpza88
aS3GAS1i8R8h6xf3+tz6BVwSsDdLaeGxPyvBYTJa6oRJQq60iQys8H4vb7T/bAprixAV1gD/7kPP
FPhX6lYTS5DCW+fRT8SYs2AYeJ4H04IKc2szIy+R2ViR+4hX84KaMCbm4+z1VKHr+7juGg8YT0XM
4ihSDGG+hO+vUi/NZhqjdYxsoz6v0LlXKAJIPgI7/zKkluF5wo8JF6awVmbDhf8VeJPDwhsNb360
blQbQ6cYcXso+b3fb966WB81ZTMEYoayDTIGm6V8Y4hadxKPmaUX+k8wghWtZ6Y4RmTnrDYmMSgD
VbCz5qklSXvdpnktgaFnXNKw5zd6HvNgdLwEMsuwHP/rxwBgNMYxVp6ERCUggoZjx2jju8XiacM/
tOqXACIlLqWiNNECXJDYHUIUyow/ORXP5ZqdoKBZhOKIGbmIZrrkdx81fNATw9t/WCM+Zd0atoaU
a2h2ZXdH5lFJppjKAoy8qxCFlNxXxvwsQ+jIuGf/lBTo7OhInHroTBqjp6NdCYjj0v++Otnu76Pz
sKQ6PGisAP6nzAz2/NM45H4ywT+AcyoWY8Nkn8O5ax0jtqOtNtfGDCzMeiAWAjTmCwq9D06Au79B
n3CRkpHrELaUAAxDzIkdy9HbWpfQ1Zxo0Z9S50So5CeD20JQhOG5uC9KooxaqfwZuhdXrh6YzF9T
5vF3OLa5+ZQEhW45DoiLrbNczOzxm8tiEH2+sZh96JV1morwgojy/02F+PowFU5NpVzTpYWgSDi6
QsLt6qDVLuqV1GaYAkG2au6TqzQuoCaa6n3a/Q0LkQcWM4r/9GhJkYXopGzJbx2oq9D0+dGDwo3O
5M5ulbZ+50kiD+kKrxYluiWBhWQhN/WZnUDObrNI3s2knt66Z2NSjtQQbXRjp/kaXHD0TP1pgwsc
VpJODVict/Eis0sL7pfmhpfs8tXiCaLdWAGaVxbWd3veNlUZvXRzUu4KixfZiIA8kMkhLVUhEpPc
HALD2Edy4/xQa/cdZ5DTq8RThMYuSmh6GncEGx24Q7bHdtZbrjslcbI+wMPED6//Maj1OhE6WVeg
qvJoWnQONOu2REvSUjHvR/n++C5fQ8Obx1PT9c8qTrEvT6xrbfvfOMWr7Q3vzUESEb71NvoNzpQt
2AgHj9R0pbvf3xIt7Y8okATYWKrw9DaG9O4EQwoeEMEm28cjxl4inVD5lF3LrTWmMT6MQssWlC1N
+2/TcZPE1VKsmrAvezIPAB/Ms35/RWbsMs6Do4pfVCqbm8jAGeWEHzYPmMdGkI7LjF4+V89g+GU8
wFZqDCI97aQHrBWrhxgoRfWmbjSLsRJ3MD0Foq7bpb/f15QSU76OtPPHlx6rItl/roKqLT8YbM2C
bLOw1K+2CSO9s/ZesF6wN2m+FkC4fJ4HapplYPQYx2yo5KkJpx10lfBRtmwDcdY77vI5pK2dKQS3
ll9ohwR0gbuTumQWZiQCBuKF7/NEF+IeVmZrFelSxw5XrJCYgu0Z3TXM1cLVRiuOmDmfbkIPf7nX
RicMkkvZN1u0a7QEoswVi0Tk3lnkPG5Y/IXMBdW/7KT91EtOskAjq/k0S2e9yUsY7vroOK4cN3Il
Pb/8eFoP6itB+R6tvz6SmDL56fNHeLHux7/xDExKDi+Fg6BzZT4ITpsVdjZrb/fKBnBzFv4bnYkC
Tf4nteCIrZuBQs6dNAAoJYl9WYesPWPh0X11eiXdduwZxxVr8rvcmvRoh2MC6lH1E2dpCMVZhvkU
c1hA5bfQhKrzEVTjxTIArG0T0QcoWg4dJBmbl3Xsufi5dR+FuGn+hoZdZbVlNWKRqjXspeZkYp53
+95cxuVUdgpKDh6+fxpyOyq9sIRaAlO62xB1sdux0Q/iaZYX+rQWREDzKHL2IWb5DOOYOowzgSX/
MQVbtZ5aYqxhCfrVq7+AfEdcDOj0JNlT8iVcqzCLteTBaIc7szqvmYaXYQsAHGOkkUG8jJ26L1l4
rlCtvj2Ikl/FZB5AP1wLhPDEoVncWX/svzi+v+LANaMHMfCXy6Hx5LsukXge6H6flhJGo6Hn6lQp
gnX6MWsddA07FhAei1szxbVFOWqIZa+PZFYYAhoIIIxCB302AUZK1x2K4rLmSX/ta892l5zvGc9k
qLj+o6IUWGDWX4Ekqf7YWs4FegjxgukdszI21QK+irkUZ/1FEBkRE9dVADuda0HaWSO5vey4w03M
0OWglNzL+rB4w6YEqDd3ZL2EzyxQUVIIxpkWeIHBVDcpgp/7FBF8sbi71hQdj26QWKmmoAdDFsz4
fV9utkKMUzd1nafC8w38uHdRHRGyvJRPrgOdKqnedYMHElJ79nJj+T+mosQcvNS5oie/XzrJvxfS
83wzRk+2L8nE9xlTUj4o/BM78AjhqNdRdxP6Hc1A1+CxMMJXmEP8RG7LNn/fgywQCr9Ic5EAWh4h
BFx+4xy+dIFY3frnZeUYH3u9Ucwg6guND0GM0/K2uwG/El1lImNGtEtKLHXQoYeo/GnErHqbaueD
gZtK9x7Iqt6S5SAV5Fi/zc+5VvfJgNASKcy60DpmUroLrnAyYH63oQfy6cC4ggQjcAXt6QV6M4Uc
bbRSbgEFdfAcsO+NoaIJiUCtK7yJwOJIaQBEBT/UQs2JshVoTuekdLFa3s1auJsQKk36qko795Jo
WJSsBhX86ECM4EqoKQ8bsE827UGUq2sbFXI9QFSSjLpzlXs8sgY13SEsh8fc//wyGFKPKSwoAOc7
MojfhtWwXqij1dbbOAKXxsfmDJOHpdK7yLvcO4nyYf76yqG7DAea/kog4Gn8DtqNhsa99R82gtso
rt16h5XIHLGqCOFXQtfym9AzLXDlDdMaMBJwD2xFPb9YKelp5DzmzTqCXQlVBpdp8gun42QYiicL
ifg9HLHSgDQi4vej7Nh8HtvLXbB3WBB9QJUuK4l3JsluL7yAaDhVWRbRuVmslWU6wnyeSmrhKtdv
mn8fsGF+1lRqBy3JqZHtHgGt6wLuOpXwE9NyxFYCp38Bn/p4gUu+hwlc77R5+hbNXUJpvAACDNYK
lLZ8Q+MNSs9PLIGQvDOyM7PR3RNjnWXrebEijPX+AvPscxKbZe7oBQ7oVrCPpQUUsPmFUQoLUMJi
L/0pL+FOU+1UxpY/ye3m3FyNU1EC8Fpg0KGLoaTNKCcZ//FnQHlytcR9e0q6flkrczHDdimNouSn
XqmNaG3KupJ1AEiDBDkZ7xWULGsFIQjb2VJwBthWn0GbKehLQJA/IINJ25elBxRToRPAfTH74nbE
NB+X5c1gMqRFOGuiNhhLclLXLnKpPxN7OiHy1DgLPFxu13+r+Q4vdGBWw22BCWcieEOq9qr9w8lC
ozLa4NzWGKZSlPHwB6mxfgKSK9r3Dcyw+iQH8biMsVIcvjUtU/64PZjK9PM1RLiG78nD8e3f/tn6
IPKwX7IyvFp0ha9OsvIv5NAOF3Shtc6Rj73CTQZPFQKtmXqHwXKitsxEJFHJbPos9PnSDuGTh2+8
qEDi+ERwCobtBERLzREQslOWjL05dsFHY0CpdaXXwdwNeDZQapreWbwCJHgDqr29FOFKFJFU/v0x
GNMdGRYSx1O8qMM7nn+gcM8PQPdG2djRddIAUye/3jOF9BrIlHwKmBbdudcC3hk5PB3MUbkkQ+tO
b26biefmgq1R+4R90LwdUTYbRxF/hX7VTksYFCzQ2iimlgf6ixLD6TGDY0UwpWe8lGtymUnzgVIw
bkJ9Xrqo58fAmUKBcnIcaaZ3SB+K1lDS97j1mIDV+uEs0vKScL7+YukQ91+nJlB21g1/P/TF1YFJ
FNO5SHwFa/nFqL3IQFIy2iNn9VQVHGseLXYfsj0jf4YI0wTwr/owYAO6Y1YWsk64NMAmMT2zsPJ/
jLYC0s5agMSzfzTsAMZtr4K8NM6fJ2ioyQQfsiCe2obRlm6cyF/vclDHu17GOuv8+S9cj+ci7Dwe
SDCjKzILDi0dLQziIr9IkCCXaCsAkvJWWyylj/1H1+dJr/bd3OKYgsA5gxywxAzKoLWRLNCDR2rB
IqubGso3Sj7PmVL3ktYUKZSUJmSMY3SF+HFC7Ik1w4iMHlHM9xImPobdMk7ut/0emFQ4ekH0e8Tz
A7l1Q/7RvennSD1cazD5/sjjm52vFbkq4Y+9HDQdEEUne/CGFzMg4CgDvsRF960tZkc8rKiCGC0u
Vyd/BzbZBUXTbk3vKgKeVT5b6ACmdHjO3hI7UDgtRV1J8EWYcQVdQkbUP1+Y8tA64mMdLDy6Ky47
XpqMw7PxlsLIJOQvMXOrp87m6mKErMTSX86AIHwzZe7K7JAoO8c7p/dAOegB90rPHzkQzhWZhIpo
YR/VIIlF7dzgpI6ubCDZ/URD+6dZPHHb/0ZB+3IP1/TTRMQjnrfOwzafegbMwW1LV+tXVGNHuD0/
pqiO5hC2jCU/xg5py2pe6R9wMdTskLMqVwZtsGnG2UTCb0vhAeyNUwc4I02HVgPV+MlY6zJLYpEE
px1m0WDJuzA2RNieQ13IVwiYCFmTFiaklFEOWtKBTnQ4TgKt1hb+Kj2LbtkHFNilC71Vd8L1oAjZ
EgwaRMy5OF3DF2gyhTLxTIIVhXzWii0jfYM/xuYJpBVbD+S4MprAxvjnaCxHLsJJRsw92A2RYdV9
4N7UKtyWp29orUdjOzP8p6g0hGjs/vE1UCij6eKR1843yWIK+Y0FTGvPo+M1P78xAU5IfMqNGyT+
WdNdT36yAXwF28qWK7NRNYJNEXQqu2gvSd/g3u3YnP7gBeaAbNJMAYiDYQxpfjTx3kARePEQAamT
CNX46zETkw3dosqubBLxBezRo4kUM2SD//1iQo4G+twT7KMyh0ueDhA4Vk2CLzBt4efc9SQXD065
F56f1UH4ldVmLEMKP7OBZwDPIucaByowwFu47gNR1sPOZv6Ox85zxUIohiygDvbL0oLMPCowAWZc
Z7BLh48iJrF52PLac4sR155o+S7nKxrNlinLtFwfhS1YWHXdAzBh7G1+rjfQSaHLbUcuBcuDMWcm
9yL7N5stU6/c3Jb1K8zcth9Nc8BfczVoccnJuf0yUoiOH278NeYXO2lxWtE+VbpP8lREVcv+1avK
VkVtR4ArlZhwMr2iJcwlSGjpmPsNv+aJkOQ1OtUWGg6OCLSyEYjxvc5Bt0HzjkY1oE1oc3GergcV
xMAHMfzzhdgWlXTes2rGbCjWN/cplgzehEM3ou8JnB7P4U+1V0FdOrnkMt8mK1wN0Kf4IoQek2Rq
XL3JV9eVLK5bNfWJUJzi8aPCKwECnuGfBD5Pvw8GDXSPiTxO1MkfeKkn0kZi1os/wMeODzZiTT55
Jqbwlp7qd8JZ5FvoACwP7kA5p0H/GOX6/sFXLzs59rCcSV8SO8c0dojC0V9+TQ8wBqTESv5GUKbZ
RnUJZAc8kK2n9WxhGB9FI3NVs1JPCYzqVxPLkZ0r+FNEYwpugx5YtZ1P6lp6Mabs6j4cEzilah9v
sfMohFht9UIHifbrNeCuzJBq5Kw+nDNpJrtPyhhQU/h1GKVsju88Xj7PVumIca7qH40wuHbBmB6J
HOkqtoIvWRLvJe3kyGX3TEqT7dip1qTiH1Nm+06YF2YOcZ3+5V+EicWJ/1s/rJfzsZX0lJOsOwcj
c5Ob25GATYcVA550xGeV5IPeR3WMHA0ndsUR1fqBaMyUbSexkJHod+XYxDtCJgvyLzzoXQwx8R2v
+e5mHjfDgqYY5VH9us95kKtAOHFY2abr95xpbpEhc7nZcRdQuPoVS443CehXeEabzCGamm65B1VY
OhKIL/85egpCnaprLHnkxI0oo1d5jM5pbcCN73tsMAw40B99Fs/2v9QDNDQ8E2xeYChpNDpKi48U
fkNkq0RpyMOxvPpogtfDHgMBV4P01VDu1v4AEId7t8K1Pg5Zq77Qa0qads1Q8RSdhfexhoh43run
W/viWXsE7UCAcqKnPo8eCs4T2FDQtRA7Ffxb6/SN/HaE/vZT1hNLjh7VeS2aRFot5PJr99iE6OPB
tYSqRmyP8Wl/q+LO95GclLMSSRNDGqfnk99G2ph+uB7n7WTPwYs3Vrj4Q+SlIJMaBamujtAo5oEJ
Zul4fHPU2vq+AivOhQ+qQnZCsmlbvXYNU+EawQjH/YklrUJFuOvj8TaMVP+XuP6dL4tPNkPOa8Qg
C5oi0Qt6J3dkY6qqbpQYalYk1obc/V+7T4COeQ6enQIQzpKJLrV8Q9Sbke+orfPzA+WHVZBpDcW4
FhstR3LKxnNeWQ/TAJYQM0OFkQQZn/QLWwhqkmNNfyAQYEzo/E6XyfQwgOb3bkVcAVL9VOpprreN
KM9NApmssSRL5rZatGVqdg5zaPwltffTvKQL4BKYcVqtautHnbgpizscolnDjUEQUbwG/FcdalI1
ztK0Ss9BNAhGXy2VQoHJWRFIJyAISnfBoIB8wjRYVRmBbHgnlTOdrQJKcnftzB0DLdEPw4RS68jK
3orRV2BeAA4kTQhIevc2R11BuEg3HZq57tf4X6VxGHIy5aO1q/IdUjfvixOhXZOJmM9DcJlFWEnI
OfHFqd8wXxGgwr011Px/K4R+m8soDFU/eXYoLR8Ybiv8XSPYsgXmgACo9WCpfM4sVtMpzn/Pcw2S
n66OH4m1ftw0jLI7u5XGuSvs69mbcQB8qbmhZMuIcxGDKSmQJvhrLxGNjcZnPPPoos5aS3jwVUGl
og6C7JRy7iCHVFLZd0m3RsmDIVJ/3P72iMk0pDXBzOVbIsyQ0ZKeiJ9SS83R1aGoDQ7qTPR8bc9m
Stx3wvju5zN6UQYg0x+knWAiQuS35Nl1JkTj1jqb8SdHX99sHjzrZVl1Na9wW1pYuS8ccKzoQdTa
KxkNQqfOUUZgk15zjiJwVqYNRynFCdxwcBAo2BgkZXLc7yTSI5lVxCXYfHngM1MEc2UuS6+yHFG7
r5Y4k8/bY4rKDJRfcZdoCCNRI1LQbCddux1DpSYA29wLwXYysV0Y/0UUb5qgV0VzWhEGwYOBswQW
WYPNfnlnLytiLrJvQ2VIcA8K4e0VfdBKyB6MY6bg6v4vjVICd4pP92u3/qmQkkc84gVrIUgz2d3x
dO/M0/28+ebHUf5nJ2fjRj/KbAlFrDf5RdmKwI3qF/b85DocjRQGwM13DYJQDehPhc0GEQioJFo3
dMLjavOTXpoKZ3LMckwtZcgtsnTcFu6xqoJynIdZuctV1goGw1v036EBc4iAforLZIpLk6Ws31by
mNTs8JVvcvRKFfSLbsSVTmPIhnvNG9csymsxPS/rPK5d3K4ODRKuwUEnIW7VWYSv/4Oga2cNQceU
zALYDpvwwH4m/FKGJGn96E53BcP5qddkrwtqxnwEofn5GtByEclU5kfTp63/14+kyx35IPOvoY3D
Sjw/JcwV4MR7BxcplrHjLuHJqc4cFAqt8PwJz/YKIcWicfWrjVgB6NWgmxCqBFEnYy2Cg8+PYGAl
Lo+UtHUvJ85Hf8KZPQsctSh8EeCS0jjxqrOgrGlbH0oDscGAHK8mTCMtcXRE+uzy/CMWeNQmsxN7
6HPwkvXOQcBved1AGVjN4YOjkVydVpILIne1BkkEIbKJjh+DTWs3dsaw9lmf9NvuaFNwxVVidN97
hgv605t+Z99f9yyJ1MXuzw5/bT0Uh1WtIVywJ2LRcJt9N9Z1CX5x6vpt0ZE7bzZGCqTBcp3G6uTU
reDFz+aAbZ6+xx0oDrR4e7hrF2s5pYoj20WtVr/0KSozKgXJaMvvRRbPwEvu5X9UqjQVuEQ3SvNI
qG3GRFX6yTyx2pQqg3/1OTC+ChAYaYGsuTB/KlQ4FlaewQMlTJ3dA0Yugl30zNrlxFdkJsGFwNME
mrmq6SNWEqJl+yB4xViaPJNGCBE6ABtfBDQgkgXwc2VaiC12/YoTgPDbVXmraDTqpW5IB0jDv/te
4riNBOdfvnKGcceZGq+Hiz3HsNr5gJSergn1WPproLSHqq1ATfUmLkhLoTj51V6XYB7zc9IioLUZ
stTuDj6odcA6JgQAxO/Cae5+Wqt2Kkk/b0kGCV8IshL/D85BKAO/kvlurZXIo61+FxKXiipN6vNz
GpDTilIyDO3FtnAjilOoAzhxB42yaYd6orSET6TR8mo81Xc3nmMRN1PqaykLcWLhP5xLLh8X5XEh
Lnh+A2weI13X0oZPQySvwPaAbSMBXQ83A+Zp/7Kx8CTdlE3i7C6Cql+Z2LnIgFo/W6HRTv9Ea/f+
eZcjB7zAp/S5xCy5ptLedX8fSLlIE0pv2Mu2D1N4r2Hh7he7+eyAd5QFmpHHXwQAiLtaTlFLPeuj
Lk8cf7RMpNRxy2VlunuRzesTwO7DeNGp5DXwYmUwlNkinqG13/ciZQI3tzOGTaaYVNMErASUCU77
CZC7IHRhiskONaY6z6WY089mJbhTI7vs+9rQ3dU8lmWx2ty10pkTbhYz5qGs3xDr7UL7VpOc77vg
tyisyPZyKOWGwG+xtConDFsQ6A95Ya2AEGC6oHylaWcyAyns0po0Nv3HyieFTjijIVl+PLS66K3H
P+LYZwLNWNzHB7cPI0JlfoZ1WaDKCZngNutyfvCaiu2LXz15aBmgvyVrkpepzxvEkg4UMmKvVTIA
75SP2I0IE43biicllsZBSqclbjc8ZIhMYlfHaexPUCn2ijpVmoRYHruaEXYHF1fdIcjp+cQglA5c
hJTFjbBSjFqfjJn3zNj4tsRBSPS8l9+HjRD1K6X9C8h7+vP50OH4f1al0/HnOo9NGORLXXmBu3vQ
apEPGE0ajGIVabYdMXdDNHdOSZ06oFNfPCihSI9c4hXNLHHk+ABj63le2+rEC03eLEdSSEIVwdny
dmqspXpxX8uJOHWVCSeLGWRh6f9zFC/yNP+Lu7oq+Nm6IW4V88PB38zEyOz51zwimpGNdIewqoXI
qJ9LAdC5DiBHY1x6VgOL/MFDPVuE7cp5kSby1whZCj+7jH57lTgTwAtFBrOrbtuzbHz0Tqn4Y4TI
DPFM2O619DMLLu1RU8wYNzfCq+v6TR/MuWwXOThIh6zYruqYqiPp/jJNAmMvgMTiaSdhJ4eZ6260
H5PNVH25wnbmRQqyyBFQvmrv1PGjG3BSyuYN6E1TxXXf06kzMicUret9kPAicKUUV3Tcv53a2t9T
njmVlkJIzTjY8sqzRNI7bCF3Bb/A0c0mQRn1stSuvYZyMe4x87qI1FjS36+UHZpZOSLOOU4O6Jhu
a992XtMmVhPKpEsPKDn2DhqxUAhAGrTjgouWeSMPvEKQ5O81Tm+z22KYtqVKHBLpvwXAiKNeU90O
+OjF6+gahJyxZkhz3NZqW6PE4V6JFOYM4J7t38ABjJ4y5CYRwVUJPolDXNWrCrTWtUfMDQWDJqQI
30mNWhRCFg6RFsezdbTA1gb8ePCsCuMSkYNx8gGS/nSXQQM0y+8pRJK5Nst7qExjvMEesq5JVK2h
pizU9Xj3i0TkZWsLclWkKarRervMzjU4+9vCs8jvrEplUtTPRxyCHBvbauXC6uorlXHoFzH2En5I
mVtLMQXqs8UTj8ZB0k3EESYVc4VTGfeT2TgyB5Si4tBSFqQKHTdNxrWfZOjezZEJlsJUbD6fzVjg
w0xwoAQ8B7uPicpKuVpWtiIqmv5OcSqrftxFnSA3F39UnI2JFtKJF88BC3kjWknigFjURxgU5R03
27XGT4aUwOJUpi/n+Gf/oqFzdmWNP4hKEKB9dRwR4aT64X6hbCp4NgQWeAThkuCHmUq6mGlaFPBW
P/XmFI6HCczEDRWIUOXFRSYz8GGi1pTrPFO6j/lbKXNI2msI9IgH/MFqeohTXkMFXaPeJzJViHNm
9GNH45CJMY45UmlqhCjcb4kifvxCu63/vUv0rcDaEfOaI+QKBSb/orw34bCZtyjdjw1NgIutvM7K
KsHJM7M3YosGn+znUUrYl82QEXDTz+gfTm+h/4XaMElnmlaxxOgmvfKLLb1l+CRBYX8F2yt+r0B5
Qr9WV4LTy/i4YttUIxqH7Z5d7eFh7OkAGQu5Ewg8X7Wl4Vai+klo/dYsfIBcznfGh6k0fUMzuDIs
k3f4FOWRbmKjh9MNtlpni64KJYGug9ujczuA/HIdmyAKqM6777BdFkdNvWlf5EckGATKg6VRZVZ1
e+NH/efBN2ITkEg6XeSM7m0kaDYgh8/YuskoDtDiyYut2QMPDGhSa4LHDqQAFj2vM0E3k4aGnr1u
fUEypSDyRKuQ7EHvslRgijgC0Kiz5dUL7UjtNVIt7Pw0gELVMx4jYms9VWB1ntVsHGstrVNzEF90
bMYaXIsAy/BkkGZ61OAls+qncOzXoEJXyZ4SBQoVwuF4+TPYzzRT3DaI5epEMDtpcVzJhzth1zgk
2XqsKfnLhnmkKX9GHFTEjbDkRY6yRq+x90mQFckgG4KQZm7a9nlPq1oeGXyq2e7tB2i9hFVMuuwR
79L9v7DxZz+AmFHa3CV+dICgASsAbEtLQxkTCc6GEXr9CkFFGcj0TrlnnRN9mffr1h3wBs7r4etn
bsWUvTwPgy5Z5L9gv+uiLoVroldyw1B3CZtGkje0upUavCZN9VtxQNmlVEnqgaH3Jdp5cNaghr7V
KkXwEPOjWvU8KmkjNFqpOS+p0mXM5kHWcsnx8a4HpPv5ukZGuae6Cs3oU2nyn8CzrufzZwBTZO8k
okWGfyGOv57nv81RNfqSbwiKcxlOep0SvWnSHjw7iRCPyt1eYBVzFOAHNYkQ0h13a6fDJAnoboiF
msCAiY63m3uMXt3018kgg/kPQxXgKRjKu+7EGO6lJKBolO0QaSwo45TckR3MyxR26/UJCs01lcix
GQnZnQqQhtSyCIICJFVtAPH5fNsQGVMMeXgh9O4lmM6NzpTO6NhgcWcujEbGB7V3LwxAm8Mn1SQu
Rjc4j3odvvCVPJqg6wLvDQyNr53UcjVcIaV2LqPB0ntmh7giRKBL5223DPjuGefZEeLbO2pFefQy
9RB/FwFyyYLkNSAqgpY+PBUD2cfsndJ3fS1B4m/l+Xn9ljwysBvu0Cv3w23WSS2G8QHqW3FKRQHv
FvR2BKhVbYkZ8RKidP3eBdqTuD+HAFkUaw2oaGfK2cFDYavgW/30XZD81goQgm25iWNNVOzjs8C7
n3DzlcSdS72jWCmlsLjEqSz34qRlZcNLFaoYmhm9zMgwEyecWSkzsQ1XgdkMAvLkv+NxR5xzTqPt
2Jw2R7aMbzJeqOzzaEjhwZxofQk66N8fnyu7F7F25Y7JraoSlNi39X9LdlEGsYFHU67DuYnr/HC1
jfghnUnGZZxK2qXMFZV439dFb4VTnLtFgX5Q2sgXnnvYsSYVXCGnjIGYl+Lwcrje1FqYefL9Hfnu
5c6Oo9i0AdGUhZio7YB/xKdZis/2t46Wrh+iwFHeK25BnCO5WThsqaJfMmfdjcT0aRqh1u6Sz0oN
L0kNkeqVlHudIwIgVULGPzUjO7txfqyE+PDllS7tOOMkQt7LLLAbNfLfL/WMOj4YvWPAUDqT80c0
HiHVbqPe2DSD5h2VSTY8OdYzGA9pYYlAySAE8bJMYIq8l+iY5tpPqNMTXNXIdXAKwm1JyEUBMC9z
ket7/ba1B4b2Zs1Z1M3KTOzhLJNU9WeX949IrHdH3/uf/7RThLi7wtrCm/M6DUDth4vhJcYl/4Vz
l1WK+mNnBa4o0qfNpcE47Z/BLf56xVBktNk4uhJR3LCv84kPY09MJsog5+za4QwTYubsWZEfNuct
9wtBwEPQWYZqdN85kOzzaYBcC8Hv1TX/7N//N7tvYCxH71Yu+r+HIp9VUP25UU8Tpx3HD5aP9M2Y
6g3Dpt4mn/5fMK8seg+zM8rf0Fw7A7Q8G59pylWMOUX6rTLcX3/9vN/ByRsYb+tYWTV9G3cm6sxn
mAJD79Q6v0xFXsfIdSlukTrGa+NNqMsO7GJEmJ4VBiOlztdilnwmB1S98j4P9I6Ln6ADOgBzyrT0
6iys4qrvRZLoOk21Q3stQ4LE/mbmrUXQrCw1uv6V0NjEtdlNjOgqeIvbSrtoJRHxlTJyOHVPodfk
vrJxmy8NNea24Jlf27d34VQzlJRZPaQAXZSjkcy/YKUlEzA3K1+iOtk36v6w1GapyDeZ1NuQast3
7+v6Ut7UUoeIeOqWGIkgkB/a6eJs3Y/0LYbMbgpmf0NPE5Cke+ySHHNIM3BXzQ6mILUE4mcG5B0E
iG/TB2EnENJQOhau5GM9BYToZZ5hv/ATQikd2CW/HEf4ejvkCg7zVsaSXAbei5M6fCS32y1EVSq7
7jor2vZF5KevhZDNE5GcKuT35IKBZkpicaJhYZvfZdbxuJzpU/UTXnjCmr2x6RgUq9InNOm0YM8+
QVQxo/SiwmOve6uBYQ4PHf7wj1C7h/GazOiikBMQdCyhGvHWVvTcZybw9P+Rafza4owWRoLUCGJT
P/dkZeu3OW7KVI9nYaWeGSjCS86Lednd06mtliO+BsY4WWov4nyYCQMJnszfsOYB9s5w72LjUWdG
+R6VLddrFjBPypCxdPW+rQEuXf7vaV6+P9nFOzIxPdc4VAFyFZQzWDUOL5bCPRUjxn3mdPqcI7fr
jQcvPsLfqfzZJHRMf0TkHvIbFiAKCopeLDSFgwRE83k8ddbIUwaZNCQ/iY09SkMBtai9o26Ddlv9
6H+sds1uybVXB2aZl1EsPp1B7RvC6JzjuS6CgpK8ZByDTx/9Umrd6Pws+fOLTzcwNIDX46yI5pli
iSZmFfvCrqf/tBPY2TPEJE/GdbDGq9mDI0A7emzFEOJQhIC8g1xVaCYYpkpoeOHTJhJh200HUlW9
s44hWkbZS7v06joVczwjaSuUUhzAlT9ya1QXdSXRTN3gHbkLgomYnJR0Ssk22IDKdraNXeKBNoCa
45kozvEOE0eJBXDXk97xcM4BN5fNu2bPZ23zUAHeKS7LVddiqMnmUC2Q8fVFPzgMdqLiAouqGit8
ReRyL5k9Y9YOxRzsuulNP/9ZsmKvVbxSH3VCtE3JdoS2Qq3WqxXOM8C50J4RcRSbSjzRghEaLWoo
Jl9EBqSt/H84wDczdvxiiX8oFS4ZqxtPQMZOvDGVGVWTb7J5jzDVGM0zf1ntw/+PxDRD4oteGBYu
rxC1Pukbu/4G3GIRO9jgN3NMOs3AlWI3wip5zvH+yK8k0nZEmPh/vYZLN/dUWDB67P7PbweISdp3
9BFzOLlw5L2qlWequtiUCraHO2cuuiKRsLpFVpij7BVYeEFJFc4Tj3IVqohTD9BcXRdSZFTXXzHv
LjRmLi94nYlPD46TDCjHo9qj1bsYoFbc/RHbY+LQR4gln9T4CUj74C26KjgzUQIfn5PfPKUq9lse
RFCjslqDlB25fHm/57ELBY5ccAl/ve/jCVx+JTgHPQo0zoxJmrFrMv4pbSntV7H7BLO7EyTODJ1K
g7S4ygBgSjOL6bM6qAVKCeKmeIrLiWEQyidsEf50ONmsAaCoYcGC/Oxg0fnD56KfPRQjdyUchvkh
waNCV/yf0Gf+AUEGvM5u01Wz6bjqrwzwRKfP1y3Vk+Y2S3fI+p4o/L0F66Y6Zn2krS9r2bJp3Iss
K9sPGjwFA/WWfc6rh1MAPhUskBP/H/1If2Pl88wI/HSQSIwVPH2VAK7vewz1CjwENufngxyXsfKu
nC7652lbM82u2cpn2PLQaJExJE2wT4IOI1pDt18gPSWgIfHbQP0S4JyPPGTkvVmlpVKOV8lelzDL
ku8vUosxDcYSuFva0JTqXED49e5x8Fmknzspgg9HOX0wWSH5inFVCeGg5Ql9csi3oaZnPzt5kicN
9XjX59dHwa+FD2b2obDvIJY8lxMAZZU+7x+0sbWehwws2/z1g/gN2SsrbVa/m5Ppo9Sg5YT3r+Qc
YapbV98C4x5s/vLB3nDcujeyBzXTMjkPTgpU4APGxdo9eXx5GiBJdOcUWVDzLfrZu0OY8JJK48kc
DJn5xDFYdWH1fi90nlSLMJgn4zR3XSrrWFsiHJJAfIdjjKQrlyex6LAK8Ug3hoan+Qp9h2UhNw5W
a9inFm7VS/2ePrP118R+YjIFBk3B8WxbeGaBxqRHhvnbVmQXc+0Cst3o1Ewczr566m+WQEIHWjfw
tj6AKf7RKN7xkvaRMHohsFAUHXmagYaoQfKfbbdW9+CSvI78Fgsjn3KFLJpM4iw4fcaZfA5AizBt
P9DzkIVrKZWNjtbYoUT7fb6rXmjjJLsl3MKXuck5Hu+OjVNoFD8EZjoOc+FogGe5lr35yRdOrNTJ
XN4mAHotvdI89Dt5neY2dMW5aKvr7wjI2n6oJka0D2NTioCbOpJDxxlDn8jozAI4jFSrCnRairfB
Sx0q0nso6iqZbD0kQLMQW2QpRPaY3yjXHfZODIJjTSQ1FuFHfixWBJbyPHfOEzp5gN1hzH0T13gr
eACL3dPOtTkENBG9EPXKt+ARpztPwKKx6uppul/XSryW5nVSCt6OJTWasGp1Ldr/Ltu2+/JU3C96
AiLrHLN7QsAfwtc50ngo7bGCS52iYXCbVn1JtAhJiw5nk35WizL9NRG7KJ10S0j7CZlTthXjkqcy
GXjXpxLxvEwcOiHxAZxFXx8qzmZK6mVNyRFdjh9Bh9VQHTaZpwyROuGDUmJvdXpY6oe548plKUAd
kzQMMRzYwMfYmJerkRZ72p8p5i/Aul8QVNA8URL0EGI3NByr/0jU7Pe9d8UOqLDS0UvFqS3N/g2I
vsgBW3uSECwLRIbgCkKYdISze3B/reNFroCB68RHuiXzuYRnc2r8viEugUpJ3ovv4g+L832GItLw
L3Hfc/iCwM6Vx80Riqmi6lzTd5bMNE9VzSZbDx1t7a5aNU8U0VTB7tzMP5nnI/Pl0Ux73Pxi0/xk
FjhigJPY0kx2ELd69hvntaFFoIO/vBT8BoITR0UnHK1Ri/Qw60jeIztT6KKOWtppJK3lb8b7XLlV
gY0bNiqLDYhDJaQhsM3w1zvb6BKzRLTwsxDpvTGnkF2avKyp+IZ5qjKHeKPKTHFqX0GnPSNk9KYp
rEWJxs5ew65vKn0HkMg6UhDA/M6D0tl6VufgskOhqL9xqOCmeVyMPkYJrPHnn9Y2To75vwmAxA9a
UAIowMufhAyXv3FDepoz9iYFwyyiBFoXtVlmqxDgaEHnFFV7i9ejHYg0cHteHF/8a+S5sVBVjIou
X1LLPG07PwhxU1q944h1z1QcOyWe3Zz+pc5OWWxmX1tmGkPuAhxFykATI9C68szMd2Maa+HUQXfj
HaOUAeF0AjEFkanivw3apgvwvfrXCUQaIyIPcsP/mmYPKBf/JPlW/VcKHzCvrsoKIIcwIne5lYxu
1dc0IK6ddVdRlCUdR7zSPzDLA3vmq/4xqAXQZX9BRafavOQ4jrQpQPYjJ+z3u/cSmxFAE6+PG3mJ
ETvccxr66n2APpvnJPTBpuFfKzHGzmAcIIgdnDp0C3tDdgtkhEdHoc7M8v0bZuaFreUgnjhewnbX
rW0WIL+CwxBoYbnPv1qrA8MT54yG7sx/LAfopnESLBYArruSVZwRJA5RWAQvQO0QTpSTUUnjCM25
FJpxEBFE0nF6TccQxjW8T71uJV67IO1lMpGQ16BC04glx+xLHsL+6rgBTrbQaze8LFwgDZuy3lKi
N/RQgyYmkz5o+CZcFeFwri5699EZVvQarX6uGdVK2YVFQAuaE/HuMSxVNv262yTjDhz+7SYWedOK
pswDQWuf+2zbgM94hKhj5fGsE3EsFjMopG4vpos+GqUFjjFEeXvEKloiARESyFO2p6Qjc0BLeJND
XZenmrdSdtXMYHY25i9ETTv166fjZPvRXTA2WLLnkbjnHHWpCLKPOcPzf32yncLqd6Za3W3NB+Zt
pacNTIAzqizneobSMcyPeaKX+If+jyxXCGAjsFmppTFa7/BXVjXszb6fQv7i93VxfK2v8DsLtmM5
Z9eqTmvzczVdqO0Jtp3mavPejyWFBnLgB43GnXZtqdybAb0Yxcl3abVwkuLzOvpdVUdiSWC9Ujul
1sBvfNqB/GMWJ9HlP5Fh8/CXaKgOLxj8Wf2+dO1HqyBqnECkG98F1fjCQlQqkRNQ8YRmWHmdQPb1
DKKBaPx1lZjzNolZYgspGGj2xE7zCIIsPTVh6bdctjfxmNtTyRaHW92/b9CjUTyV4ifma5St9uPN
ruDhklWXEfJ61yxmnZ0sQn/HM94/XZmmT+OnlOmnDeYvLaX0k4cNYejxionCt8fdbZnI8UzE8WP9
+9odQG/0eQqXX8g+vt31ty/n3cla2tuZ9gbV1DxxJc6JuDvz+zs3rtWNo9UwSJK0xD3D8EjsN8Ys
ba2g/nVPaJdf5XUGfIyN4MSWHgagbIlzBnpuIDn2eEee8OOzbuU3kks3OEsdlS5D8V4yt1c2/tEv
cYbE+zdo4KqZ/U68XT4p26sVIqq6ISuOoIstDlkXLRId9ataxDE9xijNqru+leV9cq3nCTXFKSUW
bNGiAcmCD7aMdJyw84WIOfSSO5fjA32ycMe5IYU5cCrHVnWJWnLS7HZFMzyvLbzXmdv7GjkGHEfH
EloDFpxfxVyA1wpJdM8t2UA6BoOXjEZkRHxwzgyrSDZ4WvedUw9sXs4DHtYh+sarQzUZ/GTQcfAJ
YhVnZ5o+gr5SCrRFmiA1ZDSxx1F+XzdZyehiNSAC5ZZ9zKfkfkhAmFgutDWHXKiHVnaWTGqO+cSJ
mu0K5lK3lUS51brjL3D/u890IL/eoXVGaci4rVf7uxJTT1i6tUwwxRkZNtMPMvouPeehQGOlsVWA
UXW6TmoNYnIrpkjiG+ycngc6+Kuxn0LJfWWqc69x9S44/tJbiQPiPLSmHuuKhLZqV7s4Zdsh4gF2
ITY/dCUI8+mszdMFNaEwem2YQYC3GWqhyLxRlfr+XbXjQxYhRUHEqBrVM735GRTHAJP9fLiktHXW
IdQVT9hAFEbANGk59qQUIuZEJSfzFybQOdlEOY2upXH/R8vzJBIJe9+u572NmzfgsWZq2iVKZr+5
V03A8L+iBJpSr1zRei4vnKAfePbluupeEc5BYFimGR1qVvnHvKHBOZCNmQhe4xKC76QqhdQ8i7HY
VB1WsJ10qGizjuHKSRwIl3iss8+SLFAXhYlkdelJZkYfH4gsllHtufqYeapHa54+kNxCeIR6NXBf
uPTm32XxcbXqcym54lugiHv7V035bqXBet7Y6ZTk7sXdos3i6qTdshk6m4RhMi6vSFufa6YLmf6j
wdJAAGMkTxjxJCvkdtpYiNhxTMo2YTj44pdMPhfemDUM1zb/LjSaDomNYWwjpEJUvzN1CpHeWLel
UMhth/wGr6FhsFmHGD3qYu7ezf9B/GmjGYk6wmkKjUkeJ3Wc1yS8Q3kEQ4/8XhKI8IjHH2/HIIRi
LYbc++DYXEhGk+R1GDuCacGZpr6tXp0QGAzEC/Dnsukr/9NPYEqijPY0y9PWouMB9PXbeaLMUsMc
hACX5bjaq3/hc4QZlz8nsVTfJDRVjyPerlCcumXVhRlNQi2k0ZVszMLpewrurG8Zw8penyGeb1WO
tDt1fCOYPr3H8LBlkomU8pHa/0hCEMJOVFE3VEvYXkkROJ0pL54prqnP6K12ccbPe0zfyJL7wMk/
05c3+ymwMCTajph9yEQsbNmQCoRUoviZal7l/sPOkrgTyAb2pGbbbbGYfQOwmgHGdaKfTmHDqg8N
16Bzq+7yL6OAv7H1sXERmfe5Ml96nMf2EF6py8fzJS+aDOREHPLc/3HfWs0oT5mkiF+W4FJwTDs5
duD5iVYCP/xm310CIld1j2DFkmc16VC52lplIc4KmVuvInFmFYeJrJ7FfKitNimig7s7aw6FdMcG
5+8671WDSAMMBxe/24m8Cov88XNAd3cFe3GyywPQVceq0Fw8sZbwWWrXi0N1qfum7E/oxlurRuyJ
frRyiNm16e7g60jkGr5TdGKdvKAKA3/q6cMY+p15d7JxzJIZNtZpXg0nQ/QjyuctBf6M82UAitfX
QNg5V4gqv7Z+hqOh3RGOs71hCx5EFOqAh9oPC+olDf1fV6TfPxWAc45mFmJN23GzdZqSM61FSWyK
4Ejl5WTCLZyPDLAKQiDlEUujQsCWP0gZLdM/MnjozjyR+0COJ3ubvZqful/j3vahGLwh/RJeIyB/
mDbiJvg3hA2BGIgS6GlXePYzhhc/EqwUUCFY2TNJle7pLfnc+Xay3xDWDn1to704Bmnq6NwQQQxa
p9G9UgEEwY9Dh2lM3xcbP14rgKxT4yzZBFoqC7Ieu7zXyfKsxrgMM38Pgmit8bwM0yk/drY2D7zf
L3teU94GI8CiehAAlaqOUViAT132GxSlw7bnaglssPVEPx/x0FjZ7mq2tTU0Lv68qjTwMkwGgse5
ajt4YXh5uppB0GB+S4Z7H2kKkgIpAMOuD73wzk8qeIrGPsAPivFZItt69x+Crghh9ckYkVHN/gW5
N89wrkckW5h/Di32zgAUL2hQeCrGbX/oT3DVFOCdgtNI1ZJH/074ItbSaewqWKx+NiQ5vdbVG2t7
jVx57IShUZj+Sn/tY1jZO3rYRm1xHi51N3MHwZGU7GwZA8S7RxbDHOWmwEQf+75f0mW+2hx+D/TH
tvXR03CWzmhHq9HpJ6wpKhUknFJVhSSNdW4X8VnfvDuvA9mdw3Ai3dXdQTugQUJzdxTshpb4kI2O
zE9WfrFmY++exzC5p5it8oRGthncZytb10ei9N9e22+ajlLdaOGl2+48DrYLW1Rq8mtoADQtZvIl
0CAnMufwTImCk5ESGgdHYq9GODDjbZCru878cEfaQApUmdG5OzqXheTo8sinTFtTr9BUlwGV4Xvt
PorQj5v1/THijYdQPbwgpel7dNVHtRGCjroItcjLB9nQbaYY9GMTdc78CB+DaTQeh5OC9jUTQ42Y
GaKCk873iTD9yrg5WR8YtQGUENlEYi7lpipf1cKWehObzgthdb1tSBxPP1jglbZq1nLl3Y6rDZnA
aY1c2OpVsO9tbQ0ikBOJ6qLvbXANBsGCPYkdajpDOXyYLsFxb+ZQcNdF5wmeGRrZKGUICTbzYx52
Ef+72ukjcPzQT+hCPqHSdw86TMXKf7G5qAjC7i3UBwhgaFxhXeCbxSsjkNiBmx63Z9UVV/C1TEch
LlNGVezakLB9lZI9O8R8sNxYW/9wLTO/YnP1dwFFD+PuNK0fq6mCoslqHItEEd942z6byBTSErWX
RMGN+mQTdVvhytgxmBOtvKV14h227ZEAF3DMZ/oG/UNIzuH8EOq9W47g9+AoctESSNuL9LtfXpyn
QOwGLjsF1btEneiyamXJBx8Bp6KAkKnnuxnijj1Nn4BaSk596q0EyNzwNJpZi2dFpCIqv+GVruxn
tHXmxQn1i2IEYMGUWyEE7UKZcRiZTyWEBd0cod/pE9RyhpVvvjLttGrD7ZRCO/BcWxSsEBc6nNS8
hUQI1JXtjeEpgzSrMdChs5GQX7Tf+qqr/+FOL6tBWlV4H9tg5uYKwt88+Xf+ysafJ85woVgL/gvH
Hpm2YwTS6TJawqVs4kPMtAaBKv2q2JRdQU26NROjQ8u7R3NpC6uy6wq7raYbOwI5Gy6DoVbLk4+1
k0mlKRYqgOCpXvaT/8cf+WWK3xQynnUk+DS4zHEToD+InD/Yras9ghkUgu0ubWYMqzQLOn0d/8rh
VYPLfe02xksxKvqD5CMdIpbFxxKFCg8ZlLrPZD6wd/mxZh9tg2dCT5U28HPNAeUwyfrRfH9PIlGf
tCg3a6nS5oRnDX4tuz7nqMUs30bpwMYVNBXoJAhm68fgST/ZGfeL+ZqyKuukamm+lUdIScJSUl0A
MJ1BerPvl+hdiYc6m8tA96BPzri0laj9CXybf9OuGF98hjpBgTrRdIxytJPmXo8IVEvv00D8zTdA
HrS4BLWSTEtbvYdxSEmO+Cfv/L1wR1ybX3hZgNb+VCNrTjPdHOxI5mCtLsN/NuZlJKgXG7Zmez18
JB5VXxwj3aAR2ICC25SVcTRxJzro8A0TGBNvCSNgWsoAlW4tX1UDZoOGsIDogJf8xJQF8W9wzlJL
eVHrcqgjIfaOXqlY2y5nPJIlldwo5Un90FRXU48aDEb1zxOvpDqMqkqorun2mqnDIwjCAVLcUgXR
rkzIV9QlgRbwg/axOgvp96NO9oOj/SUcVEHyoUAD4OmvoTDyonDX22n/Qau5vu84nplU1Vj8ElF6
7m6J5ljX7oktut8nstHlw2BTkFDOAtFRXZb9HwDx2C5peO9zaUXzv3n3qp1CtjJBOA7a9D4bxyu0
joHR533LYeAwBp8aTIBHYd8s3vkqQ/zk4Vs9WmEkhsP+3KIWVhcPwUiPiUUVW+o4A8NqeP5wN+FT
Uzk2faN9FPOFSbUpjh5Eo9FEX06/Tf3Jf2WKi4jX/5zAPA3gi+LKyNIZPmY5v4wLGhz6KoPuLXxP
2TQUijxjs3TuNsBPoROBokutHKWZswD4HVA/Xd5HRxB8pMtVVcC2Cj6yTiKkh0Rl6mm5bR6LVjIy
Y1T3av4VgfaRytjA1RLcOAg4D8fKdfyUuqMEKuj8lAcDEXis4vH3R3HmxtXwDigQ52JdjQ4ff1l0
wfogwc1Lrj+6qXXuzHNRbGfNaJOwQVj9aacV+FjD4FQshLKqdUP8OQw64UHEO/yqmCVPaezSac0P
bvVeS9DqLdy3gG8mY6pnDro9468Hfwli/fKWm4FEM9O3vMI0jCjG+hI6dVjA3ujjcp0gRw2UiPxc
4s34zA7suHzewJTUc0UTGSx8mY1cxRS1RP5kxhUWx2eOo0V74P8jrukIYZlQ8ssdfDE4I7vm3qad
WKpibcde5fq8g5csW369eWpitj2tOyfOwMjlrsKj667U910tHtZnjeaIoLWJ1Gvsq/kiNrguS2+e
azGubGX46MKTfa3KF1s87BueSw7xl9jAiwrOktuzI56quBWQXQ7sqGPC7UJ73F7qv6ynjhU7PJ40
lVIFtCHWLhHApYx2KAqJxpc7pMn8aqfTtgizhnf2RKrm+V/QWcvQLJ4ht7o5DZA0NRooZaGi2Hsv
aFUDfHr54eT4zIDJuPUv5YRK0hXBC02VW5b9xDKDRkCR17dP4w2IeJeUa2xo6viA1BGu7sO9WBhJ
BK4eLgBmKThtJo+Pt5p2p/c545ycrJolDv476crPoNihb/cOPq3zlyycU1uij38JA8b4C2DPR+QP
nAnogg1epHZEl9F4LC61rUufgvO7uy0QRiic1Tae02ySD8aGSXQAUIiy/CHfmX3Vycs5MeojtMzA
ALi8bcZAHUcep0rV4LNvlc7rOiICpSdNrZan14Z55TXKQ9VmQYnx31WBa7M4ujCVpjIkcYxJ/cOB
hPTKaHtuws7wlAmCooUjU7AlyzzT0QYd0wdzwyOlmj+6l9Un4u5zXBHNPwANoGHdDz+KML3RAzFt
ObXSZHQYvGOtSZYkCee4z8kxQITSskz9CchFHOy58nwOOrq+Jys25Jq11XUFRBYB7WXEqMDB6Nxu
qFRnyN/bPulhAtw9p0NZq3OLg3XyxJFz7LKC5aoXXVbYPEnXzl2iOat4CHdd6o7ALMugjcGOwSAO
WSCr1H/fk39vCVvb+pk0S45/T8wlFGYdjlTUYzc2IR31kLwCEImlwfNk4fmsc33JLxXc3eydlQ9+
TBS+UDUuSjLdsizl+ifHqZvHymojL/w34swmY1s5hKIC4xa0pDsxvJOjc6ZYPByHD2kE409pYwWd
XrkYEaWGZaSa0eygfwV0XCeVvp30DfX66Xu0B7cTp8VjMrz8dck5Wb4VolXQPhsLZNnw3gt4K9ca
t0cbos6R/3ip3cQcJGUZnSSIwZPmVPyBnKE5L68PfOQVjQJNsisZ2aD0W5HDL/5m2uzvgnLvqnDw
nP4CQ3jJGj+DxiDdyRB3XfaW+4QW+LMgG4FTEQDTdmIMY90TxIrHsCQvPoIcLGZ2ng+QjmaYpegb
QG7F4M29LpbfUfy78k+YpDqOaPbR2v1XrVz6fJDntZB/jmotClfzHWXZEEPZG4nlEi3xNLdmkf21
VAZkUx3QgmBpsITuAlwqE1JjvtE/IyUVKxTtINpkQu/1k4SWOHsnF4p/UiKLys9vxaKG8vUNsPxw
Z7Jaa247kz9o3WfO2Lq4Q6/x4eiMldzQweQ5gw/4gvxkdDSbm/ZLU6LroSW9Kxkhizo9/MzSZ/2T
lOLvlzWw0juBEWCsVMctwrXKrF5FrRgKZ0QzwbICiqrOpOWdoLkoacbt/isCTUPZ7Wp5eUjTwQDm
2+evoLXXbN99QK6OFusgIve+EW43hut7y8XY7XChiJMXWUIacuxel1rbp+pbgEbbVavwKxlVm6uf
Gk46hIark2kTpRMqF0Ur1Fwrgu/+Yo0hZ7hi0qiKDDDYlY+m/osrlhsmtqa/VOkvFno4vs9rJgOB
+3THOsJAcCTzF5xm7VBc8gWPoJrNgyWGeKTJEm22zMsn5MIYAc0Pj55yeQsUe0H+bKMFAF+wHFIE
w3yYrBCmINvSoWgDEgOHsVrzS3/kb3xqMazQX1YBlPgpF8hADtO2XCk0NBqcKIMFhPpJ8O0Waak2
DyvafrtbYHKwCqu63SwSbhgVqi24+8kHqCfysnk8GCuZeCU/Iv8lm2CvKXLjNol6JZXK50PyBeEe
usJMV1UrBfuLq3gF1se8KFQpX1eKpB2YyOg+EkqKdIj9y0tcRLVEB8bKiNpvMmUWgFt7vJJIVtJC
T5ih1gSX7ETzi8wPEdom7DvmCACVKNDjxeoreM4/0b9yUgklFxX+MO8V3lo4g5YdXsGLT8Quxdl3
SCwFrnALib8aSoAdWh47MsPg2B3j75FSqp6Q0jyCjUb+SPBDnADv8WihZATCZQFGX4hk5mUQ9xu4
9LEy/ZjYcq2ktezEXrABYlFR0dfe8Ggl/6wnyay9Suq8EFxkH2pLf4SVEPKEJ4/3SRAEORTweCiI
GRZmkwdJvdHWiwYU3Bn6M0LXdvqI0fv4hcNi648ny+abzJDc2jgsVJlhmNFN6yA2OhHQxMIqQldL
ufP9UH5Y9qXRPmOTGzM9xHh5U5skmZZfadsHl0y9tzfd5toz9UvXmUmTrcvkeVBcIPgQoIdrOIiX
TgeMzaLEG/6LS1Jwh6dM71IKmG4wh6fesrOKDo3x4QWoQXX3vJcIaU37cPRvcwJKl8/sA90Q+5iv
3iW6yBoZK9RVLSOi3hcUBH/Bc/uUjCVyGigE8gYw+IyVrPLR2qpP5OxNdci/aOw86oIzgkz5sSfo
n5CEG/ZQJI0V5FAJhubv3ahR8mnORmFcMTltyBLeRSvW257U/44yq2tnnHssSfcuA6lyhbOoWfVv
ECP/l1h5n77aTqSP67z8TVLG0exzrBpW7OPVOu67NrVRlICePNrj+ZaTRyNUbZ4tAKcYZUdRNQGj
SI7gxBtuchq14MUS4jECwL25aOOTDZsi4VOPnfoLFscuKFhEJezYmSsOSseeJweUZVJ6YNXBRhMU
Xh7DjkYmLFDPESvXFU+qgxNOkgEPjdm0yppFeFahhSVWvD37TvdADHim+53tSij8jnAonj9BazdV
rl3Tw5+R5G+XWYspAw+7RQm9n42qjvWBGuWMDHvnAZrVgJ3dQMFAwjXnEl+sEMlg8J0ut5XZLssM
oFjVf0NVcQJL5tv9VJ11rOrjHYKl7F0OTFR1klY54059UtJlC7/HJUNpMDd4rhv3+1uOMp0sCufX
lLRlQnNqYDjOuUDN9NBV8eEmv05a8g/uMF9FFC9jrDeLFcjji9VO4fw/AcADhgmNL9XJ873Oartr
pJ8lhdTGQA0NgyUNHB3SSm6KxPy3ReaTGVUQDqqEcnhZeEqllxx9EErjDBa+Tlg57HSe/OXrWWnm
S27obW4x336txsiw6pTUzrOY+G+i4Z0ORlE2lRaSHo9mUSGSCk950yT5lLZmnX5fMBR8PtBNIZ9r
mKDAjn2jJFpQrnLA6rshhs2icXpX57MW/7Oo7thsa0FqLkAIy4FHwrE6gifeownmlOGZlVT2EYVu
9KrnJNgXs50N0+hLy09MNxkN3vETf2gSAsK9qK9jhHeAudy4kwabwCXAMzwvPvGPNYI7eokr1BvT
Ie3vmQaVwJQGQssM7KQj4OmP6lFkpnHdMLt0UHNgowMFm4FtHFnWqDPJino8ckJRFkmO6H63ZIl9
lm9+uDCFoa5Av7qRCsZpalW+f4Zc/T3/LUTRPtVp57AXrRAvAHMxNohZAcaolMS8P1uji1QY9YPD
V4ukCGzab4xAkOKJTk6DO4nwc85oBXoEek+jS/2Y9+Dc7+Rj5+DwPNAmhosU+FPLmccFW1xENlxG
MJd5JjUBUzQBAtrCDw5ZeGmScES4nrqLvKXsiyeYv/Fd99DnZDymitpRBRj/JF1f4Qlg32tHFWCj
0BW2nPXQcQimnySlYvKJWATnT+LBsQ2htEloUnTdYcQ1CUl6jXDXJv1lhxtkydogJtbOEMdHcl9I
daFZH5q4g9lnpHUKfdogefw5tONcWwZF/YA+Qb2GmNDsItKzzxJPob+fPINDc9Qpzn/ZW9Qo3WkA
fTPFddwSw58g15Zq35aaugImaL+6tZPYJcXtsWNPfIWZCNpwhWYaWKay5EprQqZ/5JRPzunPodir
sZK2UAqDFyM9NR5F8lX5lV4l8iWvNwcwdskmzJCpcSjzv5lTWdL0s97oPJlwhI2JLAnXOLd9vTEY
rdV0n0gtvbZod4voqKs0XC0EVQ3SM6i6+r3m/sIfwVirqkNLbn/emQHWhLfSs61dQ8mav+jJmf7N
3hdId97RlcXG833oc8BrERUsRSKFqPREy+esMxmunw0ByEhDozy6ksGO9br/ktm+AmtJ0TAfiprC
Iw2nIg5yLr4orPROV9jspRMBc9PUPhd4soy2Vf7KXIZ7OJCvxmzUkJqVwA5tl/8+KbvOK3sbyk2e
Imk6acLXyJboGy3IdSQ4VX0ahZiVgsQhTvx5J7WBR3eHy00Hu1WMRrbsntNWG0jEbd+jzD46lvTb
DQYWHOL18uEGLeTWMEKqw2vxaT0k52e0+0vx2kkr+qb2tFckEUEBaODU3C5jkOvkX2icGdsdS/19
9onrymH6o026VETLx7+tl7yMq4ozibhdRm64GwEaGrJDazceL7UzA7sc9DKJdLRcPCxfruDiqM5f
r9DPytMfn3PA/fvsZgj9rBbJOqQiV43pdwl31Be7lmGInb/siBZo1zbINoi23QDq27aZ6u2itJAV
5ZTp3idxvLI4TJ9inoFZLfjKwKggtR99jhq5Hg3vjLpibIE2xb76CNAw5bdWb8/ZNcDFYDB5N4Tk
pIEgnbNqyPdiI66bILSn+oGOuELqIbUn6DpKsawmGwEw1GznjSZ0rwGWGSNlRUrcW5VCozGyVTUE
jDL4nIaMwWym8H7jogcRDOUCpmDiLtYFUxRadxT1yclQeF24Y00EiGHfAHYl6CSiWa3Cohhh5mu7
BIUwvTsjSMvd5ZqA5itr59BCb8iyoZQC5l3XFVHkoMnbUaTl7uDZ8B5Vv08+Q8rDf+8pF7JroDkP
guqqPruS44H633lEXAzWn6pN+Yly13OY8M4Q0hJ4wgLCkhOxz0ibNs6XvadJT/xekHtqjlgb259F
seiZORsCezxLMMgLwHVHI8Gq+svu3uBMDF9FlTmdwz1L/JHnMmEcNPEjKwFM3Wx2KRs/ulkJxpiO
SgFn7CR+EbMCIXDA96ZhHx+BfIKw+ja8UFZ4E4LiKDBh2+n5YFuH3leQq+bGIgtpe46IgLQ/Wk0y
oXdyGzdDWXGzlaaQEJp9cxdkuZX9DanDCQw86Pf65KowH6ptuwtp1GiF8ApiFp4WtuUmg/ljdLoZ
3ws0iHvzsZe8gwmxY+dE2wgTTavNw0TJg5DZQx9Tz6mdjNlYKn+iJaYjVSAR27e/G7L+px87u7Q+
Tq1F8QYi6aWSbrT5+z6AJV0W3GFSxOfUDB7St3lRuW4El+KVSkbg2OTlAeMi/tLivp0VbkZ8wzrU
hCbVNEbxUhfxNCVcEwZs3sr0KxrCiHKld+/qDLJ2Xz2tgAuW7xh6GNAgt/fu0Kw7soQwHlwjWjPQ
ZPr/TC9mWKZqBTeDWicCY15GFdVIgQ+R5YUYMJgumNnqoSgLhRlPMP6FiGxugVlzbKcwxHdwz3ih
C7GviV68oVDKkSqdsUIGEERA9Np8iBvFAOLpMQ6ZlbWzOKGuFcY66+PMygDm60E//FuENFrbfNIF
iI3NYTec2uC0pHTb4+JukMdpSxJnXrune1I+LZy7Net8ZpT42oh7gUgfsc8CZjLMJWvmiDDRn7fr
ajK78SCEeMUrUc8o13xy05NA+jf10Z22UM2Rv+mgHcN+7OsjDuzr2biDvtYP9sTCaShDn2gPR8xY
/o8QcGynUNPs6ejsk8yO5g8+P7S8fFglc7DiYic471yzT2AMLtpAPrca8uVR2CDNrsUORfJ88smZ
hvTcN/FIgGqCHmyt5c1OYTG+g9RzXJarMFhVExMJayd/8zQmnwLsBS10DiW0gxioi8CnFWXMKAMO
Y8JVtVqAzfXPP0M+l0uTHlxxOtuA+aoq7aZWfYKQKy+DY9MJFA/Dmo2mLNhO07xYN9NP3olVctTB
wDl4NbtcXeZirlh6SAv18SmD40TKfBuE72oTvTO3o3oZfAKE+E8/OYkin2Wgzm3vVih1/4mMoRHT
7fZX0gtU8FppyPkrJ4nhKuZqwp9U47OYnTMsimuxvRy0ipzVAYVxI7WMx36RJzw1Vrdz/M8fNeQ7
qwsA+NVv2FJHQBJ4Clx1bUCBfzSX1zMj0ss2IZkj+zjsY0jUCs8JQivA/hasXPv5Fw1X+5i+6xOG
/qAZSy8JpIWeKhuFeozbFBdYz212ssn47SkB5HEKZ5yFqw+vTNZKYuUFIeYL2p3I12G2erJhekK+
xEV+s/pWgwTaDS7/X35Bndz4NROrPY2RpGBk0woswYpJZJkJ71egvQw4+Vw0fNona6/P++iSWuGK
KWlI/ZRONucPpxXEOP965l+DDa4P9Li0vt/zRpl5Vl/1Y1WoIc4i0ZLSKRaGVjfxBC9hAkspQLdA
93z4fZQUTW3r1zhyVX40ypUHWZezi6TeeB5y6qO3eu5tYnFmNMedvMX3/eJjqY+fuBKWQJABabqd
W8sQkStFdiqPD18y/6W5SBwlgBXY3/Nf8i5bj9zLpRTW+7rrPvZGcSBMy1rr9miRM1d4D+iO0gyV
eksc+Rf/4nBkJznqVHr9nWNwaQ7XVkSL9J9N3B4Vjvts4uL5I493TRTv8K14Jlt9rOpWcUPVseYA
PlYfdD8JCRgeUgA/TuJSR/WTu9zaHenwjcCv/ZrgzJsxGEZ5iPh4yvM5MD6r3PB0YSvPhtt9xnHG
bqHCauf5aF0ERum3pnq+a00yhehR5JYuxSS6wfzHSYFBF7hgcT98ypp+KBxOIGClnWeZF+1FOXzg
EKjEFCaFmPIFdipQcoQVOxpQrszL1LyOdI01TiwWUvkUdGsPrdRguXo0sVZVell2xp7uDpWFO4dn
BAg3jfylkOOmF+6QdKwUoryNbJooVBgmUJJ02CIa8Zf/ihxo4Olpyk9hm3Pvm6SRKf6jWBikli3G
MqaFDsLcISud3mU4ngUONaIM6JfYplYJBoYedDFbbgQE0qAs2NUxuXBXWFU/ib9DMfCJ/6+7qP4f
i7xBccbG/ZWaLPnVEXBKcYJtXvcB855OhQ0Glgx1SMEKHrq1jcEDGZHfXdIxpzZ10a2C4/pHucs2
1+pMP/jRYILnsPP0kiPdTMrwJjxCV9cOfHvUmhR78GeForUt6xjSsq4d1/q3//w6j1Lr5Lx0tGV9
wPuT3+IEYrSEAyr/11yQj6yTR+VBEjyf74Vt96yoQqjNCZHCptNYXXeV6TZ8oYk2H8156Lxzq/Lo
U/+HWhP+0Cp/sQyyZ7bCWWT3L/s0bxpCVlOVP5cTQuSnuPbm25UO83L6s7S4uUHZ7FDYLFNv0oE2
dLGFZdWrQxCpd6NH0fITQ1c581TBXyNP9iLZMxF8c16z2t8iySB5qaHukQA0D1PXDXSKoxMM36jf
9T1gYTUQB5p1z/lDs9IixPgT8EvZSpfpWW392uFLRe8KV6plkQgARCyr5Wd2Dppx1B4+mW50DAvJ
kLv6uTDnrbrcxxETvU/WfpdTi8WmOybYq222ayKbO3UzQ6d6LrSlHgS/1IBwHApJ+xIWD+DnzXTq
SrBZwHoMkQXu5YFBuBaRsXE+UTGOIJ6hJPbZHSQ86Btt/q/wrRtvAjcm3vOWAmTJcb7PLIyhucDd
320gX5L5XzHj9umfEy1W1kVd4oNwfqeD2LF/67wDZDLQie27F/a2nFhEDATHwRFNpbE92XpZBGii
AzfVNPkTk1X5WT4aa9xc+pgYVbgVPXFGKgu0mImGXU9VCSCvchJHTZxmSzi+gymmc0SfkXdQ1HNf
L3CSreZY+FV4ADf92RYiEgTU9F2rSq9KYJYpU/cK+Q00x9a676xVkN10Jste6I2ADyhzftPgK+gf
QdYCEKjpPPsz98BJFa/6FET1femJgLyZS5q5xBRGAJTTNk6I/i6v76wYXDVl3DRNnZgq/PWeSJOn
ZFTpkZF8/0vnTJN31zG1S40Mc8eZ+1CpIyE4MSkM7onoRMPxIwNgkfk/PwGmxvuDaX+Ru0rTSkU+
oLqyQyRcGimNqLC8Qc0/JGB1t6MztgJcM0CaE9/v83woQNgr/L0pXNzANOlLpL/EjHvz312/8/Yo
SPVJRr5tfsBOCJSOZnoSlhpQPGtdrZ/3rXPpTQWkIhok6m/nbTeNY9i6w7CkmmsplcXwPsqVLCSJ
KJapcK3nIJvJ+mg1iiir0lWumoMPAtK1sNQYeHAOtoK5DiHybIJbnhqggdBmKt9dqX8RYgweqNGt
sr2HRbwAEVh+jhPobZ9MsO65RHNR6p8HwnsMyEmBDm+BgTDvLvY4frjbecKLIdfzXHLF0XegqeoT
H+hAmIZjB4Ld2pdvfbHjaFkz+IKfRp+ohtxZQALW0yDQbigb9h3n1GJxEeUEvdTLGxa5lQDd8hAj
v6xbNBHBl/ncm9oI8y47AKR4lDtlKsB7/+BU95TO6kekStOOSU7xg8DK9iq7JffAFjr1VyOrF51L
ipC5LVzGRceBnvgOFQRJ8QOKkcf0/lhHad5KEFYBWn5qFYpSTVhjGDmbgB7OXGwHuCgNdwuvotoq
2KP64ib7tn0uniD5DuzqZJ5lHO3scLFONwa0pFr4O2KzoECMzS3olZ/oMiWFGAKpJ2Sr2kAahbKf
L5uUwJyinbdPZt2yhQOVGbpxRRCcjQxJu1s4iA9QBZy+tHwjs6z+OHwL3ZcmesarK0woB3STLGr3
LBdzm5hYsLeqEbxoJ0VQMAFhI7XNicHbplJVrGiKY0nyaE6hFSQ1zyqqqVd+8oDL3SGeXBUFwkcs
5KCUbb8zxLrW8zwOG5VOAR2wOJXh+k2trDCKsJIPMHbxutWNl1ZhwAZpvivBAvk2p2iIfbG1RMEL
BQMw2ve75qMHjQJe4bDTb/zoUG66KglrllPsLMmZBsdnwAxI+I3hUZaGHs9HFAzTnkcIytoX94VE
x5wOnqcqcOgSbQGu6Fek7hpRjueJrIZfUpm/4ljwR0ync10U+rrauZ+mkP+rJz+qnvUQJNclnNTg
l9OTNLvj0nxyGu0mcvcFsLxNAnsiYK3FLdL8caWBv7ITIFId1ohb1qJbDM5WIQBeIQ11Ll1B3FpL
Excd7AIPhL2f57Jb7/cRby8J15JWIb80SyHYPXaA++pwt1I18sxl4O92MsK7o9uZJzLCG88mp25Q
cRdTt1DchNoCCEc7WxP8Oolz2oTQMyUGca1mKwjz+5xoiYnmfXiwV11AYYYkBEA3/Vwc4k3BVcGZ
Y4nxTQYZ7vfquCoC/er1rh5txvieHyJz1YlC577j9ulDkSGwYUDdHeFgwuKfSIKGiakuNrSyiUT1
dK5o4gHUq9G1bYlR+W1BMV2LBA6bynMiar+ogmzQGF2C+zmlq2akWUDb1aFmdLhAOTe0PbCQ2sta
8v1nY3MVxcx5r9YEzdPXeM3NVX3Ni8jfAJlEjzAu3gsVjSnkV1SzxSahNOcIYounjHHW6udcdXko
heOlt0NjgHoScS4BvmI9q3GwjHdZfMnGX77LTJwgfhBvskCVKiFUES3+nIBEoZMvj2wh8SAJNcWr
/JbjUxUtgA6lJvEycm1y9mfeJXAomV0M5PFmXLP/+4sH+h8clvU34uq1kFkjwWFF/7lGd0hkofok
ujtvFy2My/lJXaknchEwWkHuPE5810bmxDhb5cwa1nfWy7yAAdQLlSccBBl62ichOh6bO0j+67tG
e89JJ0TGeMHhU7vvIz97xV6f7MU62CoPS04cEDe5SlQ9BB6hoOt9UF8s/n6ZTE8/5Vs+DyHr1h2F
1Xvt2iyv52ReBO/wPtaQcsdcNAeDvM7+p5Y7UkdT4RAfViudaD/Ou7Z2nDK3yJX/AW+buSFSBVv7
aFlkrcFZ/2pSm43f8pIq4Y7eJf5zXFhH5/AexflbekmPRS6LQSR0d4lKwnoIxbD2s9otmeQ75zFT
6lk6O07oL5m+DV7N1dgnNmtSzG3PiJhiOnTg3qiJgQR41+PJjfWQiqRCpeKXGHqqnirzejlVCmQa
wtqhqPc3Eu5YvEnulK9rc5RWGg8deDuJ6YPdxnSEkDlbmmH3D2w+8Np2uju/T7jlwQz8hB1dePKx
cbi1f7CB7uGSNnz2opuNVcZq6U/UdhatlGZ9NlHsJelOxNxrH2fop4K3a/uTnAPtfyXAP72wcgzZ
kR+xgPk9PhID2kav84z9zgiSOCAhqjqiyQ9HhAdDMwahMDAuiz3OSJgHFKQWgcDaPcCYBRXHfRLt
Qz3qXKJvDZYVvfzj7BSJ0xe5RYoZnQ+MDp7APYOSIRMJUMEWg4aT2dYM9qGeqbp73sMCjGlLtouE
IUF8nlcF/7qaXX8FyrMRrDcqBVQis58nPkTFSAuiNeZr23YVOyeXqkC9CtAcELIM5HdkTp5a/RsL
SErauu+uM6O85y2G5JDYOUsYvQ/ane4Al3gj4jozGIf386+zmJTXDMJLL56MD+Th59mrMqPHxt5g
4/+4A3euZATSavXJrAyYrsJLDPklxaF6hxuocqlrfNurSmddVnauXeCgZlu5BG3Za2kSEeazyo2h
c+kHSPM7pz3SRpBqlh2fGQbDHsMMmuFywnSslu28R2Wd7Vo3RB2+FeLooFYvyHZBm+YkXUjVtvBM
W8ZF3Varn3Zp1Rjr2vNeT1hrx2X7S7ZqX3msFW16askTSWUvyxTJZHm5KkTUiM1J2f4kGopsJ0XD
LtLs9dMZNaQb5Q4dFlHS3xZl5+ZQ04w/Eyc+UWsAf8vTg2gHGJzQqkMhj5cReu6TJ1b5xNc/p991
JiVyW/K4f46MXLeLIIc4p6LTgCpLFyugEeFqhdduFJaGEd7w8iEiQU4gQlZvDA0LBI91omV3S+Pd
7v1/AZB24Xg+LK/A+Vh8L89GOYuTMh+IoL1N4Byvx6+q5ceIILYqgIOaZ4uM5iqolPXuOGqqQzUH
QXrHONqXY4wrRD9mQC9Qp1J86UFrepDr5t5Dbmua5RwK0BzzolSeSI15PAoHTU0qLoxNvXsvBjjX
Lhg3l6/KA+NYOqxch98w4zg37lQ1RiWJZuzUpxaIpH5oaL1wR57+Jfp9YsHRtBD3CWct1qExZIyf
RtwyRmGcnD53P065UT/zBvT1XijNU9U+T6YFnW9dx2+u8AFgGfjEGtnJwF2SEL8BSf7kVI/fHCTN
1bKPttDRtBAQNo8/nTx0HGYlKArkOV+Mfx5jC/I7Pqk89RDqWzi4hHs2Cm8owUXQqUOEJ0rQYoOZ
tBrx624EeOrbMFAjop2H5G1IP/dg0tHTOOMRM5je9XNrNIiQ2EOaugWncP+Qu/xjTfZwVJAODt/4
FtTSxCGNJ1rfC1Ldnpy90LZKhHmqQw0BXoUwJigzn2VCHMRQHgM5Dt1PpFguh0JFp0CZX97XqMjv
RHBJwzzWrzWpKlV2SP1zE6smS8jR0meKkPmE3lAcPW1135NB4BBIUkuMpEpAeCnTQdc//0TM+wyP
oJymgVOCgoP1TbvaX0NSCrP4KwlB0RhPJYdEwWkR+cgEP2LIRBg7Q7tVRj9fUPFzVrWiEairiiFr
q01R5+YRFvtr0B0Q5HxYCUxi1uPNMeoBQJBl8u2EQgEemlYOwQ/Ji+iCArBPpeOLsVbgytwVH/59
NV0cTWIP6nDrre2VAec0OfZ1aqjqCohRPjZQi8IlpZgO8UsoqeQJAyDPZEO2v1Bk21WQBJt0qyjN
yEwhpqrNiS+ve6EokJ7j+Cz+IpE1mIY7uKj1uJV3KgQR1Z3cPNQLTv2x+rOxujm1DE+1DjUAceXM
Z9BsX1avMT23Uqwqrj2zXR2vZwSRSapFt44rblXPrxRlXA7fMfczPEaV15FQOpiXxJ+FE/2Rw8vb
j8gxdIBKfxzXYI2UwLhZtEbp7DCHSlaZ0s1qQTjuB4pnFcbTxzSQoyjA35KRw/IZFx1U/n0WbIiJ
BZEm/2SdV5OsN4kNJxtQRe6+C40SQbuLXo8OJwfiMyVR+pZALIoPsLv2/kNW+UUAIBCQ5HBsJeG0
AAPG4zyLtxUBTncaYe74EGKqEfnVxGo12Nb1e0/GsohN843+ONkYT0OEYNsWyUI2uI9ROtpH9q4u
+mpI5c98ULF7CsSreb26wfDE2FEV3kiJTwGxUCykt+EE2o1vUztLhC5V5QiFwiTFyxfZSwnT+h24
33RRkrDS2vX7fnn4aY67x/1lG+OSiuaPRMcnHKfCW0lmjanwE1UBApKCugPs2aYE1cLtOy6C+wwO
eebQerBiouK/9bHzwM6zgxQ9zbx7dC+GMk0+oBxVICY2m2d4b83mO4n2WqSRrSYR+3Vn8vL2t/ep
RoQgYobyOGaqWWDq3KWlFTyde+4w1YUiiJ2bCHPI9A34SkG7jeEOdPEktNJJ8GaFTV5ktnSuvUD5
eqF7MZVtE+QUyWsc3JCeuGS+UWxOxmulvCxRcr0Na3YAsJhlfSXAoECv9iSX+CxjNXioyOOW9qYj
6cz5iQKj9bJUk8wMCwvinNNpIzEKXqy0Gv+9qQAKldHbVKeUTfAVtJQGdWC+l+6b334gn0Ts6Bz+
l6W/+9VSgWyH4oFFzgIhhMQfjAHl2miq+LiogvhuKPNDlGB01FO3wEpnjGrGnmRrk9FOPRUbjH7k
EW4PuHM3Ht8R1I58b8UulXACsJrIeHrPJnb+Cv7G6kbC0vedeNNbzWx1TCLQJgmFMDm7/vrBLAVI
el8Nyg+xAPfnAmWYvY0dNP+Ysz37KQxnSt6nDfn+PUz739WMzMEsPmdmy2i7zkrxndaaqfhx8GDY
G+RkB0FwMsydfJhk4tLyeDeZeEOzOyl84USf38Noh5sR83DI51rSz2eQUGw6pMBo1dz1R4QS8K2C
ElfHoERWKeXEf+aMSBTn3OoIUUJigrzuZtWeRuqyECYa09wHW6emcyokSpFf8Hfqu86UfTVGgR6P
w0h6fLlE7Eyvsmk7uuPqnjtxzyyMHjLr7w37IBwBfA+0sDRpLlyYPZj1Mno4DsUdWkw0WW38utTu
fLnyt2kQr7IXMKdlE6NrYOaXDICS7SlVvh1eDLxlU7u9aJI2jdgZ4x2Bm6fnxARiSfog43a+RgmI
E4D4lG+LM9G+R4xkEN7OtpzisR/ys0IuuraTikxg+He92c34W5+at+C/qq/5ZONbqZRMpPTNBhrQ
VRP3Nu00HR5djbtDs9bCQmVxLdxcXMVNCBarGHB21FhdZPsSnmUVfNkBX1gFLpVArrOsRBZwcuZM
lGOANw1eH0Wu1GkS/jNjp2fAEPaNq0byKZjKd0IaTrerYpmEz2lPPZOucZDiOmvzPC3Q3jAtlmgX
yEzSHPEuUyVBDcGDChy8q2EYAhyB3dJmDR/c1Nclae64yt7c1U8EzRVsRrWHhAtQc59BIHwo6MAv
2qtWiq+RDEepWIkWVYb+9m1h6waTzzT+FaAAsqnH4+n9zMOK1BrheRQ92hd6vLOrwZcb3PYKRfO2
dZ4bB2AUn0iby8gQbZdlSxIEVl5/2rovNgbSwYhFwrrKu+D0ke9thXvN/hNuVFUHPtOrPJvaoqSb
8gIJKSdi2qPdUpDnRTCNf6qaYs8OYouLSbHe3kH2rM4rX9nbbfYS2uPvW2ZtrcgeF2m9kHhRP9to
sGG5/juj7ZBbBxCBVsvT9ei3Mus39dP2VZXFOqIJxBBvlcXYZQTCKgUmwAEuaZRO4cEx5cCh6M88
ex+81Q6aJNpEKR3Cqa75fmyJC3Wna/fvZVS3Uy6mlgUWTiw6NqtmmNs63DOMtJYa3Lc+ww6nP/dm
5fklv6P7hKd7llGz1oAuh882T7U1JPestrGxDQcKDN6c1gNAaFC1gLiwlJari2WQoLIL/WXEkhce
DV6snC1aH1mOJ+xqaIpIxxeRyhk1ltgbB8zdJLM4BdAeGoHgyFZ4Rmu56pQH3po6n5wawrEG1b/F
pnXNi/LRF7vCmihadmI5KJ0EjSPtAhdaLouae65YQ4EuhRLpzqnO4A41q/TX4jZVQsm/PFDHDQA+
iVuswQZK/uFTYw8hvlITpxOQUFJ1uIj82QuILSIIBBB1Y/lpaaLm3DXlzKcrdXeX8GsvVyoGLJAL
QMdv0ZPnw78zkI2YprQb45ekN/fsc9Xw/MZ7WU4p0WT3/nIIT3dbRZOHZ7SuAk5Y0wlfBHYLEP2y
jkXqU8TjZodSPiWFHyh59hsx066mTP5cRqiUXrNCVTxUdSccKdR/oh+WF4ZJnwsP0Xqq9q+5jXlf
1y+WwSFvAnKTw87uKyf+3jR7lc9+MaTcKPenvBtvFYH1U1YyOQUlnNQKRaJJFA9NiQDUBpzkZIKP
rfMjyTjJ9B2T9YT9X6QCvVveeNAShwk9AKrdYcsEU1aBrThxghksdH+nOkR7LAXUrX8W9sHc7+je
JkoMoqWLfIKGP4jCGFY3LwhPY3Cq/HeEA3lCYLl6WKsN49QVL1V5gZ9DphHe/Rre8Bwch+gOE3xS
bUvcW8XseEWOhsdcnwOG4qJjKF4WTBEeO4mITeKa18HSueXauuqd+XTO5YYifn1C00FobZ/EBdxW
aYj1LCUlF/vo+K/y8wodhsCKeiqGiRl4YuTvwRLsLP9B17Pb04QUwtbTnPwf95eD8qKJSkVsoYh4
xvpki1yjDSYE2Qh9ASdDziSgKC3nzuDHQ2g2NstxXVMVTOhz1YuoFOG/MRKsLLYz8PxMNPJVPgyQ
eW3k9IyVQtutAgyzMUXtW13j3Bj5Q194W9TeCAkyBrWKwtWAEA0yz0CM7Mj5/Mk3NeE5U1a+xxKf
+T60KDWaou2ahyQy66HRCa+TA0l41vypYy/s09tMLMwsx4msL8edmM1xGycJNZclkUeJ2S4iGwV8
Pr2ZGUp2syPE5Yd/admZZkSz2uosx5CxbIh+dh6fBAK1DgvQYYWKSA8CysprfkqDKn/acm+ffDLb
peJRXAOsBDw/TD5CCPvLTAFskCX5KSrZQGkwxPe3+iaIiqYu4APHyFYxLEsSQRqgZKDQTouj+LIT
Wh1DT8LyUNdO1rmOCoEX0WLlxzsCm8o19msRDlHW5v7rV4wRHFCueCwslEGNbCyPs6kBWS8a7FlJ
LOvfReZnWloJK8cn7G9zbQpNiY9tM+Om+JOJUHAKryXF8qVnUp2lG4RLX6v3/snjHhZ+jRCI+dgm
TIxW89E+glkXNO2Godiz49R1b6Y/MtIdqhmJS7jU6WEMQ2+Sc9sPj1c34bgnfIQpar2uhQqe3bxY
X0fed5pg5BTQqP0yMDoFGm0aLtY4GC9NEJtC0gp1RnxMTGJ+xDKkiaPGOCQUtWX4KRA52fWo0nuv
v0bVNxe1Du9XRdcBovo+Y1YSJdgnaVZYQ0sTj0L6vRhmj1rC/+nF/zYQ2b1KvR1NLhZOzTshNu9k
OgLm8qL2g/HA4yccWRfh/TB3ePycDQ/5X26UMh4zuywCT8ZiPQXTcBbyDy1YwU56SYwvYuMM7yRM
99bw+4kCiW3Kzdeni/RMxVQ/rLR8sP9xulwr8aUuIHKVRK4IZpgG8lvs8FDjQW+7qb2QgT34Lz8T
tbfk3V3WP1SQ2JjaPXmfDhaz7tiJyQ6S1v1xMSbLXAmlr9VtMaXdHPkvLFR/LlEDlx0SQeQyzFb2
1TmFn5h1/lQflBa6Y4ujqEWNwSqgvHi6qIY1TmkmhLnBRUGhckuxq5Jn+4vR0hlPDzlk36n9H98x
NIEd7zGcavHlHZqGg07wDkdV81DsfJZUCH7H1oAMDdZmVH7ROq+8DYudCUeN+yqrVZ+7c0OjxXYg
FFIT4Iz5cQwdNWI/PMfrkdYuokTzGC0I/I8SVJwIfupvYCEWVauKLShQoj83i7ADV7CV3Bbn1LxQ
Cg+qF3ERjlhXh9hWUHNoBjfXrPTFU2/cCu4DDJB1MNdvNT9PaFiXunOWp9e6DR2JE/LJ4Jctw9eG
xIjdmoHcBk1U5El4mkIAkeYMExgGUpFS92vKDFzTjDVw4acycR8VtZ5fazXnRVs+mYcXVD6zz777
cMpl8E22p5/r0uiVK2F01mRVavi8Awi5HwUhpL/tiTkjIlO4eSvcay/Ea56G5fnXRm2GeynEfTPr
98+uJVVrNEfxTCWxXh6Viyg0K8sjJiOLn3963eTBq0Hhc+/I2rr6mbLYvBozA/Cyf/kESTDQRikm
oWkDV2jRvow87vjYOt0of0VB/4uELfTts8kOPC/RyX6ZzPsA1uml3MgFgImD365iV+3SE3GDHZWG
CajltQBy/ufAKHIg70M4qddohP+PqdbhAXfv+J4clEkVpgbu7oKggPHlYx2lK3zGR6yYaIu8p3s2
j1dHrknBT5HW1BAXIRTUqBGXpOrcQvSUMfSmIPl3DdB7EWqjXkfWKpSGS4Z2sqHh4/BEO2lRJoBf
lYJirQJBDXy96UwPYlmVfa+sXTMzghJe2DE1ddUZhMkcjVgPJeS+PNUDUrAi6mzidS+V9f+sGMk9
5UwIrxHQGFrpE7BOJGSlbOjGBV7A58mLXnlHA5t8R8dThxdFte9fb1jEzV3qtN849oqsGJtXXoib
5BKMneQNz+fAM08KU3uopSjl5Api2IYyYr94ULZgf0hrgvJDAlUkr3gWP0OeU1evEuiOKsov5MKA
XqWV5CTjYeBmKBirHmiAb3ylOenw/8JpjPjEBDmiKcwaCCtihZ7+SU9Z9kHJe3FTxOw3KPGABvyh
JkXMl87e0t9cBQK2SH3WyfrCXXsWWw71Qi9HBmxagsY4gngkre6MpbN+v/PD8fK/T/tQUpdOMXVN
g6MXO7BwhJsfDKQM/QNXB7BZg+g0LfYjyDMnD+fU/RogbfGrXD7t9v8S4aExKrLrK+3l1/0xSpyZ
R6tSxxNyxvb7Vqv2/YrgaEDqUdTgG7c6bY/YyxMNZvydP1uitPwt1f90XGowbDh3cIIeiF4sR7kG
ofSylNpdsgVqtcGj70h+YraQY8MndMLwY6fHFyusj0mCNihKLJHtJIQcvhvv7+uy6SWkfbMm60Ev
hLBK8TiVS56KWeMk/ClmbvPKvH075lUHkMWamJRFbylV3+2PzSfzs3SHA4xclt+duYkdYzFNzyX6
0QLX5/HxNplyPVLrDwr+vL7Zf4BXwhrnrPadjvQpJVKshjq1Z6WyzgPlvhABkrNzgDDgsnFM8l85
rA7kkT9kZggqVuQnVuizcFa5vb3Lyl5zO16Q6sWscsLbO6KTN18WhIk3Y6X6jsbUCZi5OCyKSWJ1
wLs37sUQArxLXUWO7LBM+UzNq4MLkqkzTSbwdI7607jV2K9HOPKHh4vEr3eFaEeQELpZCt4zBrGa
ZnQPo/tWDELrVr0LUt0yLnLpOiTRtuOreIr3pBIDzELE/da/GwRmF2xGwpOisXtpfso47sRjgcGf
jU2QSEGFMIhphaVDJq8QbsJO64HmgrBLsQxHmnQo13HHhgB/+JBUErBUYyp+XmVAcVME9VoUrJ0c
o8xBkVxdQaMifxCFJRhMUlh6hB3pgvKBv6ERENTzKO3zI3MhXnAyWhQFIGW3Oq4wIo+0wMD3kNfK
WR7U5N3RENug6RVHJo9f8Xa4c47xIYboow7rd/wCd7vGKB24UMEn5itOp4N5Io/lm2X1wr6KCE7o
j5VFgkgeHvIysSjGEJh3IZw53XBVSlxVoig3L0wNCeeKaWZCnMDCLSgruaJXH7ltPpE6mElncwxM
45OFJcvYKi5wErVFiEHHdbwUbXtK/XPNkQlnhnj42FDvJQRUlthJo2EtVqvite9kw9r9XvBSiBVk
is01XH1f8zODBQScAghYU26ZX9Ky/jdXHrQ+FsTO6PG0aDO3sIFfPphnNcrUt0iZmGSFbKZFWVze
W4TytlI1kh2KBZzn7vtTAWVX0HWhLU3i6zNYhNFs6LvQKdIiUzqUH+QnOxi+NMbKjSurrga+uhwp
5YQhm4Nuyubrv01XpiArlRnO2ChFGb4DXcfk6pLw5BsmQMwujc3n2VRlslR5V5mwy9mvDD8t4G5w
oQfF1O6HW9WtpdDA4DyOhORg19pSbWdaU0Vz0771P3qq11o5b+uVoUrmNIlPkmJpvdTFnq1eyAob
pKtKOrbCFZfn9ZR7QjDa5PZ3MCGBNBgd1vpyP/rjsnE4qBxgybAFlyQVYFRL6sFmjGRk7IGUXI/z
wXX3RHRnQXE+TBZPtjiVM9DGf1+eZ4aMR4AJyjuBU7NXm+u135ilmjZw9wqb3sTz5/DbuH8TOCIq
GZWLvHFC7QBf/bkZkETDDA7WYquczmOv/iTod+IB3Gs1+w2JGEhYL2XQQwGcz2I9ERqC5TK0+Zng
jCuc2moqlwSsCFUrVpJv+XLrfSurQedWxjhBdMx0S02saiIiZIUGPL24ACx01HS1JpaKAsQUq5Bg
XoIj5U5e28BZmJuAzj6FsTHQVM2KgV1qWgWp/ECO8RGSTHTTcS6ZhoEkgUAPh0KWHnHBTqHSboHH
utuC6qYEOm3GlDg9IzmycKpK5p3vtPeUGPCS9xPg1p57LDltP9tTbu+WLpbDaumJQQSy8azEnHja
Y1fXXqEIn5jtR5wIomzq1N+8EhPfh/rCWhp+OV2NRdlZ6MlmkH9US5SFn6ARca2fhQUzUv/f6sMi
5xt5vl42PLSQtxoxFPKjrOtYgLHRdR9+XQfvDQXRiNY/I+rNpG6KJNKCRKyXoClEjuPl1Ug3H2lW
5RDjXEOLwAEMQbGc02jMRO7mbOYRHZ9gVrSVMPgIMtIQV0+Y910kzgesY9OWjgMjJXwEhID6s8kM
JV9WCQscOaeBE5HRnK9Hu07QHZmj0hn/n0b7pyHhBq9BAFqyh2CQkhvMOH9GMGAbWImgwFLfgdSl
apCbUaXWsV2sGfaZHSTqhhOEZEiMfSv19VBPbL1x5PnpEzMgEXuEHyUPD+WQCAqXBhhQHrvZNxM2
FSaFjkHVFVGgY00qs5mnFxiqFFSdjknptymyk4F7qLCsgcL3dEexcO47oWLU/31Q0kA/Reqse5HY
zlGq069Cvk7EZbztXZekS5r5kgfido4pgGiYVLe5gJ+yaCmy3Nwma7GKq8XfkkSJI0s/1OdxDOiR
thbPvteNH+Gp7l9Vf0+nXex8y+QvIEHwxYXfQl5cHqiWlJEqzm5k+blZd9wKOAKo5Iyj9Lv5mQ1q
FEj2UmcNC+TZHFG0JZXPf2CjW8Pqn9/sWZJwwhLr4xdiA21CQcbiDRxTXbEnE7WZPxMellSTuPcd
MwEDDsqhfxduJ2RLIPAzt/sF7k8k6gWlJ0ap9Vn7ec2UqlBuSLUh7Qhe/7Rz5IezyZ+UOcJ6KEFp
DuOS+lfUAtQej+EvOHhLhlM0bATMP7sjGgNW3DPPRxh1R0jNp+KwoqbwXPL1FPvByblyeo2Z5icd
xu98HdMj90NNaOTmI5RYAoygxhr+JLFGo+VZ7xQ2dqFOZWtCeeor3wnFL8yH6hjQWggVscBwQikb
KohKk7bYijO5hgO/Cog6Royk53Gs7TmN3pebj7yTBDB3GQ6NBGbQLa9jGVJkjhBjHtMNk1wiv3zH
8OOfPdQevFWMotWpAZVrkQxV6I4UsyDVUVyVbN0o+FrBVA+EslYB6BZyWUP9gnt8lEHZlh6ekUYq
T44EvNfayvQWFd+ox5S2F3AUQDB2HJU6Kah6vILBlftZJoZTYpNXfXiBG1+q6RpiDst7jnBg+WHE
yTiK+AqzZfUwZeVbEsz8WNZtkh41JJNaDH6tU5nzB9xPQN8Q3rNaROhxq+3vKNrG/yH3UmNMOBXj
zn/FsZl0zDAdr1rb2riBI0EzTiga9x0wuOrAN7gipWy/kJj0/4KEW5AQ6i5bBi9byuUhwoxs33Qo
HzvxqsNd++SAeAh3jfMfjaOanA/OnAxcuv35rHpUa/mDfwgToKoDheqSqu/1c1JBFRICLO+m381T
jLwga1CfeLOcRZd62MUvHevzYtBOBxJ25+Dg+kveetBiiIIyGs+hvYBvp0UKEW5jGoSoAYIWyLPv
Codys1Vt3dbslILHyeUueN8XTIaeIM3BV0qAeEdxN2xDJuXsFNjMwDzuC1S/m36esxj+1cPtgZhW
dToxmQf9V678ZMbW8Fgn+8oQT09xFgpDXqo46gjytXTIdPkFeBbplb00yZIPqr0LHSSWoDrvHXef
IK6gWaZPzA7qwUdvPiK/Jzi+OwLNafxQuR/nHDF/mF4xy+BachHvI9kzup8zMnuJVQWnlBtd5EfQ
T79suPlJGAsc/n5oZM+J8jmDUvGAZawdh1fs0wtCro534bHDJGoe2TieGJkY/CVR1DpLaPGF4Lio
m0cl/psddumpar+ZTEk4iyvTPM4ZLs0jbgk8OjFJMx7daVz2iM1bUc658WjP/lhrN8YYIuWP/kce
lS6A/gjzxIOubdyxnHyqw5T4LAkLQDDuF9j0yiiaHALBp/kU2deq0DKMKiLbWGAyx7O5ceM9VK7l
Az2R5aRiYzE9gPt75feqLDTUdtxclRJegKUopN3kb0Wm7+UCq7u77tw6psxbsvUTobH3Kx13hde3
5EC2L92KLmQHrW/5CZntdkTG59XQuD4ECMH6UazEruIazIPiEm9bAGOXp1SLQYc0cd+ytv987fDC
Jjyhy438SWKBXYGq1Hi+/TTGKh0DcrQBbNq7rGpO+rCPQje6WVDM64p+wD0LO5b9K763RR9BoJ3O
49LR2tAOJk7C7lsgZPn5Ip5ukkg4nSaMhvANh2rL3epfreJJLvCt8A+/qG/hM25Fg4b7Vkqmtu9g
lozNjStBQcin+mnDsI+xnIE8f9zzAEWp7nlEWPN0YEpYv5PbFdhyl2awasLYLgWeIZzRoM6FfbEv
u0CbW421TwbbUoLkRqntrPUUbwnrpQrZCPw2v85N0rGfmBbRW1YY7w2HchERHzlq8dputn9Xvs7G
nmuB8l4lgjesmqrjsEjpOhpdZTzAbQUU1eDv4vWhVdu4jHBjpI1FLSpNiG3lK/zdOrk9I7mF2KuZ
9t76Obrs+i/iJhchWMOtFAaQVw/M+wpU1NFYNGQoFCwi3GtPuQAAu0MUiqm/fHiP9dhLYuYgrIq9
hcX8F8FH15IeZFIGvSOCC9urAeXlNy4VNyA6NXUlzVsvb4TnSxpApyLACmtg28D4+XwlDW/ZqFNd
ua5EffcO1e3tBT3Yu34cNbiGaZ1+tUEffMLqTfX9rAj72pTRY2sG6COYUVM/L8xoakgCkIEAHoz7
+dZFFAnIf3LqYCahB+niMka2+vtOhk7c2RjBeeRwq9UOiwr/W4SkD+s/Oic/ieEfPEIMY4LHOpeR
RfSTaldJDhx8D5WVKO8zVP8Djlwly+gDGUbNHcEJ9KUSwsGVH22ndWwzmVp1O1Y3Q72utZcVh56w
ZPIR0DwLNVqbxxH98v5r7MWJByGU771xNeOJr3vOME8wwOADjuRBL4/M8aeyCJGYPSz4jHsqamxe
NrD1/IVNfZ0k6uoKegPSUDiBr2AR+WnixJlVMriTC6Gv99fxvJqZa60JPxg5JQxEAZYdViaZd5tA
MxIDrEyli7Zx6IAwGvc20Ow6sYx81nzCpsH72868IMauk4oKKHg/GYRlJOZjw1ckfga1y+45W6Ze
6Dkj4MGnGHJhFzJFamaz0oNtjYUs+dmeQulYLv8JnZ4TkKQ02VUxL9/10VhXmAN3o4wcp8Ca56/Q
03xNS2Tuw3WSNKUSBfhDxu7vF845GvbnieLrHatrj4UueqL5232AwHyGMvQoepXN4Gesrep6NRx9
zVrmCoxUmilfbfvYqSO2+lpl4nXFgclfoDRhvl2xmcwd5OTkJVoyvznekWbHTEcPyph5kWVARuZn
+qhF9q8Mb5/bfKNgyy15e8AjogmGmFGGPgJXWerom0ivC/jfOXtoSAZ6nORgK6J0dE42MgKK4K3I
sPDeaKa167ZNmO49f+J2D8/aLSPkcmV/ZbcdJFT3zn6Z6nXhGbPH6P4Qy5jBR6P7z/b4l/SNwoQ/
UjkWe0QJoTmTTXZ6LcY1CPgXVMoRoMQiieKCnHHFwB/s2fldprNV1oxEUnu9rD35C7gJOchFbTul
WrSyoCGoZvRz+LpQsWrpJXlbdFp4sYdvUP50XMLqhtDGYyPrQmEmNW7ZD4W6tQ5omPautROpuet1
Y6gatgDEw48/ipeDQc+f3a8W9ehP9g64lf44EqkPFaJ+DLKP96gtyDHFhZh86xaX3RgKcjQshZrg
Tu6ZUvnsdm1vv0wWRvDLhzgqp2nNKPLQqAFAlaJQxrE7bXw1v7bHHJZqYDE4FfZxewjPiP3ub38d
yxPcHNVRbMbdpH0qP4oNBeLRJ2fktArth8LROlQ70lEnRG2JoVxqc0Z71HHebBQioptRhS5moIdl
vp36ti6CeKeI8c9f223UsZUbhjL85ZjNsW+b7P2D/AQqw6Wg7iH+Tsqc8YngDDnglOZgcXKRm9Es
q1hLpAHBtlkk/u0C2u2w1j5wZVA6bmvFT8d76LpvQ1Md/07+VbokQsH94gxsOYE65pPzGFHJBKx7
p665XqJ/GpHJu9hG8WRn6ewUpEu+NbPWISUO8ld7diHEWhfDHkN2dWiY/dXxuhWmO2Yh7JgCC4vp
2e9qJuGqb8xAO9NB4/AQqcX5AgOBodTbzk7hvlT/NpINjYUIUgQoNoo7tZjGXcQ0bXP5K6wFEekg
mcds8eM+A0a5zvPAzYJdPz7EWsMiyOh8iES8jb3fwrBeT5X3xlBS1aYsVwOyQ9uKQYo9CwZx2QED
paMUPiOllXkekpNENuMJWgSasKze8Y3jlXidBitnlHoJiG9wQJ9TneT83cKaQG2I6CaZHMlqVv5t
uYtIYdPT6FmjDB+pwFb30EcLxFP30TCxV2T8/H0Om7PuEM3wlRkiTw+qK/9g5nzQ1RoS1fj5CKjQ
P4RRSTLI0GxQvxKaVJ72CeiiE201HiaIVXtfwphHJian8igSDs8yjal1oTsEBgv1WtzvE3/tqDoT
S9OHTq4szXAIC1MVi8/S76p83Wtwtbf0InIWBVGIXr5b+r9x2LVhogZsVpxm+yTYxuXrC4VDprrQ
ok6XCbE20wXi0rUvH4IEKmf6rPU2eDVj2Jt8Lm8Ngrzuejbkp+EdMJddF088iusa5qzR5fO2Avmt
NaZ8LDebMLGLCcwcNidxR98r7tGL1QcNmlrDo16JtZLzBig9lqpfOgOBSaegXHUPuEJMN/cGYH+N
sBqYoIZVO2B2lTagfjPPvCaWhH0uRRpBsa5wBX9xrFuwWuao+R0QSXz9pz553RuzogeR6E/eyCNf
7TMjC/VJ0HHqzwHaEo9obw0Gz8y3eeHtjNPCHTPxjuSpIsUWCD06GUEjvrn6k3iV5qsqm+c+pKdK
cP+bEfUWjFSkb4WXAAxijs/XpQ8zKK6Wm1u3mniDLnyOo6nnanm1ufs+1WjhkrB7ziRgdD8L7tnQ
LDjQYszdRtuIrvgMDkmNhQzEN/oo8BTUVIxtLuTUvgBy9CBzfIOPkn+GgoJuOVrT8qOJMZkyVF+x
grORlPOHHXrbt9Lhj/MSDmOG09Dv/u6l7fa5XRd/jQLtFOStARJTvlHEcs9PpTh8maGpEJMIrYES
vUNRELmJzvI7cJeMurSdbT9B0dFaoPXh9XEINgZPQ8Us4mBp86xq3uENNE4Jky5LKrei7MATzd7b
GDoZuXNoOTzZC3yithKQMea2bDz9TsPOhGQk9zDOu/rlJGp2ftNnzX8w7+dBr7l8utQnviL7qcsh
4DtLTTa8jM8dPlPFaJ8dwfv9fXujTAxt9dGT1hrfnoUUcGEbdp2tawWClWtlsVqTLlZqwgTD48iC
kunXHUlaP95/nl33DQxHiHOJZ830gNFvjS2u7SB7pjdfxddgVRsfRRGl+e+j+RzpktTkKvHp1HuB
/fZvRXfSWsw5wiLwo3y+V6acGd7Y8SHw5IvIjIe724AG5JgRfW9pxbzvDpXvXAV4FFdAwjPpVo2M
dIpVxemjjW6JrSSrLvbaH2bJeBzXnPJjF622pFd6vtvTWWP7O1KSW0X/IZjXO6BdlWQ35FnVaqSG
55iSHxW2SrA99GZf9JCfy9QwtdIof5dklnqPuQYJJMgyGNjVNP2ubbCXBayi3wfOv9mZgliTYJcH
Rjy6NrqRpeFSCtRAOTZelCeSuJdajTFpYZHvnSS5hRqXMYcYQv8sMKusmq4sivSpwIT+ioedibCr
fw44qrFgzgzCoLyG7yc+7Rxse6ziCKXmEDCUqqo1BoUd1WINB0oseifT6dcLQD3LZ//3FsGkBDJD
9uv1yaITYp/A2e75xbrIDyI0Df4smEXoHrnFQNTCWjXWMM7B85j3VC+IH1eiPDlcIUf6imubWTGg
i4OZ7E5NVkNCc5hjwOFYHn+FQ3sDLYHemfb8C6VinmSyRdLmFOgaPxz3NhVXGMlwk+5FCE/oPYr1
h1nhmO8LU32swRbMKHfTh63pPyoJH17xYe31JDe32o+egfQ7pPfyJCwSKLddNpyXYeTz63QRVw0Y
4s47eY9y4LP8Ibhh2XoaPqlyY3E6sO4BRID8inu6ukBeZmk4TwUqs0Ya+Y9n1i/CT7f/fJvvxOIN
G/L/Rp/EWvsM5JwGfb3BHSGK6AQ7s1Xcg4I/fWnuM+uPrZK16o1M84jUaKfxf08wBCw4kDRx1vsV
swS8Je3pmMv3KvsXndcnKpwXep8EAHMsdXhKyhnJQjRkGsqSO8ltCzyY/8opRFHVqmKGGKaoQSYG
YbahXW/s6pMz8MDZgjwRsktS28t4/4i7Ay7UOaN2RlonP/mUCjEgL83Fb2ip3UUnNuL3j5x80zWb
mcTPOfMCdgQf+MQRxXDCi5+wfW278H/aBUj+q1aNXb6npISABjTqMQ7xsZu2Llt1GIxclih/nPbJ
yZeEJ54fguXsPVNbhJw5FqUdbyXf7gklwf3ekpFoQ2gLDKrDupx95q+NGRd82FEbSniHtJWAVI75
tB5tLCeMjTm9j4phGZXrJWF1zGkATK8DscQjiB8sS7lrLYIqwYdieoW2lai+amKrCuubJ9KRq30N
nHP2Oi3PBZQohkL+1fWPpb8xy9AdhzsL94l3dTjGACExajMG3hOcyEdlWajNtySEedn/cDBCYLh8
/tPJOFeN51xBt46D4ar5RnOibfBo8SQledUTnQW8MtsO0aErBUZ6sNED/bH4vTuidh0/nGNPfz77
0E+ZGfotAsVSdYfDyDRjXw4fKrI1tyFoLY60/owUJ8q8EvtEjgp5zvo6AJSYgKUUwW4XdX+lSaNX
1LRuwT6emNDETQafSvHX9Eo+OYSUVWRREuJ49A3lw7G9vA7cwGbVJjsZmMVv1j5qpGR3Vp35wPWY
wi2iHcYWK3RTGSRmuIBEcwUpvwAoH1PlyULtB0u7hyjAlDLEGJtx3sP/MeHC0zEDE7X6DHu/vLUW
OCPDTI7xN18KkSPcz+XkM/iis066/snh7fgj3kFaUx2CWvuTM1F+z4lAaFVGR/+tdd2ZFhvfuV4l
up6Nk73mOMbMvZm6RAz2uBZe31ovpE54/rOyVnlRWHW12THVxXEoOkfNXjkYdAg15idGgB7aopva
advSqfSe9U3U+6EZ25SeIiQNWDe1l0dfGLL5V1DIDS5wBzg1RG6rAeSLbVN52iUem5fIQVT/MeCf
ljSd/55LWRXmmNWu4a6i/FoosPK+Kx3hQFTkAb1L/C5+8FR1GXcTmb7xS5pnkQm2VrVtKSdT3UI+
aTy+1NriqAA2d4uF5mlTAY67vbJgs+9gWuOL/FOeA8jl7PmPfTi2EfP97cKfFnNEfb+/i5qQoFXC
NWq3H3m9z90LY4kCQ10Yt0XoFMTx1+0jD41155XT3hEpCvycubsjJ8NrblpaVe2NmVYsMNenZNLs
JkrRNXmYMf0XAolNu6vGCZr/VGpJzPePZz2C9l7RUDJAR0mfADmwtlYK5uz+QRZEVVupjELh0hSn
zrq5pkeCGTJEXIjFnJYvSg9uu5FWhuSCrbduv9OSKqcOHHkuI7SsSM1QGjIdez8Czcon4p7KntmX
ec3ztqUgtCGpm8FUrSLWQGB4QM5UoyDal6s63FQXpJ+nHfSRhEOm8vVWNUGfMIB66AkrxLnbSIjp
HkJH3oiAHOVJRfShRHqCFu+crr+3CFKdK/ZOCphzn8xaYY/vDsL3ziuO+aV5LKcPCUbi3BioCf3M
cFSChPbxYuZz3y3L1jTcUXsCQNHo06xcAnL0b0jMJnZqOYCJc69JIL/5RjKWLB2lcQYmt9CFKhq0
uD/Ip2cwehXORTKFV7LNuENKXHgEQIp/wfLefmDyG1T3VxKhv9a8NmV7NZJltV41YSv/swoNc93T
jrz8eza+ar7vOLyIccV0fVHsu4NKtjf71iYkWSAn18iu3q11YTWqg8O78g/Klpe5G2RH5OCyFt5n
9Mqxmhvqskp1AlAYRgRHX/zJbV06P+gezegX7ewN9v8Ld5PAO/RVTexI0fVOtQ7e8Wyr0omUNUL7
zisZnSxixUXWHQMrTLxOa7PM6sw+/IVDOiLHm9Gw+xsc4sAn5NwRzvDKr670ZDtREZ+ArTSXdZmt
RXAG8wpuYp+2hPfEu3ZW9AOIxtGTgT092eTX4fvAAvpIIwryvdr0Mw/ijhHQdyYo36bLTWuRGNV9
Hui/N4GBVvr/5IJkT2Hd1taC1NHv9c6VhpL6qa1U4/merUQpMlq1af09oWn3is/U/w5/eDyH0CeB
bQIwkpp7wjKrtEJo8eV8ZLTGyQrwWZL6XSHkfn27gP//8DQQhK5ab0x6i4kDPO587m+wYg5EVA+g
gVErnm9rcEPN3fHVM3an3nONo7QOGMIx1R7ukfaQbEaRiKXbiaNqQXXGxWlZCvHzhskzcluv97Go
mbXuDKohvs/IjLLgF/qy5f4amr0+/JJeHI5fusLy6K3qPDc8DqiaNCY1cgaMuVj/jrqdgkbd4Hi2
uhAzsBehPWEi6CG+D+e/8Sop4PV2EKSQW6toNIKkSF5GQP3kDwOQEaQE9Ar1FCFvbJ5PF/+Vm1sR
qvP4yYZWLli1HTvX8CNO7SvYtgEv/747DSXg2zpsRW3dph7Ly+KbqStRo37sOtdoK148oDyr2QH3
xaw3aDIKDkCm4hf0gcSSsQquNeS1tWj1k59gt+2u209X8GsJpJUR4bZb0L2rxw68XkJNti/SDAwY
IwlhvbTsBCrR4NI9PUANhQ//J0sGLwPuQW4zBR4VwiKLfaovdEPfmMZOYdfsPLWOt1VEsnmJtDeW
Okf+uvHx952ZHLejqbvDQk+xjmpD+dz98v/E3tCB+vR67DbY4aap3JoBRamW0Yf2+YjGi25Ul/cp
j8+00SJAR1Qntssqp/BnvWXDRuher5rAN7P4SrVukpdjcIlhtZUg4xkHcymqTmBBEvXPEVgPQjYU
TRh+TWkqbuZeiw6wNplgyYe19znXVK+YITZWplmWaFnRyXZQrc5Y2nxUEzyWPzgn5jTGoSqvVx2W
6jG19ALURCz/b4TMHE8ne4hirGp1XwzbWxgfqmbVW5Cs9KpREUA/b6okkoWM1pXlb2MsW8e4gSGJ
gAUOAIZmdASTHpc5zTb+HWHDioogp29nYTFTtl7JBp10+GCP7MkJ99aah3U5HBqSK2h0O6L6YjjC
cVD78hwKQr0b44OxfVnZEtaQxRrR/qyfctQ7tF2sl793zClk+v27R6a0TeB4RH1ms7ik41eCSSv1
hgLhGW46t7PamK4CCrrr1rl26qTj2LLjChprPCA0rMQS2QAoZ7tJ9STjFyabgeUU23NYl0MTTj+I
B/XSvDuXdBJJB2+4toFpEjqWTUzuM47ITWT0xNAIXKgFRlyC3m7AkQXIPy05B1JsuU2iyx/dDTL7
kjCrLnWxWAKmAeKo27FEeJCI/foER/FogQzd4iSS6sgAPv29Yj75r3xuN5VhcG4IA55b3DbJP1my
4ZGe8X3Jptb0tu+Ifab+veqKsGctoJvNsw5CFUtdmC225vjMBJ3i9AC8gchb4M377THbFfkRUwNG
qCuE1yr5Oeo0OgfovtnAYi2wiitDEHk0mAFSEEsoH+od4rEqREBjQkKCcQvDJ1vmucjDyDi0A2Si
V8vB/+pSIObtN0Ju1gIdezTfBvKZ7RUdTl+SBvwjxtFuoIjZehS639jw20jFYdLqSQr1MaOS//oB
DvcZqgpLCxcrUrPiPzFfGYr6jPH7rHzJJS/d6U0RAD5GviptVlkB3BK9X8iroxnMlcRSF04QWcLd
Q2iICIK94grY5/cjcdWLXxzdqnvD0km6+aDIq9glFiKcz2e8dw/rgikgZKmrzIeuX2OA+76ubRg6
2O3wY64tPOYzPqoyR0E1vCOSh4pnN7H1xZ8UpbXy2VwkuL5jJf3AxpRQncemji3qmp3pMEaWbfRj
gOO1AXz+xtMkxRoIMzshXyQVlKTUCSUXhlg94oWN0d0DY2q2lTKigBQv3ShjVd82TKVMPMNAupFU
M3ColkLpu/C3Aasr0oXhW0Vdr8LCT2Eq1rpDag6iv+37KGul04MO/HHxk0ht9oW4O1egGPjF4NdZ
RwW9EHUc/D4cR77iux08Lre3WgWP/SEroimlJkOyBD3hsXiPr5SCLkR7uoQFEuzGSf14eb6tfAq/
PptIwcxDAhKtQ1sqBFUJIXeInFHvYQb4gQWjaLdRjSPz/uYd7J9pxWD2KJMO7gkzQGHZEG/tI4c6
x6Nk5IIpRrqSaqES5lvNz747TGnP9YOxvcX8bmXt5kqMB8TSF+gq9V2fvKQWgK8gOF0RVj7cVsOZ
drx8Ac2+dvHGy1GMv9UCUvOUv5IoPngvLaYoepyYRNFMbA3jpa1Og7fzwYfkTWudhhjoSmRCV7A4
4PGfSCOjuIPCaIvlOuBOUzlsxtE9p1ImXjCcDJGn+9uMkpmD56alVcMgAMYH/1UY5mjZz0QsgyG/
y89Yho91bUK1OUEr4QjhqAa8p6JGAtVw9Xr9IdOJuKIj0QNfOqojJy3nWUSyv2DE/juVar30arGQ
kxyFBej0qL1jBpkss0lEmh1s0gojb0WfhzRxRCozrBSpsX7u64IvvSxJ7UEIXhWTYmG8hZkhpvO1
C0UvMmjc6WJzxbuTp7BzYHfDaKnQOR0JSnBk3wtkxe+0yvAMFvy17eamMzQldUsBoT5xvCpZKwgw
C2KtTgPQt39lsd+ym2QY4lrb7QOqs4li4tAiNb571mPuLhSGEPHgy9q2bwoF2WMeZ3nuH0ZdycqK
ErVYRWi2C8IdyDyBJ7KsTatW2HjdUL9u3y9/fghJkX4N/L82p8rnMesmBE3uC034P48+9sT1wtpf
C+TVuVFQ5ll7vM6UK+FDHWG2FsdkYePLUmvmhy2Ml2jgy/gNvHIQz7VykIawYE1FyYEG8A62GPPJ
OdNsraptqYYZJBd4JynvCY8cHJx943SfYAlA7cvy4WoWOTgWqP2bqH25V8qR33tmfexLNreKaYFh
5pELvPQPD9WsErXqyRMJfLcvUnZ7YN588XnxtE6AqkeGXyE0wqAOovAepgnHaX3KSZyovvg4Zs0x
22+tCwUCXonSfltap5XNW1+wrJkvzxUnce2dg531RfYwN8+iaKiQL61N992vPjnxroHB39/VH171
iwzm6LehB/zcNewJTFV8V2flB/RsUEuX+OoOfTYwYbBwG3FIduHJV3YM0GQfjSierrk8lO4wvxSL
IsCy0mDDDYsv4bM8AON5fyOLikgrXUvShKiTeRhXjd6KzYUQZAxt0EB8/xfT0+/y9Jf7pvuuAywD
W0bPmescQlXuZnRdBFDgIGUfbk7JDQ3g7aUi1Wu6043iCITdpQbTxJt7FpMXfxthHopr/naLQoQo
JnOiJ0R4o6dS1KlizOXzv/dPIJIoA9fATJYCo/cIhc1tyDy0dPpPxKGhuEbKhZeUsBU//8bydjqo
q/ok9rKpAeMa+8BrtRvYP+QrYt+GYvspmA3dg0p5IVBrNDSFl6gu5QHaX0lisviZvE9yPb1RPkPf
LjeI3Uoq88u6g2IvgaF4JlK+LfCj0ddxqWuFxJ1yWRHnoZdAPImm/mUtUiKoCqAbvwc2l66dSbHe
FQ+2TNOTysWMvXFpgdh0AX4JDynR1OoBqnNt8TwPj8Vws961p2jgXX+NmScWthv2OtB06TbTNXzn
dpBeX/OGo9TzyGNDCy8ipFUv6l/6Hq/IBzK+nMHB634+tSslmnYW/h12nZV0OAIf7fnVQAV8TxVf
iSblrrD8wLEHmkpB4H0sAQGB1OJLaHJhQr8rfO44ipA61ty4AgFP8NZXxA8oC3xNxzyjGICYDakU
OzRBpJMAlDaYt6ng4QeBt4hFls7+MlpBN6qhoqEkP7YLGOW8t+TtQgmhjLyB4W4bwN4ap1Nl6ZTL
Snc3R7ooznTzM2cccwJJBfLDrXZd1XdyzUi18HITI5IXMZq0E37pWMme2zbAuOQV2V1eApg3EqDV
VTZ+zRny0m0NqcMbFVRawjI/qHzkK5VUYFuV2ck7FnYPosD3Y+A6bkpnzypYQLzFOaQMjTp5Vvaa
kz5MLyo6UqosiFLvc5AiHgj6dllEfcde12iyahGHsfsFTz2hBosO+pGxsPG5l/oj+ieXdCkb6AmY
2dNdq46xm4mpHX6gwssB965HU171nBv3/T1VbmBeqpqnf3jSGHBr+rdIZvYHZsBVCkpHh+xtvK7d
E5rR7KmC3gk+IhNYOercCAYSVIDQv2ACWFYtJm/hPQMm999SQhqXn2D0QcGAo/YytYL8nuJUHMqT
RvJHm9zfePLSd2eRc9a/M4z/1gzjI5L5c7DQ9pytE02GtBDzX9XVpS0IQ7i9AqqoNKUkBIraU4Xv
rVUuwSHWHoN7d/W6unfbdl7V9HlpYMXwT2KfC2CEg9qGQ3Awr9RSpvi0tI1AREM7/aTAVvzg1vT9
q66VKfHWXCkHgjGF+woaSJFPrCdGeGEopgaV1IeAUzNnk4CmKrVOH/+AhQVMIh2N5qjJ4NdhNewr
2SDBgvMgb9PuRgHDPSMTqSIYIJAILYLfPNyf2d6Plkd/SV6QDSPCYI/MlaAc06z2K3gsMb4ao2t0
egGZ/D1UlN2Mg8iW8m0YoU0W9sgqHTSxpb1kPV0wxClXmhD5/luGGh2ucDD+hLbt9jK2TfDyTsqP
KR2kgl60dsFc6eGbVRUTl1QlDxTC1pAgJK0bJFU7jalWrSi0YUkkK9iOl6WUBAzgEXelgoeClFVJ
t7cuv4U8IdxcJ3nkhjIUpByEHyWH4upc9vptDxQpFNjqIg22pZ3v7C4RsTrZFw2GFUjDWh6IgmCc
g63hbmMuhaQGyR0sKcXe16Kn2R5nPohfUEkKhK0iXH40kDr4ZBFT9ju6Z8LYLJ1Q/fIILpDsc5/P
4VKHqdIpbUThBCOv3FG1vPCDYWzKq5gBeG9qq1Gjvxw8J1SqtUO6jGSJrLMIiE5FvjdIuohT2s4U
7ylZqqlnb84550Rb6YJU4D3jcCXeI97ChGlPRPhJ1JtKLga5b9aDwChfuLkEvCzqXg3n584WbURf
rJX9qu/MViTjo5H2+b/MUXsqUb5gbiwoNuT533SoJxeH7waojfFQBtoDX8LBeVDW9os8o/WwsnWg
9lZ3At7Umzaef3QsjgxfGkxDpw3WiaoeCoE35leQhZ/dn+TiBV+n2Nv5CrvE0rf21kcO/f0d2UCd
7qazNMZdO4VFf9B6xK7wVF/S3DxpUSGBGLrvwawOKAuYkC6GP7n8NK1PI5apr9lcZIul4TdMZgPq
16nuEkfYIaoybxvLN5UTIubzm3TIuCkqCw0qEHQaA09rlEa1miZFwgAiLA0LVstZcK9O31mSgjzG
u2B1WcFxvHbQ+zGy88mBg0OaFomoPmUUGanJNvVrTZXC0mAx3tQSZbQvfXLsFWeEFUVXP67rcxOD
AE3fNVj/Bhks6wTQ1f71f/bjTsxzDvO9YmQpA3zSPpi6/DSzTfEp3vr7fSNd9+tmsGbDSko2smMy
wP79n7mt9kzlmZV7EqUiGTivrJJGG2J72G3bkpLQMoKOhGO2cgn2DVOJQHb8scpcdyckJRl2ZJrO
3Z2FNYWRfi+xxSpaoGs97ckI0b+yWwQNPDQwkCuCfId3cPi5xaWS3+ZWNwNnenseUDVZkL2Uuwe7
IbWXzPcEFiEzVMxMwBHpUtYkDlN3b+1yyw1sWqSbC+O0rvgIEOIPzuOru10tnuJE5mbq0SPO/bmK
BHHCFf/KcUaXbj/xWeD97XBcwrPBvzRvyLrmYCXJoKCY4x6ihbOG6UOuKcbNjaNvu56AKKOYw/WC
l3dAVquuPijfS2mK1LlmG6uKm86vncClydd14N6ww7GePqADnrmjF0Ow2AzzUgzcpQ7eMs4pACDM
sxeQxdrVEWoiCVRiLZBSW/1BLkBs/gxLrRYglt+jrus+urwx247Wd61F6JQkHIyXYbGur8HSXYZG
UExE4YDPgsPe4gRYGxHShvdMorWCWGtuxFFucQYTM4nHxIrXvVPO2uGUdnqt8j5BlgP0/EUwyn7v
62VYGXBwcfuIGcOBYz5B5EYY2I2bqc4vHuZIqcLm+/GkOqMxB7dpN3CgB9rBjECLD/66G8dM9O4I
mf9PecI5g8FmFYF37c1xo5OkyQ1YvImd23gT3DSYNisGz/j6pjDvztrCAXJ3+k7fjV2JdIzopt2z
Q8j40C81dQ16N21V+/Fm5SDAAEoYc1CA9WOxzzcTI4ggUvspJujzsZzQ5ScjKXrnhB39ITFVV2YQ
n9P5o7ENUu4rzEnWSLbaBxwLR12D02MswJYwR8ha7M/KjOOVH2VfKk5P1hjUJ4mtUDPyUcFlpTUZ
OzDg0Y0A8CV9JME9s/cR3cyb0johi3TKPumSaqFlZa/BzzklseFX3aLgUDtQ0G7F2e3jCwilT/I/
p/lDCrystsFrSB+WAhB9XF+WvqIQ+eq3WpM/k41tK4q2hn0NHKMBSKOR0kpce9P9i6Auc/rhPpc2
//6XUvtu2ren4ky6f9eQpwCaHtg9xvPaj7HNfwcuT2DWgc0NjppUNuX25NHrRqzSuLx3bhKDAbsH
9Q8JmdzY8ZaZ0WUNknuT7DPmKIliGjtZMxxvqPqo65y93MyE+AoBAAa0tsvsl6pg7TbO7mfRITnE
eAM4leEH8kaj3lBO2991MzJNz126xDZTolE2CBX2KLcv0d4vYHhPdfh/Gek810nb521Uq5uHbmWP
S84I4zNxEdySGA1auQwJhX16+ZdaltG5h6Hk3jTlpVJiPM52ZhTd5AXGPgvzR50g8Hqr2rS6lpNU
oP7oH+z9b63vIgCiLbvacsePR3G/q22w38B88A6TyeBuQuU+C6fT44GeHELxFFqE/3njI4WirHzk
/J0Q3u++A9yhCTqsX5S3P1Sv6bgsABjISrMew//mkV4QWTSEromQVd5ZyAteNI8VbzUfWPVjh46K
W59y4N6TyRZIj6TJSlUdU6E7w3g/XdSDY6M/4tPByv0J2/1dYLotlDM3P7oO+3xoeq0HvH0YB/wD
zIuoiR5rsc5rk+gNOpGh5VNkvCoosdOBPXHHnKJFvZiKxPfVPYnx/u0ZJR20QD08EYYPaC3f/jVf
VuxAcbBrUYV1VNn2nRUPnF0iTHr4GqPb2p38Misvkk438q9Q/9VAqI1LVzCKlVBIKWEDRQ/iUfox
WdrQer5aK8q+M8TAV4eegW9Ck+WbTFfMJsrDrvizxIrUuOmxx3HiSGDW9VVkWHSLLWLyRTje1Quf
yDbD254CAi0mk+tGI3JTh7qiJTNO089uU/QEJ5HyRVZ8zch+sUzGeO26AfSPkLaw7iCWeJPO56PJ
ZVzgToxHUUHWd8BHps01JgW8hlwrIc/ytl00/vlhvsA2s/b7NNnfhAZ0DXmkgREELKhZ9xEJiaSz
ZNrtr3vax25WGNarEaqzL4TDLiKh+3lYbzoFpdHEBqszbibnrLuZfBAWgKPklUqUX9vKaYA58zPz
EgGYGhZyb2X3vhbk9m5JrrsbdRN9m9oGKeZvn7pBbbFkYkQe/tUzVEuXpNcYWlrC9n6HpzHNMa8b
WBH/1Q//f2IUKXh0D/IDh1GUJiemO7ZwGAttJHuCethQED6yI4/+mGVmqIzAAvufRIuCzuZ0aVvZ
UMslKWN9Yu4OG08++87r0MZa1mIXLvzU5FP+GY6JvBKAH+NBw/BdZeFHifWUaEA6pNhJwh5KZNqS
lfb8cwSQeS834ECiLAmqSS5tuYOQ9WLSYKJfC8+cd5lci/5SfSaeGtHM5sfTiD1qtHlToVY7aY00
6D/+TrgOyKXLqGtFo6zlzw3C7DeCzXtqyPR/0n4f6uTrmfFxI72MiDvm5qdO4OW3BeeklaJlElOe
SywR4FqWPgT8moD9qxxH6hbqK0VM+4+qbrMlBWomL6tJNi2wb0vsWkhId9LMURx5G2mVOFk71Fyf
+hfLiBLWrargGx30T+9jApsDE+xS64hYFavjcvrhoIh1dSH5lEKDXczLa4bNbuae7DZW/HSkxNRJ
ZyH6+9+EVXwVN983uZ+rDTA7qWMJgnHmEEv9/JDQYOLxN99udbHUdqyaNV6huDJSNJWfv8WgyDoe
RCsy3zjSlcxqgMMtuOOdTarFzcmnvAcTwbfJsjKl4K7I8XLZ3nAtTbnmxDGZ3dOJcUDHCmRSGEOC
c2RRyHOwdBMa65YczQqgpKH3wOwIr3dz0h0S1J0KNymqwaDrjwGc33zr4J8D7ZSdQU7mwm5Ev4P0
cgPY6T8yNMTblfFiIivQR0ZG5rsv+NsqwSPX0pgjcSCEiPUZZUBTozOToTviXFNAl4M9sHXnJv4l
dQ5Pb0WWdx4uosWFSdKX6gqBxciCE2L7l8Esq4kcBQnR4M46jNJNcT8lBRDQt914xzKopxwa0RYD
k+9wcRaR1XZzeN1MvUCPYF3YbTYNc4vY2iTTeYvgUtLxrRqfdlDTJ4vEt2t8vWlxIxkd9EULaL1E
GCakLZT7rE/+kJyyCC5QP1yEiTyvYW1HuTpZtOrC4irngqOe+ORHr7JGViuVy9H8hm0RRi8Lybwj
jPdijdjh5nsIXm+DuQs65X8nQP2wQqjn0Nuza0CcGRj0VhcO3eDYwf4vHAtLXy+SaAvLgZ6VjoNx
n+XllovNynPCIsT2Ef2sB9eXV14yTlEQvBQjo9O2xMMSxy1K6NQXOa3VVyk6EZwrdCIgz6nWn0c2
1fVyIm7ErujkklEdAl+4nJlisZyteR0UzxD/KpjeuZ+8lt1+L7DjRT/2HgSWuBQFLUxv+DVzpMj/
dhTnqTYUtV0kKbX1/2pJbg1aUa7m7N/X6E9Cf51ExTHKHKWeVkplAXaHbvvn5ITwABNU/Ma7pCrG
+ob5XkvW70FCehrLppx0JfiREhbIgZTaEYIrzwK/yi2k5FTkWxRw9IUbVxc+qUE3/o+VoiaPn8hQ
6RmRzYbZ+TySibt+DSjWrw49QgSWdkhbF5yi8nrKH+QFsztlnpdC9xg4aQ9uZR5hZYphekULCwzl
F9D9wrbb0orvhj5LORsYPlU//memhbCZh0ppB1Y+khgf5wqMYa83KGKcO8Vy5w9H/qUuOH6+UKWF
Wj1kZJE0iHU7uSHHzQCtfJvEQU46/n7GAz/g3NqbxFpToryR9QQSMpBB8ZxheYYdsqmBjMkXTmvo
Q7aAj2ZF5DW7KG1BgqlhWcwIqRHkzJQd8bQ1me57YbyPFSt8TBiib7EKBs1TL7Q+bkf5kTrO0+cJ
Uo6SuD7KY9KhOSIfqAgeaDZwLz3Ch4ls9ND+P6pVONopllgCPi443PPHi/vAMloTbZ3S1SYt0vui
RiWocB9VF/ehjHEoPoXHsKQr/8awZwaL4CIq7rYa7VhAfUQ4U1zY5yIdwVOGFxLHL+cpZQ2vgI86
YKm6gntFbt36xi7tBUygzLurMfIqT3Cuz3RDDhUn8SlMdxyIOA9mZ3ffP+XRTNdkgpPvIVKCvTYF
+ShSwhduNx6JvdlSNraFsV3WU+pdWOWh311MBBpZ2bTblzzoAEHgPuEYKCrUb6tSWmj2IyXBxlB6
7YkikkyPIPdiWlvD/rquGBk0MsN/xVZaW7q31FWTItNSxQBCtG7LY9X0aaWOxOZONwhKZi4yadMz
/34uDnoJGWZtbfLTjhA9B04GsQ4HMCz9tleEbYIrSMZXZu98FOLlK7gyJ6sDynkViaT14tZ/fz/I
KjOb1qT77Wm0PbVAFuMhh+WYNE98jjTzBZh+SXLsuac9bz2WvPIA1wLgLUSly834agSwcHbstKhd
4i6TjacMBsQI67YDJcpaoLtxIc6Yj6JHGm4mtFibrJH8Inys9Rk7/kMuA4XiTPMDeLDBFvzk7cjZ
6PUkjmy83MoB0t/Rq3WftLLvxR1f7j/J8HOu2EaB5iFaDhBXu/Vkh/6Xdhl0HdsmUieQk0Sek0Rm
g6X9v+wjk9redu48UM+4d1FpPmW2edVtyZCzMYb/Wvm8OA2iaKuddN96pOyeOHMcFvXgj9mf+AMw
mdVzJMNesRZoQbW1kvMOrYqnExLGF9LiHrWs/VOE0zzSc7d6Q3c7aTQBOoK8+a27FviPq8p2btN4
w8cheHKeQZphHXoFQJPRou83Xfi7glrs1L9z6bDNBOyMgdIQR01QEpNPrUES35cSTYawYUbRRZL6
lV/W3SI8Y7HfTrPGDTn7grkq3UpcQ8s8lrM73E4gMsf0WkCoI+kAFqsZA5inErBpauVwjGUa7e5q
6rgPQX5HQlfh0AXe18IYpLUE0kR06ZrGYo/zMus5Pi1NKnXJsWEs8x//K4ewxzSygzFykIxtQAFA
0tUcA1HtWYKooGfumiu8qapfj0VJdhNnfgUjr5vzG9x6/V4dnQoPNUxJtDwBWVl/BA8NGjAxMOfe
g8rqYvbXjKi8f7PYA03iYOGiAueftmYug4n6liOjMYH//lcpTJ6CVRVwDnWiKgGagEV8Uyig3X3p
UDSAfox+aUpQjKQtPM12ZIMWrpgmw4WQ2zGoMoHbOq1Zzo/qJ9meJH+ACJnUDM941HNEtr2l8z0y
wDBsylzDgEvRs3CvWMUizx9vz2yL379Tnre3x+W/SwVE0D5PLaA7XwYSReuAmwASA3XA0BY+Mrmi
uagtjXHV3x1H2Gy+lEuCUOei9AYUWlxCcAS1BBfosu4k/GvQijMdD/1LyW+x1+6TwKLGtjkrheSZ
0GlpLqHcGQs3dnXZxRPctoCZ8gR5xbBHxAD4QDRQ1bnjdxXOQVOjMlrRbUYIpR/4/qinu5QiBU6e
mSXlpiyOQrD8jaj1hJeOFw46XdKP33CBNNC+X1BpnxWWKZi+R05JMRF9DpGty3JUzguQB420YTL/
cadM2WnHDtPfXbPYd0wGwzn1Nrh41AnKb4GGSYCnBfZ9niq1iCN/UaJlTIwrHyCPLgG7Ky38rmI+
0KNcrfB7w/ZwLslQqzSg0/0vda/XnoSJuikQiYNGRfGg26o/caWLgMt9DZSXZ/Ci+GsA4pv8BFMX
F3L4s/QgEZ8V5rIp5SqtznVA4RDdm82LdfI0mIJD6OWS6lh4Vu7bCh4fdcZsvu4W0FWqRPn6Kpc/
aW9dTT1uKR+Y5VPT653oWcYl94+hFVDu/1Q8Qg9b1s/+nniWVU20o6JiK9ZniqZdR2JonnrOj8z1
fASZ18de4zFhPCMmdriK0bGbfshi6PqUy+gOXeIsXuXQW/LA3VUM7YGKDxEnZaLG14VSUN6Y2wCq
0NeqVX3HCgmgPhmN7wHaZq059Pjc8wuIsO+oS/iYMWD7YiBAAoFBmPuZudllSrr6KdxxKV6sob8P
2cH2uTIqOZ/+eSXiJa3dEj+GqmUgS/BIcS37Tc52Rk+k6A4yLgzYla0bgITygd3T3pjxgClmaD9I
NJIpX9mY7UDwwsoQi7gTcjITCOppS/WFi5abuGjd0iZt6+Huyb81YBLKmcEZ/RbA1IwAlcCS/QhL
AmC0s5+qxFCgIwmPT/DM/W4by4KId9G6BARLm/IvejcSjdtS8cjmpXAPur85pP5Kv+I20bRoxaB/
xvbou0qLewbmorsQaWUAWMzzGFOv7Iygj7LO5uX0Z4NB49Pblq/AjgIv46G0O46bh7jnRClyNtSV
20Ej8ZPwC0zrSK0mmkM0bbcjkrOmPnpIsaUQ3w+IaU7zEhOr8TpRD8A82sK3Yp1xGmDSr4geCE2G
BO/idtpCXez1sbyjTEj4TT/TzCXWFXHE4CN/tEMoWFeEI2h+s4TLar1O2KTs4M7uHPvp6XRvDX5/
2/PCs4ial03M+ObdwRijIiw55tKt45+kGTvmj0LhU8skS2bj5C9Yl85LGAe6QuFMP7GP4erxgpPd
W2/trC4kIfNpJlR0p1gs0JL9O0ouoiDtes0W1C1Ed35cl7SRXCCFj5R4PgM7puU0oMXzffnbIs3O
ey39h/AA/pFhJhWtZkLEYONjq/F6qhhcL/bG6hhBk/7cQt4LmV0UUWHY1J1nl4tzWh/v/dJ2JraY
1L+4p1gOkruLWpzo+lXHlDh/Cfj63abF36W3uidxdZH8gG4X2z7YNhAZdhZzUaO6V9YNf2F0HWaD
Eu6yJTaNb9jLbsHuLtV/y8GJeq3N6YRVO1LNxaAFOoOh9Cxoh//cE7cNNHOm8X1AXxnTn5tpDS0g
8TOP1E5mYbUrPgEkBXfARtzfCvXsNfQlIl6SqPODrypcSq03jiTu1fG/AurJE7XN75q44jyKQycl
YmhT+40VpYtBv9ZCSslodjZGnr0ltec6CwYll54O/82oONy4PAB5tUMsCsADInC3sqHs1iIupCMJ
pEt3hBlgYG8K/2dmT1B8vEqi8fIO8hjmZF4YK18OobSWy1RrAmvMEKA9lFpkAxrV3QEkTBXjG9eI
ieOq4Wanocjp2LE7xMqY/BCMGQg+uLstL/MHV2O4/sjKA9YJmcsoqpcyEQgWjOIJWGx4iCANHdW1
9DTIRIORGOodzjeiDJav7YzphlvdqwjAJPLs2RrBe6UnRMkj+qx3Yy9Aq0DLlD8L/guKaOmonkIZ
l4npnYW/m+qnIfnHdFV2kJ4WFnkGZfe8lng+5KjVnjlECid0S9k+Rp03g5m9+YMVtBodTO53MAGa
7wFmoG8HnidF19uKiDyf+7U0NM/2M2RYQpaeR3cONdSE4q2EiODqP5INaqgPB69Todz05GZ3FQFh
4TgHz2nHfzc7oYMh5QKUyKa+FsHda/FMTcD1XofdJo3hHQFvWAJy9sPROhesmRwaj6r2rAdA3rOX
Oiu0jtuyZAKn6asyh32w/EkngLIWtQXa0nfZtAx6uc6SyzqdM/jCRzFNNx/i/NtGgL5drKMCM8AK
SvetN0n3cOAZCpRidkpRWLolkITguRomoUq0+GMW6U9uUSN3QFn2BhKFrfbq5K/0g+/0Hi/awkzy
yxevevG1kRx2BAmnMD65CoecTLbE0PD2ZmxUB7B2lRRUUfpUZKt9gRmo3a46DSUlKejVBfRHA7f+
FfgLOM2YzGQKZHCh1rWpDzjtGE1fqj1cpFvAUq0gGSW2M59lxuzSn4r/XZ19dGeiHjG8Yj77p6gD
iU95AizewkNg5T6EiiK0A5RsGepBfa+U1sm6zV522ooZRndRTmyr7AelIsh03HHERRqnSXiHZ4Z3
9cLz+Hs+3sg6mShqxc1fE1Sfs5nnMTXpnWtdHtTxmxC+YOCgMclns3Nb9DuPStxxU8XlwzBL1vvy
pcdMEkJIWOmhSIBhn1SwdTaSb5hQAhx+o3LKGqcY0N7ZPMRJjGOtrTlINQy5pK2JsA3J3RwhPo8C
inELR6AxsJ/yNJpNZsKkCq2h0cTKvs7AgfObWOmTAxkfurGHxJK/EiUIls7RJWE7K6N5uGxWUoii
alPvAs6oP9cfZ4FotcS0XQq8kHVLwPoEuHN7nzMtrck1ZNkI5aMh6tr8i3ZSR2PYh7Au/8Jt0Ogg
eW2m2mJEO0kF0Js8gpOcQXYm8Ia95YHu200Nz8w8GX/k1ddDWI18Qa7kw+FBxq7p5qV0mHVFyXda
4T8nYV0xqlE/ErzujIYU2mEC5w1Mt+3jHHSji7CMYYPdFf58pyIbEqDPBuRS9CyHfyjdoBj8Tp5F
gdip/5BPJa3TzyOymHey8pmhRlZgMH1OgIaYzuLjPnZ/IVnRM6i6uXDhPlCZMMXW+qBC5CTvrDxW
hWR3pEjeH0L0ra3ar/obD2IKmlorN/IvHLlygUTEkjCQuWbawy6WWqa5SoLW69AnOOI8e+6JuI/W
S5TAepISVMJ2EvsmmOvJHCfBaFLClssohEE6mquxiCeM9UJiAJcl5PhR/Sl3efYtLi4CrBpewdGH
KlgjbnaXBfw+IO7tL0VKNNpuWoCMCGcOC6vDTSWPjDeddSVkkvQSW5Bm/qdjVo9ueAUQnskvWXMM
i/M3/NzmXIedos1zXSkXN9qjZbHqvUfKEot8GMUNgDNqmt6BB+TNjP+51uiwxcgip8kP3oPaQ4Lr
X63qA8sVGplVPk0G2pkFYAKFo4acnSqA7gFBN+27FNUcHURutZsOPaiaIW8VVFGZrUm4tasj+q+H
UA4xcHvtadcwif3lXngbj3QMnYSI6crMohHqJo1mLHfT40+U0/xRfaXej05iZEbZgJcJimVA/EIh
kB/beZQCIpKpaQ65+YO7YkQDTCML1IEBiYB0Vs4DmekDK7fth535fVPiR4EtIcLAMatRYe3pthGp
i8uS+lnPJhe8AzU0aRJxwqTk+RRu7RYrW4cubnrKVJBJfXbyiJUcb/zU4DmCNH5jSevZ5svyQ0im
OvT3xupDz3MXH1kAB/wNHSlMKDxyS/va+36zLqHQmW4PHvGEgPNtEUBxOQHnGWOJJYE8sJwEcr7m
6oyNMjzHTkLRzWA03yFhlSQu83KsP+ox5PufHVmQLhjOE3yro9mTP5hPcYGjeoeY0GLvft7dcyis
M8/lC3UigSrNZo7BuoPFCuGdniHc04MKpqKr2hG8C65T9Vco/CC0k7zjBe77xWiHXh8CdUJDFKJY
0xAyf7BrGYEs5zZtg5a6Ph6hFXcF5w3hwkdtEaHDg9H7/RDwDxZu1deXUg1cxlhUfS1Gjko8H04J
i4+ViZi5ySgIkzk7asdfbMS6u2JQRpVENiphLP31VOD5kP41H+Nsdl/uOqwKH5OVyew3fwMkCVbe
DC0bruW1g+lIsFI1skGPzdi6Q/kL7RVY9Um4WTkSoP4xbx4w88WK4KF20VdqHvH+xsmAjXLVisnY
lnCuzcBGnEXO3pZ362pJhtydvpuBzCLVOPtQIukViXTG+0MLm5J+mmRQXPM+QuRCC/ZEk6bfVyDd
mqBvBuMiG2Znf2tEZTGvVMNoBrelFNKifwNvZFsIs39T4QFWR6uhgcl9F1i9t8cqIWgdIUaPjM7W
xKx7gCIQDRjulzDUzZfO3E5aZFMJJDvEtTJ0Df8cAax1Mg+TEzzOa0nlgAtZ+z8S7KBsx+xKdbtb
DJJUCZHZ600heoKLWgGtGa6u4xyE/Gv5rb+05ZO0k7G2nIcwpxGc7VUG27Ned68FuS92nAPMo6Xa
TldR/nxzFlDYCxVcARZ6t3LdzA9FWyWLyfGQpWZrZpl9WyNwGAqgkMHnmZgg5IQbbiMb09fg94lt
mJSOj4OhWSk6d6tJM/NTnDZFuvu4a5GhwzU4hEwaQ1NNktnqCWSUlDysNb9iZb47JKF+kSkOrlFJ
HEvne1axd/fipF9kCmwk83MgZpQIxinCy2x1bIS6JjYxsFD8kEeLPbTkhRkwYItOWd+SPeKhjZ6S
AokUXGdLqQswj4zTRcTEm7G0ftDTGW4182/GCWaEDv/Z++r0EY97Oie7HoEv9+daiNl3Z+9Re/S3
CH89Jk46zHO22UfbUYMTUhyLWV/6HmNSGHngL1wRCsu9x3sllgsCmFzFirDU9hANY/42vBOaSvL1
/YzKi0rJa1GCfmqsRLRiqizGtp8yg4CpnKtHJB0K9QGrGeLO0N1knmm3lCxhgFWIKawM0o/H2Xg7
NpBtWyJ5cpUkusepO70Seb1sgulQ+hhQgdwOiU9kpOaNxh9bQ4Kr5g6MXT5v30ucMnSgZ6b/bQfJ
YeDPQOcqYjWTnWS17RoytmsdBSnBO5ZhhbaVyN8vr4uS+ZWknrDXlVjjQ+hYHshjSkLm/noRkZAg
Sig/BTQFxFeAJAkJtDtkYJSbPKWdCwYL++keHmUt1WfXm7K4XPdVGNUs5TIUgD5xXh1RiYRnJ0oO
u3GxnPHtIOUul4vsMhX5uP13+8pqhMcY9Qfx/zxoMLCwpUEes1r+fWbwxEdp5AzkHrIcyrVxENxr
BcfJdCb9oHQqUjYpRByASPav5IwFgzv80MG8FNgF1xIX6qnM5ypgl2CScBZem48Eu5g1r/jcOypo
tWciJyq/ZN5u/Qfk7FcEcThyUMuEds8LeRzR8RaaCtyo6LM/Irn2/msvmyU5f4uODY6NmXvRFMY6
kpSN8ir6dUYZLAxHt6+wxDgz86vt/H1KQQNMl8jeyCg54K/DxiOmKfxslrvfNeZZGUNrhILbycuI
EOjI2+y4ycUUK5V1Yp1riukVtTt9vXvby/DJlO8KClMkZqR+vPVMtktn43KjnlKF/mDd2Xvwjsz4
HOs3MTx1ZyBS8L8THMhxVwi15X+07BfDYuj5koX8t1OBs+Jy/cHb4ilxZNkiRG5RfVRHRMQbvk3z
TrH8YMovFrZmMP+2kAy2eKyZsmLpDvSMcojzzK/g3cmRiufJyU4y6PlubNk+1wtPe5ryBcQ8rLpz
VdCu1Yc3mi/t6a5Z8RltXy0Grx5lyQgTB6B2IHZzGUMNh9eq/Z4pXQmK3UfKgchd8F9QOMYbCAZX
61hqTd5ey9sxKYKu6cMm1hyokxJcaIZZnpCV1d+gDF9oQpoZGagMm7gWqE0hUgO31Y7JxwON3OTN
edu2YpLMdQzEmOmLNBADiRDnkfA1OOJnc/Titgx410mNBjOF/EMVn0pZZgfxhahmIDW/viCKCV7n
Y13+gbAX1XOd9gLKQZjFrALZhXAo0wn4wr3WPgiWHoGO4pUzPeZwNfDbG6CCoo57NSVWolosbbSQ
T16iG1dq+EYuTdzdwIId86GhMHp8z3PBIWLEt3sVLYkI1WOW4EUMIoMQ4kAzfrdISXKiScoX5QZW
TUSckrT1GNz9PyVO2K/K+CMLMlVYyAJAMI3VoOp2anYrgMdddHiom2qD4h3jUvU/Xz8rESe7JHwP
8lXjiJaar0FAg0MYv0y53F8/gLHeFToj6RPa8La0mdV8j+DAQST515H5vgewSFcHS0Ghral02Bta
TfTVnOJiYtYin6rQGLnRk1ebxABR89H2xOS/BH4MBJe9cTQm+9PtnZbaAos8Rg9DCDBZLqm/tDuj
nkm4h59OhIV5+ltpsrAaUody55sHR8zHt/6HPK1UN5SJmyD2wSXRuA90bk0c6osmfG9F6QWnEGuD
JpHsEvrbAZ77l6jtpVnSVfbp3IXsN9+n40KXU7Jk8A377N9UPl7NdOabS4ReH8uepaBoGZ0g1e5s
lmafqrXxYxrzTOJNSdY/+u5wpzUSXf8l+e0tI72gS2GlATlG/hQVVkfussk3PBOFHhQOOr7AazAs
jxzyzuY45R5slxD6dalCw7B2Y1Wz1AyjWpeJLTrYk6vZEjN9htRNDRe8tkwDgNvyJgv9hqkul215
1sJEI3HzLrsgd+ZLomUDTnD3gQ6FD0HgcjXA2OajcdnUWVkgAVSr1Qtrw4Idet/YHnd2/GCSryNo
Jsts5ahi0An8ln3UGwAM2wp/j6sdNuaaD1POogjjXZPSKUlM0VCWsQDSBfh9g/JMPAp7E3Bxbgr0
yIqS4NNJd6b3TgzqEg8P3zTMfPxtSmhSZ2hWCSn5fDHd++gTFHLBeEhaklgI3KwAuilHKFeeBPo1
e882dpYwRekbb85/PNLEuQDygH2jaJRixBH24VZxa5pzcLUfkra1EFjSGbzOvi8sNtcnCZ8nQ7az
9jW1DbniEvMF3xFVh6F3QVz5sNIJUBwdB+RW8ZrtZzPHnqbr2JOZrypQhTFyrnittIS4vgWDUBFQ
ofu9v0UQZ0bbmu8KrUU4AZ0nvICMEqBpBfkGfRQmmcmA0PWx2AALUS4PT8v0HGInMva1LLO/ufUj
QEqMaGBIoEzarpgQ8BVuRnoucWwgWNeOGuBHSmvTtQZJocPJzw7liT4Z5QVxriwXOicniRD9/y5d
ymi5GdOGYA+rbaHByY2Cud7eh0mFroRYJc0ZbUxxjmShWKNKDQFM/cOQuOaRx8HeNRDCDpfItJQG
kr+u2lV4DXH74QMCZ/R0SM1UR5X8x5avCAXQeF/TFeJT3ITvEdPAYcUS8nDyiFKxUVM41TzKawjO
8stOW3FQ56lCrT4aoKoUPHsbMtSlB0Ke+QPbxINbMaNgyQVfMSeuO0pgfKPUxcsfELmGlDX/bE1U
a1ZYc5FpePtUcNV1T3vjRItyMFfMmIKdS18aDA8/aUfZdkNZk1rxw9uXWPba3QLSkMS60LBUXHyH
tSis01oH2zhvfstEDC0U7rCMgi00xM0U28KMHFeGCDzFDQ3vuqHaAX87ENxrTO1hyv2tRgE9p7/8
j1Rg+So2Ie1fwczYCFh9kzBMaC+csbXYj2u5hjh5N/D8qpfsKl3GNSHngacWHZ2eXa8v1m4LB6G7
DI9h9RNGiGswHazxKktrRq2RKq1PYajtvSY4xt9kXZbCAnfdtIwcVAnf1WcyJ+5npRd7s8dJLH2y
OVY+qKY9Pz/aPmh3THQIOjik+uvZY9b0k/z90CYvZVO48mnzkFtLOA7ha1j6dSUX2Rjr0SNCL8xQ
/nquhJX6cTb0qk161zlYCd04c/hsUpaZZb+l4a7VklmZJzdghhHA1rNibbN5gO26AJocq3R9vJUt
XL8dK6/6otwMI+yyaVJvO8lGyllnmsvBt51gOzAniZ4FFBhCpYlDEeG+MNY1OgthLr9w20XM54Ec
mG7+qAB89nCEmebacQUguS9CJnp4Nw3qh8tOAp3v3YZMETvYByHNyKoG7FV76PydDiejKsa1X/Rn
+cXm2zNoupb+VfYjJEB9qWgmSgBL9hV/4Hk09hGbxGiyqhKJendcA4omwMvKNV1JssInwveQ5QKN
oBeWI3yIhfbw9cWPb6r74EIBTighjuSqiaG3Ra1jkmW7Yeq0Rw8msecGlRobQRKdcHy+5EOZgIyD
pbJQQRtdxRBqIN3GUFS9w4rNlwjzHw7KyWk+EJ4SEPtdy+bDgx6WKl4IjymQ7b4xX154Xt5ZedMW
ZV1pb3h2Arxicz6mUgPc6ndGk3e8fPYPAIxnst9dXHxxL6+JXZLuIvtQ2jlesgbXCMYvU9q/SiST
GYP93MaM+uytsbMxDLpmxAWJRnOjetShnmHbdQoohGWp8WzATB+dVd2S+zk2f1By7ZX3ppf0xhBP
EdwRXrWZEVX8nv1qNEyls1hUeXTLbI9uLH0DOxl4PkZup4nGxZJJWKme3ibuTSevgI6MMOKEhesJ
Y/5A5h3VypNfWJ1pYg1fE0T4trbWz4jdgE5TNS2sM032Q+Y4rRarFGSa453HZWt1S31hLE6iCVrF
HOoH/TJBnMYjD6MIOThWQnbwCjuwEVu90hn4ckgc2zM/yXcJo8OtzuRlCSYtHo0xHdnLacMvmRsF
t5n0eO3yZtcWGM0SS8CaNoWC9lKcCdW1pcup3LNP9IweUfPPJba/Qb+zgeclbmccwWfv/V7H5fkM
/LQ4z2dLN4gTPPp9Pw9DekX709lHt0IZBllPQL5NknwpuBOR0us8v6UmFL4dRgXW2mN8/qZY54B/
UmqKzmaR+1awOkXV6eznoAnVCok0NIUkSuh60wLXO3F9WHlMFgjHSbM9uukfFOdIKimZyQerlaSJ
Hbz0qn6cKbSmfmacAoZ3u8K/9EmYs5vM0bBMtmSDVYy2uZbkeQWPP3/lQp9ch4vwcTNwBDzRf6BG
uQsgaDdlZUSJhaBlmc80zICwXb9nV4qjdb9IbYUuRX5xYrQ5CnW2yVyy2b1j0Yt4KpTW6/W7GMwr
etP9qQZEzoa92oHNpwTe9X2OFdkwF85SDHGKqHmhfrX75MFeSb7wtvzpFju9vp5/gPH0YQgI58Cm
fAJ5mKTNf2uNZKcPiQd/2xbRr6T0OYUHFvRebK0pjOHgk5pwYbwJJv6zGhkcUCEtYJrkoiB3Y0FX
eXH8oUtU5dU09ayKjK7M6ouyqeZVTVwPufET9mPlihbRFT1sp66c16yDspsJ3toxVzc+6kgigIAl
nQtHiw0cPceIUhTWCBYe/36Qiio45mjryzo+kC5JWQKeltR4oaUR3YUcc3WmMtOAMzzR+uN1xBzq
X5khVSRnMv9DEl+DdParFm/bvFWtuKWAVtlGXFO2rP5N+FA2ZuOOY8HYOJHF6A62tSY+VT1jCSGX
U4ZMXfCWDAMi/FhI/lbc2yOupdWinSru049qXjEIO3uHRcSgqPZIvxGvmoYJi1bwc1Lx4V64E91+
zz7lBHj9V6nKevOAR5woxn1hqgp9q87wrJSwGZujxIJ3F6t8PWeTZiXcIKonKy3lEJxZAhV5U8RD
HpiO1BgJtp2J2KBSnRG0Y+ujBVWF1bcAjfl8c/uIXh1clpIFpr/kdL1cQXfZgVXlIHj8i/VLp29v
w/e+XEXUaeoImqt6d92NrOugseC85EVEkkKFrjQOZ2MAWi/8NQryXZYhUaOa24XbP9h5xrTMWgwZ
VcpHm2tXP1YVZ6c6IoqMrV6ORu3ksces6lcWt+TwmE8Af99JgrwMkJrWEXTPGLdCM9bKacGBgKKA
L4IPFZZMrs7dsVVS1SX+4LNWdLpFlcwFTh6V2U3J7PGnUFZwBWQsWIkQtklLh+2Hxmn7SuZLwcfm
Ief1SevICSTszflBsENK24ng1uWYG1SvzRMUIajIFY5cAuuSFCvGR3P8/NJyIxQMA4YrrytiJWOR
uWDzTPqqXeaaVlF7WR0e2dwBZ//3Wh+pH8lwWamzYiSnBgfRH2DLBVPOm39UNw8b69PsoDR85eSD
g4osfYL9iG6k63z5hQCJbkVUwa54EOPtBzHov9c7IwMd6tXChO88D7E25Sb5weslvcD6ZZR+BQ/c
U6+lYsK80mnm9fQdo1KegGCEp9q6MFoP7AL2UdkXeMhf2ozIhRK9e/BEw6tY9m59yXooKtiyZhOM
Hu7xMgCPR1XthZSVhC1WcbXF/EJXGJ5MVrk99Cooe9BbJURNhj4odzv0zNP5MrV910zbTpkvQLl7
H+3BYpDPlm+4C1hh7JlZRmHDegXE4hw1CcMwuBW/VTfHKGPXvMWvsqsy0g8NvE4nq2fQ4Koyr9rj
e7WgToztbSH7bN+g6rs27SW1wF4hgHsVubMMWbgcuuEX9oMhoCT0QVFyevgPK/aaf9EB39TRdK73
rYnUhJ2f4E59NFM3VpvlMuTO3aCSGYwekYF8C+uyZLbzuDtkWcizqCeKUF0qstdwoD5xPC1L+ycH
QgVEF3cI0KPJBHbU0uuIwvhB2LQtrEHX3EwyL4uZWBJsWPjlkMNrIVAJGI5Plqg98EZ5x0LYp6U6
FpId3zkWYKXbO1h/ZmIpXYJjTaRmMhXAvLgSYYatNcnzNXpTNzuG6whrjcW39ILneUzN18qPITTz
97KBx626phfg3zqyp33ufO72BSTYLAX7pAdUS2BzLSZniydoRHCngtrGt1rG/DfEFcdah5H3zkYC
n+xj6RvmuXuD7+nYUuzidrfu2JTKWWqIu3N9CjgHvcxiGaTlc9/T1VAKblNTgn+CA3KL3lVMS11T
Hcr5qMyJnHCOMu5hVgc1hmdTvAJEkecKZLS96aoxMuR0gaWX1OsS7qdrpwsXlRGa4jP1B4U79QIo
lubJ1pWnos/sME6J8TBmew06mFrDMBzbd9rAWco0+u6hl+XyQr54JGCfsxU+353emD8dWU5YebpK
lJbHBDKPFdoMRUhCIi5vRV7h/hE1PggoyxdEeR1ukQleXAFgWKuIZk6uCvSTXV2GhdaQmkD75a8Z
w2vNfzTzmTiV8LGoxYr5sTkaYQvb6zJFuljzAvxA1CCUPrdHXplfOoyDKiuqeXy83k9laEtOHZhe
J/0DYLI+FPMTsVU7F8kOd3GHiwTVx4xuJxQ0KaYkqiEG43lBt1iS7NxQOXFCDJ4rC3ewIGj6zb4j
Bz3ktLjQVXR4sShLO0JZIASKxJsDowMdFcWDgYk7tGeb3AGCBoaufueSIMxYI0Fe25k9hKFNaZA2
z3IyfFlT+/+73lIbsmYB/B/Whndn1iUqlXP0rRJV0Az7M+2EcfCnIieY/jds3pPKe9AhuY5u9gRZ
3IdH/3HU3yFn8gRy3mq104KUDf762Gz+mHjxj35eE+wEBvY9myPiXMTFjBJCBepnp8sUg47I67vG
jSqGziBd+PbZOp1G81Qnh7z8QQ/X7O1A2V4zDFz0WJQIsNecjtGyHE9L1WQ/d/2e/2xj1BZG8fAA
HhZAW4sfjAjkAWveOwmH6qlGOWs+QqxT8hItexgFbi3VzzSEJrVIx2t3JwU9E1/ddE96dYTMjPVs
1fLabyvRM3lzNnOxIPylKoMVEEfv+VGDRD6rEeO1lyZhK1oPfdGtexKAc62mJkD0UOqD0j/1shh7
9wg1Y9e8reAijvS5BuftvgVU58KSKXz3IR5P4ZKG+QsBlmV0E3KIaaHsqgwW2i8fkTKhBs4DFoOj
tng38qUWhTS+AgkLV4Q3DIDu1u42HyKzfpgAo4UQ1f/1PI+j8DAcuuwFXRWgBD6NWto0Ud1Be5z7
KaN0YVf6Mt5jNcXAgDxi9uY8bjwapPlMDI0bz00DdsKw92H+Wc7QbDJeSqz+WXJVPH/SaKqZhWRc
M5LtVjfmJPqQ+xpbrqTrkvKjZp/yFTqMdTF46NmX+Z1e8M89qQoCVOcjaqgzlL/23m7nGZ1gi9E5
tAkC4Pzs0yxLqQdgiMiQz0smjzG1tCRe7cItz/G/nz6TZYgAUelERJE4BmSXG6Jl/ObLGmMHuMGS
92RLoqqSioJleUvIhJSCCR8Vo2N277qPuiCLKbeYa7H1GDVh0eJB0MK6ZJmEc2PzhUvreC0aZ1yV
EoISZMJZ5nnoii+n9ru46B2EWF/mGq2B0j5BrF3SRs4Th8m9f3FzoV4YyheFQk+JkLBP0X7jVPa3
XE8LBdPc1LUj0OPuUKAP69e5MWzEpUcf08ZgF6BqZCM88c/+PnTNao+iA59ewklsK7rC/By7VGZV
OcFktGd/9BYrCgOa3RUPjTuXwOBq4uyAyvjs1mm6xrpmklk24879/8dO0pEiaZMnT0FH31af09Ll
VeltsgtZNRdgPG8aqHCKBXrPkbipY8ySBF133UnzNY40HrIi7hBhNwlcYVoywSY8yK+DVOOFFU6v
h99C9qLfauJP+LofcupsDQawfAI5+5fMNzgjxB8j3xNgGZ98P4bP8nu7TcPc88F59sm8D4nxCOKK
r1IpqEN4tvA42NiuKeNUO4ogwJrtpQPzxfSaIuW9/74Olpd25ufKYtuqiH9+AqKuzc3nYQHOI3ab
5jEHiqoNdkaJJzF/Hy4P1ivTfYRumOlU9ymQljHuxyF5GkQYT7HKuQWcQTukqcNyqCW2smkfkb7Q
37/xDdFgqLzojSdeo+4tPlc3tLtFkJcWWkgWaRNx3imWAVH27Nhbb5q7k4ZMRCPhdUnjpx2PYbkq
GvQFf24OXZ2q07w6Wdn4JEgHZrzcrXj809x5FTNw5RwIz0fWORVOzG7OCOmT/imr2DJZfC2MrrCI
AtIryFOHtZxe+7pI4Z7x6KVXFLqQfh0dyHK57uG/9ONh6jemFsgMEiLRTltWVInQTQPGRHwqXIk9
NGMClLeY6LAP4zpFducXK553nc9TA73HEB0ea4lkwBH0/KcYNSh0Z6Ums/GL63P7Y/YKJgjrcKd2
S7VG8ChI+g2trVJX1hs/PSMv2r5pA9WIVyVn3Le0RuTgm5bOPp7wX+1EHRQ49Dpt2bwWgQlNZI5T
786abMNMtKO9iVLdFYn4qa3FvCRGThWfxi6MtkOfUQakDVoOD4Y9zoytlT12vahZg1NHZQhAWamS
yDQutVvjtSNZx8QgTLwlX0SmcYzOj8GiZB/m9iOmj0oVYulM4GmeNOlbpXOJ45MQZlSKmal2r+Wq
XXqglZwLqAz/9XgWh2/50/JYnnKIDrJH4lJ1v1lxwuMFwCzu3MygrFucR6KaXuf8D5Hj2h5a2a5a
XlZmSbDSR9N1RZdSdei0v5l2Y33ySQW89fcpWXHFq2WNJ3YKcDjSNatIPDiL/huNjBSc5elU3qH2
wbOV07KlRAEet9fAemx6Ft7Pb+riuWmDAnkwq+D2+LllbUr1Ag0mXHkRUIw8hvZxKwx3Uzw1RW1n
QUmOnrNglCbgRPXnmae2ELFF73EGT3fM6SY0a1ohBO1WUI+YikkMwMzzyt5oB92lraHdIu2DnDN3
CWeQ2/P2VhAo7Yt25Kn0HyiRvktfF6693zMcKgEJmyaJx4gLCZFqyYVj3ZN0igGBR+QKHPad9vuS
Cr44UAWl5ewyBmXGHEUN3z+4SbWyqbDs66ynpudohM1W91BoCdiHxGlHPP7C0A/9MBP5Uh6HeRMp
+ewgqXGlZDAfxd0YRTRrTetYEzoDvPIQqsDJ94gO7kDbOvT1ob7HuM9r5oAZReNBzvK8bijp3G+N
XI101RRtIdm4Ztho6aG58Nq7EmxDOlgkFjqi+vxnpm+1jFKWPnIKctBbu+nb/g7C3rRLZMD0FjRl
apQSeMs+h7tb2fvtHEHvPsi4GoKToAmzx8DtHoGIhu6MZsD9nNCrwOMn35nluaCNRLMcnN3ws8ta
zBptTW1VQzD5YVW1Po9FDaCLCHY32fBhqhAlFSd4eio7RaAJWjvbqtsfoS2Jj3FRlDRohfL45tNg
nnqcqRuCIaDOc5FBZBnNeyj+EoQ6Gq2EtYyVELSXNNRc7Hfi3F6vzd5pJj1BKkQcIQ62eAEAe4vz
2EHc3t93D5KSTH4bNJ50Fg78bearAB8KJBqDLVH//uMhc1lfpkUUWxGDovO9YoBxQB/jvFt2842Q
fPytXtmsI2IkG1WAam4F8Zm0FI3FMrMrfoaKhOG8PcQtFi3dU2g9Vzx/lta9bcw9QwwHIEVZ1mpj
7IcB40NJP36fEREBop7Zg/5c64kBFhPmJNQHwfEk9dEiSMFtFh1Bd1PXRcc6KpeoSU+OMnO411lF
TTEISLe1tN7Os4mEzErVoYnIuqqa7W4N+8qbngYopcaYyQrKhJZJm+LoYHkV7TPXC6pHG5UAi+us
xJtuaxyjbdk/vloHJXzIGSZ1pEgtgWH65SwvU2vHwItjD5IJtXbUS4zWiGOEgR8Yj3LSVphq+rD9
1qq+yk7jql2p3t9OJ4Wa/OiLnZiLNMRheFhXfKGVDQUWjvDnyOT8izh0K26jZlsiJuC67BuvK1NF
TLK1X12lIO/oY4pytVHhm12JYN+59AOIeeOokylyB6Ybv4JwC3u3SY5s7Ts8Io/uYi2jcCmI1Ov8
V+Di7zIsYAhmOeqDFEI4NfwN8+SpEgukHz9N3ISXfld2ywf+CxbugUUTn6PZ2bYrZK2vcIwlBeu+
xxcb55w6oNPfrc/LVBWBiQkQnQsMmtARg6m+PqYhimyd1iTznPXCZHMu4VVlibcXaxRNiZ2vN/XN
y0J2QPg94UevbtVOOckhPY61TJsyycoK0L0nAkzCFjm2KTGD7NVZ8bI2OZ1DhADQuyiS6a7LgPwd
O6tUI6IvhgevLvoR3zDVyyS4GUxLwDcUVEAoi7i1EtZc8t4iQt1V8bOqqwIf0l7LzDwREZUZqW7s
OXGqdznZX/l7dKmp/PzSSfDb5eyfY6PP0zGhFYkTa5ZsGbbd573CAu9eFSdN+9vl6wihddF2PPyx
OGZfotA9snl1UP8jkvU8g5GIHc3L8NJNQDKos31A4ekKgnNnRmruK5mT+fagvBRxakvjdzKn2CZL
uc8062hXMP+7dT4xE1z7PQYIxIvQSa53dLgYHXo0beTxzhS3mwy2iDDxPlvldPe0Fo1m7pE2Mz9y
HT0FA0vtivPP/KG9vyaYckuhWljvpLkRnds2cNfn6o6dXK+Pler0jqmM290FDhHQNv4BexNOcAed
Kx+4iE7CCmlMZygdG+7Ew9whzAoKJZyvErwWtrTWVNZjxqd81cOsi2my1IbBmG1hx57kWaX8eehI
fG6EigZNghIah2QfQUBplHmbpQ5a2xTx3ygGWJhwH2xOAhL5U6eeMKPD5qr/vIO1VoXFXtftJhCe
hXjBURZlMJlHUbEiQ6yNLInI0DCpu/L/kTtXJck1ASLZEFD5JT8QoztZBdr3NRqzse446p6idWvH
wNhbHOnqmPtqk3Hi3ezSWxESEhj0/67Lz7d5oCMoTV+WR6P+JSG79j/BPW7ZoHTRNLBKE31SHL/G
6NI6dOXRi8A6+9M52WfzqKzEV94a2gSUTwuzDN7pUkZ+ptmWZnEG2tRT4lZFwWB1lGN2Veske0Z9
9gdiNwxjr9AFL+eyAqrzXtOpaxbEFkPgirPDkPw82ReTOhg8IwZxoz3tKBJIW6xe1r9jACGtoOq2
5tHvtLUhWMge8wKqPmN0ytqbY2meFX8PKUVlm0tbOGlbxSkm6AcDT0hv7ctxF9EsLIU8+6cBVU9Z
ZOd6rdWGWEnq8jfOLFCqXxVNtoHuj0VaiVAm7WWqlddDlgN+RR5ZziD9mFigeMHC78KYiuKpP7uS
0reS+xHermx6rhruwgfFNag3Ubw3kSpFnJS4GOXzmj3Do3uxXK74h0BAKb1DfafXeqqkpZnwklBg
47J8cwK43Rf3++OJsxGNeyLxfwRBIKJofSBGeqtpS/ySwksFmR8fYnhconOXZjmkr+Vn206y2zgB
eJCQ0XHg90XriXbWdtlf28VvF/SQ2NKn0It09kf0mit1THqzjFt51awCe/NOZMQvH8cHA3nLMXwS
zEjKI39MoaRbftt6niPtOWjmrrqFfb6a0rg2a0t9CocBqqQxVSLd+Vlu8HXjarnhTgXh7nCU96g1
N6ro8LRoyNnV0O7RAcQb058J680a4JYR3OAoojdx4PqK/P4OSjXZG7dNDF82EySWe4Huu6/N4k6n
iFYH5Sl1Tm1d50JU6B10BU6PX2+5z7hgCzS+qh4jUeo7B3+nWgi7pwjvmM/8cI/9EBvvPj5ds0wp
XM5Y0PiC8tiBjQRpo/2GBv3/0k5LXnRQYdJzxcWPtKw7xJraxYq7XORYJ8Zs32KtrGPzHI37ovAi
7sKZyoHj5Iqgiguih+zqVw/d11DozCUzRLt2csgCWzjm3XHtsIoC3qsBBFvWGMeetT9TrIZ6EVvQ
lBflmPWBDmf5W4ROUva22Wa8XS3YZydVqwRHgq/m1zdapvq8YForCpLGaX3yl+SUrAS0qs3s7yEm
2MYVRV4zaYfnQXGzDGKwvOWoNhKVBs8j9ANFz+B6Zz8rN8Bif77Ql5LC7lGtOTQNniEZmu5ZUVDZ
4Q6+RTe81cvqTBQYK7fzfIxDIXBsAOyTO+RvCRpHmbCICM4x3XWx/bV/ztjvUMNpfrx8GliObHyw
P1F6yjBzYsaWxnWSpi8YAAAYguqx0h/+08IO/ctSlLb26FjmRcNPezXd3amPjvAvfK3n/8iragYh
SoLiwNczL92WwKPFh4+MgNlW3brt0Vo7M4f2enAnyOD3pL4hG82ngaFn+SQFU7SSRc5YjeCBnddl
gyAPPAtfSHx2fReJSpe0ys1CsLhf1LDQ4r/IB4TPmaZNxvSQkgYLZZafu/F7cdsO+QJttYRhqgvB
2RVswrkuLoeKGYgEwJm7BrgtR6pZLHAoBBAXbkIi6t59TuWn2uBOfOSH9WbRxBKiTMsgTnEYnXQG
YDiLK4/6loWVW4jAY5hBGRhj87VA3mXLPUoGSMDRj2zOfAh/PKAKsxaNtTjV+SENeQTCACAUOi83
YndDbUJ4A0Z0YGzbHIw33LZj13/43hm/nDjvwzFe6BbtWq+QUV0lSQSV3ajlM+/ed+e+knVfZgPe
3WxT+n0d2hRTTEhLjCwPGhjsozMsKarveaDqBeb8I9LJxWywYr4C8qVy3JG3X6ksayasftxAVXx+
8H4oPn0vsCf1r5QRPxX9SxN1TSvibz4+tuUywk5VB6/L4HkxdKu5HgQhMUtgHszVHd6t+4ar/6KI
DgB3iVye2sOb5fTeyQTKFoWKPYCigm+sjLujaDGHtUQwmmGNaBJOCswFmV14FNMR+kfZCgJVA+B1
z0aPJZg5G4mnqx+vdKdUwX9SFibkdMT1FKIad+clwefraNTAYDN0LI+OpzTATcRRoFyHJM883vcQ
wlfcGrOnsmWgLY2DtcQb2Qobc0tk9xLFekE4hLsaIH6B1L3HZwKDFVBbsI1sgjmDiH9HXFtzRLCk
qN0iaGY/yy5tKQ+xeQZshU4RFE98wxlVCMJ+0bh4FzBGmCJZL6GAV345nvSWBbNhZbc2p24eQToA
qR1GE3QJsQpyNexl48HrNREdU0HmvY40CMvvZuPpC0GKkIyAEIGGHeVYb+nCj1Gp/KnJMsOYJPib
QyKgwRoxddESPPLxtlFeXIFkGWhWvvlmGBgtPQwd0G2ie9+/4ZQTMDF+3OK9UBjZvB7MHj+62BJa
wIamKA1wBA01x+SM1j4rMmO7lVBl90fQ+8STh1G5oho4RO/N/0MdkERcoYLw4KFJgjso1yIjUNcs
ngYJOwAT1O0AWve9nY9VgIK/ZmNqtQYBeQQJpSOy5rNcNdEsAx5TdznRZ+MHkrWIfZCXpZvBLB7y
hMPubgdLG4N9q8X8+akiDdGw0hMVprVseOh4zmyJ9/IS8b6EB9ygeKfkGD8loRKgviKg5TcHibGB
f9t7gvH/UIwMF/lxZkkIbFNfACZXRIKaE0M4/jxtJ8oDOhOOB2pay+pO8t5CvRlH42pijGju5r79
9SLwo0j/m0bzLjyOrQlJWxSsrCSY7e7m8VFYphUH18HK4Smfa5lJ8PDKYcuct1mqMOgrHIUWXlYl
9gxSYXLdfjtnMPKSCaCD7zEsgdAhiy1VDI5hHXrCVMI33lv/ifFIJVlSK9fAnrsTYfIASYePU4hM
X44LG7CEelvh8Madq/2deKvvc1zWco3AA4pOsEgPJbXeHN8l//17+TIxe++hvWnfGiqzYKG/xJ5f
Z1UBleRVu0r0umAL2B82h61vb2Y/PeJWsgGGKcxWTinC1oVkOK210/X0cMH3k0h9zDPRIYuYb52K
fK/epQ0nS63m1WRia25hKMxhwQy8K9M5DvObxKaT6jKAuFY5cbypd5WG33uFkvNuYAw17rx92P3Z
YUoo3eQESD37J52isHeSgXvqDHHKFJ+S2BSGyH24QTU1lf628aAhbB/rWn0fIbmBKEmUZSfZhYaa
K4abb+iy6dua1G1NFNYuXnubsUTEJ1vwgRpkopesyyY+PZGOlSjKEdNfNOdfxKwGXxKxxuyQ32vF
Zoox6NCQMP6GXNW4gtyVHrE8R20JQok6mD3g1eqqeUPowMcRh3v3+UPiX5YzeD8R4btt81mtNaJl
eO+U2Q0eusxbJMNp1y0PsXj1279AX/8r+BS2pqbt/PCFpTPGdzN8X4Th96GFV25gJe+QIlGvC5JF
UeWM3fnEKKfW5S/7XzGhuslX5Qdhh4aYNOiBPhsQH7AR3NExsBtpISk5/rJJsDAJovHCUvLFzKk8
WifW5O/TrRv69n17r7/uL47jrIpovKMTBpT5r+1ANo29m4RhzPqOYLxx7Pq/YbobCL8Sx2PPIYPe
DhwhE239Vwzln1GvtRHQE/hLThr5XM3Bd/i+n8f/dadOWHsiV8xDgXOObiMedgU4fwju24WtraN5
Vd224Sg0iREw+ImVP2xf0fZEzsulK/oCKh2Th8dABp+ppIhndBs85ZlSRyWkEDxeAL+fos60bABz
qvJCEkhmbC3+pBQqLQjCiejpa9SzVqnTtvhqLMOYo/BFBuTwwJ8hnrZT0T1uGucTtlr1rZHXNBwV
ZTFcwUJjFw9lafFLE2ri/6+7o2C635dViNzW2/MDUzze/KdsZfm8ikZDnUjMX3Tew3lJ2LZOjMl7
7wPIFvZX+CBM1iMJXyWX9pifdQGiYsZ1JKc2Bi1Zyu/1AJnO33v8qCOd8J8LcLuZavEQyrZw7z/7
GXRmWpmRn88OMtzYaohxka2nmp3K4Q951A8oHPZN3/ikGd75oknz15o8uqLP5YCwmZZKuE7a8Rd+
wfqa5K5R4u2TG4WD/Lpp0OMFoA8ehxUioqNhssCxLBhnNk98Bsygbboz8yB0pHNOsk5l118YWAZb
RR2Mx/SAKwPMQ5xzyI/J5PNq5414Q+Kfd+opn1sgJGuaxa+OTMqpVBvinNImzpUFe5UbkfQUacw6
Jp96cqtU5OCpqVWqutPIJLhByOtHP8OW3D/0otqB8AlLI5Z/Dm6kQdIX1ggsxPPsums6hwVZaEw0
3qf/zK9pSWnfs35GUUqFAYF9EXahIqhEdJMdtf80tpajaprR87DjOOgQdbKVrRC5z9ANWMF/sICW
aTii3FqOaGx3FvmnplWk0Cql/v6s7/+zIjMz8HI8KkmChr3Pnm7nSJADrP7WbkZAGLwtBbe3HRHL
SXuIc5QZIa4Jq9qzrQK7e6q5OfEer1aa15erG1yARqKQIzflIKB/zgK0m35gfi3fZ3cGjlhGzD+s
GLQ++vWjZGBKwtNiWTJv6nTTRscn/OrL7KitrH5ropGz0ord3Rg3l7NQj+z1vVW26Oslo2vHULlN
NGSsnb4qeYqAKduQQT8+3gxU0JsJey8kxh2raKVZOC9kYL5JVGYp4iAmQEEGPbrJI13h55lqwqjV
4Dmc0brhvf92X2cdEwF7LhA4B6p3AWsDTJwmuowGDVjV7VGrYLCPO8RilHqrMejLeisg7S4Wlwgo
aYTyYmqcAG8L1lugO5XMZXG11ahEdKAzB8e2NKqcU9X/kToZKJhqADCJS6mGTD7BzF1666ZdqG+t
YJn7qkINg3WSCwBW8A/fHTJWew5BkGxlG8eoUx3GWn19u/cUcMs6DZpjyaMAA1raXW2p6U0lyqY4
Bw/8Z4SS9CVUGylLFQyerVt8qdyTyxJOy/zll2Z0iZbXzpXdjlBynkhhajeKbSTLPKW3MB1FPikk
QSoKD8gO4BrrCXF49AcldpBlrOIHl/4cHqeVLoDhZPQqB2VgwSIdM2i0eDMy3HLemk/8LcHrHlun
HQicGfs6Cwo1aWjlPtbuepHl1BEwZGJCVnLQfwL7CEk7bPHKQmKiUoob88tNYLBLRL5SAcdLk8su
jt7B6NXEtW7w9ANScAOpM7uFLq4uOlZ9tmy2aGG1pniWsGO5XfPWShAfNSK3MuNh/6zn/TrIsY8Z
kUJJzp5tKl4FACsmMi9QTrbmnJUYqlyrHFAqMwcp7QP5nl22+pvPjEGOM6Krms0fdZmCMJNzeyLw
9hRmV6e7/GPT2UtL6ZIsjBslkhloTXx6//aklJvv0mCVSIwGhE2+EjzLBgVU7XtQroNvSPeXKJj4
KoOaxjmsEWcniYXS4zLmOwtZgBOIo70T/QbMW9ajrlfvuTiHYsrw0Ao5/gV5GV9fy5hSZEzw561P
7nqGsNN8swYff78dc/GhiLZz254Ix2aMcYtxZ571r9h6bF8JQ7r3f4jeiw0QaaGkUHH3e7m1RAfu
zI3BtF9BuolL9/AB1tNTfeRdqL/J3eOlEbkhRAbkgDNiumfaoaLx9yPtstjwpWNSQdfMpytMI29v
wCzT/c2cK5EkZEc+UD8oUYzcgu9hR226SUIMk25cJ49UGfiJlESOD5mV/TzG90D4WF3YLqR9Pe/t
ZJsEt1foIX4kXv83EhbELargc3ZTr7MbAvJdYcHqgDDLwYLZcrEE4XVNKELM2Nb4WjpAkqq68Ia7
f2il/r8ZVrPtaQq+D6WkLMFR9GoDoXqED77Dkfj2jt86Pdvk0pWGmYf1XIyOuEQz8dzYdSMQ+qxs
Ta+YL7XcNR8nCz7Jub9R8tr9cpRAZ4jk5/M+NvnvaWFbmMsOzEyFHfSP1KSejqg7NElXTS80Crko
ygfxP0Tez22jaWapUpyKOiqWi5yOeIFpnc0AJIjCTsCk8b2fXWsYcTy7+G5XA9CGg/k1jJhEdAIQ
tDGwE/hmdOdLGwpzTVMARxL5td1+bk+CUi0TIc6a199rrcMvm7KjXBBFYDCwzncWtStmSRe89x56
lXd7vRBv+N/eseEFpIsRSqiKpQhCa6za9SjkS2+5gZ8aauk/v0KIUxGlwhLJjWwkDNGRbotPQ32+
rrWxR0w1Fg/qUI1vKkOJM50lOepap6mso9sNsChSSPuPtzDpsQ8ZBdjidFU2p30fLbkwvwE38Dmu
bdNyTfSBia6Ex+899bsz1a5egGbMKLJn8KlQQw5xh/Ml9Awa073SAwdziI4lwpXRkO0VGy1pd4HZ
+VqEYf3jEYNXQbBauAzbZz5HNPtCkYosSq9BEUwjq2U/ZrYHJFQGBtzuYj7eYVpZJUzFx04PRDQF
OPwGB4ENCMIl8ohsmmg9qizu74y8ZyFrGUjbPSLRoF6y66iJCdYECsKwNsaMlYBhs7Fmv4dFu0pI
Ke5UWxiP0QIoD4ooz1iI8zmzeoEXSzbcI08w9aQatZAC7RuLMNL9Y0BGc3O4YhFfSJrvyvA8WBFo
ZoGcTH/T/swdpDOUj7tNiOOYFvdEhtGJIHX4MP+y8vSTh7YCXOCWtpeHMIAgFdP7EciQoTSD0MQ5
7sjkadrYuSMSN2mLeMvSWiutdUuv1u3KEuu9T1CEmcngXk+scwBzfkTPmw3FGeh24Z/qphj71cRw
PR+69DrMM/s2HoEUKvSCnVYRTdpC58ANFzIyHipCag13sKevMn3Qviboakgu7ck0a3p0REQqymqq
sE5DPbbbNyJ9T+wxSDcvIJtSkE8FL7vX88MCnBANXLZN9p9qVMpY3RvyzP3dm4MKw2+VK91PxXhE
jrcg8f4CSbrHbPrBrlBMcDONhMR4MCJM33huqtLqayHeJ0F9L7wbVeDhO4A3OA5lAhiMxX43WfZA
DHehrK35tShWWFl1fJgO+mUhsNZ6Hz/skw3Y6TM0L2dNzWj8PRlSI7ZICFKLCDzgyI57rMcWotj4
MdsK991FWv2B3VQQaxswozSUG6PXuDAndP5xkVaTBb0CyeR0oVhY241wBAVOs04aKe4X+Fsn28I+
6gilwmSkzQbD7/Hvqhrt5YaIFCIWbsdpMMYFcZwBD3AYJhHM8ZyiNbFhiClAEum2gg+8Tp0o6QsF
ZACuKeVphGYp+oqdRtDinZKRlKVoldje3XReGK3bFFUMSA5DUmdV6G5GFBoE5WyTx9ngAHtI+WFI
g+PeKTJ/RG7cKyBv53gvsBXPhTxUwkq8cHtreZvx5I4HW6vcFkPKNkAsYTwPGogKHG9Gz2pELgK2
g/j5vUHBEKqrECPwCGyQnEX/p0t5n85cg9xF/146UZzTMg2tGi8UWFr+erdLzMA4chv+UB2vQF4c
fs4Bd0roADVeenOieeNM2Hr8gYXea7/jk5G6v7PJsZpwvMvIFDgONxY1PbyyU7WxutSEeKLFEFTE
E+rUQKo0a5UfUlHwBhqX8IpUlNpX850o4gC3fetwuYTDrxmpgM5HXdCOVKp8xha2q8t9pA05Vv8z
aGldDZtVvVQi3wMM4UCBZjujh4hizbO1tF9qVk5hoe6dbA2q8JgqbNvA+k79wqfpRov52GN/eWto
ZYI0Nu75o5KAf5mWr3FDu/HuIvc2rczy5480DAF2P2BbXcNyGjpso7RT7xACd+uK3XNoai33lwWF
ZB6adSI7tAb8QDSBauotVx3Eauv6SjtWJFz3b4l59jsntYm2Qv/zjsxJ0emTXw/h7gHKkBnacTSm
7B71188FGidkxdTMWJVlpgvlJmcL6D/f+gLxg6FSoydVvnX4tpMjNKAy7GrpW2zQq3axGYIUxrOG
YajvzJv1BkcwSEr8qiq2F5BYm1ZEagRke/FiwFnpDsVw6fI0kDVF086Clxh4kV3iV/d/MlmAfBoN
C5HnWNpXngwqkphk9Qyylx3DLLGGm2H7oCZ63W5jMq3Ga9OScDgCPwmIPYKz376P+CyGY0bsYagI
CIDc58lw9ZsXk18mbvhNLSiN3u29qwYrN58l6surBbDQNcGqg3cqcVF3nprFSFI/JaVSasDDnFhJ
mG6mtJxTlzK6AsaUBTDund1uQ166qy8OtW/Qy+FwuWPiMQP3F005nT2zt5L/XYodo9I0H89SOBNy
NrJicXaBKQINZN5ro/TIZbIYWHhCBIJ79h9YIO5yjiLL+N5Bl0Ii/uGt8JXZyNC1G0QMygXX4Ded
rHxsV4wWhVnK3zeuYoRalzVOx243HGtDS9o9/m4U/6oj8Ld4TEg/NHOO6ub34Axmr2BXVLABwtR4
u164GWH5rpC64PtlHsn9FKiN/fa+fomlYicj2i9FvPU9bVSyMoN0qYrYeH9LuCXoHjNT6nM4oV5g
L78MihtCBRbhsLZqNQoAFJFE80ZxA5shiFaNJ+K+iZQmzuVvO9WWsDcQHiSm6hIrMvln5Q26e91i
Zk2E7tikADBOv5d3j6M3qTNdhc8YFyDpUi07ou/MG3NRVBqb6YZLwVtsfZHJsPAKbAbGnsCDpTnc
Qr0tywEyV+UwYnLsdMsX0q5e+g3j4Pl2OOo1tHWXzlUGvfy5aH4buGGoLMdRyYoiR2iOf6KqSDbb
RfQr6bcp+3tTDqXMemdvbhAq0sXvwKgK2RiNzEL6Z9XrjLxnSI8ocGMAU+f9zDaySq9MaSjNOBBQ
388D4ue/f+nRVORVtrUS0aIeY0wBtHgiw4bnMGBb/X9WLCg56XQxIDBqPvPeQd70hebBE2jnVmyp
kLDuCKE7//VQRj1bvv1ylAGZxlTj85hfZNp0ykWewv51o8kgY94/VGDUzfuFo1Yi97Q9zr3y26dH
DjhBStviE3j+IpoVbi+Y0d/gSVZR9BAfqto7tewUJXy3Nm1xHTT+BK0oiJsrAFSse4EYRskkEG2V
tOLCys3wrFAXr5zY2RbI6F2cavJZy94T6fuM5DHyCpoj1MPlc64Gx+WvfukOHIFJOnz4o/gZaN7i
d2rtv58fogCdYBZaX/7jXcObX+iZ/4vzYHdfRBVNpAgAYzHJk7E3pbY5ERzR0eRCTUksmlfQ8NiF
EO7ZBrvRQUehFOOPqRm8korzzyWJp9/5HFpbz7+FUHo0msDOqNhM9ZKK5LK3DvGxqm/SyJ5qmw5+
9hNKQ8qCnbN2q8SHEWnhn+n1DWmfTx5Ncru4QUPrPvGB5STdwZz/leIfHO+KkkbnZW5g9P+YqElV
sfcxfgKPF7XIRU5iVdjiE8ZubKZdynUQpl8505zFrls8zDJE4fylf9yDyEeS/kXcACvQBqguaD7Y
wa+OwV0pzK+R4w7bLHSci+31ejnoGIhtbbDSvmjLB7x9oJDdl+6UwIGyGb/v8WvYtZh3TQ61ucK3
pxhSvDZyUQ6zp9O2fMLJmIpA1kan/cPTbul5/uPtPulsq9yTZ6t36YW2RJxmjaae34LDmDHNC2A0
+YFqrZALg9ycNwyiyopcr4N9X4BRXm7JeFHZ2Jalje9bXS53T4eSOnfLpxpyKlz1pasQHnWX/51u
Z5I1ahGs3EbfwC2wBU5qYTNIO9TArSMJg32/IvPttDDr7tYvB/hkosOq2sK+tyCmDfdSdvh/0+g9
OVLIJgfTa7X2R0PPZvPD3kEw98n2KtgYPZJoc+B+gEKWSgOMJral53Emd63LATay4sNyp83WHBdz
t1mdt6LjQPZDGoE5kv4KfXIWM6rl5zHg4pmZtlih8No9YyKswln79iO2/ystkVbsCLR29233+S82
EfSA2duyVPhu9Vzv4qCiZ7eHx3oawVs/ceIqYls4zE3CUqn/Z4gHtU7LsE66MOaoJAJr2ZzvYCad
FytuP9tPeFwcJc71o+rMhS2QJSalnTMHUAB3X4VMF3Piyk1G8EbKkTEUvFOICNuXxMJgPQaIpKif
GpKvjmcAWz1TWT96YlMIjmpzDkmRd/e8O0WoaFkdlbxV6nyu7pOgNzOWWUFB9RD9K13n12Ne+R9U
zsA0cf5/94UH/zaUFyBh6fJsbAPp9QoKQnFDvhIOk5M4lu9ybKwzxouheW20tgQYSfVb0+xAeK/e
H6/W/AwSbsF5w664DBAMyiRIgsSUJc839F4VnwP6HkcjfwoOigr77k4pBw6hrYrdgElVwfRowR6n
gxbMbITQtHE7RBXchdoRABD1IpYH2c9x1aevkNmMULyOak2kYoI20id0iyVxcTS/nOHQ8uWznkxb
k2SVFzw0TrXynxyqtd+lRMLnWOMu8Cu/n6MOdpMk9TbHTGdsxBooigxIzcbnW5QfjmAPRXVv2bVX
KfOFDm1/wRTrp2CqqquvaLbMmtLvZxtPn4Zoa4l5mhCfntxCF0/ctcplxjsWRpu9dh7FuhKlMdEr
0k40XwERtiMJPghjw3nnxVXQqb5vItCznEqpD2lwqhk8r6GqE3GfwJyTliDzXPqsIBvGElMD7TpR
Zrv0HKJZKOBq3bZDc7KZafi+QXi7EGDe0fEn1DHhRzggkvVJDw7K/hX8ZBxBCbdpHO/tPRlBhd3q
x8hcsnlzIs/mQ+Og9HXYckNpDvk6YrtqxTEDi1IQDXxBxeGFWaoU1Ruf23quMAaZ0g1FZVB7/j5R
GUCJWNzzl0nD1MsxL4K4kiJT03ObYdT+fnswO5TmMp7VC1L4qpIBbX8cK8FHWde7GkLjnKLTaafH
N6l2OOidmIeee1nDAvVU5lPEUBZGku0tYTSpx3pds2yuiNEIxBumLoqKi/hA3OzKmitgPAQix5iC
INBXWLkU9oz/sBY+HC5qAbA4TkkAMvaDJbhVq3Tr/K0HopvgREDjvuAMTvfLWLRjUYyZ1lPBejCb
BlIXbgMzQjunwviGh8ywFKAMKR0PHLsppkmJyjSomuyzFGqWhJ9b1XgqtCYG9s/M96/tA9FeNoS8
yiBJnu3yh9ixJaEhFMjxEC2zqduHUpvHciH3uFMUwRYR6vgTlIvLf7GC9i5MFijDGbZubu53Ze6O
uTY6yyQf/oZ69KVzUxL88fb0BkLtksxbs0sGUpBuWIW1MzGmtDzRGPbBzJZ7/aOtvK9eg9SzwxWn
1Yb3e0MGL0OO3kApM77SCf3s43SzS5iIkcjC7F/ImsXDO7IE9LPN7PdC1aPQKURDOWba1A/3hKYX
g00tqGaNS4behTVONFQR90s8/sGFPPenYANXlDCLP+rYx8k/Ru3KUP5JSPIPHkJj6Wz1yVOjtm9E
QJ+g6eUWwvXfNpMsVMm73/p3EnQFa36qMCgPojEUyNmDv2sCn9qMi0q2KifO/5jeaAC177wig/s1
+PEog3ax2GcmKUMKfyVgbDWYOcC9AwXTNl6Cq8nGOchKB58FRfNqwQPaWT7VgRz9g5e3UlA6DAE6
5Qrupv1F5niIRiUDF6y4L8w7C85ey6qeaY78MV+olN9c3AJFD8/7nPYjcfHZClnaUVL11MzGPeuV
74Q/VfAm0qyCDSIY1VvIfzVNx8yHZ0U7VosHTUwgAgdqdHoFcnXFVyWxIMLSzd0dTqfmG/ykPUi/
vjKx2Wg6+z4GflsiIyg3XgK8NFyQsCilYAS5umkGwUa574+N+PlstE6rSUCarWTcQ3Z1/ghDtPrf
C0vzM4m2eo+LKvvCV4mgiOWIBX5G1TFuPP4gBoaZiao/if7XOBZNfFjWjETELF0l0hMmEVVXPZrz
fSrtSPAYzmAPCxjGtC1hmGjkYpFiv16kUe5wiIxyuyjMFk1T0tQ9HIqWYkf/rmxRenUQm737Yo/z
PKZE1WFcgwq31AjVCiZ+LzuxLaF4V9P2uBjesHDR6hiwysuNqAPS5f10T3iIuu9LrBbLngBngXlf
upqL8ZIBF7UttgJOCVhDnDSvnGAu89ZU5+opGdU0c1TiRAPsHxMCVW33hg7xWJLZEiHkSmKPhu2o
liZbbKyOM3StB+1XJkdK8htsWTD4tlHDCioX2NNZmUAV1FbAhq5RBbe9mDcAq4/abFk8yivmFdX8
d8Xry96nViRc2kdzvvpAS+uILZWK7VyqChjx/i1E0n2DwVsSR+77HKxjvNZiJU7+006d1oU80C9p
clNeXl39U8KAtGyuhtoK4O/ihleTOOsR97iKwZ3F/uoSHDJeSUWuOw0SWTiWilrBhRXpPQDhud90
QbXxDKcSJimWczT0EkfZcNRvLcGUhllgxWQsKSQgx/FD1JqnkNoSR6WRL9q0UVHOArUy0eiUmg/x
/tHrqc6H3kQVrzaXnBMoVFRlqxmWT01X0d+e0fSxwnBp60ebFf/5vqDtOFyLAeImheG88Euose7U
n90GIG+T+DQxcmM9X3PNRqb16MT3M2nOjo/lOoWJqFzvfjc02IY3tSOMyPi+wQJBmeT6JGiOND6w
fF4jsWFLwhzlKAYBFNeXnarvnNvqLGoqhLXYHxE3uqk2RzQKuQ+JauN33YdMQLzuPZQlgWU+V4JB
hP0EMnyhdDe/cqI0IRzRWm+q7PKa1JZv8mZJW6hrbr4XV/P3V7Ses+nwME4r582MVFBvjArcFoXX
so5pejgF4PN6Lq4TAxqBzbTu6U7AbjUYfIs464Xkj3zR2SAlMaX/AiK1eTRWAUWtv7dwTPQW9LVh
1ZPcUJmxjXOMEsGnhyKkJ8rJdMWz4qGkTLmIUD37dHcGlp7mqHZWkakP87DRZ493yb2JLkx2A+Ur
slM0bFoHtbQANfYqKbbrPZygWPDMRgFQTIVWOfAr5jFmLHXJmdMjtPQCBRJU005UxtAt2a3UsPBo
IRd4TuCzPyG8jC93GGe+CR5sAaQoGLnDIiJI6jln1+KRD38m6KLGu5wAKT4vap0wdAfg6SWtag4y
CItYJk6BGaa5KxDmwMFhCafbLnnepw9Hk7KuIVnm4oNaMPATgqEMsUIyMJxrWl4SdyZWy2gVcE5d
KTgOAbO786D6b2ASybeHIRFkjtWA8+/LAudp4TxK8CTjYo4xnGoMcMPyu0IEz7fJ/RcsszI5FlEm
/RtCr3gYVLEDLnDH7sitI0Jkg9bGDwBa312SgCJci6f4UAKzmpMNcLLXIVfFnUA2aoh9ary5cwlA
Ajx5r+q9/CsUs+uKxopqTKjQ8mg40w4AB0aIXnBASoOkiDArmXLNHGDmanD9rIV1BCqV/9MFUzbj
uNc8aojUU4QMw4f1EtCPNzyTtzQ5ks+w2K48kqTnkM5Gvqgm2m/hpI7IW2RlOW9otBrEVYlu2lj0
zh3bjJxS89uF3WQSBQEeyge2DMelMkjjZQtUFVY4k5ROXtBpbzwm+Gde2OaSfhcsqd1p6d/YZcUl
HU3Li5Vf+2endneQM4zrTBO2DPg4QkOTMFX7+Cp4Y7HQ92G45WnHYbj7LyoUUToRwkhQqNtMm3O9
Zf/nWdal5TnHbmD4SnDOngtqgwIgEpw/MpF1T5K6OPiwVm+q5HQOKUUoZPo7Y9GPx64JgSlFhnZX
5d6Fo38n5UlFOaZBWln2ITledzrQJP9k/xcWTmT0jkfz8Eb06BJAeej4tbC32lZ8k33ofkZppJQS
S+Mo74TUZ5Rcvad0uxcxJf9yJzM66OTE3Jf44DSRnpj99E9N4FyZhkNZs7aAWWpnIOT1bbc/NFZJ
mjvNqVU02rKu2Lz1Q30MUSqL7MlDp2x7mLEQQvP1s6aphSMrjujqC8vzG/NAdxuXzjCnT8Fageo+
WzeS4bBqpoW/oa/9VZLnNndwOECi5Bb8yHCZieJAhGtVD0LApDYuLP5lD1tGqY5l378jKpmmK+hT
6JMiihEQYPwZV3w4dN+SVik/YJ7Tf9LYZTedEwTStE2x4++ureJEfN+FtJFC8u+dGkYSm2X1SlNz
qZWG9gXICO3eqcIcIbFdxJ7zHpXNogWCWuNVuwA1r7vIQB7JvIGasgUCKWHLGuM7taZtoZVFgu1B
Cy7QKvU5rxJFyP68Yy2J2aXW3L7pO0oJWgol6pCStN1gW7UZbiDwHhWsVEaVtYQvNzvigLX2cz3T
AyxlgmzZa+URZBvnrC9aXBQeUlTGT4jbQ8ozkdOr23bwbQh1N0H3lkQFM+psfYZZEUMyQ+vMDKW0
scsJxiI/efRRSEc3h3Ts04LlKg8JLd9AugBmBl2naGCKTfi0ts0cEUDU1STgVAWDmmCHfUjCEGjn
cdMzUc+w2dgSXMlqhel9J98+Umz87F1r4kiXBF1fc1wFNID2UKj3KPrevKbp3omPuRAeRlY81fWA
RbHQknE7rVBRQUGYA6oLmURbB/90YaVZaJAB/6EAfRA3JZuzyTMldnCo6q6b+sh5YeIO4ER6bquN
1w/UDGvYwvw53t0rnmKgdfk2u3hfRDusvqVJxYxuA+4t7sLI387IbadNJqflwtyXNNlUQMFKBQB7
goWguEZF8jWOF2FQpoL0Yh5EzIV60MVCX3DRrsvWgHH/7LhH5PEX7LPrfciLdqxhFnSkRJuLTel+
U6P0D3Aysg7pxKnmN4y0URK1tlxOATTxY63ZP0imykQsdWA8ztL50/eyO0ah45u6dCJcpUtCmgbG
srQ7RtQK6vMTTede663tFJ/XEqVUieKNk1i8NSJawT9yVALi6TBqjyP2SCvd2DVhx/AyDX36tONQ
E1BoUvLjdtOAxXFmG7tQeOta6TbPAWm+nHX+C/NYEGu6Z1dCukT6chzExKTFrp6FGmSV2k9cQENO
96Drmx32TfmIQ408Knz7OhzGOLwXB8ZxLN8PBcZbt/LJqhi9NbpcmnryKXCgOuj3b3YlCsdiwF3o
6FGscDWFT9JVxHUIe8s/5vB6j6zH5Dnm08B5N1/F4rzi2Hep7p2+687E2jYX+/RTwHI9C0un1u7N
hNpfI8o3MeqIeawwSHPaapW9xrix4UahaHrwJjfXHoTPtxQDvoaqER9++zdFrWI2EOyoS4g3f6dx
6XCAFnyxEfM0WJReyxwk7SyA0/zNbrPtxdl+cKPI17VQw4IxCnQu829TIcRXhptX1hQuKPoyCZD3
kVQJQLKQAebGPmZCi0zyN1P3LjsKrMMnfmqUT8zGJbkYJ0hUwIpvQz5OPGc+LYB8sSMpc5ksrSwD
l/8w6k7/0DA5gdzJ1Av+Et+ZmYn5alMfurFubx+SdPMkbrdHGROpMTieA0+/pAVrQj/OxSzkX5QS
jzi8XhbyMgTi4rJrDMNvwqJFN9FuQCIU3fvMoWyJNENhOBlYigJHRBZh24RGMaBNtt8H+gU9bo5S
0OqX2sVsQVlEHsoJ2lwmrDizm09h9g84w8BdeP5OfHE/6WtJZEBJ5WoEw/j5wNVzbsr2l6rahcTD
s+cy2gI6wkL72weMhWSJb4Jw4+hh71j2vG+z2KAu9WH8XCcqZ0tShNJt+ToPc5FXAPSAAXE8Po38
O7qWZeQ/USjUmWX1gDrMgHdWy747SpHc6AAx4gYZ+GrVQwU/ctoWNJRnQ3VIUkzhWF6UuygYbinZ
ftVsAjwGjPlTYLuHKhWvnEN5RqnTSLbADTjg70wRUXSt6RORGh6pA4DabKW6zYmIqy3BkWopxHR0
2+IJLHwG0iqtU0AvHSjmBNr9o1P8XUVCYFUW5Eka7K+DW7RBh6cr7DWJYW5CQy9A6QI2+YGqK5FZ
gLwNjK4cDAcekKB23kJrc2RwS3w45Prk8QCA9Pitd46zc+5ANRof0jjn5czEz1wlkglQtLy1rLlz
RFWInpQaRj0iJ9E/HlyvunoknxYapCn4D1sdDkSF/9u9hB3IHKmxynIMkTyjjftAqvKU0Lb893FD
9J9oIezEbdkcfd17TLSx97AOKKxv+L3iCfceVmnDjZjursFF7A+QpcFZZkIe+xjaHTsryEbGEwqm
YO6TpFlQOErcsfsrKqvSuh4ID9O/dWHkzO6JTFcV3eqXXqufEXgmdiVtOnChDqiWGd+jM1XpC0rl
xNzzfQnb5huFQLji2iwgMmhhKSufeQWR4VP3aGynGtcI+XzGV/tbFw7ILiTHfnGcSYfDstNrGd5z
wUg5cTuVSn9t18bwZQUx2v+qIJWHPseaKS83+QhLofe84AsilVewXNVW6UaH1vb2pU7wEWxzaw60
83IG7ZE8R8UCELwFdYTxHBU75e0BGQwkEY3xeJeUns9N71Y8nTJ0htAnfVMGhx9FOwOEHbyBTDwm
iKcTiAKlF0ZriJIFaqFOUEtvQIIFvwCtZQmMScaJmMwVkdC0jL+uFIQ0R8nnLL6Ud0CqE3dKr4Do
GvuAFgz5hgTX1DPx0McQWX5+rGHUcc4jw5OMaiHNNjy7FPN7X/LHQQm4YCftWyqcXGEi1kLBO4ia
GUPcyNN7wDzYAkJMX1DIB/rgnHbWP+5X447WnhhxRoNZH2HhVHJfeQrLdp110UjnSpOaXknQyoQc
7xkGMvySVuSGM6Uq9m+T//5A0fykURdtW/GsVNgQ/vf9pjMNmCE8e6zwAG31RciFyZ1QaX5F2gue
K4UgecbD/WsEcTBVzM4TkcHG0Hl8SeuIiBijQrfi7cj7qvbXI139aywGZBl+Umt87JTymfBbDqFY
jjg90Z4as6esBVn2BkPfsxoAtfJFqKqt/kO0/dkEim/ps0XZYn5IAI0rrcv6uHctpTRPjPie0SON
pn76nXLnW1RMOPKXsqFcwwPElnrRhQ0/wT//AHh9BYj2l8UNZWA+6wjedwxserQ9Q6/YH5HlhY12
Eb+ryP+7kMBidl33oEzsxusg9uxz9tje7eAWM3RTVwaDJkaQmtRmLBtIeBpOwRIe87QweT0+KdZp
wfdQe3aabMTVTMUlU5gLilN5etw+BGZKTOQKaLEOkIaJKFzk8PL8ecn2huN2DtBYpMzdNopgbPnW
6tV/Jk1FHXGCNi6UIKHqaRsf7dSgJhEy73x6gagm1PTB1MGPMZRgOIJreIHkdF5S7C7ONU7dAuVJ
KS9q9n39h7POTjfoczUOuMAne4jg+ZJ8OHXHK+AjW2fAik9zFcRFRkw+Gbi3dAED5fG8EFYFYjNx
Em7Q86FUknYuwITrg/MB4eWU9/EzpRJbM/WVY821D3ZEsz9KuWooKSwo6Kj69mCZhCHTPtrt0s4S
3GyWPPRSlSH/vGAk/qCS97PmmUsnNuQD26YJfSJB309jJTj64TYXvZ/4EMAUN+32EqX1HXg4Gz1R
ESyOTTDJGlp6awqOkilh7WeuZKSlwQa5T5iCbi/aMIhfUGtmf982eKv4u+PgFnq5GUasNZBBqCy2
mCkpYo1kkiVCnI8Ce6/U6+Di2v22moc+sNNafgzZexEiQ7o/CUuJop9wwAhSDngxqNJRAxgPv43J
KCBczfkVyZYgmajcJGKvSYrKX6+puxj9CCvHEjIW1D1BhhBZ+OUYEo+RyQZ4DaPUO9ePYNZ7/SNl
nYmUnxsZA2ooJoHaUdc4HJWtfrj5V4p5809B0pP0H4H1qefqx2Ja3ZIYryLjWAo05x1xR+/I3v4B
cmlVF8nr65EMiBN8Lh8XoJFfZKy+rAwjNs2DMWazIpnVLkw9gaHf/FCW8KQq//CQkQS6P4111s0U
oXYoH6DtszqGKQvS+u+64V6pTXTnfbl4yy5BQ/Xyi/JZNX1qoTnndjng55oNIkZv5WL9T7UtQEHB
Gyu0bxzBdfjf8zt5lxy8DLF27hYLOJw1ieJgOjb1XwSezpzNE83OgTJ4FUYkL4eQQFDsNsVmUJwW
ZalzzL5+HHe71QfQpsISYopcp1IMtnD2zYoqUv8zTF1W5dE0j9aQjJB9iKeXb5OVnaUsaQiBw2r6
GLX0KUO/yRGfDG3ipvngOx7mNIbgeA4SE1BD8fmq1/aXE9aE7UBwgHBQgFtO3LUC6eTUto2Sykyu
IaebGmTLfDY2aecVZ1CZEemhqmRLLXQHV2yNvtHXhvnQqDMvqrYzMIN3EXSj5YtWDLv9v4vn/NCh
GqNoq+Wb4m9kC6Pi4D2APs6Zh6M0fNMhHsiULzapQPUD2qq4xSPCTgRp6SwxE7acqIu/nszL+3dk
nHkxMRb4ecgRiakc/TFcLIndGb+huGL9AObYxEmebjhZQZfeX07W+I0zT3EWIRK58pZNLr98Aa3y
UWVbByhROnQGyqHfo9vqA/weJflFrCaAZ66erwW2wkFr9qkGM85z0qSb1HLVX5BIJvKpd+2K9v+C
rNYV/AO/z8iX/CDvdWT7m9AphsHHjKPKmtDWA/VpUdymO69z4xkY2PHy5zoEfoGJwHfwuAX04TmO
TzaF/8xJJoe0HjpWcbiaxM2opN8iiMaaaSUJq4WZWSGy5iK1vc8MRIJFsVsoUqkEf6aGXk2EFJMB
dDuKUqaHlcn/Ce8pj/JEN95jsNIYwH4o7g5kZ+hcKLuwuxj1FZ7niU+CPEOo21lm4meRD7k39NkR
oFRiH/aFnG9zErs7novJLrhYduocSUS4oXVpptdbgA9AHZfVotOXdSmYUndYt3Y1qcqRDIGCLAfi
/aEGJnUesfQLURNyZXXjJafQN0+rockj1imrMg4IPWDxH9T3OW9pPrGMAbFLboOnFw0cFMqkeHJk
MZs7z22n4J0CXMq6vYcM73HQcdCwmvcge5vTFNOS76x0Ih0J8RL5+op/iyOg26+28CIoCv2CNHN+
lucpkA9Q1X+SXNGMr/Kon3HTJiVNhfSr1nko4wKRWXy1jsX3HX5E65NuJN4UTzWDGbqa2u0eXrad
HMmZnVvvxT27FVIm0j4OBGrquViuZJwPhQbxD/uZWmnZmInaCBENeUhIjYfSDB+GKeruRCCTaow9
Nv7/UVSvQivBRjmB6D0KH3b17rNmBPIqQSJntHOwrloYKZnaJljOXyQdNlKlZRSUTZ+5vqMH2bOK
tS6GXnt8CX/KFWNdQAr+uGfHJw9AeOkhfEDP7k7DuOjvI2jztuxKWBhorV5Xi6PLEYL8Ui8nEmSJ
5MAQ9sZCnqAaaw5SE3scjWLwI7OJNHcUw9IhgjE2w6GjW4woCRP0FT+TG5pIx5AjGAaniSHgB14O
EEhZlL4aibqxL5P9P419sQW2Sc7pCUVWtaQ+Oo8PVXTcnnmB92BO5Z+LP9+HUF+u85UL+QHkl68X
+3dSWcVoHfVawo2tLDIDtCljZ/3IZzh5I/OssTQQZlEcaue73SnxpPY7SKUCcjL3YpuRqM0KPG0M
HrzdNHlbp1GDZyXpTAeh9MxKWgBjcGWAYOz9gd2pZkKH2lzSuB4caXyLehTZeqS3qPjloCXUMIRF
Xl0wsY7iGr0AbQ9SO6MC+PG0JsYGyKtgzbFktCCXVorMVkLRWXCqavRkbS70Bzwu7qNSoK4G/X6q
iU3B9UrGPf219s4yY2A+Yguiuv88C0vPeB+tlEn8XgSw6OGpu+zdbg8t+D6VmbYBawp6/Y46M0+5
m236447k/K18MVrI4wdgudz/bTNiK8ndDwbj/YyC4YGnx9b7PmuM8s/nmXJ6m0DbhRMUEh5zqwg+
zJk0SixNajyojLeIv1t5QMRz9f9Fw1vLC8ytYqdzKYgz7B6KkJyCShJiuXoPQp/p9nNaUmczsliU
TacyP216L8RvJGXony8egPY6Iu39NSSBZlThSlrDD/1W5sWEFozF/1Pq2OobfLsUn6JE65raN4If
znxMkGtiRcDHEMAePoTIHJaKRW0YD2cB+YNZX63yK9e2cAhfhOT+2SuBClXEO9883GKc1Hv59Nsx
dmZErqP9dKLv46kG8q1y83ms8zzzOSM/uBRWIt3yc9S/O8whMaJWODpeRypTp469crpRMtVGPaOu
fisDjQxjSn21jkt4F48q6ymeic9HyJ3hgoZKZi0nfH5iixsi5foOpK7xMkRYZJc3P/6DM71MWIfl
grCwup8zmgKVg2OX00lFFcqmMu22jqLt1CQlPKJJ1IAgrIrkZwXL9o1i0KKbGaEjSaI22Qocj6ds
4Xt1QTr+9EQFgZhomhogtoXkZ76Rx+oVIgYfMh1SZ2TQ2whryhis22E1+7m0GJIvCnbHaA++SzAR
6b88eRzTP22U5nf95OWA+hj0JD2+to4IP+moakM/4CHRuUuOWDayArFny4uM9As/vNqqSk/s/J6F
+x8thUEdJj7yruNO60OEkcmqYZZGbrLudo129LCH0oE7ElX2+Ra60ZoqAdktr/+iMg9J+Qb1q5t+
3cId2qn7LyWxr1PYuJcoQ7PU3TxA8sNnqwRrNtrbrUD8g3fnAqHu30VOcZsCDVierJ5yIlaoo6m5
Q+gtpn8NShk5m/MAzLmkfRfBWu5X17sHGxq696PA3MBfFLsO/1RDdTAaI0JfJ/jB4YHnjZ79kSVj
0EHk9M5cBtuFnG1zCdSchDNfQo3aRe4hmTWqKtYsr+b1Hd3XPcbFPvdI5Wo3sQO0T1CRURfgsTI1
+XNZgbeHU8oOIrXcE7ICipnlV+hbrmh7n30H2TAc2FA/7/82IaiVrD63P+ihetLbMLVdQWtaR8Nc
r3TQliIC4Ofw1+Hu9U8p5GElog7w4N5Xa63CJdZtPuaO4dScykv2cRFdoncYKLi3Uv4U24TkT8aU
p4Smw6oocboZY/xuuKBOwUcL6IO0da5E65JQDm4PBBq4CGdz09jwFB0ML9rgprVQDQwUbYOg8on8
rlRqFaizVQQUoEaRiF2IILSByef2jsUSzLwvCLkGMqeK2vXWemsxcxuhbySaa2I6ltSyQmOp7ii1
U4DdsuWljYOdSBY0rm8HwFcx6ILS428huPUFRC1GvmXhvOB9YuTxrd6aHeB6P4QZSB7vDh7iTRaI
05050MYhiYYyP7k1DLGMxdLN4pIVPDZn07XZtgOtT4mz2IzX02pZMZWOCxeOB3dGLNxq/sQzX4xA
Jr8SEv3qjfzmSsUAlailX72QI6xF9xTmAwUAV28p/bYDJ19fiG/dyzrK4fd533bq/HVr4mmsr+JU
N40oHE2UACWVJMapCCOdg13WbZxkd4wHEGSrS6Xl0I9ddKB57TKRWZXnqe6SqIHQ4J8yppvjfsLY
13cKUiACW1wP8DmmI5cWNYQduvZXoxDGVEml9rOxYssfNhdcyo2r3s9/Kq7KSlkP86L+KDxLriJN
ajwxte4MOoFF0wEEH7Hr+ZWskPexq41UiL6AtugnP4G+liiI6dJ+70l1zfuSOO0ZMIYcQVlqKq3o
oMrOkO1YVK3XlSPEUxv3FFgoxs63q/rm+T/ArQH90SQ3XY6CWEt3aPlMdiIq/KxwpI0AtwyFSiPC
jJzsO9Vm4jv6WvbzOnd2/meYoTVi4S2ycy2ftMuiKju04WAw0/UvE/moHQt6wTZFalgP1+K+U8tH
J59+qFQR7J0BWL/IXI0ZzlO79NfdPTQZ1Pb83uN8nQHK41/oJB1UvVqHImRfA7CiZFpxsRliqUsj
3fC8TBQ84121O8qcJiIvgTkOIbbRO83BcH3ypAqtPkqHZbmuZz2zSbfVqbQNvYiloYm57HP81lGt
1ZS2I9aCLEIe1pI9rmUwtZjq86Lws1ihfTo6iYdQudfTxLe8mCHQYQlfW+4PUzMtii3EP0pcwcPe
gLtx+WZXMz8Do+HvxGB9eyyNYv2znQbDdZo6fQOLPJjH1pTzFSENYiLlfVCqVTYQbigJsdnItvP4
/HllJaLaMtxMVSyYD/Orihagf4/1G9fIfPn2A2KrKhh7xMFNeZgGnCT5vKc4Ts2HMuPmiYNDPiEg
J3K6cAz+A4WTpLneX4+umzb2USmKPnzQx37CWf353H+/AJ+uCcGat/DxIy3FcpT0TAvhaSg2e9Yf
02KtPTUQ477ZxcmFftreQPigUhyFYRRbW0spK1lDaI6GToI2NtwfR/OorzLUKXX0z9gMiuBPFu+d
9Tmu1fyHhZ2hEym8iyKYnVQoauE1nSQLQw6NOo2MhAZH/qWkBoUHXj2pVrU0RGM8CRkrOYyEHjwp
jsXGZjILOGm9CtGolnbDhznEmUHLiKkwB7tWTZ1eOLZT1rX3w6exyCsKDnquX6P8gFMvWFedn8tV
AJ+kdPTyCBBe9Z7vQBEMWKBPqzBScKP5SYj7sDT6NK/RtTyhVUv4wFMv+j9haFfuWhsDnId6y8Xr
NfC/Y2lzeHE9JGtgm8ifMI8FyCkie2+umsMvwNV4FTeW8mpYW6H3BaKORlsyuYF1wOKYtGcOraiB
IS6hRgcMF5nm3CclPQ9Fj/1+cOj5U0oJoT90PUzpIJUsTswjs5aKk/4IsbiRMtbRGKwvWyM+Xlnp
VEqvL+1pSKo5CwrJ2zahErkGkNACaPFDU+dW29Sbh7izlrM4vOCtzJ0KqELtlsUT8hbicoTREZPz
JmSboru/m7/mxISQ5Yy3a8jYCRTVBFyZuJN2ExdAUnmu1T4NcGOljoI/8/ZzMgAiH9khRXAPoa7S
b8sNGcPKK1W6cMzcCFOS0o80vDjomfu+XOLNEfbt18ktj8OuLrywXjD2kN+Yt+3MVHIw3aXUkAK5
xyONjSpNG3wyFnshZ7UIDlS8b7yoJyoBTxdIrQYEgpUHAZ4ey2KKVWJ0wmUQlKiDCiL+HVJIxJrI
7kl6bG8b/PBtkfqdlz6KPdMy7DuadgvEy2ozjEzQi8QdxEWwSGsgOFHfD9azkuUER5XL3SBtu/ch
jZOCfPBjy6DN+RM6q7IVd9CchQDdO32giWrM2hz7QXk7thFHeKLy4Hc10h8MhXy4yOOhTYZTgUcP
V6IdGb/JPNJseoQwPnJf1f9mi8TjCPH/IU5/kdEruXhyQ5xoWCa0orCIBtCVFeMCIivwjG+5i3O+
Hac4f1QpdeGehZeKPj9dG0iBi7x6rbSAbj0pdRaKrJJE4CasmPyf8OTRiKMk081kC+0p0/IgDiGE
P6b1YrXyeBdUiohA4GCGvxGxmt3j589/7BGCInf4mnzxUU9hpZSAWDuPgsORnQrIsMRI2YXKRGAO
5kKxEnZVhKNxr5Qob/kCRCKLBUyxYly7LY2jrQArydVmgsxigubsom8K8e6htFspDMAf7nlFhYg3
X34rV7BD/4eCB7vsqWCVAKuQom7g+LgtBUqtDj0KY6TiSH6cUL0PdQReqfQ/u3zmj/Se7ZJ0k9ou
nFls/2ggX9YCiEdZ73g+DFyjP7mz5YaZBV8pdl7ihlaOgtx+7i/uqDjqo0dzMzHM8s5051tzuaZ/
ZjLAOUTw0kW59nO/IuY6gcwYz6+l/IAF6UREaYaO8RfdFNfGdF9ARGpnMlojIYo3pxd+Q2ErP070
i4CGYCEklbMVlvO5zsWDbFAAB1frRIbW0nSQ2RDRMRM14tK8O8gyBOL6b7sr/pUAbWgQ+Zq9NiLb
lzNJy7BPJCmBFdv161vdsRt91hY+ppuIXaWsP/tzCuyh8k+7hVOmyJQ0q92EcedBi9hW3DdsraSK
EjOqAx0ZB2e/UWNht0xppWDqFH0uoXiQBo7d3a+BobLk2ViL3vJOjC1hUQ2y7PexOUgBJjBm9s2U
Z2O72iW6Sg8CcynBxQAywOFNRP9JRAX7RakE/ANF4Gqggr34OMkDzKMAwM44ArbdjjGo2AUqo6kl
lkcWxE+mWTcBT1sOR4FeCwjkZSPdE+gpOgdWFK4xGOCZx9ef0ns38G4hYLIFNc5r7D2DATVodu1e
JMV+DNNO1ljKZvNz2Kut8aSquzu0UW2TkahmKbBjtQ3DJLRp/GznbqWdcu92FQ0ATzsp2G4AJ0sc
g7ZN7avvhfvZr5T6Lc9/Vjh+3jGCy8by7rqifJohFkDEmOBT6MsFuQkkD11JwVUiZXDiANwo8iSD
xmDGmBcLcfEh3aSrHNLBh3caul+C/S+QRsGHYcDdX5OBlVFYfROSl93mehbgwY/lfAcr5NeN07ir
axrlKRbaOPDxvC6i0fqcMfFbx1bF1kuiudZqALMN2Ml+y+Z+pMrCWckR7r8X9+5GfyTRkrwJEute
AECkxkKOuPx29Avdb4qD8PQl/jT7GofcvTaGP1/G8T1IU97SuRlk4x/fH7juXDh1gN9VpElVGYBj
xyoDHCQZ6rVDx+g1c+dAqLGQt+D9GYf4NYutOqMClsHmNjSLmdDGtx1FYXOBluqTP/p6hnAhX0Qc
JyC9tvYRMKx+q/zQHL3kwmjJVppaB0ndKvMAlMr+HQEWAYg45sJfHlsg6ChSjS3XeJm8Gm2IIGyN
CAz0M4wIksbDhhMbZiJdf6p4+sA8Vg5AZfOqvgnKV768yDQdk4/+TYy3XAitJc9C+BxOmXCZ9FjG
W+ILsPce6/YlntmW23ATb8pt23s2sPFkk0BCax0sJUxAL4coESCq+/vJgCbxjcE4NHqU01DObkS0
SHieXawV/e07OmeUqYYX9CiS9GR5llMOD/+TCI9147xL/kndagCZ9S1t97jtKLgTSdma8fGeifZH
Jm80nJgptkvaam3NdsTh6NhIoHy/CKc+1VL2r58HrXyzGHnjbgQHtA7WZ6xza/CB9UjaJn8CmiJo
pxu9H/DcjIRmAcF+iG5MP2qJvDhuFyjmlpZdJToX2QjtoYaRpyzSdvOGBYpQ0pIjF/irxQjU0epu
DvSipMtW0LOre/SYVE9bABVS2eS1O+W/681ts7QKsMZJpsRVGQauoWITRMzVaQ+b1lyCfeKIdfA8
vL0d0jmsqBOOkJTXh6dthqZ9Lfkx5xEIRhIs5Vcl77MQtFroS135zlJvq1g0ShMe8jotQ8txo2zw
EZiMiP0ke5PA6wPwUIr8Fwphy7B847+D/Ga/CMq84UUoo1gzi0irTTi83AyKwTn4TigbBToLYNDk
HIrWDEf4FCPQxQIJqoLE1J8whywcafA8kFMnakARkf0S+g/KzDwjDEtIPaZhgE/SkuuUbT4SUSid
gMc6oKc+EGQz+N3jrhpi/HLXIbebDKh4H3GTVffUR5WN2j2wuyQImqPXPAKlC7Fmox87wk0I8GrC
pcRPSH07JUnqSvC7SgH+YlX7M7GqHVrEVmycCZorxp8DqSAKO36cVnXzg8jfu9w4CuuuFP3W7xi0
+7iVXRJ0+emmQVd9dmBcYmimXYIR0oxpSYdFbRkprXJKEYlZVequsiFe/plcsgRoITF33jKYY6nv
BS9awmyA9z6Er6cQDo0y7sC0+eiTBc7f7h7qGvwdemSTxK3rX+w/ZkX2IUY9vAaOlZyQeW+9LFy+
4WvYjNJMlGepV0s7/p+rP6ZOs0t9zkpwEvWbWtMn6GERGdUxwade4uQWidSWV91QNKx2yOjxl5J9
/4NtmobBZbNdWHqIvQSzRwW/2axt/1kJpzWRkH6iyG+flKRyHp1DtJo4Nt7UG7hNFjxBVz/etFcC
9698+dYi+YdbPzH3ySO5MPQRnn77MN5NLloRzza5r/KVqC3cJ+5RcwoRH3V+f+YFPmXNZHvzd/UU
GDDWb9RQkyay20bw+OuecoFY4m3C3sjO70VUMW7p7FVZ6zDG5ih7+sIxJhBYW/1kZT+4NwsNRLPL
KaRoj9XM0qL2b88hYSdJK7hhREYKQ09xgzpQEjiwSrNKvhDSObYcz/TKM03qzUcRiIXTZDqwX9xD
Y41fcda3ZMNwCaeY3zOulVk0ra4nDiQjIup/hBusZ0XhqJSJ/CfKnQGONvcwUObJDOA9MQfBE3nr
TrG5HuS6xbAtePC0Rxchky5l3U1ORUH2ctkSdrE5YlTVBs0jOVCTfmo0aVHWMWyFghHpteDgWZY1
Ii5Q2fW7LnJuXcEIqpC7AVYzkFlhdud2iViAi6oezuuiqH0wt33rI/IWyde6R2uNw5PXHCE/dfCr
LbzyTkSsha9x06uxaqcGREtuTBzz5sIu7o/C8pJ/KiTu9LlweJKiOfDghTLiL6nFNJ/xb22BcfgV
rSX/FmfvVs+IsRo+n5RUXoDSCTSyZO3PQSAc5ER5h+tlukJJhYrpkdTqbuydkmXex6ZjpRrvvCm2
u5jEpnD+nJSbMVcFfmJRKSCKWY2Qt/VhCkt/S/SB+T22y0jLf9bPcCYvBFCrDuJrqPmKLO2zor0A
Nb2QqPAp3b7QxtTSiHsnF7MX8AKUiS6YrMwOvdexRTz/0qAYwY3UIS0KpOwdCVcQVvUx/Y23YOab
MtquwR4hJ7bG3pqvL3Emd79xM+GuTRFrWMX3RL/CZteVIwBFzdDkRW+LrRP7wc7mWLtoghkX+MIB
3mX1lCn9vKZMmOUWl6tAVninfp7b8NYX+Io7VXsqN7luYtbrveWZpoUsAisLWjxNfcqgIeFiM9if
I00Kd9DhULdSZAQsBQ7p9jvR1/1tIRx6cpTPgSt5RIZPXCl7lwiuqS7NczYB5xWSdIvPbr3Un7zh
Y+0+znOFfWfBYLJ6sFLhm2faaBxjxIwLsTYsQ+G48Y3jyCOcFGIqHj1iSxKaN7f5EUXVJpZ8BR6S
oVHgf/myuPWmuZP257mr7OtuZnKmTQc4Voq//3X6uhMKzuSr9M+aq2+FNPIC0TXVPh50/9ufqvJy
6T2tUmGQ1+w648CbYODbiECsxydHhAyZpodqcDqCU9B0Z6UTl0R7dR81qiZrlkxutkMkeohNhDI0
UZYngsFjYciDiDRKqDZvftvkkxB7fREB2RJkomXOGsCqDRPxyK7LHVBeSOyw8zEIDzGFwSoc088c
4eXxYI5JzKyhKOS31DUq/qDCi+FUO5gbwqQYtGIidXJ8+vmc/ZMXycFHaG38DSeV9xxvWhkL0Ero
tz2eNLubNOM+FvWgFMsXWM4LbyfercDR+ag66HhsN3Mrt0rlHIVbr9icK9dkQxsmGbcH1H5UQLjF
9HNBIsmKlGXJToyl/E6Kv/c1/nxIrZwZqWmIpRc9dx4cngGC7bgjwmaHKKgmfavNjxmaKs2xn2Kg
zW2rYMdz4HjecwSOWYyYpkSYEZbZV3Jb42A+Ii6dx7tvy7iLtnVDZgkerR1fn5DAYLZec6+RRCmd
n6nRys2wc8bz00+bf/nJ/hoNQiCGuyUvbBbl9Kd3ajKy4/A+nWzjk1xQtE0CgSG1DZNJ4Nl1EE2H
Lv9njqbDU3mwpbRNR4GFsvKBh34BtCsv42FOaYBIFjeJxbrdbCLuMBFEn8wo9yicE4VckPJMk8B1
/Tl5FVnvxhQoHbZB8ZseDnI83x9tf4wbl3H5SL/HhoEHIsASYdahZPsKtH7ayaXGJc9Zx+B/kyNQ
tpu0LCuAZKe8ptZmVCNwWfbcASV3T4wACaZ2UJ/9jwswH+UsGfONNq1uVSdqkTIgAEvR+uCLCJij
vJpqaQhDKvPDGsqMC9U2V3PC6jF4h2tBAJp1wHOyt2pgkP5Z73NqOizsRAevYdhD1OlQXJAhitRl
4+URu5n/Minh7Nn7veg2CI3ebjl5KDSnfSBo0nvQEXb6wcquGJ7KJEqfL7W7M7Ny1TZJmQVwEUrZ
JHqZkRQVOmAgQM/vIBpxHZtZvBiub9C1ZHK7mSCy5soN75S+nKeEY5J4mkJciLJBSfKLB61o5B+q
D9Ve+rs6HPYYNjtEfaQYwuzPWm5XU1Ne6A6n0tl3G4hTx3XFUa+ogFxaeV1Sm6OOXWOYo6vEGzof
Sfzj02NWjlsg0btXO9zz73fYB0wRdbXaCCC4AOr+w/9xJkeA7FFhzNNwm2LV7docXy1l4i+j2di4
KXntAsnmtPapOaiBXdPc6t+F25D8Xny5bL9zFo1ZcsZ2h3OmyTdtjbL/Ln94fAePPuAXO6QDIZ7S
dlxXbkItWinTrGWLWj2oVlAmcDEjTXOzscXLNzCoYAvmLqiuz/lOkNnpQDyEufvjo6E464hKwohj
7vBY7eLomYi5BfXO8Fp3X0TMCGCNu3qPdD5v5jC5bf9tCptx9dkSv2LZbh6UF8lMl69c43Jl71mw
HpeWhp7RCBtsxaI7VJxgdDhskbVtB7HR6ol29Np7FumbEyG7LJyYZzAG7a/j/DfPzBDxePcL0lZo
ejYTcRixqrIgnx/RZ7oF91mJNAN+BqX7WKq2KrRQExr73iCfAmDegsmAt1GgkS2d5lGlgl54sqAq
8TZ9OR3nhU2JpKyJEvIm+RiPfLm7n2lqkb7bsInW+sP7d3oWvIFaOW6vnBXgq/pU/XzKHVqgkCG4
y8/SGvbidh7/2oBgKN/3sJRQYfMKIUkSAL2kfWkJKSxLbd+1bSp1brSjsjKzh6TK9K+hwxN9hJ2C
8oflZZ5n3zH1PX6TMm6fi5lKiav9eefoU28G4jXvM+iFti6eDbf0oBO+6iOr8gZyx951vKpemUWl
1hT0lhSYYq08P/vxrIgXOantkn8ocNFuZ0BfGa1Szrtyh2lDINdgNJRNmLJy/W0Eb2/+ZnMdB7PS
J9r0fwQf5XJ3F5qKageZzNcMKQQ4TQspeKa1MlHsXnaijqgC5mmeGp8c7oqXfu5YqTniKMushyV8
qKZxUR5PdYpldCVgBSKL2kqsyETGUMY8B3f3Yskm/BgL4eJOPpC/JWpLDZ5IVtfvGAJuHYfsJ9Z2
qxjYZ3L/sRDOFZ9kv7eEkP1KcvoxooIf2GK/C10YK3EXNw9Ce2v3YPzXUnlR8MszFoonVKKscklC
AeipkvIY/rfYdCJDY7/as/CMfKHHheLLRc8Zm/XRLLwuvCSsS+VUF7G/iESIQ8mlfxrd9F3QtrAB
E3jaXG0B/3fGn0IIlkxAuM0dY6qX0PZA4jkPrHWObLrxuKLBGCpwTjEA9sYejBriiHm0UQ00wgUD
SDE4juAd0jW8itXUJscU1/ag2rSVk/ix0FSmWYspplc7AcPlzVrPOjD0Tz2JnWjUER3FMICiW1b8
QoGLecE647YCsbAzRooLL2VGlVGVdrC1PUD4dwvns4BA4pCaxqvnUeXPOqZ4dDktEXlOEkm6D9C2
fE20rCpIwqW5qFCH63qqGinDHdEcy/rpfS9yco3+MCw7oXwuqViXNgK1qBQ8E8WAX00/jdg+0gxx
NiSEN3dypa2ZVtwCrvUXuvyRmht/T4zyfeE7XK+XAWTTOo/HZACvTpMfvWr9ZJuFW2rJp4a7Wfg1
YYyF1UYCwZB6V3Rhhce/CKSU7mYU7sPUrgxvF0esJi4+H53z7ZZ4qTAKGaHV2y0K6XqouM1wyV2J
ZL0DQHwvW8yRfAn2dAT7NUUM+tXmr8MktJIYm7plAob4xOzHKGycz5wHux74nSMca9bG/TADxthI
LBrGJT7axHZaaO5XYmrlBOv7MknJ8ze06m+27QuJn13G3qrd8SgsrMloWiEtJBYF+qLs8AUuzy4+
aGmojhDnycDtpAJ5f1etQzU6+nPNZkgJoXe77p6GwxvLl8gU1NDzoTswl1YHcOyi51VN8zv/pVs1
5Cf1NnqFcoA6wqZeWCE3CXf16EKLgY3NdsVck1pPGn/8nvYKke+3qRbhc/8eBtMwrdUuqXdT08di
PBAU2KoNZnLJPU50T0aHnTUJeMrd4nZn2oaqdrI4q3o7bDtGh5YMo7HXWSR1FeTUbqZFx+oPDCe1
GZFIR/sPlTOXfBzUWNlNg00MmLvFz0qoGtuRzeM3XrddS16C7GnAkYZiwShPhd5Un5yqOBggm6bg
SsOaFHJu9JZSkJcRdSSnViH2fpul6l/4rpwjGjg3McN3WpdhwFtc9JIpbOPFCFXYRpfzGnmBx5UM
nN9gqICDXZDEiaHSrLRu7XLRhkuQIbU13KzAf9r9wmPJvlR3HFaxsaghph9BLn1h6gfv/fOqmi0G
pSIP5/7nPlu2NEjTqf2lAldX6wGJ1ts/8lMm5czZI6tU2kkO9plz3ntLaTuTZSjZzr2BINC3BplC
e3nFzMWhzlWm7FdLob83k22C1jAPuuQLX658U6wqD+5W3GATdWock315QbnWZKtmuzdChzzVM30u
nC8XagNBqxsAZ+Oxhgn1W61HJZWHdenNnx3ys/o2lNkjHXTrAzuqga+SOUOHhOtK0SbpPGRTWXlD
OAz3EZ8enQYd2HpS6S/d3FnH17w7pmp9eU7f3YP/3AzBpJyuC0kY3MO0l4SnZ8NxLhqbVRWk/4vo
JY4lyIjJbHw11rsjM1LKIVWswZzF/BY7eLkCxyYE5H3BMnaKG3ZhYYJn5lXl6tdiCdLr5Zh85kK+
Z4lG5H8U23H5RMyLtQ5M4Hlfl1xxejZSzRtzUFxpyhCqC6/XhEP72eCaRpXYvxF53D/wFGfl2+Ym
kxPoVy9Zq4r2eBgwaUd4hcgnFltggSvatXtdjlPxODKRQN8VL9uIUvMU7XXFXM0SXtWAbaucuSmR
Z0OGbjettBXsmuGgg0FRXuxRmXdiy7WcBAXDAFsQfCwShzkTAiSFNCy3g8MamBQprfTwiOVyU9dL
uBBm7OyKLgcuO4HWLy7dEHAYjWQd9ubt4IlLHJ/evkFD5K0Ip9MUcE1SNDLKasj+bFrEKBtSW8E1
GtW3G7p2b9R6amfsqHl6UxqhSPGge88SIl4cPMarx7/w/YweWTrjKSXHWuNYUohi4iGc4R3xT4xc
rhGVwWtOEpuFPbjuwh6HpVdzEUceOENXHCGWxze8a+gLyjwaGMBJFxKcBMDi5JFCdUNplELDKhjw
Gx7/4Exm+EXNKnu1jH/f2yuM2i2OSUm0ULuZKe/XnlYylozhwmmtvceTNU189rSEQd2lBpbPw78R
aiEVBOAIBoCC0wR9TM/6UH87ZNx22uiZApVwudIthZph7CPv3BlK5FmcKJyBEql6VtuEcEEsvEM2
2lUIuCu/ANXiOcGqvAJNhyThIhGZRaRhFHPT1cRjIVy7NeVnv0O+n4CFfulXaOHzzUVC3RmbVsGh
FbBhW3vKwsVj1g4Bl0bHBB/81nuoiw8zxcYLDILhDahcVpR/MD3r0LTTHyL6Kt5t4cM4WdYjuAfW
4z+HGVitp0C8aE71Z6hz+V1m1P6oecM7DL29eVnCNkWDfzivZdQ8K3ErzPuV6IP0uumkXv+RcjXi
92fJqKNfq3+8TYlyWNBKe8CWjFDgG1V6pIoMi+WGM37Dl8BABi4saga0rzl/InIkw4ja+U36dZK4
Pz4AK0oNqZjAsNMuQWYFhI0sD5gPn5AzOTTIcbBV/EITMQsx/QEPIQdPyoYofKcRTOtDyUPPLsTo
GIFsLOe2tfmmwSaDzjWiDH8nLtAsp9EkG3XAWdM9oyBOE7lkVvBkUJfXZ73qPAWzW4PW40TlJXxs
kC8H75acO0bJU8eAT5sWBRjkPI5+mLgko33HNKfbHlDDnADvYWgcmE4E4kDPL8C6KiiqVYN8JlTY
qinXajvvbEddUgo4Q7Vs1YzqW+fyCGKry96kbrs7ZimAqthhl/ueABsoR98+YY86g6GtwskLyV9F
1bOBSc2O2uWGYcqGBNXf7PVwbqnRplD5E71jXDFKQw0h4ozStgIIQxq109LSe7C+1zcnMb08ALl4
BhyoGLOukC1LMp3vP0BHUMWzha92MCnuUnbE5Xrg9mJ8+h4FDccmW7rxk7jDrOo+SecovNMiCFJz
bt1u0Gx+b37M2J48VjqyuPhbL1WGPk+EeEvbJoyIOEIXRLCnAVxk3UE6mbekVEP2rg5Kga14sY5n
anp4PGinFp8Yi/T7byvYDgFpHM8dlml7AP67U9XTlBEspHGxpX5AIBgrV9+3TxXUoP6KkJFXMNLr
KHDzQR4NbjqDXOYzIsHH+3WIqFuQduRnDrXvJCIjI3+IxlyamGfmOqr8H3BdCql0vb0r1NzsRBS7
ws9XnOm6Xt2DjIRKhgkk9+PIO4WPQ3FY3rx81xhCb2zh/LT3IO5dywBhReVQtM2B/vfCEEQk1lbH
wAjnOyVKeXX12vbFUmv2CjnFPAsOi/e+RsNNqr/DjHi+BeXXgwSfcIflpkY/YYYdCavI9oqd+pJq
Gsj98aw7jErqTnAmdVycPrE3PK1rcLCqriGLzRUELMKcBjWQe2rjNIWHQmgWdgWOfMkKifuFgWbh
UvpyLBfx9iY1f4K8iMPNksA+oCvUEKi/FX0p56Zm5mqWk8qC/ciEozJQUl9RAN6BNMhcmwCaxl5y
gd8ayeHN9EnOxrEi4ka1zBqpBqV66GWu3R5+HaBPER5tjwhDQPS/k5gXmMjjEq5mKsvqOgDVdtWE
LvTHJ9fzjEC0+anBfkxdTdnpihjFQacAYJySz+IkZ8lUeqaASWmjT0gIXhJiNxsd6CfIJoyPB/vH
bxWm3QEA36d1vp5zH4wq2jrpioT4dv0gNlKmIquvtrrnF+xpvtgRmodZPY4o5eYPDe6SQA5aNBGJ
S4t87YRAmbC3cT6VctyGYlYGrcGnlYj508PVWISteNPmkdMklNLI35xs9lQIHOJLLFy9rfmO1N5c
1JhR91tkYhE2sGiarBuRBwoUonXHRDtDjF9sZWaEORCm45AKLNby7ZsqgsvEXDKqO6S8W52POqlp
x3M/xpl0F8PnDtZKz3L1qOZRZgHC3zRNUs/L6+S5RX3n6HGDQT/I7V15s0cmqFxEqyaivzX3QZ40
EkIr8xE3nbKNSOJeje5id6eAK22AeOaHyXoc954hxO4AQk3BC+hF14V722IiqdcttUP03uBI5LMI
ZtAfRgvRIovN95wnOsWhSonSD49vzb+pcGmsomTcj91EXtFZlcqGnJuBpbvDZjH7U0Dxkkf6Vx4n
203uyUhV8Fhti5C30xbiDYjGdB+y4gFPeDsMUUMGnNeCqRYggoBfBFksHnvfcVBVIFtEHnj/DKg+
IOfwBp19+sPPic54hByjYdIzUCZX4B3D21vkX+o3gm2MaLggEet/azP0wXQE0qn0BSxb8V8A+yIg
C95ifIPhZiqC7yui+vjdevH3Ube0m1gU4PqyMYl3exZlEFjbKSorftC7FAJWjBbF23ajXsGBfLwg
SzIm/9qHg+acxRbl839TUSM1NNTEV6fjtTwJywbZP1Dl98I5bMI0F5Z5puROFnUZ8t98OElWlnoh
pJVJwUjnUm58nxIR/Fu5jJEqQufpi13nQxvVQO7Y3WOuWG8BM3x3+8lZNFLnLFp6nxBr9wP6yJsb
QhH3dN9quKwsr2q5G++wA0WyB7nvTbITudeYG3O74RQ6ppfBOfHLK+DC0luiQ00Pwh05Se/z4+/Y
KY05Lt0NpwI3KO/Bk2APYHjGbxA71VSGY9UqvNlLli09qCHmPwk3wOmaxONyqkmlDQX/q3nOP+ql
iUeIyWa2Gesii+mlWwS0KORGtGRM9vvLpYr/FkggFBd+y6t5zzpqQ2iQabNFD8k7is07FF+0S0mE
6aTi0YnkkHmnnmLNby1zPGD1I2SWBmVi5s54hNvdbZqXVUElWUO4o6Hyt5OEgEw4CdIGPnPmVHNV
kkkdv1GM3gOH4Dq+a4Gb/ubjSiZUexI1pNJI77dzn4El0sRoeLFCrO7LfO8jOxe8p+tIMgrKXXWo
FCx9m27Rl/RgQ8XCtJD3RUvXp07mn7dFFumzhel8pO3PsXNXGQ8TDU4l4OYaiTmAzbO4CutJT3VU
8TOnbtzRvGd2IgHufZ2CPJbqIp5F4dvbgEW0Wvc+B3qnV1ZActBcFBR4cSWxGODt3cN7RsiO3Ku5
kvtQDAJgfnoLJIz2f/H5s/O1aRH89Ltvrj1UOoOwTRFw82sNVWr1U3x6JCWttJLs9Wn9NzvfTkgF
AWm/7i4GzHqrsK4+UKSxdIyonfvqcVHKwXnFKe85asyqjYGr0fzGB7Bf8HRKJPjWDxwSk3yOex5J
OdLv+AT67i13y4W7TCClE9yx0yON2FPwy5j0z2n3WVl4y9uAx8Jb0EX0ZatNm4JobqkcTFHD1rrN
QPdzpXDclLAciWnGDFKmkWohjhwBGWLKvonW10YLwvrTX5VCT+5qgTXPEYgzix/MZMqNz0NN5fSf
V0OUI/rWVwcR/5CYthnEIyr3LqL73WMaSejdrZGNuLtCXdd9/C0Lr34yDA9azsT0JzetLfZawqaj
woLrJe3X+ub99VH7i6AZZ7Ru4ct2oumqYyqX4S3XFqf59tl/P1YVpefXSL/BB0qYx7STcfdUG7MJ
0WBSa573mJFi+OGrLTvPe8fCsq0ttfzZWqXB5xtxyqS2DaSyulLVORTNKKAL+NJzBwOS6jYHZ2HD
u8fETJcowvQB9qs/XRh+yQItk7QXhGOrYE/CGgAJkyeELYLXPCcZQzhxcqTqAEh/GfYNZlSzzzgk
XYY7qOVlmSC72kEvzHFoKvyaFDSFMoVmrBpz2J7aKZdN9fOhARzlGKduW9iXDftFaEGY5dNj2JQM
o/7APpTl9bfw2ftEcKCR4cTV+F/Y4uzsL3QA5DEL/D0rD6N+IvAM0OwqOnCxfm6nSUMiH7MPzB2S
v83hhee+4Fs+gH2b5IvM1djLe1fU+cp5TpWquceje5/FfHXUNmdt2NOI4SZRHw3igz/0TUk127E4
pohK5NsnvEQAuJTx/VtCQOp7Cm4vs2I7F8mXXcFPE18XjRsyEp0Bm1E4B4ys8/NPCXq66cfAQJuZ
HVaNTdt5AM2AjN5nYzVE5WkAWk+2oEU/WNfEPyI8T3qnjJpl3plJ5aVAtPV0/WEO2odIO+xLr0U8
mcDqBhNrleyQp0pLjYi2wDCxGjPzfLUoSun+bKUZoHAWBLqzgAlzIuSimbg9dCUtKmywF/XKbweu
jV+lmnzvenAj1VqWnsH8yHMd3Z94+J7re4NiSApdAq78DBNzZ7U/HRz61ObKoylYKZySXV4yDHZe
6N5TPEPMttlW3M3EhX5BwAUS961ICUIHh5QkxJwOvgJpc0/yRoijgl3LyvKEtVZgxpRXHbqJSJ2S
KP/DLuPwyy+DeyEipFLD3yNJEHm8jwZSh348ONYk1oIF/ylS2uAB5Myxqfv7i+F6FQkDfBYbAlbQ
WXAI1Mog72wezSsczAyz+GZjq3ytFCJnWjQU75hLIZma6nD6MQzNi6dQ93mqhZ5tgwKekUeJTIy0
bTAyAO5Czb9Pg5bn6J8FRY+1rvtNlM3qDPpf9+dEHEdFxcEFyaP76bDhhHPFNQPjnKK4l94kg/1r
8MQh/nP/2BSbvKO7vf5YtHMM9+9NFxa9OkydBKyww4W/1r5Wlpz94tziP90K/wXC2z2+OCNLUmy2
iweQKQd+ABBhACpXwK2JpavBOn9g5r5m2MlPIerYBT/txMFv5qpCT6MvnQeY4sO0jsoYKrKeEtyP
/XBb4GuOpSgZ1OVQ4a96ywSRift6NeXoHSoWAYYkoueJHnanSqekDpk4kucM7axucBFaNlEndXOH
8hnSuECmtNCj5UPTOOOr0fhxvc75Dtg1bty4hKCndOsvtUS1Kpe9Xt4OsNb8RgoiPD/h7LzG2/nR
Vq81ol7CR0a4WNYqfYBw1iz8nJNwPn8kAmIJsTTRVyvW/c6pfYQ317KjMTlMlbLyGERK4Ji435Ad
szk39S5uC0Rh8Nzo+X0Tlp0Mcmee4g+7GRwyziQ86KwmOh9Sv8I4uqwmv4/uy/zGYgCfDGL/s2xL
y6O2c3Vo04xi4nGQwFSwSwjAI9j01I/TluYQZiIw9DeUJyDwMpDfT74xSRT1OpXRAoyAE2f13yZO
RIYCoP6mghqFYwHLMdMFD/OFxX810aRL+hqOobJX1BicG0dyigG/ffTBW5U9wU+3UOK3Y6nHzxAJ
5MRNIHKHSLYNw5op6MW8PHJX9dtgFMVy7kmY9AbObLTfDhoRvyIYFq6XUufWtZMoC2D9XEkAK6z6
acuuPV08ghqk5pU9ZRYaj7UUUx45qXwY+UJPTgXPV3uADeSTgtZF5po6/SN7Yd3BcjmOQ0vwVTg3
CH1y8UVbAzimte7AvYJ4Fn/P1rKHi1UljABT0+VUo4MI/F5nmC2zGH2KbYwI0CDgdICRyq5KjKwt
hdpxtmi1gNRKnOyRI7BgR1cRlBIoUF38aqNxPcjl10L05R0KBp+w+xrykKITPrtDqvi/9zD/tece
81gQBNAYo6eLiF0j8z/gfd7YX5+XNUj1fF0nrDdZ2Vbynl9ssRH7Fbh8d1KB5070Rzss7DNiekWa
UsU6cDS88rbb+WcqM+hlVZlTdZCPibzDWV7h2TaddOL5F/guT8Enqw/GyMrZ9ug7dmxPE0Upkvwj
wdXg1yyqhU+rUZwcVJHXCXtnLYbXuIDC0dXnRZjOMZPHZAgibpx0bjJkUhiw3/QRm4LWzjRjkyVj
FByw+EwRLAjHXYaj06AlKwyOebGZgDxrpgkAz3te05VQ23/wNmB6ZeZzcAG7+HZW+0/uP8FVWG8Q
T6YgGAwzNxRe7IRXGJlFyLDeuyGCG7COpLPyQ8ubiw5CJSbNIImaoHYauHZLccGCpGrGbJTNkBUf
IT/1UM8DsH9jsJxvch7E4OVeTQB5fFlc1uudGMzQseVjNms52rVzFIc79LZYVf1xvjUJcvVMIERu
LwCmO7ZOWzhXVeK+OqYmKvyNtptl6qpmYOLyGH7JBF4M/Vt97ijPylMzCssAAtUEzHf2jt3rLRSo
EbBbEU+Il3pvioEPpPvwmnyYAQQn0WminxWMvcyfX+Lqbox0oiu/0MBVcpHZHlflsyWP8tgFx1hn
p3oKhKJxErcXjyZKtLeFRrp/DhPrw0Ym4WXk39Kpoo3y7HbPNWpIv92tvVUUysONmhW0p4y/Svg3
ZLnzoCL+2Guyob8V044GAoZa9jkWt6GZSAfJrwxAO4l99gUrKvezxX6qM7l6EBgNHTObj2T2hPgi
CQ4sXrEI+KbyMUDXqxyImeN9AHV3fT232w5RbQtZIo9vDoHVzCpHv6/2yr1Iq/iIJqY0IGRffmj2
Pu5JeZYquGtNCwwg4OWAU6z8TAXezG8QcedTKYeqtxLAf2UMxiQdLpOl94FPhJ3bUtPzZtFaBHM9
AGKAhLH7g58b1iEZY2HOr/6riM7avCTZoZ9XTc5UfWRpTPInJonWSXwt1dh+S08PZeLotz8k4gL4
Er1mILqHjFQTtiORPZhZf83PlZ0G0kWc/hGxTpql2cJWLotCFZvfOioUUzeEctHgkjh3Ob8QcO9f
NSxPtYWqs081IBUECGuIMTcEKpKLy/wC8D0MvMzFFZOTsAT6+hG6ibPf34Uxtc1I6MLV5T3omUGX
u8GKb803snqNZ4ROc7CTjuXBM2KvyKu+7My18Gp4alUb22d93TuKpQylMhE2bpS9AiZsVAmbaK27
JXzsCwDO5sXPEQrZ5g3RYgGIaR1OxWmBITuadmDzfNOfHmrIXPM5Zpg7Zcu4W9dWYbN+JW3izStt
B8y6DM8muN+MRXr3jstyVfYjghPXxrNI3uzpl+T1j/EJ/6DuuA0+cDaz4Lo4SiHaQ9advuqc+xvt
H/vV77tcv/gK9z06E9iDJ0WJ3rcjzPqdG4F2NqPhSZ+aOs1oGOSck3vhpB0odvEmBC4VEdK+ZCGk
iKAuuvXUVKemW13mgmC0ztnmMySCBUHvq+k1bUV+ydLRmTWsAhyE/8bMc1qkZ49Dq4remF/fB8rB
6A5OOV2jret3ywx3I/VBCoFTU1kXToV335tS06mDLm4SJKi9uwg1jzHRtzbeidyOjJvzpniExvPo
nK0oDFt5qFIHi/MbDwMUoYaP6Dl3yWQvkYs6SyB7k6dl+Y10dgtvPNVQ1Gpbcby7EcoVy3QQEp1v
+K90PxpmTShA+wAQSgxc3Z+pyChrNMTXiqphUHhCSexXoDX8Ge27VrKVd4sHdmlZPvgEuQaXWEmF
9W8Dp2YW7fxoRnZDq+IpzkvWdzB266qoYjPsREtLhukQz1D5T0d0k//sv9xKSvltH6GJRUdsHApX
Q3/BOL335iwvnJ/2r+tox6eJnNvw1q2idqOoboPQFbCnJWBAWlpjsSUC/z96fpw57XTZMY72f/Be
XJaN7dTPWspOldry8CXaT6g6lgFqMRI4MATxXRPZhPtxdf4kIKGs+vHOmgBfJUD5gliGmrLWC//z
jwvc/+Mip7xsjUUXy8GQRmIeVCQBd1dlOpwmKiLfV0lgzYYlepE0Wh2Idrcz0j7NEOXLIokZFRbX
y2ZcY70WxFmBmA/sK4VDnfVi8hqEwhkBJVQ/hpKIPVr8HK88PLc2NfPuKvKWXuldZ3WZv0ypG/IX
pcg4aaecKL5pZs1Msg285p9eu9KV897BJf067krvzsYAZYquSuXvi7aExbfH304AfoL2YLFyhEH9
oyLxanJ+0bynJZmQSRTs1Eqdas4cmOiMcRTJG46BBqw1hQRiyzXZXA5jgYC6vguiyg7K9DUbsIuz
U4I2PgKezAM+aZJcdXpPBuF769rnEhuUJmp7CjV5w6kT9m5Cp0YDkJojxqVg0e+pxsf7rYkGPqxA
zCkXQ29+IOXi05w5w5NI2ipiTJjhDDvw8IBEYwPVlFvf293Mds4DaGtEnsIKOMtgu47OQWvhH9In
9NVf2kpv6etaBEAV6IQckXIbfVcDqBI6Kv4vPwCEfzMykd2pAZhzcKTn/eHFw5njKjPqTQrJedzL
w4ARgsr9bau5AdTMw/VOro/FkHloBnkt3rq1/j+YwPzt8zDsAlAPMdwyHSgXgDhz67wQ7++Ow/jK
OwYRDd6JtaDQcPF758nMY5EAaeGTGIkz543XaSMZ9AiTun5zKud2nAg0meCXBc7RGM0qf0khQdET
duohnzNBWkHdUcJZf8nSvjZy9sxKNquA9FkmvIf5yMU/GFt1Hed9mPEjnziFinsgY9sgKup+hRY0
EL+QgD5BrsChY0qAFqbJTR4ABU2HnPphy4WYqTPQ1KvD32OKLU2Fpa2Z6IoABLfxPg3wSPNsTbsv
9PC7T4k/4UeozupN/JHOSTbwDBxTszzRrVKwTmOYRRxQPszHRo0Slg3vV75B3GQkFKukUsR+Y/ga
wldqBEawLIFcloKcrK2O4W9WCr66o4FVZ11f045+4huk3nf14CrKvf/xY2M3zk7LcK59B51LQVkn
wYipI+MbvbmdsuDt0bWrLThF0i0LhFbZ17rgjiuf/mULVcqMRrN1gLmoNy/1nJMr1cF77iJiBsf0
9HRcLjIx6qVtJpWl8BaJGBr+9+Bvbi8AsoNI8UJvCNbursmp/hXzKrKy9FcY6XxdN1yAbLTrrdYb
p9S76iidw1ynGKA82XkWxjkbeDtjxtU6izpljVEtbMjHBEw0ODKbKViqpLI4k6otZbIIdS3UMO4B
1EVIblFxV3WrMCUAoxsGDKBXncst4kkm9QHLi14SXG87LEBbXA9ODKbWCLsg2UQqon1HbZhhdodE
GaTL3qItLuDfK5+OoFxW5yE3LDuJkXlRfFdTCzVy6CBGQB42jwlNGwCwqecasDgL9XCFCpURA71O
jfTrjs3b5Oj/tdFW3DMEvXylTo0Qt/UtlCnVGNYEvVBGKRc+WU3lCbGlKPuIOwPm/hRL1Uc0HaR1
OdONZfyF6nGcimdv+i7zM7lAnniaJkHTOXcu+sjSeGdfPJH4xQOVK9x5wk2iwznvi3ffRrhZLCAx
KcmcqQWFGaK6cbp+kAiiSHbxqBHTVSNE73wvL4ShZKH55lSubd/CkyQwhPT62Q/92N3NA0ekl+fN
ogAfB36cbJmo1lwsIP6V0XIyq9TS/PVkeNncaX6KMk8fv6Lq3E5qaH3ErKUfclGE0DuHlUmtb622
AO+i7UZJVOfh26hKmPaV+yeuS7AVpSM85kEbU8ZuDyvahzWYgEfKF70+ew+1M4/2TjJXRt0EdWAx
lL/fYIAv/rzxKbF1v+ptHin2AtSmgB2LMZt5O3CyFOGG4uxGYoU9ualfvJd0PBHUx4Xs/QTwFYmN
h/m3gCXzspMk2LTHMYXBAQOom93IdDxlYCaQIZYubHwRqLa4Hg+IBaJHG4hGJrpm4QkhUppsG8RU
AY13BWBYg7B5M/p9MCcOzWmWeVV09ePocjEaVACz1XNhwDQex9JQ2CixG4qF51uam/Sb+puk1Ayx
JIMVvrFQ7NJCRtZ0XFcW86d5sWElHowDE3O0nbq5VXIgdz/eUHBcQuAiP8JkWM73aWNOCvW+TbZd
Q4Sge5HslHZaOdPx09PXH4QM1eAG5ys+B67BGXws28M7xwFbsXko47DmLPIqMqkxYUtcYhN69mFi
AjpCi/PQ0Wpedx7ZVdhizpXjWyDYPJkmDcBSIp4MM3t8d11sQKtCjCvzl5rUOvu9l8vrF/6LbefI
ejKKwSuwh+OPQdsNjx1H0o9l5fNDcfP65SGW9MzS6FyOvCf6hRbNPkwLjDoItw+fDFGjOFWsmasr
bOdS3yO4HR1kARMgeXIGo08koqRX6YeGD3PNEH1kqDWMC/xOmwUoNWcf+6PDOdrE/4C2Sbj245c5
79j+O1OgxyuIMwOpbGN3KRvH1kIh9yCEuQeJ/1m37YlXxgOQWJWOiBFh3k9Q4CPGszNVkAVwk5u7
XQCZT/TA10jBdeoyo/8ZYH5/LjgtYN2Kqv6kFBqXXA/RgW8LaA3VFKcET0bXuThuWFYrGEKg3suZ
YifzBvG2894YEegy/NsUgKEsH26JCbdxG+JSg+DmfzHp4KTxnMPwj4cERIe+NbX8muYiKc8NigZu
zrLgJa9wcLurpX3Q8U7U4t8W8rSqBttXXDm8TV7wFv9kucEfitWivuNuNU44EjVjRMMGeqAZa52j
zeq+DCypSko+Oy/8bfdwvlihvJiACboZ2nuA5JG9TcN+zvTMb08/lAziHNm90nG/gHMemU8mr9vE
AJBJ8MG4Zk/ScHXhOw3eqscvCfc4orctN0hklb0UUtW8PgWEoP5F2sZoXK0rxrxXEtuGAC/2uEHZ
mpF4EqOzkzzxAGiH9SlQKol9whAVX+ri30Hf0Vty/z/Uc7q05PEv0fQXo0rQym77pnMsa9daQYmN
b/MkR3rp/Cu586raAeuBQlVJ7ujzZy0mHJhGivuKonHIWNy+wduOtyNcEk0CFpAonxS9lbxtcgOz
ccNHoQENb2TeiwtExbzsHyIeNXgaP/knrXfTTR5ta5R5NZRHyshKd0ywojUriwDK/vD4SrTxDsyg
jlowtuzisp4RobP8L4347VeuO+qH6uRVIX5mGQwlO5aii/liETtAUSVEvJiOC+WrMiJk3OIrAAcA
uaPCyvUJ691L5fzpu1DOTDwPBSII8XuQqUDXOaRfIf6dlFqAFJPFRlLY5/6ijrzyqtmus7KCiTQW
DqDwgQDu+Pl7D+q+UlyfIzDjfSH8ZnoBriV1iqmk38vLUHCD2yLhO1fin3S9eVdNP8RDj9KL+qaV
S4Rz1sTTgaO8Q03inzoYPWIS9JzGDwr5XdPmsz8/rDeIbiGWKD1yRCsvXwr+709iyhSWRZxSZjZL
S/ibR78qL0oEEf5dEZQNlB6VH8CB1tPTZONQT74kRIKmmo/t04qpuW03tkY21seQJ/sPsWVuB5Pi
+UDDtoq0xILZFybPvueKQlsstq/xVWAhl32CdFpv7XpIg5WGjnyGg77du5xu0Ufx2FGG3zq79auP
CnWCqxdw8joROCndSxXkS5XJMavL28AlByqIHztP/xt5TUD2NH3zRlAL+Mh46P71MpuVW/TsBvk3
0BKsqC3L3W1OTSzHZIoIaAcQ6LrnIk2C9LJl1yQPPwwGDoUW1KBozk2/C8MA69vhMG8Cns6xB5pN
f/pPEML+394A6riQNPfHGpeP90Y0jl8c3nGQCiCP82+E2oOkFvQb86kqJ+iDBlIH9cUHZaghAkcO
gnXFuXn7ML751IYZNd41rlSCYC21pgnnyZafsMN6DTkjl/Fz5Xku5CBasYsPEGK6i8OJPLUXYvud
s4u+Rq5HWF0DPtT/b9iaHV1A+i+BhrjcFazKNUBUZQhlzfciba/TjSO0wnQo7Ir0qdd+l9b0TLPe
RWopgKJtX69Y+ixe9wCiwLVpX3cJKs+N4serHwW/GNoIYChmJcxdDx1Demspqmf2GYhlM6mfZLnw
P5n46GcWWu6EoRNn5BpCcqwvc37zMbnavOIOtEKLNt4w+//riFKomT/iejRlLqbs4brbZYTuyW41
s0R7Pm4Yegxdt/AzQG9UNhmzhb5RwPYAC1MnTpj2b5Rf4p/Bswga5dXQOQFipcxPW/dDCRXG2mBk
njPAz63Q5p7JlQT9AA5PqzpfOw+iirbRWtNaSrGQvQFbkZ2TF15cNuKonS6iqrH2apZ2eUfBR6CH
+L+oaW61pnHFF1QWthL4IC5wKD05ZO0miDBt/bNvlZkcQIfs3NP9fVzkPHaiFa5PqVI91kcqpUu3
YSt0Jup1AikwHA7Dv78m+EvdWKSls62d1x/+eUqIxKLNM0lYwL8YhF4Ax3T7dNeQy2ZENVh9xrOK
nwsy2R8o1lETbRxVgr6/bKjtjikJE6SMWs+NP/PUeaFhqI7bs2EJKHn/T8mHPOcx76WN1YGq6+WJ
5IM7li0eFKa4cM/BruZYO8qSCXToRwT/34ZXanaKMyJn8OjnfnHjBxQqC9rBwjCFl8/f2rZvFJBk
AxeR3H/ZmQ+uBcBVfBz8DGIqIDoXm+KF8HO8959gZFIpqcCD695XRjkR/XSTQvbU4uNwrhajiFs3
5vYmbjl6K3zRuPuVe42qtye9Ugng/N/gThEYDzGSjLGGG8AUuDhOHUtMgq13D/dnGO3hAZ4vDI+e
IhTwxI6vJsKnrZc6D1AFJRkTjLAGUReI58miuHguzE1GFMi6Oz0QAH57IRWqD4k6oNbx9lJqK/5L
TQwiIQbIY60+McXkPOr48yxQ7TCJZAUhHLzy2f7Q9SQbyVNdSFUZhXLNNQOj7tkg8hlMG+apN7vY
ABRus0UF9qHYnu7I7DbV3XkdsQ/r6wFSSs7Ng9jlRoPJOJ3JPjwgu+SA8SSm32b8C8wqqXHaOHR/
5WOHTaNeZIC1nZn7865It9yb70txdUpSvt3+b+RwACT87zNNM3JNTB0Yww+zbVOGCxT8wcbR+xB0
i9YQTVj3wFqLdUixDdrpOpJRYCUzQuOw7YmOrxOEI9ejp/bEM+SunlnP/OEBVJJAI0lRnrjaK9lW
RI8/JcydFa+dgGEVQ7qDwHMk+rz5ijlFT1MmaNsErXmHb34vuOAh8m7rfRrZW35nZQUKTzt+bnw/
t17nFTDkqT24KrfQSGJYvTBxADRqvNXZhFkMqgC8jQdpx0lSgR/IUbRP7x3xaBxga7nN6GHm+czE
aXUoqRq0vocKQdsMrpUSEYaQO7fJNzzuIWW8v+dzuEMj2rhDUYhRtiPSYvRQpNXQveU+E3Nh6PXC
GJe23ejQ94okIqqfq8NGytec0IXy7UdJP1SteNAbW1NfuCuKpWQDD+eXJ7urM1SX4zRQ3SwdFXoy
Qzv+Trf6nuAUUqRDw4P2yF2IiSSx4h4kdR1VKpIsOG042nAefwIblFeburll+EuIwgElRZmg2FgW
pHdfLjHKGLxtfe5t8dXzqjCY73YEoS99TyzLH3c6asnylmfeyeMV/dbMbNPdmWCNwRHYtxzDiLO9
mQ2o/VEgApYG971LsP10o231Q/2JKZTLi1Ac6xac45Nju11PrVATMB01ddjtkiHpi3AY7SQ09SSG
w4xo7RRjimFzw2Vn0bIadg/l57/KrNbX7gc8eLua7JpeWvqtvs/zZl1mAU/LXVYBJ60wO/ySPqQa
Z+bJxz5O5X20e0HdkepAvmTHygfMHAIKvDoN9Pr8QZq7qNJSNm93MoprmlRS2Dp2OkS7qOEWP9BE
gbr0UIWX7Ty9cSnzUkqL1EIyxU1Urp4QHC9fht727Bt4qHSv8o7vOvXgyNphEihkIf+IIhcsD0Lk
3shzL1aMabLvONVuq7zUISqcRXYA5sSVyOsF27C7vRbKR9YlhTM9NX+CQ2tgL1vXJu+m2Enjzqik
pFJd86aUnIeQVPRn8fgjyHnpP8YCNRr4JkAGbrCh3yc/LbCoA29xIAXhrThmLGUg80FBCDrGcxM4
vGR1wX2EwBXThBuuK5G9zW3JM/W5GhvJMXlKherAvCw9Iw2X7ZF8Eytkkt6bYV2pU3XnsgqIGClB
X6yVnXt+YigQ120UiK/VMKyx8EygDnQa2W9Onaxsbw7IQHBT9z06fDb6nwzQYNgkzLx9TOMhFJxT
Td6zJejRd8NsuVTYNcoV6PN+seYzFJH6L6rNA8kT55gqXKmkyqWrXJwPQp+P9Qch0xJ5X00zcuMt
EPYYRW/UL8/AB379a8OOUaCD6R+nQ5JpinnXNjPSRmC7+bhSXt1lpw4wLFBousR9XzbCkKxVxVX6
/sPSHBjmhn2rP9f7sw2ZOTxxfN9EW8+uXY5daJbSKhFJnlHAl/RiCDUStfziWJcnejaAaKDdzKvl
4zwl+eVjP0aYRrxmOAXjSI1xcXEaEksdEDqmeYpaCv97AZTmbBtDhQbxSdpd8jJX3N7AdELBvgWE
cgC061I1+C3yOUB8BADS6NPFGQnHJaeRiBOB1aLtkCfXl6Y71BOIoTAnh1SFj7kzVtZwjQt65/o1
R0JqBZm3j/4OnSjGx29HIFl2cTc6te0WNas/lj2IeQWsILZO4q77TGHltwcNe1Iej7swliLPDwGb
2rH3vwAcCWaYgHNbuXOJ5MuGmXDnjD7/2fe2nOW0iaE5TVo3g+Qx9+lzm0e4eGzq20msGOYBZIBW
HterbBpcx0wsqhP5V04jeGUhUqJmqz4lAG59LvBejWCP/s+lfx9RjETCrbpDuxjMU2TevRU3F+2F
0/g5SLoy8pFzN1DzFRzc0pDhERrS1q7SKtavv5uVWvZ8Qwcp/2Ejk+TL+d2nPUCk7kSwPMcr/dl6
kek895AEy+pzT0n+JPu4UVRmtzZinstS5DCbPOhvs3hUFBMGNnvm0eeg+XbuQ0Xwbhet/esKzGOz
onivUPZjdhCDWOKsMmeLKp+51Ip6sK+U7l583V+pk3rzbjpcSJaRzcPHlBnJ6X2iyd+MMlB5haiO
f9pNJlsZ8d2XHCDJI76C+VXNZdEMPHTxxzyNd6wFmYinZcG90EgapD+RMk8f9PbHqhggeGuz+I0P
rnVnt0Fdty/GzHVbwJQoqs9TJfZjf0XahJXgSSHR8r5i6mLeiNse2/INaA7CkCDMlL9GtSSXTusz
DHRYgd/sLWFW98cqka+0E5uryKIlEVFjsToWS7HzJRbwDaZ7UqelC7TlrLW9Vi78RY6g+MPGX+IB
pGKf9l/ia9x9ywJVynkiGFs0SU1ZUdrWvFK+SEOahjDJrnBsraGEovZky1oiml9+/PC6DLvTmQsf
YSkYfLJo63Po5wBvd64IKXw8bhvqJ96AtqOYx8sk+ElKpGVl+ANrjNpAeVc+WkG17qw3gv4gbvR2
shn5heb4/JwMbWoxnwuNdS9CERc58x3C5D4q6EI1p/xl99H0T/g7smK1hY4fsfW/YpFerSh4x5CG
clr5o1u0wCxcB4z3Nfcm9VgDCBoKjAA7fXtPyXm8AFpMyfmUSJmirxwhAAig8BYIrsngJU1GD+Rp
/bSEe3BZvcr2b/+CCe3ZQJ1xFWoBopGlU4XnJspgADpd4Hpi2m2N9/UohU2VeWFEIzRhHRunNCXW
8DqrQL/Mtqg6fR/uXkP769Kn48lKTqOnwGTHs/xDVYLNx4GpPzoHeH7sX2D1J8RDD2tNQclLJNAr
zj4NVDVk7/+89fxW8Wp2xeS+Pc6+y9GbylWrHUEZmPxXFrrx+q7ffZzXvg9rcUZu+mQaMgHMLyMu
Mu/IiJ7f5Zg4V9g/0izPBxxYU3XECmbFjn0EtlS+w3wjeGO/AJ7jI/Uf1m3PDxzL9lgIkHUA0y44
naHn4i938qhn3zDego8fGfQgasQMM9xat7N1OpJTxOjcx85zdqrls2J8lQAAs3j/LV14ZkxYrxxs
VL2HMoe2r9h1I7eNYibJ6K9SUuhPmZsz7HcXpgNaQ8bKVHJafDOXaXLeWYrwTX80+ZNEhNU695ON
qJH47KRtIXrorCvpF/4bGPR373yUcvdF5XhNQYv3NlozFFGPNhniiOOO5GEXjv+ZTeThnvBg92Pl
LBwYVvUyeQQ1roJ1ubaI5JKwE+fA+AFDnD1fAFdeyPQQUUvQjr4CMy7Zpe8bWLAfJV/usZjj1FmC
i58ekWZfRc1Do2oOU52TRZptQoB0AVJWpoqEqLzEggG1z9SYRRq9GT/cEL4aX9SZi34XKaSTRAJf
y4yoNownKyd8Z9VYSwcnmkSEreqN3dxQT7q8mL/PecbLbW4anc/Vj8rA45EPL8JUzTtYoJBhYUMt
rWSocKvCbxqqP+nk7BWAxpk54Lvx0WaRRDwbPjhrbO1S3oPKAT9At8MS828se9ApC77dSCRT2p7A
YYPzYI0jgfAl+A7HHZv2YtAAGIaJegt+OFl8HDCGS/eT3vWtfmCc0GAXs3o4BZB+BODgcFyLX7S6
pYFv9z0KeRzZe21nS5MWx+UABpKxn6xzj+OrOaPsWRT5cFp/As8SRWG/lhdE2Wq25rIZPTYjHbIN
VatIfFL2P6zPCmCot4ZLTQG3ei+xxZSLH3y7nL0PN6DruqP/jE3UPyAKnV43ZAyRUlr1PCVo8IJb
lc3nJBBvups/TtDAdFnj48zwMkHWBGkThiJ6UNE5Csk2N+bcN/QAHo5n2+xjCg0PZw0CdQMHIP7E
s8i73LysF12Bexsi5lgV2nSdtAizBK3+CuPB2CfTUTh6fA7pedGFkvmPtmBFs7CYi2j9nkIz9kp7
XDCq7Z4JW1RpTrnWObNBszEHw112ULJMyeN7ZA75gS4ZWowVxdk57XdTUOH84XPZ21GPasZQfkQV
6z/Kt0D/1K1F/1CA9UO59+bCwPQg0M4tNPiPraRPpEnsS8v0x7oheT636un2czr4DD7GNFj/c/jH
FmkyIofWmgxDa4bC1vJSeL28mmXUNc9yCl5AJP/uEyzhGRHcrw24MseF5zH4k7wxFwqZZS/n7XSM
bthqcW4R4iUp8YjwGtsvKOZTifetkxY5PJlHAYopbjiW4kmfMfn82eUVy8HulHtvI1ukRryDu6ZI
Gm37ixiglCLvhYIUzNCRtvLprVJbbkAItKg5LUWgDLK1Zxr21Y3lr3uxgw86EmcARp7q5iN1hJvV
RaBL1lqMbGY0P/ULYLoz5ngclPi7tui+zzRl54tWyM9CUuiPmBvWLKp+B6BYp/J8pnhoUyfYS93e
oSpVClkmS3gZfSUfOMTV7QQP+eSgKulZYAVsTXkk2CA/UzR35xJnqkicVb1EDCt15fj5nnKlX5hc
D2dE9dqISC5xRCoVQvyahOlMfTQgZgkhjq7kT2xqZaLg2JFqZcWfxA2GZDLU1pyp9sZ+w8cRNxrJ
D2Vqs9ZBcI+MKGin68dlnBjtKNRBfSdIjNqCEbNHElFB5Td5+A9jQB/D/U4vYfvws/5V94ca8SfF
KpOHS7XBjSPRuklxXxUR8eFJsuP50Gf+t+x7mQkvdnn1SM2aMQz4/PTOki0mgy+Qhn7hD5C1rupY
+GfMoJMI41Z7BgoEGJ06mIS4IPdS+QV6mG1ObnVqDvubhHEm6fC2WDSS/EeKM6ZZhDmK0+ySt7ew
2g0imV8YaYKIGF7nciXsXJJ+5SZvyctxcDIEjqmseIl6yNcVs6cBYXXvP8+g+Ue2w1W4aJURsgtn
WcOpQXx9cGV6f/N4PhVC4G8I96801jU6P3+zsSkqwKbzbKwkJQEmo8CLvyND7LkdvslwNalrTUhE
uyind8ZlYN9VsLhP7H9TEsBQWPZOmw+0WA0cQax2HXLjjOa79CnyIbfpQju9fOChirHbVjGVJpPv
VxRP6odY4wUz5d1HOX/0r51HMRcPYDm00t41nRGK0PJRVfp/8iflbw7Q4WY7tEkKHQ1ZBMVwf+kS
h3KPcVAgZXjTh3W5JWrZPuSNYsVpATiLy8MNoLP47KlTjk4tYi16vmEN7yGjYPUD5qTTQ08hdUJk
KB9yUM7Rxtp+7NrXnl/WGXtgaacZVc0eT/dSfl+o7sv9RhJLnSCgeuv8RB7+cZWMzTyZz6tH6ERJ
itBuDEb6NZDZl68iZ8/F4v55FoTIx3MKWD4C0hpoCwJ5+2OVhSUVJS+ht7LAj1lG/7YVR7EITTi0
3FndpaowxS8XbkWaZyboWoKl5Obwq5scdEiJMROrPK/fLJC52Ba+cvV2Phf1wvWW+KRP+GMTbOIM
DHDa5bnmpXFV+9nw+WZHFmDs7XqOsyXOZEfziJhERpq3c1Ga6P4lUg8B0k+YjlEkb8a9K/2+8bmo
uKMkaHTmGDI6o8A9dCMHgESZA9it/FkquG8VxgNDrh9HN7xQXClZU9oG8rFuVRQKiMJb7gWyZs/1
EmwsyaoV05D9XJOT/gL4bERJrjxE7UoRZJWKtUbL5xuFlRxixC9fXRaFwOsb+k8r7g5eOFDEtJlg
xBh2vkPGB/N4v1vfU76u5hTpTapHV4ZbaOxL15U4CoVJr4aBD+Ov+6vh72K7mB4AP/9GNsdIXMWC
8oAjQOfNpQk6cGo7a9gN8LTOXHCFBK49+FJEZNcdzBejwhKS23w5bZkr6HU6wokXj4Rs9CMm07n5
l+8YWf7skC6i30UgrUWjNmm4t0i08IEvaDWVw5TxUKah4VCuuaU2ichwvmA4rSjfzUA6fDOlBSrZ
luWHAwRkIhNeDs69tPFBrTezLuaJjBAI3ljEGpoHfCBFA62GOS409bQa4Cf2b684OBH87/prS8yc
k4azh/aoBml1RvRshcUfQChVjOM74udinEg/WXA5WHofqnOS/ZYWfInL1HGQwIp8y7GaHW5/gtLz
NJCFAkjIFseXMeKzBMEwy1lPXgcPOrAcAxgyj2HMZKmndMMk0RQ1h5eLaOGWOfMoORaSfHQ+n/Sr
W/0zsqqS1Ks9782lMcfXmnSCIu+PgEpSGW15BgopxnEgJaFHJBP2q9GlfR4DqAu6aSVbHpVj4Jcu
V7VtTVZgXgO2bkoieWKVxUn9/GiSA5tzlUXgSS6ig2A2zbdIIhldBR0aLM66XsVpAMneZ7lJCCiF
rhK0Wche9ZmGHXZazUr32xzCzIOJ+XaSgmkQmTPKf2PJsEz4Ozk3EcdAZ3O3JH7EHql/FHse+o2d
EfOOcapP8i0vWoPkI6XBMLaPiLQCuyK2tsnWlBbZhSbEbzqoUkbviv37D9F/1ngORXS3u1Z7rS1u
X1yWEO+jfm+9hB7NcIYHGXNGHhMAZczhBxEo/nLTQjORY+HBn51Q0wIM3VzuwF5cASkEesI5axdv
RlnH93bdOEQKy/SNtHLY3dOwHBhuZibHAnM1v99/hGLPNhpk//a+Fv313PRM6kLvfgbpc11GNzE+
XiBizBHjVM/ZCU2eApKQAzAYVObGDSptWh8m5zjIkNujtjXiPzJcGubvetm97LXF8a/tjj4YtpmT
A146iR2CsLy4CCrDOWUQQ8fd3UU0YnGtWa27/IDOVL4UPhsSlEt9iTHfV+gvlrbyvdM4tPHssyzO
EY8URetODC3KUvKEnGJgWCzsCfTDqmqKAcybx/E1dgwhImrMoGu3VePPVSdsA/PcHsBMGoES4txD
dyinToGevWO7dZA6oXtASv9B0LN6zam/Ge2BC05fq48qfcUYYAI0K9A/N7PQcWVU+XxwlEMvehM2
vdhXLJEHemQuNMbkgEvb/yuN63Cw/XDwMJGmFEohFnjGHjRN9igtIeLd5THF8qoHkSCNIQdPe6TX
Bmdaghua2t14FcNnercnQSo/5BwVtYNxj3Qehl5euv5NPXLFABf1lkIl69z1tCwGaIPnki+C6qQI
EmMBrT1P0lgEAhq84HbXLABetYjJis56UPi4496iEhIB8hS2EsIe6icxKs1224nqeD6W5W5I77T8
ZjYtFE+m+uhmQomW6RSs2SR36f7RpyS4uYuTqHaZhzbnpsIDrYdO/oYWypZSjFQLjU90AUrSOWC/
7HkUfalV7Zf+7B60dFingjejYchk8NictNaHPTnjUTPsuAvDU1xDk90A2nHI6gqS6BEAExodvevA
Z/XGVif3t/N2Tvdwfyv2N9QfxRKGVCtiX4UsG6Eo0VYZsZO0keg0jTn6A4E27cgpqJFhOFmzJiIT
TFMmSLM+J0XCSXERoxUwZ2eiUzhRRkAyHrHoZ1BxI2nyNT8nXtj61UJNkDfbUxHYviQAzMpKjchp
qZEDb3+C5GvzXcC5H945MekQ8KfHa8pbiKNBugQW7Hv29Gn1JdNlgzeEoqrlXDKbhaYzYHJBe1kz
VGFCCWJpiyNdraDkas2AW095VNFnSL19P8MnHmUQ367aOtzNRcV88cHCs3JVHCzsObepTJqvgfcL
pZj/8cHy3HD8OEeUdAzTg8AJ007gJqNtp1a9GH5cXlYvtUUJ2sSpGLeI6QZ4ks3eg9BmB5z5AH46
reXw0Uv9fVh5dsSw2JmPhYsnZJg9qegA70n3YXzmv1TK1YRVlY1MI+l0sbbOafMyXAJZWhSVXtg1
MdnnNkttMbn2HRASOdBnObirAg+2JTiDPuY3IffQCC38SLVfXNjrvyG0TjeKO368gmq4DtuoYXr0
wC+KBG24wyPzUu9SkvypdN1ktM3I0RG5EMO9lcbC1NjHWVe5GaxtMWUWEqXv4FvFZZPXAHWsKjAD
ZZduc6FzOXCgMQ7rCLcwC2GNRbAZ9HMxjnkqzY5CZxQR5e8M7c/gcOfWaIAWnr4dsmpXges5KxFi
mCQYavq9/G1kYpcyVAxEOBNTStE11SsVuQ/luRNnvk2n1FoOE79cRIn5P70wiB4EAWpDnvYfIRIJ
STDy8unwnln8nFHNKDRfheRRkOXV4NbH5Vq1pH5eadboVtRqH2ux3tg7sHjFH4wpDeq+Htv7ggbY
4LPFpHN0mWsA2yau4bNlK0+bY/bZcPk+4ylGGalnicS1QJTCU05v7BsyLd+YbO44717axtBUkkLI
UvdItc8Dsm/celsVCQO3Qj74KhLgH5apJoXXwgUq3Wrr0FLM1ra6TdNUBEkTw2xgp/Jk6R/YGq9W
ZR7UA1vdkksTbLi/WcwR+UoQK+e2ZQYx6WdtjiYPgNfs3OQiWMlIC86A5hDMrbzfTgTfxgmpXMFT
JuOVuuIb+6l70N10sdUV8juZjVepwXZpSv6KkE4r92/GA+ysaEDr7ABchMTSzGn8+Suj5jFf8CrZ
bP4E36/ayTT5pao2vav+5ue1RkdD/LHFTHCTq8ji5L6vpGz0OBS9RDuKyJM7BpXcwSo5DhCtiVdr
LNv4Cg7CufBLqvdmHdiyaFrR+Os3hb8JKXa76owouHiP7f4icXZr5rI8BYIpmfbkyyIJ9CTUVfil
3Dgn8espae10SFPugC/fWNdE4xSw3TIiovxmJ1lr4hCPLZDzpkRt3QhT1zG8aqNAYivwwfV0QADi
AWOoHqUhKBpGbR605XAiC1zmxy+VIiN4L6hua04km6CimrlXOGBKOnSR0T4S9H6B2rKfbeG3Ocw0
T/i1jgccVd49M538LI7svOc6DZLGvYYJiPb53cw5S7KMLv7/af7rwk0N7+qNz4WEsMdC3LHcYjHt
wpMoaY00ql+Ds5RX9KJdIpqcja641+8mJVyZjCtdWZvEIftt5f/7/gN0PkoYgq/YwnYO9r6N9mRK
se5OiRUuVTHlYIVoox53JRA4y0ojchiIDZiZM3ixzSNQZVqNJh9xp9Y4U3apkhR7MrREyL7OfrAH
16swqOKqZrrYNuP0gkEEfYfhNz5N8TFZMwQydkC/RHVZSUjJL+2KMpLvXzL6uEAQG3Ea1c71EJo1
CmAaiMmTWtOoWsJs3Qx6pD3VDHVlG6V1+hObrjRUwW9R+wkPyV6sE4Nvk+dE/kZqhAu2Gy0u9e2x
5l7P/dI8EQiwdvKEbHyWlrNkl00gXgstVfi4o/krwxDOIBoKjosQSkINhTS71rp7jkrZyxrkr95c
YuYAiM0QKsJY8vvBjrH7aYXgLot5cjezbahJV2BS7vtPpG86zTCmAXg1ncCQVLYsIxn8T9xLWBo6
io7X/NWokvgAAbY4lrJva7etLVS89e9Q3vabj+T9Z9RC77UTYegKK6L21up0w67Ktb7Eafy0laMp
dBWs9g13TZgV3KZMDb2WE0XbVTSxJ5pzqLwNpPbZ+qSGdPIKa5Hy7dGmkZLOt+ne7vxrpYJqT+lg
SSLNMeQb8zTbFNv6X0IfrLZZxW6iiQan1zXkGz9ItUB9vmuUnCwT04xsk148wliJOJcWvf7KDu3x
TRiNslDuy9YTfYTR7njYUjOfrHkG0uTTdSrdPZUdYchXEIcfAoN9cd2GxVWNvoD73F7IicgWmJuu
sSNeQ6bcFpfSq2GZP9wXbm7xN67C5Ern+EtkrtPt32ZVkJcgYQOKKagdxe2HrYybDnPVtXCShhFS
X/BMVu/zuDeOZ0bod/xYbJ4p8veuDL60DdXVO5Y9V79iv5fxryJjRBFY29aV4JquhfBc14ERXzVk
gNyfi3RpdPA7f3i2LoXSC4cJpqh9YB2MRH6yHpJwn6dVGp4Bk7CIjnC6ugksI3Z3gqX+aclNZfSK
2tkfM0oDJmjcrqC9eTdd1C7zV3hYa3lzbWni1L8K9anvGD4wVprmTeh9Yj+t7eBglYzDDHBDzNdi
7l5y9KzOCvgsdCUP3MJuMBV7DAXHSadezX4yJo/1LcwQJrfWEbg4a3H9yLxXvTTaHl2mTQNPOCWZ
E2I4Tle7B02KcY6UCpW9bIiN2P0H+c/VllzVQMVA2bVI7pbTz2NmLqK+IsEyarw5Y2HnHb3F2cy7
M9SO6fWzhJHC0mgmIuLRNgMAarJC/5H7+DfNcw5L4nttd/C2kkfxu+jx14UTGxQtdImOExOyz46l
RM18lOQim6X/ncXIstLuz4l5bNCleix7PPhC7sXm/AzW8Wa0iWzc3M5LkDw//Q4VzwzQny/zRKo0
1jEpuKovVwfFSwrbNCcOoTAB9wdqkL3Zxr/mAQG1/f/HSkUZeRo8qLVhBkqYZq/2qXWnXg6cjsfe
PHvGHFlbPA8ojLuOz7F5sl6OTjLeTNl5pjxA4rI1du00Rp55aL2J2krBiH3/D6my6g7A3Yz9fG4d
RqN8twuWup/7B4/Idd67n3KwaEleIHP10sA/ZKjCdD4sWeFidToa/lGOclatRppTGRmyvAjtpKx0
2z6DXn+slPWoZJHCPk+V/5w5MUmljSNmSQNz/B3LQH8ueQz43sZ6pPAcCNf6ljGmZUEVKQ7v/4OT
tErjwDrMp/rdFvYO/HvJCCpXAPcENpwxfmujiKx7lLOXpJkh5GoSNH4UDnBwpIVnE0qZ3dgoB3hF
ETE2njQ7RP7lcsJslpXoffR2xItEXkpTBccu2aUlJN2V3hjI1z2vs0++Urk+fAUIFqY4/iQos2tG
kYScesdNv6f/eSDnlnL/+m1jPw+93kfIWy26vS8WcbzjPmoq8xXC3PEt0hSv6V9rcFxHre8nnaRF
X4i3yAJKTEK8SBbeoLXVZdLl/srCc7PckSPvzav8xdO60hpNs3Jbs0ZIzS9kYWo01zK/BE1C+Prx
jy0uK8gAnyS1+KB8SjU6aEI6gocwpbfbAr66K454JeQC+AgThQdY6GHdHqwwpPSE2Ks/b5RKkOZq
oovnjGBrqo4b6AkU0cB+K6LkIHlgAq8PH+CL2AFfnpxXHkzWyAOSWjJCPw2E4CY+oT0SFUV5d6or
m0FHltXh1YvudoucExhdwtbxQ/PihbxhtsBr7ealjrTP87TKHniIjRhBtwJnBDZn8j87kSbDGptI
UZArZe2faLcofJZCtQKY7OLXCOXk/cL6s9OVY9S2fB7m6EfL0eyRt0iyVH7v4AuAlfgQUD04bCtk
oQp1lESz44auoh6U57ds9WuEtDg7Ygq6lENiJGyM8y+zgKzBKUBlQhIRdj0IGgMGsqlemmDKyYhF
HfKkMT/Kdg2nt9Smh/5J+ZCFVr5byZb7nZF5nZd2Fo1dc5EMVEZj7WcJjvhTK5c1R5t5gh0SQSE+
CS3MvLGWiQh97Jsc79ntrdevrg8gqu1HICDPlCblIfCzgpZfsDdrYq1LUxTKXFC61dAoJ9aEj/HJ
g/25HkwEkCcMhGGyvSop6BGsvvWkqShTegQ/GkjqVtS80SoWLqX5xuzwEDqdz94z2pnqdrl5WQvP
VzlNikaSJ6F5aNO2aGU3UcGqrmbdeQVsyEEio2eH0CsL3kVSaepDaXNpXLa0YrjjrWm2kA5/sdZs
hUbhi+0Mt2L1M3oSEt9VlxXi2BCxae/q3fd9lspleFHlUrTSkRutwlg64j//Q8WM2jB9NYd4B0Jm
ffvMWLwWy4ttHyGRSNAVpmr063SiEVj5ycf+MgOk9XwxvT2dB7FbIsF4yfbWZ5oeVJGkcNZHG2zK
T/OPGBkQRoRORizj5XjitVye25O3YK060YT2XU/npsB99QBMrAQLaLtaHtdwUd40cbgkWw4KlfhH
mDNwUjdxI61wzMooaKVOiA+f4yOV9BCpCysx/+Ih20UzPEGnAhjDoRojdHsDwnYj1h6LbzkpbQr2
GkE9AQMyCt1+4c+70K4ZH19pFcGklt3kmV6m4LbkuCtoYLRTwhsQm4b2hcvNY3rWgYb97oDVwTvc
dVNjcNXVqq+WEnutA3K75+QG6ZgvUuHok683ZjqX8tVxgl8J+O0R5taSckgTPY1rnsCdWRVHsPjk
mjFFzsNLNt/ZwF1B9kcTd/OpGV5Pczk+9Ws0P5bbPXx9ea6pFB4LIqvHhGkWOEusXfXgV2+Crdt/
ysc+7E/FzgSlrBjIpFnofMzrrKzFbtuh7p/BmV9+FyeEgLtTIkWnTJxywdh1w44EMKR/N9A5r5Aa
HhWNko9Zh4zGyy4rIX9iv1Qc0z0tsDbnNkNIJUjlip6V/muCrIFObOWW4sEaf1BUXV4SxxqK2Pkp
8CqLAQ8WdojqGerBvjaSB5C2JpvudfTaxEYisbhgtAX2teYOr24AbpT74OO0lZAMOhDdTQ5bmHaz
5Vx4fbPLHQODXCy+oEuLbSOgBbZFFQmYMltccmHqq4FfRQIPKixxlAwYWwVlqy7Y/D9l2rkubHIZ
GTds8EeBmKbhhYISRsx0/ALSL4OBd5OdKxLSKV53cqyhzrhpNHSqNpv4KLuSov3YNBxVz8Gq/zAw
YtoZ2gE5XJZxaDEaQgMVq1h9BSsXJHfl6hAa6H1K+H/MnTuHJYQU/teHy1xWRZEQY0NDhTq79w87
4Sfz29pXYmzqfzWOq7bAmR9X2GhuqyO5jtPjXv8ctTQAlLC9TEdjCSNmOwSpYANKEEyy9GtWZ/h3
bAMcisn0RtHWxw04QDSziuAiT3FkYTulwhgEo+LKbaZSgZcy/C1E+nHfRVYNNvcjAdnQtJaS3c0e
VMMPNIixW6fN8lmziz1/esvWLc1SYHOLGe/viF4Xi77cGk4YsYI/E8Qyq+20+kewR2cZ2zubzu60
g59e3vgf8LBoq2USXnoNYaYiCld64yRP/Iid2Qyl9VueAQ0iuqFDf1d7f/iXmQzDOLijGZC3tzcd
iOBI26S7wp/AkV3l75FXw2b18XIUr9De/jJyglCPsOtv0xIvOwKi0O03qwHnIg6J7OKSho/I0F6d
nCUe8+pOqxwiGVMJTGpoBgxAkbEUd2tB/QpoE/DmhZ/e17imghvfz5/HQiaCVrg51bGEftC8BBXS
ZT5Nz8OEYkiWmBzuoiQzNIy0uBNazc7Y8QmOhkcHV7FmjmWmR1Kf1r171/KlB628SXP37R0Fct6J
j7Ss5G1W/iuCCrPFwwOJpTlvkXbeRpof+cERIopftxvK1vk0m0PaAg0Z+CZZZPAFruMMVICfcmBX
BVwD6MRdUU18g+6fhZVsZwlVviP8SKiz/QLqVWhcnUpSvXB2slToZo8A2+kp5sCubcZFdGtZDNl8
MxrFxQCqwaISRqiJMqXyzFXkOhwYW/lFPstvr54TnEWQzy9w3AO+te1/5S6heM3f5q+q3jVAE5X8
UX2e1kTCuarL/AiA391LPNzSi5M2gk1pEj9AL+bxmbpkB1cl2UeDnRvfUJC6uxUz11kPts4jsooI
w5/YHmJmjLB9JqREEmAekAz5vFmNLa/sLz70yVBBOBi4VwWeOMO2CP9r0Kr7eIz12Q9iMXtrlgAY
Ud/l1/KzioCGk/EM23abBHw5UfrhfK8mVVgim39m8I7tnMTDymQz7Ki5SXZJbS8yU5ZRXEdpeMiZ
cOYz2WKkMSneMencI11IKSEAMDl/IXpGkItgbi4oiW24+oCNJD+tbm6nK/gqLBdvLJEvPpacXHcI
fQkiloEfd7OcoyrNsAkWV51BPEJ1a7ozb3zNrG2Xf0ElrZCNv4YACchWF7PHW9HzcHcW7t6OvFGV
GOZO+HwswG04wZAvWN/EM3SSPZZ26/c3hITsi+VVdJf794qgZSpQKF4ICZ1aSD/zZdS9OLuSZnhB
pOXC4ykvn2JZoerU1CCso0JtQJcmsdoqRI+Qh8zQoI4ga65LdClegpYslMWMt2ziMw+o3hw/f2O/
J3a/nVuG5SiXXz0NFYP8XjNDJHSk0cdCwwTOtDN8Qcr4+0n/sntLzysrBTdkEq1N0gGFpXrQ6/v0
DcJXMNLv3MfiFsHuR2WgK5d7bgcDfDZ/7DX8WpiSzlYbwoCbYjv3rbQGScYhClI6ElzuSAAT8Od3
v8KEc/qOKmT5anwNRxr5baW0v8N+9yzxWBYaiYSKNBv/sgJ8Ah8S/TtZdB4QbLQ5Pvws3zV112St
RALqjkFqb/4O58CwULH5uqzDAnZaeZwZ4ID/VMI5nTrB5XGSEYDJ8DDvS/qhayPHeM6dCSIV8EDV
sUGjVDNnRMm+5mBbegcnVbRWWkx4oZV2BjkLYM8WmRjxkqFIr3hvc6Z5oVAeE86zAJFKL05pJX49
jW1yO5rgOIUJBe4+yZHcUQXQAL5fcearz1izKH52xIVhIiK+AAKkHwzTNMF0+IVYcqxHhXb7CKVm
5LaBP8QpnzBgBInwnQRX/oAmlOn1NqNXwxffGeXexdPm+QrNb1VDG4ou9FeQWF7rDY//mrE/KvJO
Mz3VFzwmLXlotv8Oan0PAl6EC6s05R+X4ACyULxJ+y0upCKDZathCn/etlPjZ1k44K0L9hYVOtHB
31QUgTYb6KoxrOxiJZ2bpyEriUgwKFr0FA8ieZPtsxZ8zPuW2EcZ8xBzErv46z7DlCBLQAb/1NNe
0OXLlksKWlHmhKquHFSZdlCuZYBoa6EopcVhtTs9LXldlz7I9PFccycNXFw9l7ffOJxfXSNSaJ1z
4lRHf+YmyBj3oGhUmIJ6OZVR9eudWpyNgC9y1ClApz7oKaoyUwohiYMhkpH/2L/PKBmD/a1jdisr
DfV4aNkUg1mSKjXdmk+0a4InkRJGxDrIlgUo9QZcNEdwT6E8cgvvhQCW6bQutNveOvtMquKE+cKT
ZhN+Q2SzwQD1qerIYbWl5A+RS8LB/5rsPEJHjapJsshfRhSJcUeeml9+wk32SVXZZOsN7UiGYMKF
GPO5M1v99K93/8pidurf79lI1Q1ffp96Qm0Xz+h0wqw7KJoLnc0XyVq3tElA/kaiQOK0faCA18+y
UZPhOfnFTkILl08G6R0/bzULaHGlxx7GsOkv7kWlhyvTapOaiUXFjlDDneeKId7j+B3s6AUwTNAX
idAyiZisJNs5t4lEZqahvmN/y4+ulT3zzJ8p8r6dLIKNkk2uvXxX1Fe9mf/BOQBiXkj4RKC5S59P
xHfeh7B4I4n9ZoOwuFrAdXzdMTYg6mJQ6/TopaHbH8HTvXpbyfQeeYdmQ8+bSZUdQM8oPi9WYpjk
83r7JpQ7gOUadzIQZcmKtC9Pw0VKDOZ5Ieqgc4CY4zoKslf/6sMQs9pUTcS4ctb+KJZ81EB3ZPc6
W4d1t3s6QxyGTcPEI7AQF77WVmtQs9HShKNcB4niXx7G2TobW3+Q8fhmOh97+QZ9vivcFi6LTjEE
R/5bFOb+8Adxi4jvrgyQVIA9246vSQ+I8sUIStMEIuW19YdOfolBQAxgnS6I3IahN1ilff3KQv31
9IHkLkvlVfRFIY/8ToAsO4k6HZCEtnrYyJase+PoOeb7M8kuo5qGnanWyeXdD/1Gzxt8KIPPgbwx
2FwcMgeXyvppkBitW5snHMn6DNe+ZVsx8JA7PJ1s0m8set59QuzKBXlAOK1e5Ep+r7uTizYn10dz
grqgooId8tXfNDQSiF68KqvEM8MK4ZtaBxHa9bVYmBXvJsR4TTc2JWCu/y8+3WJEp88MS9fMz8QE
RR1cNFtVbxeYiaSlBpg2P+l5wuyC4nwdpV07yS6trmcIbjFnrKLCHNYAizOQBaqGhBPX2hmPswvO
GBbHlx9Up9K0TzHU0ONg07vtKFiAeQN7boQmzQvBNEYJ5V97DcoCmlY56zQzJpURkjsh9UnYVe88
FSYodDsG5loqTA21X2ZLUTTeXkw8a2GJsKuunaolQZLpzaBMLcsJDY/tc1bV4am5yW7hSVPHIDbW
CBZPOjksIQl4/tVEsImaZXa9LeqiU95jHDBDCxu9LuyhbNXhdJZJolh5XPsLiWItBA4eCnfyCXZr
1xHsJfW1tp+Kj3FakyuKXavTGmPm3v1JhWUK/h8DRkrb6BeUpgC3h6AysnX6rfR6x/WMqWP4jm6+
c5fngyIQUAjXmpgeLLe3N3vZ098vHQ67EgJkc6QV1ZFRICC7aDdmVY89NU8pbfDr4I4I3WWpAuU5
Qv3iDrGK4Crq+cU7cuYeAzpIxQ6OQMC+6ULa1IwhdPA6i6bIoQ0vUt3Cj5Yn8nMQdf7qfo98MlMQ
DOZRZzr9SrpXjozkdI1UvTjAHNcPHJwz9fN0Vrah4etg2ffP9hqaSXgkM9zKOangFQ+09Yik5ajw
aRZkx0s3kVDeQJligWoavPdAFlVvR9mceezDQt0umNqVyqDy5LUWjdHSogoVfxNYWwhaDkFP+gSr
f+FL2oU4PPGs4OP2GV2A4jfGl7RlSEzq5qRcmZpA86R8DPTRu0OTJKreRXU/kPI8JKcd42npwmnv
4zEowSPtzLWDEK8zR0d9/1TZczStqCUuBcG4BQVpu6/8SiuRLs7VuJSCOJTDM6kTA+h4Yc/RR3hk
EL86vIa1EVlwyltrK0lt7953vszWyi4EudA8q1eQdILXJS25meN38cXvqr1wEAT2qYOWxEl2WeAo
wSAMGTrjZTgtJWsgIm25GCw1nBHQa3Rt5MzJwcnRUORay00z1kctkCfPXb+rko+bSWKpUlgjlMVR
2cpU/c/piB/Rhu7JkdtSfLaEG1LuzAK9WjwvRlFXK23DBRp2mZ35qTn2XjDN1JPienGDr9vWvZVN
OzRMnJXmWhmaq9SvFZp6MATebtoigceOCDzMdgVAn4ZYcdrGh9MOWWFbdwgB/hrTW0gSjvfeliE0
cOSMxi7b39OTQttlWqE/Ghg7eVF2iQVpoI4zm2p9I9sFvAGFAv8XOM4ZYQlX5Orr1F0krR9TT7Wz
oclz0TCsk8Z6mE6WHUARgG8BThO/mw0CU8BrjCqq5N09L7JgTHDysaPiLm2lbfcIA/CQHadJhacS
7FH05AnOADJteDefpoEh65RP0A3bUv9Xn/udZQ7fba5vO/BjDBmX5E9LzFzT+yWp5H1Xoxwngz9w
e3N8WX1AeSLd7G9xyMYbs6UjkEdy4f4yKaPVTcnxBscRINBD5ghO7ORlPalPYrGOkH+yEA0SmEih
JXK5E0cwclvg//WDpg8XAwPU6QJgLM7gSwZarvWQ1kUOEJGpCh3ogSTIa0Z69SkRbltMkCaLWZGO
bQJG00IXmCoDLmhMB8Wp3t8zx7MLBrRxLv7O4/OE87Aelf5r311hivsp1bhm1H6xmdSR0b6p0Zda
C8/bJVDtN7M4Au7EEk6kUcltIHintBGg8gVmx3xRw9uy3mpD8zKlPPYc37CeY7bYrQ+tInGvICFV
1QIMDPh0n5WsO4pkh2B7Kq9bUcrJxxmqPy09sDCOmv2wNkSGkBFh5PsWfUJjFI/Skq7nA5NnmtpB
Db+GCY0+ogY84mdIxkanggd1ASnesSKOYbPoGt4Pi7tDO8YXk9ADPY6yyKUtevQB66h3OmQxhYcU
f2gXAvmpLkuLhZuO01diml5AIJ+qB6Wzdd+3KPFu77NcQgJWx7CBrP1BLHHPcalE/0MdKPcJdSg0
M7NcW7UJzhz1S6Ig+r1/4/GvvMQLyQ6lzyeOXUsI/Qg7qi97vT2gWNUoWvYj7n5tu3hqKKC5M1MM
5r/bDDoTp8a85I+nnd1j6b2qk5CK4ZLdTfRIDMtGj6Tv/TaxrdKa4zIDieLtcTQWIeZ8NchHhnUs
A3vCg66b7erZ2zEZm83p87WtY2soIqZxC+A64KR86sXH1DDb69JJOJR5GY59/7AGs1v0gntYJuxQ
BSnUdYugSz+lFz+Xif0pACLoQhJW7lV4IYyC5P3KcnhZChQmBtw4zVDzDRqhAgDvmeS9yf2an+O4
B9oqldH16Esx20ZL+vmQ8gBFZKJtUhzW8kF7V5EI2llM4RnwpuJd8YxniT0xslsvT9uhmlJBmivJ
txMKdCz+Hcrhm0ZTaKNaK5or1yd45FtxoqR4+dXq7g+CSMZ2n7VMZ6GsJQMQ446xZZuxKb9hAWMx
lCU5nmYp0sZJW2C7T+hrcUU3EIoNa8JRLDWcCO2RNiCybrmuUzPuE+hfwVWDFxQP6NhM8h1nAcz3
g2U98tEwMVtqdAx5JUU9o/8x02WX+Rx+w1KzAvTsc/yYJMid8x18togXqBNLq3zI8RrpVXI3jI+Z
dSZ7qe5dxmjp/JzFjwneVxafO/4VgEL3FnMYw8RJ2H+GwZlebLatmx+MFlCfWYf4+pCJ57mnv2xI
UhhVzk7BwPt+lWgv0BrowcsmNB9V5LBqZZKmAfoHU1UsU3CR8XlC+e3Wv2j5cVK8XeIYmmtwwydu
dzyAPktsUBjHrMlWud7YGYygS0xugWEjpWW8oEp3oOeCcnchZV52aLg7jVT86OibpR2OGRTWHTfh
NR6ZBnmzZgvyaQCrKP/T4W2YYXXGwV9wIrnnjUK8zWh/qJj7YxQY0dbEXEqtz4Qp6NbxWT0ilP5A
AD+ve75sNJkWxYBCYmNnDpSLS0m+3ArBwbHIMLff6ipagmp8DGd+PV7WL9Mmo1mVH7cR88ekH6Vh
x4bzGEoIlxvNzgNkwrh1C24ThTu9S5hH012M5EFXSOhydYAQrLL0uwiDDSXW0LwvZYbPjQ2TiKJ4
GPVgmBo1CIHexPRVjY7mLxLtTa1zlm4hOc+oH9o9pSxLAYj4Ea2Uz+oYStuFT6F+MsRstrBTkCzF
SOrvkccjuYFXTZV5XJnZAGI6pf0XaMovDcd3nmbmlFgC9T0LuIu7K6WvOVFNvoGR2Ak1weYU2f3m
4cvyQIm3jGXltoCttmFvgd9Fl7yVqFXEaIYPpKvA/2TrAE/A3lasHVhuKcSDQqyXwVxSeFReUedb
glvBZYpHZq0ctvdxliiJqPubfLw6PT3PpgoQMW/E8/O3ZNUChhoH+TWi2UbNFtjp4Wg1AmNfrVRH
tTz7jCCllW6rcpOgIjDZrJAHFPv4sSHUiyknPNZUFNCJl3T0lJVF7v7D0mK61UrXo33KjyA+AQAV
8OtBK0Li1+85T1GW25BuUIrB8UyS4HBH2A/T24MPlLLcpQKTQhJUG3YdeGwlxrez5oaAE/jGHwk3
ps7psVJ8h4JPeZF8fpr1I/GpbiYVF23LwxrfjJf59GpdWgflzoSQoMxvpoA4W0GKCzBMZ3scs4+G
s2wRRiabdLUjqhUQSKGv5N2JP3wBK1vZaHeDDu1PvKUxXEjk/P+2uJbNBOfnXS0xgtVbSq++3aew
2OIxwYhmhmX341beqs9u1oUHKUh7xvfR1AwVwqgqQgpRCbvMXULe8F1raooZRkPFrTe7OBvqyZZR
nVO1fNBXJ9mOhGJNKlfjQcauxQK7k+iUkcryPgXm8IMkmqzHhoIMhM7BDZtvgvYJp9AxhFXgiGWR
G1gc68W4vJddUsACMgnrm57MacMddCg+fXC3XB/XxFci1NSyRTCIlDIA2cnTQs6K2bEQR6AxzB3v
2nt/P1WU6WO3o7buOvoPy92cPUKpCWatA+eFBgaAA0kS9vPxFo102IQDcJlLarNwzSdb+aLx4+Qt
5BUf28El5EitgID7MT3TxjuSC7Hqb27qyXSfOGZ4rBANZlIwyTXye6V3iGgx2bsHhsEBcdhN3woz
jI784d+kb+rN8AJxl54wlsWPaBu6y9QOLRwV84SHF/Gj5CxH4VLTEJUUMtyNOIaFX1PeZoi/x4ov
EP+m9HBKtyTNZ31YEI2crcyKBN0hnispXAgL6xCc+nGghScyVZvgHBu9/UZvp38w68x7T10OlJk7
CIdY7oEqvyGVYRCOsqPAPwZxcwFTwKlHAXKLCBG7oB5RpsBs0r8A0m5se+tO61RgGMtbOtf2BbiK
O/Rn1qfWP/KFg8Ab3mkr/UllfyCBQPn3l0tZtyBZ3IovVQTqdIKXW3xhx5lF7QFKM4kYcX28jC6t
SbPRv2UAfLR359+JsPzNE9qbD14bDZCi7NKJDb/nI5bPPhvZNakcEu/ejOQ976jG/fmCFOAuzRWs
YE7H31DNtHRAc1pMGPJW/m3bqguIRHSBGbmzVkeP+7VrE9YGnrwyVzPpoxqWkBxlYspzQz6cR6nu
wpyda3dO+14RALZq+9GtU+azR0S9gCQcZcsRC4IshE71hGMMHFKhMWE8k0SpvVBnJ4KWLhDzwg+e
dQAGxShSErdyphey5C31OAjwVN4i+OG+N/BN023ZntOZHA89156EqiKmK88LSLrMGOd4rVvZ3B7b
9uMAKTzQlRaAsCr70L/aI0QrjUbFfyGEjqu6keZl2ZkQn+B0KxdMiE8GZIzZBW+gNE2vTvD73YTo
pl9LVvbb14LvdIT8C2p2M90+K3JgEH+RVxes8teI81i2Xpe2ntxfiuDzuIboQSjAHAP3ueBjrS1o
N1KxpkCAySsBMQpBVbVouXJBipxoYP05DZsJZewIw3BVuCsGlioCG4sMBAlNLcFFzfB4G/RQNZo8
wMBhZuAhwe/UXAqYR12GdltAyKmJTzM5eRrrCfYB4JQmcjVnjUOHrydgqndDb5Prwxw/v8G184cN
lcjFpm22c8WFf2oIHRR+GDPq3pYirDjqgHSGYnA0Fv/SK5RodBqeAXYICHbqUR676634jShbmxWB
GJxlEx4hFKHv81qv66/SUqWCDhRCiw9TK5E5J6AL/BkMjY62JNflcRhWx8vfnIXF6mp0RMryNYR2
sbSmqT9VEzGTUySVt26vfnDcwqAFUG/max9744sJPTY3r/5uu0s4nIasN2Pgd+MdQ/3F6ZLa+2dB
lE2wcll1X4Ls8UnbzJA2pJCggiTAop631fXqAdZQpubESPWnu9huP9Ff+E3zsKxcagaRE2MTJQnz
EU4gCdbU6TZ0bfzEH7AzLyAgOwqc3Rp2DTL8m5UMebO0M5YXYQ6tryr/9zu2evnWwR0Vgk4rZzhZ
F7ziOXE57i8J0doI3n/+A6RXxrHAvv4tJawp3KT/WNsnsJtJyrT5PSZuoNd70MiQbVPo3CJtQG2h
BRtQCVExhr135xV4dAtVDMlYi6TSxdmnVIt/LhXNLycL7H4lLFdi4J+JtFnZdOr45DXZvEawxkW4
ZhsnSlebxTE6pPMeehSTdHntEx47mwkChumL5D7muEQzf3XF2nvi7gv/A1zszBwKpLc/bwIFm6xb
jrVRHBtMts4Y62Y4XhwLMIk5IvMozKi544jRmi13GTKuBFXa58SpnMlF/6hgSXlMva0G6hBMzuMb
3IzC/SHxJgqrvWJBK0UfTfEVF4nMPbmRLctuOPAP0TqIK81QBztbxub/jDxcNqR6REia7bls7a6I
sAeQtqCBkieJgXCCAf9RssEcV3IfJXjLDIoF5RKmyPm+5kRVy+uKr1ueEnrDCZXIOLDlTbZEb6bY
9R18kyVGMuPlZLx7w7IeQ9pIoTlGtxugG9twrzJqOrIj7alYCZdI4KOEhm/jEBnFHgmHyd+6e/3i
OND8JdhGKaGTy8C1S2OsrFC0Vm1OX0iVdpPsvVSjVESv+c3wzZL1+sVGVqWDvyeZCa2cPD8qAtl7
MiV453FnXGcoGMtUSWzIIW0oTrkAnnhBgOzJ9uzC4/vWzFuXsxUh2dcc9Vn/m+NuqK30awf0hoP9
ViX0UdgqcsoJpZpuni26ehHV+/N6aSzBnUb8VsnrnNo1Q8SxJI16CLkkale3ZpvlBp3N2BEORah8
pYI4LTntS0GZPHvgbYnAZNX7RtzlG0XyRDyhOQI7LEew8GTvFJCEDavkbvvVLLOMC5iksxCS86US
ojBKQj/3sG5Gxx2OUxsryg1sUMWpnDQlOxSkBHrTIEwDWxKf7han6pbeH/VZNzV8TW804LygBmvv
pbVrk6rVMWsovlxGcrdyZtaswdB2meg0ke/CIkR9PFG2+GAVp2OCCIjb62zGuJYEftAGIipLZBFn
6kj89oEdKia1ZVCvToN7tmM6KefN53gdF62f0akV4O9YWma+06qJMEhyqv88gyBC0QynxPgW/ssZ
5OWKn8PJBI7I8uXt+C0eI12N0R+AXMoudduUqIohRzdxeYALQB8tfP5VqlLXRVB7qRWuiQ+ByycY
ICnbrCbhB0nWksZVGvItjIah7AmrZRtmhWZ1DbQ9L2GppiBcEu/AaH5v0qKuNNi51cm5JGfYMrl5
f6Z6Ni5J0gkgrjAeY2a0zhEloDrW2mVeE9KeHol4S1hKKUH4deuKBJfXKftSwYdcZ5HGUbuQNcTf
lMsWyXqEyS619n8q+yhheAKSgREjwakfvHg2o2BGOpjdcSPUX6yo8AoJ9yTE1mrxi4n7uy3AcXM6
ua609Wf5+MFdOClCkGq5jFP/th6Vunds76/wGNHrPD7Xn/ITGVvtUO7nB0WnTuXt2FLavQla3HLV
1Yni8oZgUg4Gffacw++xNQT+mvmgXkbXYpIddr7Ar1p2tYbz/lwn4o2bWR6NExD0TZZZ3AShya1h
5XDF1ymAb94X7ugObdDt5+VuQu6zQPb6FCfszq2dlWYiJ9n9qLzaJgg8+dcxHhJ80nkl8UhLoZzN
i0UiyH/0yaqfZh9SRwCKmBa1FskkJKIMX9TuoGv2zgaklPUJ6BCgUYN8gfW1/UOIYD5sP+MxOEAh
UZfKQvrxeZHfHSYBdwn7/EWAWQvYqc4Orv+zTiyxHVMn9Sh1ryqiFNBo9EIQlQI9rBrGz3FOWGk5
KB4RUGaSJDfCujueBFO3Ggb1P9X12i1xNWpE7zkkOO9ukVGbuVVlDjta/fqzQZFHQkK0lBSgvVUv
f0vQovgCgSu1Hoh8AhW2ZQ69WbhqCCOo3CGIqcoMetqeUTjrQt+4KqBmK/7eeYf8SWHLPCIu9xOt
HF7bwwzfDNFX7a1bGGZKaORsFYzzaZeyWdoNCUQM4wWKdcrKN0QH3f4pmqJC/TGbSRPz/MkY6tkc
qW0dWIXgtWUY38bm54GQJtsDaf5olxE4YtsdlEDOxzEx4r79igSnFkVKBS7/Log/sQlaIRBxmd3F
C2bZqD39++SczwlrmF2RR2G8HddarbpSPttYIHHkCqFWy1Oy8gWzrgKyr1fAPTgA0ngpx+clWTMQ
bsIDFQkhnj4T1Ebd1O4hq+//EIDw3b2kjN3IbglZuABTheiYr1LqsEUeoB8YYUDLbkwFY4vL1yZ3
NF1Jcha3RMr6bMoI7RduRA9y03v2/POR+XuCTP/zJf5tChFMibS3c19m6EKo4Vq+dGYEoBg2dmXA
t6VgsCFS3kfE2EiJHZ/DfI9kx7hec4Kh8hwVRq8lIq7MQmmjdGhSfCL9Q2GtCE72rQlEZ7Jt7qit
050AEAoN/zxLwWNJYEKiHSSAP/3jryyL/z8TjKB+K+lZ/XwMjEstr+NhWMJnH+A4iOT1S2QAi89S
fi1rMO9fQy5fzwheb1kspa3AmMZoU6k29JTKssl/V6s7GUrqh56Vlxz5kMLPzbyDkJzFNT2cGDYi
nOFTRvtr/eO+DOQXDVHfHFpk2sRYYn9btOy5iclaKxzmBRyVkIaPnujNl5RIi7Rgc2sy2gcYRuk8
HzHaofKahu8dSZw2Kiy/jv8xo3k5OhqNJLoDOfQIdwMaHSxK2uK39VPz36zAdoMdEuV7gziA9q/z
1FLtzA6POaQfmsEIIHvqE4oqPoQto2r1OrH/Z5AyCScJbvvwB5dTf3TGCkfT2/veg4+021l+tMor
bTgoU2mPINVqIJaPI9BsGUUjC+FNRGoMu11J32ZGVwlNDgWmrIOl8SSPGDmLRmjlWef8BA9My+p0
sT1X3MMuXsLqkHyLD5tqsfWxo4vGExnvfSNkIjlbDUJw7BIq/X7OETZxve6CxTGGmk53aUlayIUb
rpVcgNhcz34130i7gP5mDqds3P1eZV7migNqOgpFdjArGTDKEf0vD+wuSBZu/jerkHKiXOaoTvPw
HATezG1F83TB7onvc8fjcfnlQoeQfHLX2zG0zwFcSY6NaeM6oERheNOUU2l+fDmbBAj0jfYN9yyR
+XQCzJL+rezqa/i9ucXwUZed4BUcvrorrVyWF+ljLsfwYmJcJBXcpMbvCqtUwVVmpuo1pPq+0y4g
uhRUGzM8ADWkESMLZ8lE7Kv3JcJZCcXhQQvSQsXqLliE4czrqBot+c6daQpPWpNxIefzvO11n0iA
c5PaR9kQw+FdSElFGKAEwCmiVYR5FbWipzGI4OtFRHY/FVGrrlqRx6F6o38ikPiqn/06eDExe+iB
aUJa8BOsb8FLfaXPfGknlQ2CjmrYYia6kGBGPRPqkdK9nCxKJ75QkLAu3xYsNRDZEtTc/4m2smfa
PeMiephSrBiTylNrFCg8HF2qYw/bgRISBrCXp91NbRD7qcETlhLql1gNlpjW8WVKgee0b01ZeZbK
vLzkL3OquE2FXtmsZ/1ZDRKy6IGvpJAI1+cQ0VFuZN/tTNwWyrsxwLJiLr4FX/tcrn0ojSEea6l+
ZLQHNk4i6sX9aJCo/bjeTvA1nUAW+4t8w0p3Mngrji6ZKQSiLfYd/JH+nEC00W65yFjK57Ha+yv+
Watcyu1uCcKlgfsUUEg4M8oYFzou81fw3wOoFKLAsdRz5gAOcEDIhvRVcmK1kZClvpQ72t3fUo5n
7VJiRj5LBXKCrmgUP0DUBqtX94G5vYzgIJOl4RCO+IrmCkIGvkCow6YXY4zLSW4OQcI/UBD5oAaR
KL/IsSvYR2atRmNA7UJ3SVysaDIE/pUvIgBbBRKK11A+3EqL7oF2XAQGLrXtJuEAYoM+9eWMsF+q
mWvSTBuyR2G/Vm2F6Bhc3VKuvqcD/HH9hDXFLku2PN7CPS34hkYyarsX4p6LjpYO3v/Zxso5jbs4
opmszidlYszHTBUsc3mzakV943sMkC6wEftv+YqikQThykftlwZcbcMAb28IMOa/MVlNjjaVTsTA
r9gZtcUIfDug4yU7sq7O8H7D4IdvZqfyoWrTKrJ4JOkSQzXPfRwf/Ak+yzcfpgyRfY2/0APpHhm1
UZw7KuxPZQaJioOtQ7n6/fzfKPWowJtZ+VATJW6rlWIMQR4Lt65ZYHp8PcAdSuLPpAUyCQXvVEzy
ii0XOePZXxAbiBltOE7cpb4/n4UNbPdY30eoywF46o4rKcLmsUnylAKL0Xgl0FGOjecSCpwUQKaP
h+t13iKcnJSq+RBuDCrccOyiHJ/StnWkMpXe3aMlwcAiDIQgOs5QOhjVQbxRqufPOmiZ+q/vfygW
+xYdAX2TWUecYgXjADBqe+ARlAoj/nXFKFxvE/6iBK1SyPpTst2FiBFS7SQAWs+WKHsFSF6RjuhB
QW9LUgEwFZc87YvU6yOe9cTjmxDNX/Al7qxe+oqoLzF32d23lmDWI+0OV8lB5RC1K2BJIZ6/BwuC
gzhJHNvactD7m9h/PzeS85CY6SZ+D4wbXh4UBySdW6szyrcgzzoYY1I19g3lhkEQ7RL1SOaIMNqd
UKVcGczLC28DChGRm7ky5Fdhu9Y3jtt8/4HanDTGRC1CjgAD4bK7kXNHGyL3E7sGvGg9coi2Pl13
ytjCtius647Z1oG3qBa7QJWSPq4NoMmxYZWh1+7VXPeQvr56vgP/9vF8D2DYN97iy4hNNF8uYzYb
KNT/pBAg1bDsilqnY4fMaDU7wfuLNtjG4tkifWc5t4UysEwIW2bH7UcLLwMHNQ3rJ2GLyI7uMWu2
BOK/pRnBeaFs2WeOjMGu4PU7BgD3T5m6Zg7Qna4BOjvL0NBEwddTjscxlz12PLEm32Kte8c98zBv
XisLQU/LQJtzrWJfpBwnR1BLeMEA6HOS/VXy/LnBACCQi3z4j8Cpj7ms2LVUxZy7edX8j9wzP5iT
+gYbGXJbVaI7CkRAWkw1zQ/oPDphiCo6hHh63k+4qt0tjgtWeD6u3wiZYlheUIfwSt6fjG/bH0tZ
09a3wEC1H6ym05+QmGuDGgg0ti4zh7GXAclKl1quo6zbU3VDGGIrgrG+eIVeLWj/r+CVRg3BuyCz
8kvjtqKp7V6trU+RYqbLlW/NsHaoRhSVM38DyNkvbM7V5Ds+5409Petydxt3U7cJiFZeRmGq4fL/
CRNfyzFwePB5weqaOtxhgI/t7KVJ51N3WDGrfRkeFWLmceoksxci3yXzsvRHTHpeUoJ0c0Ce6W63
xAqJlFndz0qi3KdGvceySqLq2cKP24FJwJoDLBvkwinEjfe1H7UlDlZkM4LpX4cLQ6grJkkMeIPd
WuAiwrwnt7zsU9hP/bFnoF6wltIbTgUoEoN8ASm/U/b8BBMMrVM438s/tCz8TbDRtiLxgrEnEAnC
sf+AiAlfFhqhkSNcnJg4Uh4pM+gfGnfQH4nT8nPU3nrC1g8xP08JTALivYBLejO59yx5wx1FuRos
mExRSP4ZXQBH8KabP9eUzZOdjfjqUFf3C5tXH3HAjAGHk21XvM49sSG+D6IC9Y+0RuiFAdDCIRsY
2UneBRQIwHX1FkKla6l9z9JFtFPd75R5mgiY3Uoa05OzhJB3fArv9Ww7RS351Il2C7b6W3ZWaMWN
JFe//+QtS2REHrxy1BBuqNrJCylLgP90DzgCvsZo+mt/kGrvK9uY10H5X2ksGnIJW78fYYj6trAu
ATiIUq+xOuxDMp96VTJlYkAkNlPn5jqHJ7Yqr3up3g1T8oMorEdk5pDO03sHGt3AKNn0GyxopYiP
1ubscwnojEPFfSG4h32MrPunC0W7vAZFMfazk8GiVx8dBQTYEGApp/xfBaG0BVSVTE/YEnVnN9WC
rIkBVC1sIBIHccwHeR19Tj8fWJjhRBFrTm+YpefxQY1bt2LxeHHmt198/n0BGJtUJox4yl09UxRr
OkLbSnRbJN5UvKRWGlhwG/2NLSDQV3gSH/m+wgBGwHHXRCoiWwNuZ9kdukX8ZkjEzVWg2uiol64M
Lq8S/ijsI7PF6WzX7Mwue9gvyaKb4pB6BtN6nTDDoD0Ui5BjN94Ldnwg3zWI0HdecoE6TqOP0LTr
7SPGh4SOQj7OmMczo4n5IW5+90znCp2sWfutx9pN6FJ9RKiZquzW7tvfgN5k33QqQTnXJ7zLxuYt
rEiJBW2y95LZW/swZ83O9lUC2cSbsYXA4BPvQDI6/RLcbgCqDyxil/AmuRBdiqAZuXQm7WkOpKHW
mMvJHHD/9RPl39UGDbW62vFnNn9wPT4C27POwLqnOAE2bg1/vquP0OfSjUi+cy1sE/U0eR6PuMeI
eIfktsAm+RytrpsIbR10dTaft+R5I/XjR4TTEQBGg/xAbJ3jgS1kQHdhpLg0Tkdxc+m3r3G6iEd7
PyD2f/QV/opvzQr4vaxVpDsuO0+2ePKoGScs6MycYtx7nQddPDIxzIOWBQEukCQmKNije0jGIqf3
A5+RxGYYDZij5IxxOWPCY/Y/mzOsdLBB9wqoS1AC7pVUR28OlW6+XvgPEY425YDYpoUujbsR8eEV
5UhpatoryP58S5J2DURUMOINyFf+lJN80M/ZRNXTAocnGqk93QfU5cK9DRQvmjiOixskxR/ESuby
1+qpWxMnFmix/CYZg3B/ejZaLCwAefeYugs4qN0s2YeTilJUqTu+XnxqMrOe2F4OviFyDKyuvJ7+
s+s1g1NgOdt1k/xGROT+OIhp7kNiFeBgnV1yzMXveNuhsAN9JlIXy0lm8Q4ixgSuax3pqx2quxzw
MqhklwxGqrfKvFkmuTOKDnTDiRAgN+PAjoKnshi9vosVtSq/ELtbDZmu/fCdpOTI5UZg5FoLubXd
xXCEETB6pcFfAh5hNveORy51Ryxfo202lAcJNYMh9oLAubi8yK8NXfncZIcK7N85SvTcJI1sX5Zd
x8Q/Iqa8o5V95VqnFqIuQuxBUuVBkKlo6ry738aGfuqtvq7MXo6FR6IPxdji3C+tYNS0noRdjEB4
PgQeD6iAHSPNEx2g+jRG8eifFUEd+hvBd2v+vQeOIP4QQo9auWBGyVihjYrevDVoJFSAkmwj+Bn7
JVo3AyiXcwlDCMdsP5hNsFhh4GhcaGgmhrAYInrNT73e27Pl99v5uIO+xtHkgCQR9CiBsBJl/j8v
HzobIRd77DnTgfio+V+pMk3XPUomQtVTv9YUK/UQYNjMvifBmxYXGGh2IV+GmTnU031Gbp+eveO3
HUdlG5KMHl57TqHcF8WgZLLEpoY7/eKv1t5Uvy+Ldjqq6CvacgxwPqfGFy0EW8pxI8gdz+3ZrQHA
+VQ5qi9rRu+4hxPabxdgMut/ruqnPjJTZ5nYrJKYaarMawBsVwhJ/j0LJP57rZTFz4Kb0fqRGOpz
GGrVIPwAWEoynBZ4SBpDHkH8CF/KiLOK5vNLej4SOvlE3JxaSGTPLEAnUajrm2S2iy8Po1jLZIUP
k2mu7kTqvexs7KfJxAw2RWOYS8mjqOtQYHA20U+M56D8occbV9+SWMzq/ezsRfekYaeVayrz7oxV
Hp1winPxdSgZa1BsStKudknPs5izGnPZa8QlKTxo97xUSD/lV2AYzcOEuGdnquIOjaEIm7KRdHiT
dZfLwAeR369GDfCM8pC0Wx54wndVG/Zyr0jMYLblX/RbXXjO8HRYRqnFscuD49YOiKS6qup4YeeW
v21V507UkCEk7pe0PBtm9qoZk6VrH7vHfskiFuJOoS97aTZNzH2ZfMTibsEEk7cvGtIPKo67uXR4
1kU9qhrfarG9MscsL1q/aNKEgPBW2nvMuioqKGGsxnFJla4n8Q7Wl3pulWQ57ohm01FZSzFW+9Eo
J+NT30H5fLEhAo4l/82rJxyDDBIXhVmJH8HW6hQcpnTrEzBVVOYJz9qzatg7lQJJRi80aGHAEa8i
k0lzOh9emYNBWSAyAK37/lY0bEyiK0NrQuGUTGNKV4pKS5Rxc1+ArhCsVI0QnMT0rdhLh88dJQ0a
1lZQ4D6AxGN8Y1uuIuUr76fY6A718HZa36YmcpbMlSRcxX4ikAMaqku0/3YQxCfSbcyw4VgjV6mY
sjpfYQZBPicy20AWAy2bFC8dVhZ5s9hnCHmitJ+WA9CqRKoyFVjCujj0cfXD17L0iQjRHz1Okkkw
4MmltqxXfLqKbRK12s03sUWQGtfYnJWlDVik1W6mACigS1sLYmYEHaXm8sFRWk70duDoIfRaHa+D
xpWgW6U/xw465tIc1cntzGDNaHmxHYjWz2kKHnfXNWHtIpdofWsmXTNNO4EbfAyvYNXAd4gOpO0N
vjp1G9B+QrDf1anyvaocZwThrmQsRMCsQ7ZUlKDHR1MdxKmPKV2ws0PgUpgAseuL1vKLjLTaxHqP
s8oJ1zgCSpraTeOlvFo6CuM9q3ycMzx0Yj2A3ur920A8z/TSwoRBfKAbtY0rNYtKXu9vRl0X2Y1W
WDHgfSns2lbN7QIp0fvEBHR0vb04noSVmxZARl1Qb63py5pxt2QP8yMmiAdanKjPwXBCHBZqhZQe
hVILPEe93RpqWWZ9aQ7IKEWN2YG9d0Yu5iMvkN66ybZ0AsGeQ+H7xuhpLjgP7zAPjtKMe5aD0JHG
UEER/M7OUtd5T2LccPOr2qjdvopE35o1Rr7ei2wI/SiRukEA2bgFJ9p2tinW4fP3HdmiODz1lEM+
nT1aHxNarm8vU1zcZxfPPZj+47VA61tDrsbvybLdroYgkUNcJtm2HfNFfrIKs4gdEqXhu/cQ7Q3e
N0FYbsFLZcOKLFvCPyfISafDCiil2TUG7cDOJuqS71p5K7kBsoTIe72tB7DQZnXZJADr0veBpr64
7H+o6JetWfMPTdoZDO3T/+c4l+o85O00HohoUjoTyFODbvk4fNJ62VDbmlRq2JAmbuDgeYPFjGwO
UC2/hAIi4yGWMCqhnDIgXdVAAyXizdcL8xtfJh1VmVvKf31eqkXMqVblWD1B7m2b8RaZiavB8V+V
CnSkUkC/OXgtCgGF9QyI7JiWSO+mUv989GFp19cj5BBg44sZIP9u+a5z3DGrWLLLQ+Pf7yZV9cmi
vuuR33qqNpcVPyak+OPIoTw0lyzocoqcIp0+R67fmwf+5a0mWt5JCclnm4wuw4pFCFzxrfzKpYyD
FTARQNFk3drR1OzyIieMM75ntzLY3+iiCMrLWxXdCFUOICqgy0y1yysSHjrOiqeJD5JhO0ZEsfXK
J/Pnyo+4FjzlU1bNIVo9mn5jN6ZpKPtFNvtPbpiMlT/CpLSUiUssxA2TKk4EJOn32/gPmOQKE6xS
HWkmcBVGOVfzw55UDv6gzBSzL2aBB2Zi4KjSlo/CR96hOaSOE0hwRLpBjyjbXK2YHc7VjB/WBQEF
c8SLIBymkDUgV+icYVbxTXVYMUAUd5JrK1FYNxaOoAgCyATcuemiQnxiuj03XKihdBPK0kzmT7zI
GngDbKLQlEvaCsNt0OF1H1ClrQP1jd8omLVuEp4Lkgl3UP0OZD93u/TNoj+JjgM1kSHeePj89RTt
QnUxf1Pi9c1AimKBKvdkC6WcBAH+GwQ/2mSzTiXSUoUVI1HP51iZ/EyNAxtqwf92v55m67eazG8T
S5AaaecZMvHKrMC60ZjwpPQCR6V1qgcKu+JjG4Z8wTUNjogRbCXSWBtGjJwIW7Uj3f2vx2UsJAhX
w2rs9jB0+eatVZRXjA1/sM5e9pDmidAOK31BC2J3QZNfhkE/pmrwUjcGuzr2RN0DedSAd15lTMkp
aS5spoo0L3W+DFltj34cz4UJ2Vptg/cVGlI3trMo2MBK8mokFp0LWYLxOK7am/WPwo2TugeFYp/O
k+fGWTQXMjinB2YI2tnASGC4VjnPZ4USxjbX6eV9bWV1tP0G6C/LzCGd1kAby3l+VDoLejhJig7B
cBaMyvfeiiUFM0pq8TOeS4lfldQGM49E/siQuLX7oMGsrnT7Tz8sDpk9iNPXllayIABZooeJpnMg
aowUZyx/4E1IpgCWhX87faCyBVUF6GOICE7qamlVwyrYiqn11wUtLCgNGSQscXFO6qS/ky/vSHi8
8wjOLsf4BNkD4p6k20SU8knfGSXnCbkj7U+Qsl2UJtnRO7NnJt+ugdw7lbEaN0F89uCeQJQH4z7u
TVRUlLDH/Lo8rBDuBEqe9AbVI8HvUe+v18XK0qwRltRFNAowxzTHoCWvQkvYH48nd2rkrHYMCnej
SZIYjSIGTa8m2VfGFNKUmjnmTEL7CG0NjGZ496C1OgCSSvjw1wuqsoGatV8BqKf8drA4RtS2A4K+
eKXWOffIpbz71AnI/L7YCOmgpJGf4yVTTgSrECmR1uy2NkH9+oxJWYeCb9SdF2CUudeBxcirDRBT
9f8w9PoWxglqDsWGOB/b/+lzexAHQxEerF8fFPwNZQ1q8njGKqeGaXAZm1d2JdfMimwvVtjliv6R
af+EKGUqO3a2BCyaHwm7GTh/4Faj70sNvWy7sMjLZayVxttgYCGL+CycddZ3CqLSKrUA15LvZswN
8k288Oo41viJUQj6ZmIK9xtErJmOwgw26mxH5CQFACpeSF0ErH2BVqJryFoBH5/4K6HqYna9m1ko
yKYRmzw2yvDe1+8qX/IjNu+exk58TInxEsw6Qn5/x5wvjI4RvuKAzlqOWMfSPh2w3DATOT9yN4ey
7K8AD/gqlle8xBsYlY3gpBwFw5PQLP9cRFh0jSXwoH+tnRlVt5X5B5th1FOsj3Qu8ElBU7Yfx+Yr
gJO9QqFpWv+YdPQltV7VuP+D9qIVqlkh/V5MGoOUyejmCWz6d3wj9u0WdcsklNsSTAJ12Q1PgP5I
gtsrB4TI48klvkQ3Q9bcv4MQsOHIBe8qQ9u7iwFdSqZ98vviP1IqKKzpf0bvXl7yJnzmGZ7RSEwR
/JesNPgXJ9w6hbbjhRsvNPqCN4WfY+86jp+nn98aifSqXJDIM1KyGpfdVM9unTV0gisCF8aVAvZD
T5PnxNKcV7jKo4Fq8Mog5dOR7idMZGLU6Was4TTk9uuYMW+pCg+ioJAvm/8lg2js/hvktkKe2HmS
dKBb6hAQPjJJnme5w1j3sXQOjMx5GW1eo0tH5UhGAfPBOztSHX9nxQdwpwgRfOaAxe8vp4AakvZ3
dZJZ8cjS6A+lvKDuNCbrD++6gi4QYk9og3iF8WrLmD7dA3rxs3Gr2YYuYvE6M4rOq0xt6EdZlsdk
uxNKDWerfYNuJRAxafhfV9BLd8ByLHwzu0J6j6W1x/6LaU2EzOAmOPzj1/m3nSDnNK4XqADQttXc
04brXwhoygZxWB8ZxeekUWGFBUewpKoqyaElbUSCFofIEx3uRyhrmRFZ57HJSD0pjb7DkjWXMjke
RbAWa2e0ywKjthCn+uCdJpV6uRVftyvBSpiGRc7cGfI4s/f/tVOP+AaROm0X+tALlpoQNRN7wj+k
WX3MJhQplzp3Fp8qT7TfFmvcU2ql+ySQyME4/rmQMtp3duJMrrg8F5E7+Rqxl2dlSuqmGtpQoP/9
pQIsFioJH8/twZP9tmlWkvKQmZ7LWk4Dbw3+N8FQ9Q49SR4VjanmmETc3bObHUAea/3gBbyH9689
jhhj8MEo4k7RHhBDSNh7p731TV+Gl+GO0Rjtx6TF3Z6xAAsD4OhyrzSV70LTK63/POmSiDqWRIIQ
L7EbXUDGA8fuJUbGucYXB2EuIsArLPuoKzZcLMzgjAmh+sz51jDDKfMYXV1aMfKITL7i5IbNrQNs
rGMUvHSazAAvjh/H5+gjKjhBLBnFxt2Be7+b2Q5lKHZVaCnmJkcne1L75hLhYDzfJoTD2lGZV2PA
aXLsw/XEXzqG7whq52PqlQlWLlN5KnwgBQvT2Y1loQYQkEukQ1F5jOTyWwWvObl8V+KZMXBlBr1J
QMuEwK/gwCDgj6J3gOdHsNPrMWJ2Z0FrO/EYAoQ/lLbmONCMo4gL1accoE3dDp0JvWhlPq5AE37c
sxHdMoVNBiEXl2wvQ4Ncqa8GMBcIybO9IIQwj+pcqrQgiag4I/r080wnaWMgEOvXB5PNvKAilUdK
/3UmxyHZ9E1p4pe6T5MlyoWRA3LgIPpbFJI9PF08IvQ7QTbY+KWDoTR0H6bJslLV9hvkzEYNWx7z
pMWgLMM4ZdwAsTAcR2pg8iQqUyQKgiw0g/2owutr121P20rljIQZoclWnbU7hCvl6W2NDqnx/9a8
rK5irJSbzMDDx43BD0l0ILJB5IibYUfzcG0hWKDaV06KTKcgmAJSUHySfh21IxgG+zPhZtwCthNb
JYxuynOBnbIa5QnpjkGm6oJ2TaBHSHQCVJzavyvO6yuWbfFq8iFZTK2ZWIl2yeo6iqLY38AIJgrD
sX9mWQ29HnQzXolqVHJCTk627SrsSBfXaj7yiIES3eas9rOGMkfdC+TfFdfr5HDUli5vOo2uNVZB
Uhs+83wQ9idnjQgoKnAJkpcqjk2XY6a4yfu6ROpPVmQp7Vcm2w05hqhoF5UcMLYJzQaAuHw/jDrE
T5caqsGqYaiPuBKmchWESzL0lkc3ukWqF0Yb16sPlmgVJO7HYxU82fW19OXrHOjFhDbkcCPoy1pg
mpbOLBNgs5LRAg642L79m412N5FRkBc/OQTkq8GZYqpFhlvVO6uERQDQvradzZ4N9b5LwQRQFwKC
XV7c+rwpQL29v0yEbNDNa+183IdzcLg5OwQ+UEcEj6A7/b5Sm77hJFTEAxHrKKbTpfzD9w4HEPQi
0BQqgYpUCNaKHnCAtWk5XqcJzDOsJPtHs+axlxc7AVipsxiJ0tOooIG8zK0KtDxxlUypS+xQmXaF
EXymAvyaFOusvFeLomdqG3iKay6RF/3mv9IIr6GuDFWV0Zw701hkwS9h1+Pc35jx6/HUcfUl25g+
gaHr+g+6NmeksAthT3C3HpU1jgeIBO1shpQiPlttLgYPfILgsm57WSZfMtpq3ev7YDAnP4aUoD2f
3MxotmyfxaeqBx+8BCiE+dq4ttjLK4+TK5A6FfPxibP6vEop6XqaJQxuAfpokOBDPUBe3POSFnVo
wijTcmsrbvFQwFSopKq077L/Wjm4CSD0fnQKQ11ue4TgOQGSKOVSVZrX/Bl7FqwSPkmjIjQd3Bwo
xDWb3KDFlt9rKo3g2llqIoIdMJRBSu9HRSEJTyt5ox/wf78YHs4e6KPPQZ9scvq/Pp/CmxqGkLVe
yI6TJKL0TyO8KgfuhIO1iuzfzYBDdrR5k3hbAoKu8bRxZxBzRaHt4a3DHf9//p3SOjIe+PAC1Ipj
1e0eIIBzIBTmw7atNbgCBnQUHcBOfDhN1p6r05pG9w4GezKLpjbHRU0Uv4qRaZdAiB5ykNetAMMA
Q5cMfRZcNOXyY8sy/R5v44Jf6E6zTCngahfDonnYh+wxYvck9Jjt/hVvUu0xFKpEVL60w0vxTvD/
Y07wGt5MA70CYwhan1U+7CDzGnY+wpOuwxrYcaeRW1diRYYr2Zd6rCEkQA7G+iI3wHWjkwwiquIv
O092HuE5KpX1Gl2FnuENDv0qCJdAfbyXs2WRuV4/2gI8GwE5GzKmp4UCNFSyOoWMoh6WNA40nZHl
t45oiyxyOacIx8KVPk8uUeuSpbJCH1Ks4J5Si6htfDACTwzlRvlN+z7fIseQujzYXv/1Y4WQcPl0
poY2TMWkcnkRpnO3csGGY962BVDttFY/ZvPBCnaDcJiKABn2vPxffUtBD2XQyDoktO7q68rsybL5
mUsZXdTp6aof3KaiczUFu8xN6ka5dtQ8sx8n2rf9Ccj9NNQf+h2TnD/p46yPuJksP3iJ6u3Vnuz/
BwGw4K77JIWqplJwm4AFkv8jIXeEtD33b5qSBmrkBH5Hjgo16TkcLzwAcDu9iWhkFxcvDDD/ZBc6
+JVBC04mb9fhUi+bnApVrFA212My1d/RoV3z2g3ZKJ8v+/QZpcKAT9cD/U/kPcoiiHEmj1ADpyks
46uNdxNavHOCmflfXXzSiVBht97+8+pLq7Vkcmb1MuysytHCg8rUabtFUTK/pM+ZbO9bziCz2tTa
zpCkwE6uwWfvK37rs5heJ5jnHCGmjEsIZPEkdaWRKQw8HafzJ+fRoQ+kPGFgpwWlWxv1cGNGdPls
24q0MtLr9dCwZ/9OIVUt1UBNB9kpYfRw50pL4jq9rRAfWICUsMCnRfZ21NeK0GDQ1TXHhoFeRREW
+k5YfooR1eUuf20M5RN5Ku+Z36wqdZvDCTi78B/yGK3zZomOrRaRdZ8abl1sJmd+sI93wzsJaniV
lEO8USsEp4nMFWBQ7s/issO3aenRRTLtU0VOH2QbFMYGQhcLICUaSBQAoK+dhI06CMIRGrXHxFo+
4L+Jd+bRhx8hy905RhFf9Ua43jehQzIndZvggAV6Zexhiv9WOA0i3aq9VmmxKhzowIGu5WbOiYBH
mXDtSumA8G4u+RWtlV39cnFnwSW0TA04o8fu23y8BpdKvA2IvY8hQ0M/izxg3qdvx1fxSDC0kpJc
FrhEqximPYk2BQ7fs+5LuiIXuCK8/yLEYvHMNp/QOLbMgm8vFYTV/WkV/Q82AhbbTZ2wFgPodtfS
GsQDBl4aSUwemiGeO42+SWcOyISjAZd6wXOnxdgUqc7Cn2OxPojTZlLoVqR2c7+geJaDlZIkPLAl
MVqjG29A1rk9cb0FGRKwUIiuHmxAKimtgplDQmCOHejoVIvU5ZxrFtEFVhyI8dnfX2I+CniRcIpH
tawyTrPv/MdjAu0YuDtcU/DtM0S0qsSayHEZF8Hxg89nmsVQbUDnWMn4pyHUM8VsJTWWx/DqtbAe
GhgiTUjoYAZwCAFCh/ImGrEzOiLy5mPDTwgBRRXaWCHAR5E+1FeFGpHLBeJKUB6O3W9eX5AEvwfS
L5kHV9mw5ol+qEICM7/49kNa/vgp9B0bDBoYRz4NFmR27JsYSHMtsvngInSqhkbuxN47xMEH37H0
5EUQmyByO1iBYDE/j1AdldD/sFmQT5SqqLV96nKXm4js4ijHvDxQWMSl2NCflcqC/nJxxuzbLm0f
GKbUtp471ft53t5YOyKcxyi/XdHTnRAGIqmygxq/UfaQb/n0zKBCn7Nt4u7g3sqiMv8EY16pvF7d
G8vTwxgEcE3rNMuMkMge4NDG/UJYay11dTfJf42AW3eH9Ww9BoLP/TfI6GANoRNXK4fSZ/kSPzB/
x6uF0ds2C5+4m2N+U6F9235wNypcqigLMhz/OcUbUjnEOe8SXPCFMZwcaiFXNCgk68i5EntcufDQ
4asyNHgx4epyXdPHGUrszSCxQkEx97D7BSCC8l0NyLATAnwUHo3r22yn23D/VEfCNMO+CdyQwFfm
Nc+K91aF7lOkvCbUiD5hVIYVfvShX9ji9hv04qdh3TAD8PkLsgVT+JK7deV+Ld4X6nVy8HOqPOP0
HuJA4dQoXb4/fdOhd0m+qfr/zLBzDm/nJ6imB4QtV4xrxlkkeqoY1TAxCspjdKwaFlHgshQPfSxa
uiDBscyt9GFhejbtSrX/QJHZUvUdbxtoVCmVZfwZEELMN4SKSj8YLUoZXa8Ay+0pItVRlRNpnNRy
5GGJzwX4KrfkPBipS7APE/DvJOEzoPvsr2ZqrOatpUyIGsx3qT96yKByUQcotb0Sp+Suj1NchEDB
W1slh6O2uinjHjdl6++OfAyRy9ilxwQXabnWrRQEaq272JYmI7FAJhR1aaLaJJMxsMs9jZF45T3M
HEk0CbLynDEmAny5GVHZ+PZSoYSN8GvR2afWmLKoSUmcylI5mdd3r8Wcwuw+QMUH7WjPhhpnqCW9
7LYgrSGWcLcB4r8+zeeJWMMp7YUtyuOcoUHxTr0k3KEjpmPDvl3MTjn/ks+LuxG36KpyxD1J07ae
DGIhAV4eHtwWV0dvfEtbrISsfbMPt7yQS793S297zjPBNzivwC+4Q+ebfaFY0mT7o5e7y3qChfqX
aImCltIFCvfMi6N8dRd78W/sDwrh5YVuXnFJ+1FXYQAN+j+dgDc3X5JW7TokwiCpQePspS/6Tx3p
Lpw4QLlJ247iHT8vStJEpW9CGMMoIRkxSj0sWTvWVI0RscA7cwgzemoDLoLISCQEvnUaANP2ZQEy
IIXq4nojqwUtPzSsMjkXGOIndfJtctUybi8U/8UaRrzcEmbmf0OSXjtbZPV4P2iUdR3t2Zr0SQ5h
Midy0VVpbpKPEl2Fd14Ma9DlwaLh2w/U5xSAn9485/mTxEIDc+r2xTIgrZPDHhozK6Z3rjBAPZ1/
ImCOlYBJSITPvwrQ6Y6rg5KJi7vR0b5u30EwIF8i5r59JYmzRd+0YccHgnNYT7ybO2K9l2qp0vQ5
tTTJrUzju+3uDkg506oJJxeNkQt9oVPoNmMlkX+kPdX8KWq3LlbG+MzRVbRx2J4etPszVp7qSmMZ
DQsz17Fmm2IuhVZNG3MOWLHES9MfIiFi6TG2WYPrMYrBQ/ITvmGg18LxyyzmgDaJOOyBn2p1E2lF
PNNSIV0q8MVRnn6QnV34V+9H/HtKeloKVieuI1ajHxY+HW6PcZZgADZOZCCGWL7QxCnfj4y0BM2g
bL+ehnuGGbt+fVSiL8oOAaOI1r114tTZQNwLhMz0uR8q3RRQpdYSQ2xetAqOd24SdLF6D5xujUTZ
Y8KBdR7bNrST+uDzb2NaldLpDTT3czN5nOlSaIn0IN1jnOVC8PpwopBWmy8cJZXeY6sly6+PNc76
cCZ7lxnDku3I3TkQTQxJktWfypyZx1RqOCB1eidXy26Kom+mJF/Nme7keS258/Ydnbw6NEbNORe6
HrTDlJ5eAbZYtheMDexk/MT8Te/WGWsFJKC/e2BjC23xrWqQteHf7tEa5LqIt5MNomK84NhqL0Mx
CkU7r9UQ3QJkNPifvdATmNLmJG0tOEFxOxIzz1QuZNBHI/SefU1MO8kYLb6deQ1zXEoXdSuQYNYe
cRE9+MmwEZ6IFghYqRZoDN33kkdhvPFoZmOoYc+ska1sVqDXF0hxacYvB9SC8xmtLNIdz7uoeIH7
GtfXhOREF5oautG9GQH0ZelGr8I8eKhpIeCnG41J/LB17XCXR/x8P2pztFDLiADDtqDrm7bKP5Yf
4TO1+kOFYTWJgZMTsMi6PUjbGedjTss/cqS/9+qEzXh5iiLHdDUBXXbgN5jMLKhMJYaXRoyXe/OA
lsjwasvu7r4qkDyOEpEHIRmlnnJwfTB1N3nFXNjAnev1VBNnsrMuN8B5bKZY83hcBkV5Ti5K/L5Z
zlw8F4XoRTBo5TRTcAhIDwss75Xq01mT0TMQl0oraCPjUGBO9sOucvbK3DZf7BuOPI01vNMosGuv
xS9+nXe5qkUCAAaS+grPX09KU3wRPMl8P8ftxFEIcYoYm/+D/VS/rGmoeLOtSTemBhWMWoNvwuTp
zkqFy8fChqey2WEjPjKcjuknt1rMV0ryuCLFpXq6eRjkMFRKWxHP64yotCpMkvm6ERBKhjVL20aS
2xtk12IBgiWm6PrHY34j0/W3mUcYzC5+9RpnUj1Yu7Zp66vWQXa/OAyfOM0Fg223EmVpZF7Q7fMh
MUcSXjUpSgMPikvudJYnNBMb2ongbi+UfCR8ny8wiwJ6/o8p8krHHJBfTUbxYXj+A3vGxJTeX6WK
U7k3pBhYzuAH6o1LJjfuzPRChiH/PNlskLjtwWjimieTWyl/9eUAoU6Y+5VgDM7yh9FlS76Aw53R
LnqAmuhVhM5aLjvNyz70QTstwPDA1Ng7EWMycHAaVVNwz6ztaIw2Fi0llCPN8o294bJTuMOor7Tz
lpKzNYI7rproMlifg7YmJwSTIkm8rYmmdNI6CHBfWA3NliPr5D37lpv1rPUOppXMJumB/oNfT0vr
5aS3RdC9yVH3R/Khm9C1+YEuR5TzhxjFmg0A9gcLECU2s4M6xbircfDX9kkPFC2loDoNGdte/Qig
lVgt+gk/XNuDIliDMWis5CAfpxpmUTtyHGa9ZL9V6PWUBojZG/RmRHNLPuf9INqDc0D3qtliTEa8
URH63JQlyowlsZVjphwlqWZ4XNgC+4Riqxe5bV//ZRUUPlrjZpA+JTv/QowDkSDhUDqlqOn66XMs
CSbvvxB51uUYPDKW2fUkSi8+0OTFz559cXy9P8emAgxXxUi5QM6WMsiWt6+z8eUVeOBXRigSaNeV
zc/3OLTCxN84XGjaSt9bUnBNvAP03bCRqq9FB3icNRlIGlvX2VYGMHI502f9XCDf3Ndemm4ueBbo
uU1G/wrs7dLtr28EW2n0minnqZW7cefb4II6B26jpaVxpdaxKH0r6WgMJh3Xdtx2p1AYIoZJ8flr
hKDA7z3S3Dlwj7Kc/jHcT2vglCl+8orBdvht1eOZhcZ7S4bidl7PRyJdO9p4CXKCBPjMdDmadSIR
ev+o7JQSVMuRiJQkQ5vZogRoLNdkUhXc+dBUwsmNhH7doloMho9RKT1V4td+6G3pOg1K9TvPZJ+z
gmR+EjKzf/RbUL3b3ydVGgzN0BSsbCP3cmdhY1cKGQFPPHxf9srGDKD1fAG/J5fRYVrvrXjTLmtz
n1BVRKp+O1owWpOp7oZ7Hvr5xlSv7J77MrlxjXnxvj362LqhaXhO88iZd1zYby7gmmpWPqlEML4j
x6Z5gUxfysJ2UEBi7B/t+IziTQGfdmyxYfd5uTnoX+9WQbdfSeq2phgyeFdLRpNaIfxYhaHlNevP
7BaW38fhoflWplQ4aGUsLWrFpPwgsraZP0qC5pAovHhRRtF8vcjSe95d/8Q/O1tABMiGZj1ghxtx
RnP+JzzzCEA5y7gD4xx9NqHEKdsE141xdJ+JNUDAi8ICFFrjiuMxTjGxOjgqmGYoFZjEO901u0MA
B9QDW5JDa1WTwGURpl2XB4GCPe1d5p2Q8V3mcBnkNUtKTL5tdV4Ke1OFfx734qAtQHRcTh8Sq5dG
MTbtXLU7+xiPPhm2DilSK1YXbbEaNy5qecaVM+JYxtmlb5ek3NZFJnX1w1Pg5Onqzdb9QIgIblSL
90HfoXnREVCFm3DJHVT36ys/N+euBGmnrOXQ6lhbxwFn1l+/w3kBg3KIQSLF21PYnL74GWHs7tpr
2av/Fe99kus+VYXgfbOVZom5aHyk8C8ftX7Rd+19IN3wXZd5UCMlQMY672e0vy84ei82oyzTNbs7
l9xwzM/nPEGUVRtr++xoqQReaStpYaqH76P09na3+DEYZdnleXtxabtmB01Q/xLlyNea6GHd8gCA
qrsfEzV+4D14xGR+WAk83O7MBqlBKPoaRlng9aNLv5sUuzowBUpAETfNYSmwPrftoivJT1Ld7tiQ
Frw0iRTzgxhUDEAgCr8t2iZ1s4h38/bqcTOH7YeH3GQPRbo22idHqRvWY6Eyw8AEitbQqQDb9v+a
Ya9woorZhDNo1L87dNCoGaImjgYJRECEEusoooDo+lS/lxePdXldtoo8FA8rhE8FOmajDTJMMVdK
emrVFew4yiQinbU/XV5+3VWVWsc474p4WfAC68JkBb8bLr+px8XjmE4xzc7JtTt+hB11ZFuuKGOs
3IXfK11l4aFc0K7UKfLifQ6O/wSCdKq/JhEEng7yujCqOiTgm5Vf7Dl7dcuINdahu6Nf0JDluqkD
178NJH13EaKQ5r4Qgmr+04LwTAHYrNCwPz5mwX0mjaKPQescHntmUnbAYrGwpwCpAb634HZh1YQ9
9wZ2mW+6rPHs1Xs7gdG7XzwwLfB4/K0hvL/YuPROOP0q5CTl8piwFZCT5t0a+mb1dXLBf1ZkCN1K
JhkeGp5T1HiqogjqFcUhRE0BBPyRiQ3nvdJV9QNN8gNZQ5pfZG5hiabN5UACUbzkxaXmpRFTL1Mt
xwtyS5a20yEK6FP+46fQLRqHtY8rEBHuuvlWbd5Buus6R/9x3ttyLK3iJ6sPkY7nK0oOyUjjyihR
RffzuiSoPbjVESHU+4Lr0a+I56fLKmyiYf0JRNKbxDAHT9fKGOM2QrDQPCZ3h+UuOkkhVPV2D9pP
mzNsCmMQwqj/5cFECBu4QyK8DS3QB6UnAXLakhh+39UQM95Xt1Sop+Tg8dDaLnDktyjnJeBpNtFU
gI5Etlj0EOtWhsGupiui15qJtnw1j/BtMjCw/MvDQ/n5t1hvLA1zo1liCAFliZI+l38ucZ7wjXcw
cwTcDy4zVnQrdmyGJhzfb4hP3piUosPA8fuI3jY596Z5KJ8j8Ye/9p7HXPbZBmX/vL0qlrQdtTaC
b45bRO5Eo4ZTyUwxsJgEocx5bsGlnzQfdlrJxbt6II/d7+Ikd+nrKvyX57je7sWkUFTX6DNhhTZq
mjbRSDkbpmsb1fC6nQdpghvf1Ksit3a2RmhvoBdyS5nkfio26lNIofj+084cpewr3sC2BTGf8rlS
79D8GAdPFO+T+uZAzUyRReKUn3hZQMTojJS6sZsxSFQpgZMyxLDSeXVNRbuFiqtzCDfbLXoRZ+sJ
rhsnYbix/hqe5rUlJ/cz3XZynKqr6ijjOR3jjpEHpnlnlzvmjJtdQMJmawzojuSyHusnKrdvjEUQ
CuXqKEoVcGmnc2KRWNemlfBY2EfHRWMZ5FfMDB0a6knTdS02sxLnjLo5LjoEX7opgYexquAzHD9n
WBUREsdGL6jYsd9e6rCg6Ms+6z2/lec9myWdvZ5Z0opxzfhNa2D23+hI1IFx6pliMBbu6+Dp2cjG
FTy5AfV3c49+87OvLwXUFF9pjtySianrk2r8qKEZTXDKWcSUrnOJmnu5OZd1XrRnPIuBvpenG9EZ
8OUA/7fZOPFEgm/Nq+6nkUdgdHPdg0RJbCbHx9mm6iGo17ptYitGJ00fN7M6bbWAsqXRd6Gk8lpE
0ZmRpC7yVvr6qW4Z4MvG0Yt/W+TxLeDzNu3Rrj80rmDYsE70UOe2RpWl9rRkULyn5U7ooyKtO5YG
eFtnejSzsFTj1uW58n9M54Ar+UWSxCfWKtKzEEL/tIpyA7jMGg1cqRXcPeGXYCr6GsOqrntUDh/Z
kNuZ8SpieCIKNzvQwtI/oYkZQEVt/rkLqgeMxvH87YNtpV8ojgtwZZeQakcjvVWEbqh8Cv2v7x5K
AEJskKv1847zswvmppFGlGDWLobmp04Qr9DBvNfD8KbUgD7Shzr8aI1H9nHoKLGDRTZgi2I6lpK1
iBv9uBi94MldZ56NRYF5QzUaB1kQgpQ4MHOunmJUKgvXbJLX6Q2xkD02Ity0Wy3hmc42hFkBQ/wE
ESbnzQN32hzojGtAyaUE9BY+E/WSIRrLAM57HfbYd5RMu4Pl0FvvQJ5kHJWwY7Su8TlKfO4zkF/e
0W9R4sBq/2PW2AIeZjf6fDb19ddFbMI17NfObN98Via6GQDuMost1b3RYdK8d78OL4UhOJaaLpsZ
k0/SkB4vAeDipit9AqfAjh2w0AWs7xH/X/WiAmmplaEW7Ou3dDyq2N1A1zmBJlz+Cm6TJ0dcKnqs
1GoC+eTKFVDxHkga2vMU6VmQYpfV0V4AzLc7xuoIf5zk5MLBr2I5ekFUbwazgqbhzOEHkrL64Puy
CxSI6s6FLgFsO21l4O0XsFd80FsFfU8G909jKnjU4kCO6VUfs0XyzueqktaVLTekZTxWCRVyTTJe
rmtmosi30EQCK1QwOPRwHGTiR7Y1dpl8b3HnYTK6OntE1sE/Dz0qV65mdvxmyuDZAtI41gxsZOka
J00iWdflEL8zx+lkUKboxSe1MuPtDweEkMTIfQin5DtuFKt3pSOAtLXesAbHMdhSvnfLh5Gb+ciG
v5fIQw9FCZCZhXoCm1zkhdZlj67gkroBKudOdj+wqRwcJ2cT2S8fN8Y6uUsiCBh4pGxnM++AGUha
Wlg9x68W6peOFOmSMfQzrAzeCDpt80M58cRzkzZk+GNTHi64hHZDAQuWrlT/Nkph3a0RCixtS8S1
Cs4on45T+0TbBG/uhTSVBSgku5PHrx7axGtRk2XKLAU8MI3rtbd0pJ/SXFlf7tIW9d7YjNfpgd7d
eIPH8qaY/+j7USammhGhC+hs79zUxSrxA73Fx9/LGogD8N0th6uYddLCJ4tkaNHnnVPT90M20W22
vGX+OzlxxpjmtSWJ27iUy7ymo71zDTjHeL8X7R6FnaG9AQjM8S3cHy0FVYZhZAa/lPbdAKnhkT2W
ihp3jlWSYO6QGRWrW8RFXofkf4ZhbBIa/wfrJykBDp5fqiEFAEn6Kef2mCd7qTXyIZFm31HfthaW
NQiBjSdIhbWlqwPkAyvEe9+S7uR7a2Gh1Jfl5bEoZiG0kbncG5hLMlyqN9fd4HL5unXuY1QtieDy
WxAkEUsaKzJ+rIBkpwAsNFCvYruwDUH/u3WB0R7eSXv4tNwnlYVAAlkfDUJ35q6jyQHv/e9Y3IJv
47skOlAz6bwGpI4Ip5FPw4Wv/y/PjBkOWAFq46xIhYMf3d8ULErsL3dS9h2HcS04gl/lvs70n9v7
1qYAhrkU3t4F7vO/tJ8/Rz8VwG8/YujhOgGmEW/z8lQmGX17Gy1+dJWXZZ5i2uX6TSCvw0Qp23QK
nMdk2spt2KWXZRdFSgoa5yQfLW1y7/zOkteRwjCp5P7jwYbB6nUYTfE96h9d1zcexfMjBxjBeYB0
6wQMq8HdNoYTSNPfkryQg6tVtJ3UY5HGcesPgDynKEJQAKamsBLjzgh7xihzElLxpBq/phhssbV5
0NtPZ0EkqQvygrfqK63LDacQ2XoeF7clcIuwOSPWMjluzn1k0/BDePXH2rappp1Twv+537rHohSp
VRWMnxexwBf+XNobzd/vPLU9COEJBBNQ+FMBbDBifFQ9gpMqv7hANTK8PBZrh7GYX7lOgMqI8Ljk
un+DY9GZq7zd0rXVEaXbmGoiNBjVb/khlll3TrE3xVtRQiAIjtXAEG2xb7hyVYqlTwbEU8rnnkz7
KIHJyOnCgXjLSaLser3u0qY6Q9F32B8Bd26P7Q3TTSlLPQ+RyBl72W9gWIlhRVS5iCY9KIHdk3pH
p8ohKa6YwO6KVNAgpBnTe0BmgoRCJ94e5uSasAmeH4jtPH3B8tB6+FTQu/rO06DDLojlKqzoYIiH
ZAoGyjA60qttOlq/Px2Ys6LlrvPtacc0ZDUrah0dpHv76tBMEmTYMM+DDoWqNXkMyjOWD1jEk2GS
wg8RnNuCVc1EHnAFE40WxhdvYnex0hJ029Mztn5CgTZwWkaq93b0AK6m3rjr/KaIiTpgSMPNSwur
K999eCM1FDlnCr3SifD9Zd1WKB7bApfSJ4SA1puEBOzh+cOx4mIO/5KsHGaqWk97/fYwit+GzgzZ
wXKjhE5FZZ1x0ztWCOS9qdFpgT0Lp8wvTvjO3AuCZyvLKKelGg/8muSD17yg4CLyT2t8JT7F3OQx
5oEHiLqiq7VG2FXrZKbkMfEU4hNlprYLyNTrgydKhaxwjg8zKqxjPleG+cnsRO9tk7PvyQQ1MRtZ
NuynAL6Di0/sW8upny1usGlFnoId+lsyT5GvP8krdJ1fLeTiMBi2R614FLE+eEOZW6CKPdDDE13t
WEq07Y/ge6RKr6VGJoCGfcdObmwUw4nzofq9vHmAzMF+2PfV5yxq821ZYgrfCQijM5gF6yHWH+BT
X9F2WryD5aNwG7J1yxDSkm0D/Ctp1r1Z3WHlIVAbeuGH/nvOwvaPjGwMUMGD8dLpK+Oht6r06ZY2
p8Uw4A3/13bL7FIE6jC36ItwWOLtKXLNJWn5gD5FoCYInZVc5J/BIn584h0j8qibkpAWxxlR66tK
TIrWF7QEUoV5prRNpU4KAW5K91eIY2DnlEcrSjRBwUFGg/PV8iwcbdCJG8p1Tpmjkej/uJE+5tj5
ia8wbwzzErL9mPUZ7VlxRnBhK0NMZuuRfeT/vrD4/4HuNChurICmJwWWEl//DSC+w8fnbTpXc7hU
//d8jT248zolXVFlQIjdqvZxUK+kyLxYGMtRpcccEWB3bElzQaIhoGIt4Am2Tgj08nQDSD6RjDfI
5iuh9JsIj9A2C05Ynie9lbpeCO5BqqtrHGhC74wSVPSCIqJmWPnmvyFCfP6r+On8+yeqIVoPAxuz
pF/wLvES5zASEPaS2V/8tUrbj14wHLQeUq0OV9VaKrkl3+0jLJRW8YFKarfguRA2k28vl6Gcy+YB
BSrsJT6n9/2QJ9oWoT4NxXVJ/2fTsBsMe0Ns8PJWoXcbsr9USBbCK94fbysG5NTyRcEHiEw4JqtN
/z5bETOPi0k+v5XHc/6Xm6VwdePa5itd9WLqnGj660B34TTZ6cWBRHs1OUowJXE22Uevg7GHcDn0
LqWO4m08lFFxMyEkt9QoxHcaUtfv8KeLW/a54vuTxMdtpl/pdIHhrVjA2GqPXJ/UhBScU6sZJ/og
SLY5j+SKW5Ug8dSOSkTxkmiLzEp7h8o8yyeRq7RBB8JkqDi9qm6BzEzsBEVOoqXMsYnfvP2p3L0I
xim+Cz3HYq6q4hJIJ4n102NwwsnQ6XrccQkGGOjpuXKchZVgtQS6dp4robpwfXyXb9/sBH3fOs5v
tbcoGq3dYr4CVtv4KquYstjiJQAXQaXg1gAvkAigRLocr9v8wrfkEj8krVOGnbCfxdE9eN1VBaBm
n3h90K/VTfOjQpzSwbOknieQy7WxmoKlYizqj0ZFUsny/eq9zxiVnsMNUACYqQZlz1seZlBIlC5V
O9psody91gTqWfcvBT6gCdqwuusrHcR7IAFlzza9HLOdzR4QD98QcxGTAokDDM8JoM7FJyktHQ0o
k7E5d8VoXQ/s3UcLfPAI7OZiHcFKxyRW2+Zvhz/W1FdLGU/YYgt6z9cpu/C9L5gHPvgt3AOp/rIN
vGakFivriNVw6uhnwlKGCFEGCFe5mlDehJgoLTuqts0Vk2zPCr3Im8GweabFolZ50nZA5ESSUs89
VxRk9nLNzsaMFRrT2/2tumuBzoFRVJtUsVndDGK60kLd0fzP4Poy5QoMORFDll9SX+CDbA4nLuBJ
6pmzuzpWeWPL2BTnhSe3OerXbSC6LI+p9GLF5QPaiZF3Xupw3nTA0/8P3NUEFFKupD+8vVKb5KqH
MBKjCTS7Oxbg2ZLLwqGBQM2kkVgAPCu7/ZU+TqNJuABfixe3je8wdiRnQb9MZ6Hyk9tWy6otVSjR
hpxa8dBu3FtUyjJVb33+SeXEwrsQkO0468v6eii8/WmU/ZPNSQBXdK+aEcMNdUngOSCP9UQ9GJaC
bj+48S45pQJyP+dfJ+K6p3DotpGYLzFofyXOS9o8sUwO+jM0FDnsj08sE1m1D2nlAh9mvuNllSC9
/WC6WgwrkmgALB2G3CPjK4tWvZSoE/haypERNSYbCn71klNHB5nIm7YXl7Ptl3koUy9x3H3EhmGT
1Y1XQ9TBMpSpac27ZmgFzCL5mdeezQiBQ7KwhmHxGM36gJjAulQ/fuEBQUD4iFO1pIb2/HiAbFDQ
nKmiTR2SYczqVksvAd8Y4lvPs4aVeFokFcbIuLZCsxOQHk2CIHMxhgHPkelCT+UBwbA759ZGomfZ
Q96MF+rtKwR+0zMGfjWV0JelE9Ow89RxPrZxFtQGSpFBV7MVCPXyMkAfZUnRmpgI6fk0siPHouhW
ME/rM81fqkvmxB3bXCr1DlmgzHlP0rEJVJVLB1/gMOOEaW0SA7Pm35MZwSGHH8gakcJtVs1DJIHD
QkiBpVGgwOToaUtTcC3/a/7pS69RWoD0wu0SYrz/jkmYljYXNEobvaIHEo8pnpME/tpqcGeW8HVT
zK8FjOROmHdCJFL7FcxxvqHWlbI9uaDjL97ihaNWwe6Z7ZcUX5NZvi9dDl+MJTxJecSfF8g+vKl6
dmMDqp4PR0XUSzVlGMzHpTrSNU+Tp2mhkBRKwDlhDWP3lyppUpe6JdHvyTzLylCQG6Pa/iwvA9qB
j/+9lciR3qyBnmiYinqSYHt2sgJ10pubRTfjSSHU/uBjAURes2v1ERlsTvwCP92jTWtX2xgfCB7G
rKyvb+x5BxH5RbqVXbvXfcDYRRf/7acOtVeCvMAj3+AhqSoiIXLi/wcbNrjMEQj4K4y04JH1mesV
If+dbxZZP8fU6S5Rv8wu2iUAsbunKWUdtNJ6zCRpGRbsFCJFy+8X0H/g5rsRguMYZISkWp4dxMDa
QzVkTXNu4Cpsq7GJXImEOQgeWr7kadWlBWv4DZ+FjlYJj99HZJYEz82H9JxQhQ2hOJycxs7615jv
KB4k11dnYGNsO45OZm/ZuSrpA8qOWSdBgmLxve6U07MQyiBT9KLO1ZXnZ74d78i5zc0JOJY+gVvr
gw699r9GFNPwtG1Y0ZBvcyG84hA7py3vAnr24K7XdouPyCzhK9akry9uiJVZVnrdP6GCLYd5dXS7
J1rJg5PT3bZMHDUeJ7T04agDn7vDCdA5nZFQMGLAiYzO3TDBIsuULVRTY9iOCmsqV04O5N8JV7/t
a5s6Aj+VaAIB3CYxD4iyvEgTjT4TWyCB7Mep9PihDAomh5RuJjoJc3bIzFirCsyyjWeSEqrxarvq
a6W/EmMf+7tDC01gRpbJQ+g9AdYvvcH6eJUnAiENWTFpJCT4CUdSSiNuMr2xn41dC46o52GOTpCK
jm+Z6XOQaNEKBEI0DX8U0CUN2SN55BrGhzdRK9Sezv0g8gx3rES9go5NJdjaOPxilODBP+BS9+5Q
qRnlnY2gzCZRUGQ57yvPH3tug5ZEJNZLLctj7/bNxGu3rVvGqGzlGaOgBvQdFgXlA0pZGwExiItr
hEhM1R8Nt1g4rVqeKGn3qUdaPau/uePoT4ShjUdNf0n483ZZh7c7Jvq5MmsWe4qzPiLFrCSWXvhO
mURUMdZaZU0iJ+um58ch4gO6FvBHnXVYw5G8XpI1sfZUYFiToeMuPzsruyUdaZcbbpEPN5OKlAIG
7W2BW/7DlmSYRXTeICbecgMMPh5tvlnIChFTKERTIZ1hZICQ/1e6tGyFWvae36Mj3hht+KJNwBKl
d28GuyAZ/XZQR9qjKJXysmA1mDKZPmNjHrstjF7iKu9723G3vL7dHIUXVgAAL30HT16HfnSFNJiJ
tgaW6vaeOmjYA04H4eDH7ACnX3CiKd6BsUKR1p12Ohx/FEkt1QUpIuu+HxIDM7YulKihKRLr1ghD
A3ueJoA/nXMxiU8sbmWnlM8DvH0JTJ0ZPxBkSDFG/DEgdigppMZrl6EN0q76t590YwWm7kB6CaZc
aHIlw+HBL/6Iermk0vaXYntedop/DpBu2gZnwyllcpVLGm1xVJc1gUALKBwGsObimir+kc04ux8S
XKAzys4t2Z/FkdTJEN56Rw9lItifUZiuGr6buRJYZFnSYbkonysKQBPKaV6zygrOJqyBeoAGYgx5
qTSIQbp3Waxd6kA0TmId97SfR/tVqAeMiwcBX9nO2YDc8S48zVe49L8E9usLT7D/lykDgKTOlShL
PQ/JdsvEIO/cP6bTj2HWr96Poty1WjhB3LPxohoFzUF2Lfux7SagMyXOYUXRymazwJtvWOTTIDn/
RAXuboFEPx8VuvMQKaZ6MmL4oaucXGA/jLF0nQ4z4ercYiW3AcCQrFMlZNq1fuek+kSXwRWos3f6
h/tteLomvWu4W9ABL7bpk3sT76rbZlLMBU89nFIfOy0WI7BnD0WbUeMgzhjmCLHlY7aIOQvqAzmr
HZBQlbwi7bMCAusn7k1XCy92MFFVKBAAGE01Q40DnJ/d/v2SLH8EtjOhI3LC8uEMHZFwQxw6Pamn
jy+2XPlixgUy0Y0sqRf/olUgSL8izeaE6+fwDqsvz77uUuQhn6f+pM/PYzYlJMBLp2MusjSQd61f
fwmzdYTQFTiXRq9/zUJGmN6drxrSPj+zWoFPmvTG6wX/69jGm1g6+yrOj+P8O7wc59Zjfgm10BYF
58PXEZdNKiC8n1clO+yR9Un5XId9MHgFN/4045HpaPOqvZmJ4HIVji6nMY3+OVGWoZqEmNEfJO3e
tcuzNMFEtOEPs7foGS1GVkcIjY1/an3b+aLW1ORZ4tbOlieSRv8aUpMLsM17VgxnlgR/Ha7oX+Xv
tLCqNSH6JWZxtfg8vCzfwUMX1xQqiqUMRU56jVAYy+D9z5p3NPo7+UCEjrfcUPFJyemHx/ylkss/
4lWkWthGtHp9oL0wkQfHztRp7ejxTa/muhZo8QhVcQUlkfIQ4zzGuAkiW+N5wIka5tfWQKq8bp9u
PkX/RtpT98EK3EQCbS+kR6wFHkIj/ANEKHsBAhWukpdrdRot8yWPp9oWPXnlAnYogZx1VbNz+7DX
07ssbpfYSzbjegaXR2zgVluRAmo3tYx9gjZ95m0MoOdgffC2SPCjcnJuVdlvHfV4OWTK1o2QQlSI
hrQdk5hy81nvv+19bMohp/7VJnRJFD9d7OXDNdPcWy1uvNHXHW05vqe1nmtUxHbVluXvsx669mfB
k2j9ODT1xKOZ98h13OO5qmBhMWMpX70KHraDOGYAFYSrYlajdss6PjZptg6Y1UBODUc5SXkctP/R
glaWJX9K4uSPzO/q/5S7FeV94Y+ZHwKinxrSoiNClNLi/byGwtC8ghEmhafNuEHMDzngi01dqL4N
OO2rwCJ7QVwMM+bqyhipbamO7hv/pajJWfGURG1vN3UZP+Xx116xo9OUKn3S8iyHTVIU19c+VQib
Ii7T3zL7Iz3AWXCE2OdZgnb8sqXA3XPK9djBWmBau73aip5zYvonea868D2NyVjQdWcIgGNEY3mE
kpFeusC2rlMZsZcpQCqN4HcCrrJW+ApIWR6qlYocG0u5n4g79QZ/4S6/N2LOYRQDmr1H3mGQ9ZI8
NGX1/K6bqKZ4apRlzVm42nhcYLM23IBJtwLCyc63XtMiHPU6kltxQ2+efwiccF7AsQOu1FYd/d13
uCTu0o0fNLBx9vhqWYHsnhSs4SVaWhYCiWqStpTtC9kla1hV6zDIi6CwKW50ehIAZ9DTSWkmTSzh
DlbEy6xQYF7GgMvJG42Dex5M18+DozrsUku70vraja2aWvJTJQCtW85vkrF8zw/HSe+4Z23+lyPK
BWbeAo/DJp1PB8GCoKSa/NyVE5oe6wTDKqX269wKVrQvmQfbSQ8LAJD8QnEwRl6Ipw7+fSnHEqP3
jplwk2ogEINud2t/mXeBoUdC39RiH44EYgdin/CeQgD0H9FW9iGrNRq9eEmQE7zXBDHP2ge3N/Cl
GiGCG498xAMrD3tAPjyQTwHXVjHs7McPf6V203abWYAzpzmyGZyx7JCOcV1ceJO2HtUHOjkT9FX9
O9J4PVkmQjvJD1R467ca08FpH1E0cpX5Wxc7ruWrcEUFDIK1dLkDTsmTOj1EviUkLISCkbBZZKAP
Xv5KEjaeCxvC4n4XTADLf2wcLT6CQMaQ6EuXAx9gynsdyUh/OjquoHcJSRlYeDmLEHZ1DO+BUTdW
YO7GOMwcvNhoWGJjQXLnIhXi+iS70uesRwzCV9s9uGyliPgBYEwgd2PGjB00ZEDE8qhobgJTZ+zd
TuF80d3fYtfKotsYRI167QWiBWjJN5D0JXVW6S5ERGWayPN2qlu+gB14Y9//+Uqtb93Y5HsC4j/s
kmizmdFjbIhQ+R5ywgJWlcbA7VWsozaN81zesE4sPBpDfm8nCp7KwTcLVVFsJn29eKJDVYYDT1vB
9v0ZiPGFpx8yy2mX+H0V4o2cPvethjMDMVlXceTiZ4atBKF1KfO/+Yw3KkZiN4+tmRsJyvtLfMMf
XF/L1FPZCZSUKarB+VvJVmxcKIJ+Zlh3bKpyt2MyDSb7TUCNG6/FrgnVhDfiOcxsKf9uAMVB6MJM
TNEmjS7OwTKx4N+YXdVpP2zAB2fqMWnF0qS+hJjB4NHvERdZjZ8IcsNBWo7OP9CAenM62MDmbYlR
xNwoJKgRQ2LTVNOYmT5CAZgBUUZ3X3HwtCLbh+git8kRCnOZzq/cXuwNUuiKFSMBdVSwsNJlFgW1
iDO3ceeRzQQPBZzdvlfQ2msZ/RvCkdhoM97tpZ6H4osRLW2VNqq3w+nakmbbzD1t3uRx3RAipuh8
17mVT9SlOXXnrubs9DK1HYdBcRFS7PkYVrFUc8zxCOx3ZLgFBVZXRGJwKjTUTeKxkorcv+EbOX1Q
ipW2kyVA+ZG0dW4VlGlJ7GRL5ZmA2d9JtT0v5gHLQ0VTNkVh+t9uFB+HQo2msttFUZzqShYqIxJx
zlR9rEebo9weqeyiAP4FLghFYOHqrziSdEP9Wkjkq7zKZ/kYsRZ8Ge9O9HDiRb1bnSJAc/ygeJS/
yLK68d8h6+zAJeSFdoRScls2uVWq69ZiLxR4lBtF/LgECmLce6iF8zgMnQx//I/wScnHdGrqUtHd
Ysd34yBpfht0Zdia15dI52km8WTZMVw8TXayTrG3U3fGJkvs6V5hX8CP8vxDTo+1ugN01xz9smHj
pMxpI1razWC3kW4Ol/oX647FduFQ82vMNyfHJN6GCxq0CvXIGuhOJhyTSMqyKAJz5DD5xDPoAeLp
zMHrpHoWWglx7zgHAXgATsRMQtp+dYx8p8Icp8sJ6W9c3OIV6N1nh/thJ4rXQHMvS8XDU1bUCLJN
KSFrZcHY9pPYHLXg3AIyVovTzUpvrjToQABKnEqLqMA3cjEZt0JJA3HKLWNX1Mto2J7T+bnQlkpr
+JRpeLze2GyP/5kGLnzGszzgVd3WefBGQ1eZp7z87PU3zKRPNN47UBH1ZvYcPJ0s/GKs+HjCbpxf
rxAblzx7lUDNJRQfZOpFTU6q2nyUEj8GLDdhbqIoCORsqCUR3yfHuc+JcfB7xKw2KYXNHfzlZdQU
552Nb52+X/RnKqrynSlRdKj35Q1TWmxv9tbbCttBdSTKJMG0r7BpfNFTOQrLCj4AXuOFycBUvE9T
7pYKxEZOB+rLytJi5ULVBU4ggVJqJleXY/YCyKHyXcOPMs1h8xuY/N0ae8USC1OQ0wWkxEbAM6ju
mT6NIGlq9Dy5T1K0G/fyXs0JLJEMzQtcB5u2exlSw36hURrZw3JvlABEaB7jNu1Dblo/EA5+CPwp
jKFERxoqS3xSyF7xiPYlj9b+Y25jYSdZaRoVZ26sKcZQWQj5hlRNzNa/1vLhLN4nzM8/d6PDyDaA
TRuggGX04a3wqpHg0Tx5U01dP6Dh5vxyMukshuPRR+txJicYHJ82jtGzFPNrXWOOlwWRlvalJHN+
ipfaL2/5q7QfW20y42iUUtGTNCEBbVU/kBJbQ2/v78pDH1tSVOEaEo4xE2SAfqfFA8ddMSZ1mxWU
wjAVgJ+CPBz6M7jyC3gBhFhOi1kiDXzDIfFf1nOgr3K4twtU6RQAwQagRuRG3Xna4wi68xPAPXXP
yJfq+LscQkM4Fk9OD1LWyaarWAkssh1ZMMd5ml+wl+T82dfDwdBCHjpGOqxG2WVg2HITta7k8WC7
3zCrDfhlJx8mG7TCUFZqQMrKq+Q4VblIe3bYSFVSeR5TOAZr6BUrQveABly5VFF/IsiXaIBbjnXR
ThZWbBFERMonRdUKeoWuNXpQQmtYiyAKnxL9rGXaeF4z7sA9u1ZaIcF1acbxV9DZRfQgN/6BOy9l
rRF7sfK529+7YYNAh0A5gf3fjuGXdNv8gS95aGqakKLjhIL83SKjP0a+8uY3b05PTwjtf1J6r+fl
sPBca/QUUgOyIkSwMCI8wL2nnPxAJzNmBBm9/RFefGxOcIm4NNhC46QesQ6YPdpcDaq+K+dhBCS3
+7l2KslGXS83oBxZd+ec8ZY88UpUHBRenk/LZQBd85xYU1rJinTE0xsBEQ50anrjmsnz8T4jbDvQ
5r8SZAVKhAKFfkDSgq1hY7wANGqD9uF7KyuakrXOpKt32ZMJwKjWSHrh5WrpMFwyIjYbVzo9i/bA
eXZAggaa275rYlCB3Hn/VBsZUHu5D7UaAYPhPrDSjAOvLG50p8/pJurJmCTRAVINj+UiqDMFIcTZ
jOuQL/68RZNdMrK9MZTlWQTjHTDjKPxnn6gdT0cVSq/ZXyzg5sM6dBj/9I+lfZ7YdI+Nk2gd2NBP
afXur+lrnCYg4oHnUua0mWmZF1XAVTqhZWBT+2V8c2waE2rYispUpOMqciEkEfqiajgixjIRNbFv
cAPdI6RrRmL7UrarYXXEJ6lhVqpywkULYd9nJSrHOvLCGu/vyLwSfpcXCkImy88l1SURejvuF/bS
6Hsu0XUCsXKQxMTo7938AvHJGlWdMqGnTuTpwJbi3bBxKZBLRwEMyH6ECONL03hjsQFIkfmJmtRU
C8VjaH06qR2+3Wzck1WDWPJNRLsfmBZu8nUgnxafzIasoXDCSxwa8IdtRy9+21DZ+PxNJ/ADaZIQ
/D9O/1GNWhK24SKVHhujbCaoxhZYUL50Y0pu7K0X7IoUVU2nsdPXmrj8i2yY5p0S+pWqMsyMi1Ov
LrrQ+NH0z8LYtsGnKdc0BIps9USELsk41QdteGsSev0QCG+WokZTSUcmN7jqQfe7e8652ESJd3Bx
jSccRlrYw5L+2IJZL69n1TuQ+ZNWfvnVkXmpmjId2N+GcMlEckuafoT2Jv6W/u/pM2rs6kMTrO6O
QjyLiB5Qz8aqxX179/ZlaTt1zuLBmaXyP9lF4iDua/ot0UyQktbDq7/V+dyWPLZqafRib2tQFiBK
+NRaGkfeBLOpPuj5h8b6PJ7UR2ABFZ4Ea61u23AcxZdC+g72/BY0QQQWwHTIJta3ZZ7JszaLETau
vIF8wt3yCondJ5o4a5MYsh5Uw/Qlr2rD/Xl0wa2+LmjWTn9pP0hFodlUDg81HYSgYQtsfROesgd2
LTReKaogZ743dq7LpTS/zh3JuiEUhzeJHqbnOiAHWLjgCfug//osz1IqD5QxpzaJz5pS7x7mGJZA
RrbphYLxEurTqlrCbwBUjLdzWW5IOZJOuY5ochrDcyxT2R93c/HPPFHd4wnTFGvjgre+w7TNasKs
gR4mSExE8zDfu51ryNZ+Owm4S9pdmN0UQJMB/YQYdK8KA+jwWqHAKf/FaP2wbOYdeO4cMxd14l72
QVQQ6q49osFQoiWyyT2Glw6cGmyhC5DwoNMsnLVvv9J0X3+AN4XxVsMcyb2XtqdqCDHsdaL6wFhM
7/pTcjiKpdB0ziuhQ64fTHOh6lOBbH1HeiZG3CC6KBEAyDA/3SdIfF9PutXei0azl804WtS4ptZc
KNHEecD990rkT1KR28EafhzeUtdegS5Sp1XJ2a2SdiSRl8bDZTlKioj0h/LhOxW698dZcAfuZ9Dm
q1FchXO7S2ZHZEwacHuPlneZr9CYa81zJKcRHiwsFL7i48IXXH5lTDoCPSR46j3SdXnQ7W+Wifwx
sSdH4KGAVBb9DgqN2HW5VRZPGJP8Wp3M56jTHTiicsguZBpNuE/5ZOHFLCsJeq7yBLlFaCc2+iUL
lQ+xyQtt62xRdxF+0SibuqvOOuH+zDx3uF4MCHSjdJszaXhz21haL4S6qwQzJF820meYiCre2GxS
6XcItCx05U+Cpc467E/9U44aHNlsnZcgR9Eyter8Y76e/H+StNo265Uj35V7/dJ7E+DbGYZMqwiU
MWGj8/XOKvZVZxJ07LY7iTYspCW+ONg7nBbFCPx//lowgfX1gXH2vge+TlfLfyL06+gylZJU3zMY
6pSjpvy9eKb8ZIY6LNGshItVdP17jsiY0IUy8tpy32ntma+1SAg6DNoV2ADfvtdaCxyoQGG1HvGO
G+Uh/umFnbu5tVBPclcVzPCVv09vaBjMHOaNSaGWEN1QlufJRNFhAIMrPF6c7BqgXJS+wTQ4ET2Q
bO7R3BUfzmQKe82PjuPO8uIAiCvI2qvU5ljjTCo00HArUfQ6MUnemi5fH00TUPfsGs+t+r3P9SrX
J0ZmO7lPwUqsqteeaMu1bNPlunKB+9rdUEvf7zM+1NSbeIAV7FUOPRRbre/c6o9Z0iaCB7K1g9fu
XD1HIMJm5pHJ4anXLPPuaxCcaEoFNiI1uTMa8PE93dsM9dOI7Y+72jrtIE93PJsj+2RZS3n9Etww
+dzjj6Z9F1z+zDaSYS1rNvWTEn1YwaV0Alg41jgV2OHNp58CXtpzad+qhgHZIbAWIsCBZOyQAkZk
LLaRoZ80EmSELFPbfWKNu+E2uz87dmXUszNQVEzTSzBcqlje3t8BhSV/+0rFKyB7I26dMfghI92J
kSA6C2xaHR4aLRpoIkn1J5FJYo0ht+0Sf86GpAxvGuz/kfdJgAt5dOV6Up6rGlm4WE9kD10Y+WKT
gp6GD+pqgSHr5krpJd6GfGclYzJVCCdR6apMyetDJygMh8aV4g4NSiT9iBnsihBOIhIPZ6pwhV2S
IztsvgC97rIHRBR68vu7jNJvxo0s+FDdD1oOobUKmDOqMBhXgxKQJ27LYz2iBf8+ZHFo9UsoFAEB
SMu4rbhq68LcRCaYypO1WxS9yPnCMyMl69IqX7CEMhfmzjlXywqRjJ+TnwRguXog52O4lNmqvZli
OdRZENNXvzX2hNGqlV7rdvvAhN0UXK0yZ6SWASJwEjQofK36GV7mj0AZARVs7P+QE/AHOiDBY9hb
PyI2sXXFrsT1B6xOQw9uuVFj9uEVPIyNPBX9G2g0VvnkPzupOk4qclVmR8iGEnzidHijX7mMd07u
EDtYRmXldAtLhXzwbFvok7KG4Ey/2ARAKSAHze34Fwo/H3tFy+6O54cjyu7sieqrtX8RLuym3Lf7
G8lniCNy742xqWe7xaczcGUBnDvMLjoc4x/zqc3GR8sd+mWzEDpXTQhXEjaQUQGjypDaDBhFlqqL
iADMIt1Zl/Ti+jdsDENYtJWPgZyYKufHgrYmq+r6Fi187i1vQr9xf2wvTmtn7OGrhHZgMYF5+kkc
U9PCJVVICLPzUeHRUQrG0yaJHQIuVkaKo1LiAzwqajJG9Z0HwFlXdtgX7YHJIVr6yJTARiYlekof
OUkNUGXuHItM+b54pMJ1fYAlG00+aJIgbkhDrsGGFdkCw3RVQKHeu3U4jHMl4IwQWbyS6M1Gv27O
QwuJ45A3NR9SuCbACMtQnaA70kHyKOi5NXguGuK681j3KwQ95xifmhSjtYAyId/wR9TSKWi9Znw8
/XMScvBURo8mQC+YcGJISHstzw0ZkySkl9TFVw8uRlSMmQRNreLfUlOrCgjKwnLXYfJtvQZMlU6Y
qu2Y6b5mO2NOy/50pqRxnUOxmq2jMOc4HeQpC6gFfg+13YQPkRidasXrrXiOmfibZCEtsPs3cUQb
y0HD9YCuuFfui09BkLkLqz4bfN2Dew9Fjlb6j0QtpYKwqmA0D+05kN0NfhonF7PktSWsylatUOVM
GHsDAOZFgunkj4c8XGhAJD35Je3WkSgo8rIttj6epeUeAH1ZOQCwMonE40Kzh2n94gQEBNPJWJXu
5XkTp6YiTrhoFarv+y/kt0dTEd+wHFHyrh4+GMZLjOZNWWyE7Pqw/c0xmFK6q2XttpeQ+5R96et1
7oD9T8ntRv0mCX7px0xtT6HsXVevgUA2AoQGsw+OYU5y+czR59gbGZksBwb3qUFVMEwLXTQ+EQ73
SHza4VaUBaruFlBf3H/3r93C7Eg8/cdZFITCF9AcXOBYE/hZDQu54Z2kldYnaYJKTRqAJkwbUkaY
RLv47Vt/kNrs6f0UtBwKZYdtvewr6xB9g9+Tlx3tx1SA1zOxmQWzy0hvJWOhO0MkvDS7Di4F66NJ
YUvT6H9hEutZ/wcyp/e4jIagY80z6nL302KVHkyhn2ywpEnakHAwD+eqI12ciTrXmKcSRngxmDY3
1bu8VZPswyKbxlqxhCpudlbI2+uX976qjrGjxNT7kaiYBi6SIRYBSuA6HR/ZtUy8CvK40Uj9OGrl
1R9A/Vsn80ddD+Wg1P3XdjD2OoHE/AreHV3GbrZOS2AIkAhVI0jE9B7xjJ63zEC3Prho03kGQDuD
KDE3DufnzeEWnFBh7AydTt8LvhxFXS26sx5m2Jqj/5X+V098Ypz4DMquPYFwiHuNXPV+3wUYC6Nj
6F3lYKIVcC/7LE6fOuvMhG3uE6GvmISHE+Uq6WBDFEwVFD9rjX1FJsKaX7HZaqA3YmjzRIzWtuLw
nyJSBUGfQ6gC3AfEv/jYbsuhEInolWHP7g1lISXZzy2zoPMjg3L1nX7Y9kgY3evbiQxKLHmKFzh4
s6Hn2F/6DEcK5Cw6Kgc4xqqzz+UrFT5mJwrNIPAIu4646MlczIMG17bkfRsOYc0jcsvsY05Kl3lj
pfKKJ8bfjjTuk6OVlFzC+O/ox5IBNqozPxk02Ynn1EnLitzbITEyWQWsqhuodIwOPd2n0wjnd/ku
939KOxkbcyTX3fpul5FBecBzzWVMU25Sd2D+qLv7kzq6L6zXVyP74AqcN+0IrB/IVICfrkQhlqg5
xDB1/zuVe0tPx0cyxOSKNCCRiH/ruWp6YVDsnS00nwzOhZD5rbdUhTr5V2pV9gOlEX/a7I7FQVka
aiYkyEtxkw1phqM5O/tCKAGbUdPTC4i6e6XoxqJ9sleoy4BArsfL8I3nrpmlKjINoj0MCuzHZJb4
0JWI+pqvAuaJpOYNrhtECu+XVO2KACxo+E4VgCnmOyQ20NeDOgeXelfYf4x5oyP5qzlZ4n728O9k
UeA07R3lGVaXP47Z8z9a3T1XftouSFo07zHRxI9G10eP0dGoQErQ20L6XjGcJ8cmWfIxKKilvX9r
8HcruRIdQCOLFgIYmuo26jy1/a2kYTkf+H9o9xcbqpK7WjfqnXQANUJTUN8ZBOhJMqn4ptjxzv9r
wJYxa9U5F1l09IsLjFx6pQscAKKDU8Y3mb7BygKazZeXaB05m+iuo+UosDWDfbSWWPfH84U1VOWn
GHYfGElv15fO35RnO+OdQopfyZQrb5qqLpVUL+jY3AIeB1knL+fvjIu6Y+hjmmNMtHlDlMUKjG8+
qHfH0GDGk+jN4fi8ZRLLQ/zyztClKo4f1cOMlsJ+Az6ZCOk26G2sYCSLBg4/LasVpJIJkTbTh3gH
VwjrUHm5OCWJSwG1narw3zTwyoVSJ9KToynLb5MJ64PBT8RJyc3/LNIOEZVGTAxVtgIfg6qgNxH+
kNYaXl3xxW/n5evfPNOZAvE85FiMd74tkCXHfAvu0LzWRiil7CBQo/cnpixX3D0jm16kh45RG2Uv
5VITKcmnUgmVWWTGhDrD/klzCCWCnjnU1yLdVYRwT681/W1Rml/dsvAbJonMwFtezs2qZ8KT9zdn
9bYJjzXgBHhoTfUPI3yVIkjAIvbEKFQOTgspO03nnhbnkvv+eSt3jgClEpiXHG8xUtewOmCL3km/
ly0L05DKV86Ugrizvkal4lKaIhPmb0nU9E4PyBlsrgaRXHtWEUTyzAeJvdrZUgEmxUjyzKsb3LnH
VLzwqR7jkmPtQpzXramA+Sfsgx3Op+DZCPesUfoT4dAM7SObgNa8OhiIkxf5x+AQ9dV7o/tMF7OD
c/MFNzwme1dD7MtOVHiVL9Glh1j4MU9mag6EvTHCm84+1dkksSuaD1EGhcIEVl3Hu8ZDMK9VsL/5
2K+fhgF3Nr0zG1RXBvH4w3KcvqCyuqdhr4iC3wPa7cqjuP7D8dMLM8AACl5CUyqdHwqQ/jPEv6yC
OJzy9xgzObXIJrirR9rvu61uAu9jUKb1SEgRD73EVAZj6V02JKzP9QlJLarJSZDFRw7Wxjw943oR
Wf/oRc65TrH6/MYeXy5154jk4LKP90YrCm8vAUMayEzCa9VQs9mOrShD+RNT6QrgmOQH0gWsCI2A
qIoAWbWXbJ8g7idrMIeO0359Oz6K8zMoCe0E5fdhG5q4wOHAFmzGj4ZT1PTZMuVVbLFqthL6leXd
K8Is6VPcdQ16/jGZFcRHpqsv8hajZzFJu5rnwZ7vl8HReTTs7k07lHtconYLk5WyN82OcpZpQriu
Jptbz/CLp5AyWqgfFxRC/iJs8IFTekhRYQ49+8ho4KQKbijzXIiwwqShypKCp6+NwuqnEEdQjCvp
X/KgeLjXwzeNfjp5g7fzIInGPvhQnZj1IlEuAYOSmlmxu37cZyM9ou+6jRCRI/DA0sxl1AYc1en7
8KsLbg1CCKYdkOEtkOJnRxRMjZWL/PeyuRxoJdwhaXMdFg1w+PYdszcakVCvhRBwejMf2s7nXMuV
hcmr/7fqjniuQYMAOyvwl2+vTqRC7KW97d00Qg+etVBu1mntfDYZQhgo4cGbXtHJsZxBq/y/u9iM
Swfg9QjiV2KQo+Z9bg+ppgHq9Qz7jOW+ktvp7tZYTwNJ4NYUmMQZW4UTws9NMDW6bTtogcqu4lBG
bjh3fw41gphNBkd8IbR1iw6B4vjQfCv7+0ogxtDk4XNtTSOryEvliS74ghip2ilMaN72ou/gT7mH
Y2K8lBMDpjAnhmBKHUzt6r5W0fg7bDBWgp/04KmPPKKyowpia0A3j0D1Sxk9nrQSPRk7uX5Om05k
hGk8JkaCW2dJYk4CoFeTXkw9HSi/i1/2PznQo5P8dBQfXU2Y1/EaHvJKNAmDbMS7o/gNmS8ekMj/
27qDfGaiIvsBo0nNO35E22Hj5PuNyMHUmLY+1Sjpl3DoO7RDb228qtfEl5oSvUCyOk4reP1+fj7r
ZhkB6fwfjzTW4yhHm0MFgb5fHHO7noGmCdh9nQjTJFfpuZuRYxch+wUib1aU4vKUGP02zu9W0UmI
ZAz5U1aXiwkUz2a/YytfksKMVUUhQLTyA4osp2Vnwt++65asAIA87LTIfo96pgzaiVrft3mJ/IQx
eeAM/iQ/1yimh0z70Urj0c1hkUBs8UWMQOCaEG4Aw0Km4wOFmuKFP/M3ozPJh80Js8XDBZzioEQ3
CcGZ/hpPeAIC0pSU1cKqxe8j6fUsHDEX4GeAqxTsE5lXLTtqCXEXhD6cfyvtEVr6C9v5UeIOgZpx
lpVVz7tfpA8XLYMsPC2IqzjixnrE9zSUMBqoLEiCG90KsCGr2FiSqLtExn+uWpurk2V7ZLOMea1q
9k0JQNkaIPR56FP/Puf3hLUhaCLNeBlUkrq1YoWN9mtOL09j1IqvJopPKwKb3ghoCSgJDWmft9/f
xnqzmetZyc+y3unUFdo6k+mQItroPC+6yUJgjp2SeMdbMRPtRfdukBBxhtCLgCc2SV3fgwkZ5Sl/
Fy8JmMo7+U2mzmXG5ICzFyWt7sgYJxLgrS5ZGS29ccLuhpC7Nv3k4JUTD8kCE6vYK4/YXm6jOcYL
YAABnB8g2Z9Wfpw9dD6R8QoyUu9S8XJM7ohA7qRSt5qu7TQYy7WGEL7fbEXH7gYriyXopBQYbcJK
jOtm9x3YW5NYrqvOhU+hTp0zx4r5QP1tUlrwrAhM7cpSHA9FovoOLgEhHwmob46uKvcSN3qOOm6e
P3dqPewuuK8+ToHpuF0o5RlANwXXjrUyKTwhk61Pk5X+WXhT4WNIV9kXvrGUjlxa9qm5OQTJmIbs
t6F9i5dQXx7iF9ilwO20v7EmWt9oYh2YYIY9gdn1O8xZbYNqihjxgq3IvwM/4yTMMB6Pr5ncmbGs
hdUmQtvkPw5sC6aFRvdUqSAPLCr0hnNSIA7nCi2upVjvIH7rEz47l3H3cSc+35adX5lER3w4MGAB
QH/CcoK82Pymi+nUm8GhYxcdEQFKuhtxzRZ0C2uMXGSD0CkIhIi19ZqtMetBucyRyBs8RxS+H1YP
E7j8fOmDuyxxjOH/VpCX4PyOjIKCd6jYu/nXnhd2YFbuAmc7d+eBjmYvUGKJ7KsH3zdgVj7/wmrj
D/utpRW8DcWp0HNnOAUlmnu8R9dVrx/Q45bkBpjYNoKwfaJ0U1WmX3WUWVFwsiTvGqoNdgmjIF4W
CxFY7OzdgCcg+abc1o6CSZF0D7SoAKNIA70/Wp1e1KfJb8lWrqIGgIAJptN6bgbJHPBkslocjrVb
jpH1eIyempyq2vQcCA8C4R9HqeL4g9a9XFlHypfzZsbx6tJ5eCxaaUu/V/JB30B2ZF8oNzn+NLL4
m2iQRbimNv7cLJkl0jtmMZiApkG4Ct6WbsXVZwIKe+EQXoylqB9jzdiIZcsC23nm4kLSXeOkrfaw
t6m8jIDzZ0oxnn1XP0urK1sI25BjgEAENY0EBslr0t/3v6upCi0lNNErw0d7tmbX58aWvvEiefrE
knQdXdizuPDi+6xYO60G7RAM2Hz3iCDqqFupvEIywHItMYu3Xj2MXhFWS/WBHvlB0aJKKucTdS/3
MsiO2MXyorvgBE7NdErpcGDgs7pQJkbj5HMFTjwgOKJe1Yg+OljlvVPKSO8pBpSmcCQCsS5prFmZ
bZc15Wzzti+LmUos+GdOXaV+td8ETdIa2xZ6bvJGNFt5PsAkltIV/WHxY3p8nXeWfMmZWFC++TFv
PnIRZAfY0vpdFisBRQj6e8NNuXU8s/GBUjDBXBPVJuTvEdtxPYnlhYSR+uKJvD/9Gc/uUghAVAkd
KCHwjS82xTS9Z80iF+htMo1DiG/QTjBakvoLAatIfngYLYKe94O1r4R+RyQj0Z5JCbMbkRcfOm4O
FSJd0o8mUsNYmbQln9BUWOLYuvnL/FaUrv0jKBo/vo8vRbT5g43stdygfMz5a+TfMiZfex5REyEf
1kWCA2uA4tq44X04s4YldSB8y+c0verISZcc4Xg4DKfv2Ki54GGjZbjcbxfjU02MXyBOGgA+g3WF
PYRHuGBmdayZfoEHNI1wuR6GAHgzc7BtCJE9CpmnvKNO6tY1C66v+Hx5uCdDwnyN6eAfNI+UeBK2
EtJNWNpAG1lWZfdkekSvIGgSXTamyVoeE1I0azLFrGleYBOAibo8tG6EfAAkFVRblt60HlGLx0as
3RJCK5jzt+eA9CSWl/QdnUknMhHLzTm3is3+K9B/DZcPdGXPFP0VaxXMAirsQEJF6fKIIAuaCywL
JRLxsN7QdJsVupieX7nDdpb5wn9h3c/GYkfiwpqCDY2OZlDBVparq+e6fYKG6IGXUcOahH6jEaqE
sMkInpbAQGWMO0HG55rJ7rYs3LQBiXfoqGS4URwZVuAYNW4B1aaD3FbqciNH0dn4tVST27KRynpu
DLMyxT6e4U8N7JH6uEgXdVIe1GowQnS2xT8D/nnLg4lT069wV0+Aa1o9Abgq0ivzVq13wFnS0Iw4
Y/Y4dJ81fu7mWWQRZXZgmVif5f7m5L9vfPofUaduLAcjQwlSn/9NJVjoTcFm1IwLVwq13irBxBeP
p/lDtQyXJxR3S+2GyoWLTfOJxfiC/UDIiNcHongzvzNEkxzR0ZVhcAAcCoYY36s6ZqD0AcNfFLKF
N0S65JLgm0/UlSoW3QgeP/PcefKspXyZcuO+5l5OMocLu59hxZqOfAiOqmws9dj+FsnriKsFsf6I
+GmPFbo9mUq0nUes4BXUB+ACQus/XwrM0UJL1x3cGs6qrAFuvYc6DukRvAoSIstY3NuVQC076E4k
+OVrelap6PoOsqT0VnFFlq3gRMvWPax7PN65iLIqkLgvVd6Dxq5wRLkec8iIhKKptZg82eXna9BI
stctWSvWNxFV/EVnTLfl4evOF8t98mbTw704iCTMjCbTg9mqszucF/87i4SV/pNh5oHC3K75abnw
xAdNj+/wIHykIn/qx7+NOGsw1n0XlrNUwCHfUMfLySk/WGqBSpA/gJELVSnKykfDMwGDLG4bkYNv
SR+XVejZ52mH2Y6nYCJzASikBMsxDS5ZbsP5AYwhHHPRxwNGrS2hSRgm3BG321GppyyPCjGt/Orn
i7HawuvosZvEv+2h5lqjV62Ra2qE2+yWQfc2VHKuOGZcqElE7iuejOr6zFtXPUoinv9fNyA52HjC
L5j8ZHw4EUtEt2AlA7t8CkDX6c218HUie8E7gzjTl+V4DqhPvcRdeQn77qE/OGp61n28zg+Og2kB
V7dd5Oe8M9dO2qVtgcdb26U30+KPfggQzZ7HnIAGSFO8g18UwWPwjgwCXRQtKad19a8I9C6sWt/9
Avme5tNQRBKMvG6pfjjGrP7q4TDe32HTSRrbIf0QvSeRu5i/RAskcxt+rUzOTxE9UJgDFyqGHiyd
cDNLipo5d0rg/U0uxX5FKbgPIjUMfgIoT0RnmLOiqj2yBsFVS0FQypjmoJtTeg4/zLceViUL+3cb
gBze+2Awncq+V2EqJh4NwEDVHMRnpD1SZ0/12U4ZYZlI98yCy2FXuNz6ZAs8Q1rflMcjHkNqNy53
yudjf2L3LG/AYz/XIrJ1FXwYIvjKqqyw78juqxns9CbAk3+VRNPQXX7945tQtJqUT4ij1Hz/5mlQ
QqlEwft40XtsAabAyFkAVoL9zNvOG68wV5/JxV6r8Q+RobnPrz6ff1ucLyc0DTMybwtHCaP88ejD
PgvZt+UACPVpiBZaS7U6cPAB7pikSqdY6XfPzPakI8wJZ3/YYqD1Nx5lfgKev+rfzDs2O1zAsygA
5MsGNRLqjyQF/Hs8c9JQ4UljENOs4TBkOytrNgM1e3sqht6Dgm6g6hoStZZpZVBJGLBGq6J4KQy8
py+6jI9/+BaPCOrf443XbVPjhyOCgDnIARUs8JFKLn3y8zUMSFTckm4vZO5VwvPOn1QeJMjI19Ww
jLYI422KLVRrWZRYMm+dD3zj2Xfv5E7rsboDWyTIKKxXnG+xXnsEpSzsP6cu/bi5IZJUOoDQD+WC
RI9sWgeScnV4sTz3PyUKj0N4AJEbDrGGnPCfKHfSi+CguRKfLTf/Igk5mVJnKspLAltoM0cgLp81
0eUKzc/NJFYYY+XrX8QFZTTpx+CB+rkXHXC6SY55JRcxk5OHTdI9Eg9j/HohkyO/Jdjs2fDLFtKK
QGpd8hN0njEJ6Hhe0eSWnTCsNEITy+Iu6N7TTXyVgvHV625Yv6ifJlsA26DNj4Chrezt53Kbz30i
9lsA7o+cwjWRJBn9Jiwe4wxodVf/BeY3OQ5vR5Y+UK6jjhyYsZX/NBpF5MkgfKHxqU31a8iqXaY9
rtdDztAHUzXsi2itVzpRk1SS2ke0zB54f6t5SJGjeaemEvLx8iyzSPrDNrsVp3bEsNow/sgQypNL
ducWymHSdlE9r2p+GxBgzqk0GCM7NE9J7Dx1I8JIMV6WjTYDCeQJS8T2wkvqN8gjjVGBU5NSiDIm
mqb54knslpl9WJsftYk8oBZjOrMzZOjQyWY3Z12NYRCpRTgP3TFFBHfhsjrcx5btk3H7OkYM4QsZ
aZuvN3qZmgKfhsRW4xeGs6l3klZtcC8bkv5byj+pksirSkz1RqwFUBXilxWiYoM5pXEdwLEfCfq5
cGKI8tifoM09HuGlM6BIBOXIlErBKjes2rdiWYI1pGsr8VLqb8tI6puajVPqa+8n9KU//usX8pu6
D0Q7st0vmL7D3agh6adFmpO6e+Iyu3bZYiBO8En93AGkm0tTSstlSy6Koq9oLDDVOt7zh1aHuS38
adx5kPlJaKAWxYjshH/I69gcepCDAqa9TM3gYUyyEWq+gDEXHE5u86YQQ1SKYBzCjgn6YR7ZD6gt
wninu7Z+V8k1SqtwZXfW0QZyzmm/4DwsRiO0BOAfo7NCUfwiNLViP+WmBWaJO9slHJVyiw6/zrFF
y+ZjsrEM8WMzzWFOWQnd0wTZPXXJ+Cx6paU+L1TWH6t6cKfJ8oyxLR1ZVT2IsjoQ3RpLvekrSoYG
HdTPYEJGd17cVIgfLtgPlhH62dj9J0zRNXNVSzoJ3oW8uW2pqBytC7b4fm0DzJVqwr2xJgdJ4kT3
xLOEdU+ncx9CoY8yt639hs8g+ReoS0+uLhE2vvl96zT4sXbO6WDpnX7ejUkZhXWdoXKMI29cj6qz
s89xTQqdmM3bIsORaiaHhqUOWgK96Vz8PF+8eKeW3mQSIOjsre3mAlk2LqhNKWDBNtCfxycPwnce
Z4qzJlO7B4XegrdGoR9ZxwGq1E8QFVGd2sfsATqSXJ9qn5257oosSe9ACDiQKSVb9im0/7x2FCz/
wwEBq26rogn/BJlzLDHEYfIG3/3gnEsZmKOEozI7qD+bs16atqP1Cr4HuWQPLa2NR7iTiwE2pp3A
/Jm8TFVhIoIhUlKC7b/+QAeTbeArsyQLs7+fTanEgwuNmk+N8eY5rZGUEjJa6YHQ3AAxk4NyVHPx
znFwW43SgIDyo4pUvVXueaIUdhIRdKCE09moWNaUCA98E7bBL7WmdaIY2v5dNdkotc79+9Rmsu9K
RTlVvXRENoRqXHbCngdmATPTPfIKOD5sBlmDkjBw81MDehdpL9DBO131T+9Pv7wpZxxHapHr0143
WsBdzC6KJqMRM0hCga8RiRRtDKJdkNRyXWlNAg9MLAwukrtioI+EGvKDonlEgIr/FlLAQnww9SOA
vZlM3EbCJgoU6LVY0idXKTyZBe0pxc5FW48kFKQuOAzJDGN00c3qZHK188z7F93kW62r5xgjj1HU
a3G13EnSY0JShRUp5pgSUotPwbCyPSriS8dTEcDv4leYUsJp1ojoqrftzImQntqHeWHN6ikOPlMi
U/h1BMVRVe6df+10KqL8SvQjxVyLvffDzUlwMKCGAy0RZbuBDyMAdLUndL1Mto59+ZxVNn3vd+Ve
BDpYCp8dMuctf8u30jcxAHG06PZKDA+Z5jJs6+ZapLnodkcpVh7v3etI1LypVPjkPF40yMxC7jM3
PtP4K+rdrLSJixP6p64pLmSsSyYkSlKX2zNruZXcepJARghfxjGXOENMV0WT8A6OeMKUl8TNjW0z
sW0/wAP1yBDLococMqHL3LmCwyUj8JMSrYcudKsHjl1NXsCECFKjuV+3t7AafskaRc1SB9c6Bdax
agk/MRPtwW4oz/3OUs1nK8S0usx2lckHEFL57xm3RhMnNs5CZzxhqYqS0+6jECc33edz5mFCQL57
BbyJW119LNBoYNmp6Ye3jtQctDz9A165y7s8vGxGO+0uELMV2P0dhvOvIr50uoDbuWbyDqFBUpdK
2Wo/PlnKIYt/vY/aw1xrHbskutvLMNENrIs7JlCC3hn3857w3uGzRHuxORR6jGbfOVZ+msEkVbZx
B/02GsbRYeYLbjR9/ooxas23KXifGpArDh/i+vFE+1pmhMpCfwyBaGKdb+ZPeRoBtw1H+DSExWMG
sAcDxUVeOTrDAAz4TjyS+HDy936v2PnHzEKQ9Uu5SIBZLYePxIvkVZq6CKqdSF2ksTONvZ/ktqwV
eJJUszFYrISulDtOmKnxWwXrc2pAN4oSoZLAd9dEAdM1/ZysrRvUCb7A3bTaXJ7hDKrEBPf44gaX
ANbscbxCJCJQo1NIwaPp6nV/LhkD/VixAfiSMejVtmyuycw0YXBYC1azurnU0zpQv2iI6xTPjhkS
YhfWOfToOrHk1fRZU/ShchSY9v/fA9H1E/WbeYCh2NI+DxJDGoP2GgC1K7cMU4hxOVqOsxeGFL34
G3FBWTo2o82JD27zu5jSL0fWXs2BdlYp8rZZRso0VJiV+l2wWcIYQyUyyHOPD6vxQN2uxI3jalYx
9IQi9NCQXr65KFXSFP+ecvAyfWCSyRjafHm8/mjUDMkJUbhyIaormXylJCARWzB5RIXP0TDZxTNJ
CmmOcDNU6MRkpFyprIo8BHG+LPKCMLPDzFp8l3L+gwVw/Auupm8Z0667IH4PlTozkfoqCS4gzQ4j
DUU5o7bf7i3mCL2gsYw2QJ1B9yIQhJFpa7p2dS4yL8VWckZke0+I8WHJxZQobbk0EpQJ7VsjrMAJ
KLrXORdmUlXSEA97A7sYwtQRde850tYTaIB8b96cTy+gSauQzjNM2Qmmgcm8zAeRZxQ9X9Khk0ww
9LTbKtqxsY4Y30329tYLjyXZWdUerYIwwG5Ak5cR1hVHHNObN0gzIv5R/VxFVXk5MgE1/p03sFY5
y+/OtFEFlZDo84c50X5frYylZBYCgLoxwgqW8CRHtSo7hdwhkU3PIBT8N+8VMmKtPcCQFKXNHWbE
6svW8XaV+Mdgmy7ajkhxjMz70pnDIbBHTPAM8UN8jGazXB0uyRe/NbyISGADg7TNlWm+Pkg0n5+P
0qfhFSuQZSXGqNhr6tYKELRT9qNuIKVaJXJOG7VjINMYGfxC1h/XcQN6r9WbSAfVS4XhCKYjGzDK
8BEt5rEHIlq/6EBUlQoYcmpVQB/YTFiH4yWx6F7Nbzikrl9CM3imSqznn8KhIrWDl92NJje4d6YU
IEcgE9BVwCPDdknB3Jchw1Q8BcHlJ0fPBQ/CcRcG6vX63JBEp7foJwr0/+lxX/j+Sbzq67DYaItX
nC/8ec1uEXEU2dpSuIvJ2QkDI2JJ6bhhGrQTYyIsR4HWkvDKlFUhhewnerfISqxc4ssP63B7Ej9X
hWqdjp76+/56huBjsBa7pIEeE75S1h3g7GEzGjDXfEtnySDv08GaBx8tsRfuKAOkSi9BcFbPNuxh
ayq2RhnQViJMowYsMr4EoPsgFWGH0zATirBxQbidCCcs96pFxbH9/7p6GKRHNQVDpZXdVKIzOlwI
p9IoIE8OQUCukU4XtYO4Bjag7Zovh98vQnWnPfEt4VdHZ1MBb9Vx+UtWo2q0cRsyRQwpmU5kUJ3t
iw2VpPowYplv00brhfg8fDejAo1Yu36lE9A11GVR/uZJWdFFLqjFe2hEO6Y1ukkQnjoOEhXaYoHa
yRAWaN7ih0+LgoqWq9Afc65AVRoo6BUl3Sl58LoK7U6QQY3rwPHOKVicvMx7kNBVjQ2edM4XTt9L
nttKUCNKeekR1hVN5OQBU9QWEz4B/GOpMTGhgJcCVUXlZjFntOP1BeFHOPmDKfD49Gy5E3Hm6OUc
20fyl3E8ySLoKCVuoKN00+SPCMJIWb29LM6Uv6LosWkSnu9PzpK6n3xf1hiOFIosVJyE4v0aBaRv
YaA2XgM7SLYE2vg1myyCGXjPaCyN04ajXw2HLVNacoByq2Hi+6L0WVuanx11oRgKyty7POGa8arh
wfSjmhDDQ3AFavcm+jyTRwLf16yrJjQNBUec0XT4o5VY5YsYpMEQ+JoCH4avKyuSZHB60sxRt5jo
8DhRaig3lr6Qqhj5WwR5YlTvTWdQseE8ayxk7SZ94wpGb904mLb+xd3wYpZM5u/V27AyhwXjHetW
Kj+XZLq1kEXSeMkH7VaTwEU37jXZteq2OxKMNrVxFmQ3kF38D8aeEsvCyMBFjStuF4+vgokbUkBA
HCfNzkuMaw5oVeCuTQY8n0PEJKX5CzZb7jsn6phO4SLakkxGhUcF+20m3qOopgzn/NtaXBdCCEZS
1giZGg+5hDZ6jvB9IdbwUTlc219Uj20fSUHmMZBpgNf+zfI2wY4PooItrey+cMtWR1MjKjoEhA5a
viZTiYCrCWAO9KQ3BYUyeMjS4FYUMRFFSBzE4XnRWxao6iXg9+ICMWwRBlMxQg4mJm/CNR7DWunL
2UeT7cECBdd/xZRY0cx6ZVy0HujVNJGDQ/HFI2HF+yl+1GVT0Ddpp2IcKSDUi6++hRKWZxYOm1AY
lPDap1QqJ99l2EUQW3Q+dGksYIQtO8jy3YYuS2vqoSkFjNsaEznPM6R6Xtys6cg4lIzSkGj25RkQ
EyMG9JfKUwDAfE6y0GyqRZogmGe4123Jhf0lJvNlrPhjBOd/0Z+/7JdJy1f2pPY7KytNLNExG26X
0B69B8GAqm/2khz2PLurng8toaqCnAJO8zCayTMm83TFlH9FjiA/0Bkdjc3TYGq9HJ0Q2ZwMivBR
8WqqfrDg5qt5VRDZD01D1y1WcUwcdjZbGI9+3llk6eqfqAJb7zL4pkCBqSnOXdz5bSQ0ywrR/2xa
X7OklY8aomVyFpFK/3VNlQgbcIZcspvN5C7qUlRpYPS/RjxhlmCLVarQEWEHvLLgfFl93gGcs1Tn
34dM5slCeoKM0dtv4kxQRzkDnXD7bc8r8ECt8nhiY2kHss4+HfWUso1BUXdscWS1GFRIOEdHuq4n
unhFZ/dLn3p3NjxVKyL8thBg8ErBndWXghzs0AKEF69D4hLva8Tg14v5A//0KhyPtZxiEJuGv5Sw
7bCPJecgfiOU+/Vw2D/Y8UuECwGzI9Di6bZbYm9+KT3j1H8wSH0pZqVRX+gebEGXsJUQHRlO6MwW
9SezTP9CMLOkjQE/DfxWmcoSkGPWNb4YG02i7pO6ZsGMR0ho6m4h60AGnSjB4d5rq7QM43FzyqEH
RO7g/9emAosmEu9Keb62qdsM3DvqvJsrgPrHUUnfRxux4v2InCMyBh9s+BHBAKIglgPfDmvJQ5/e
KNyVPYJp3A5HZKK3K63xsYmPxCh4g/oDeU1QMdNbZtbyOuL243hD5QGA3RPwMz9fuE6Hp6jZ56k3
5+NVWP4MTsESlVCyHXn7XnuNoZXdn6qsikVL+KNEkUCJMeE0HRRtTP1cVP8DJVPX1EgCYRdZTWXk
13PjjPGNB75a/SQMdEKSdMj8JKjo8jW1nx9BDb5ZtzK/owcFNkfo0ZnTLXH+cjj6460lO7zOZNKf
L2wqsgnry23lFe7egNlYBsH0fpvdSm/LFxB6/mNwOpg+OItgaMuoSenqL2YkQ1EgC2EqURJgn0rK
91tx9i/q9hjLT3w9jxU0go00a829CTehVIlrrglUQdVdu8Fa0iVW2l5+AxNeIODUUK/xxuREbxy2
uCKbxYNvzlJ7SWjK14/RbQyVD9s3jVwG+pOYp13zvHSv3QdgTLqt5ALLu59R0+7tibWHpNeGshMs
BDBehLw4fP27L/mHO7T32joCVFaJUu4HtRaPLShOfnMl0ANCAMdfmbVFgVChCZs8wqb6Tw1Zrt8o
+Sgcb/SKy9RVWmKFdLobJrxgRfdGxzLjrWWc73xNKN9hKzFa1fl+n7Gm3uTkGmYVpivoDve2DIjU
+Px684d5qulMPYY+OP2KobZPlSeTVv1t2yQMj2Y5dvuV3U5RAgz32BwSlNMdwU/hW9OOjbarhGav
LnyTp+zTxemgJFv4b/Uy1weWrXKTwvzfYjgVuXaATr0MIz7GY9VM4Xue7wnWcNdB81nbZAb55E3z
e/rrbXEJr37RvxdEFDJaWRHImRHAG/pQ2i7l7sVFmIILD6I4pmrJDWB8e0Joz0H5tzTJuikzbRRA
y0eg92Xiq1Rx6TCokkrt6b/U2cykY+Y7rk+Y6Y6+ymQ+nvoz6Sk3AHU31Gg5qk1iysg5LbtD+Fpw
KqbY1lMGatEdbz0rPPuOrNj21YL7ucMU6Iq0c0kokVLQXIyeqnvzzzpODGmnRoFaR4/Snlq6piTe
qv0VMOUtlwMCJzD0fXvvJpdO6ea81QyMI5DtGhlaKrR4AAJf+76z83Xk9LExE9vKkSjc2xyHy1n0
2Ng0Ke5DocSwm1e+bZMHJJ4eQE0xQ1oOvzWVS+Nr5RGWXBflhQtip+5WOqTdRE2FRdplzJ4HGlhc
4p3HZzkEL4QKMT8/BGmEBz6FknHu6x40ymxPntTZVzt+eOX8slhHO762VQsatWJaWPHsno2VLiLQ
GlhOvhvMNAPEmyOTo/T8srsaJxr4s2LgMBeBxfsEdLJMPZpTDADPOGIIgornx9OeE+fGmPvpeR2N
ly5J8SJmjjbt3shK5IqH8fXUwheblwqqRnncHBjQ0c2DOMKH1l0rhrGQLZvBV447NiKnbarLf/r6
Gj/Edtvo2eulOWcLaXKHdSkx89VaHpNaUj+MCkvT/SbRxHTUkojwIgqW/nSk/fw2h/0GN+csCza4
7/gKU4RIRgISvQ+L53Yxl2Pq0u+2qSa0A5F6em7N8opUlswUb6Rd3scJodwTJa8XWFpgboJBDNme
aCwD8dcuVtrvgmgC9FWajPWSKVaYK5biMfRCsa9i8XCuWovZ+IPDjo6I41UzDdQDfpCKeISDCPg1
B/71EXcNtDYzAAg40FXOJCvr7WbtUY0S2KPuy2UCRVO8abMXJiAOwOOoW+jJH58tOrZvj8B8o53X
/P6ohhexPa7g4YEPVsVs4ZJz/YvEEQ8KeyjWPE9FyjAL+nGWZsj5G1Cz5QJUD+Aq1s71ekN6GAAd
H2fStuEhI59alxqXPmGjpS7hkxlf2DwLJLjacPs96tnfPlEVWkOSRLYWlCj0Wkqxq/WEx++/XOKU
ToV2bJf7GI255blw4JZmzqWmGmP2vMnCto+7jfHyKfWcGkZ0129VY9eATLTwHGv6UtwjwoP2f2zf
o76ElaRn3BuRTnsCtVUOwinhzlybzLlLNzHdUGNuljqhR1lSE2aPvhinGPUGPfa0T6hjJadW/xIb
ab2eSB4RHPldvPCpWwcEmkOgj1qF4WWD/5KeVk59OrxpoZ22RBIhoXFWaja3Xp+5LNX/+yfmnuiN
0HVPRj3VDcyuXrnH+hD0olgVNtnvJd8938MllSpB4eZVCU/EzlGNJvN9isyxm8kFR+gBMY7wF3c0
6nVw1dvztTh3O0uSg2aUybsdm3j4T0w4bKxP7ShmlzJUCe1OFNv9ErBlZWCq1leJlbksbttsfOv9
75+WwpfeYi6S15w/VGPfY4OUJJFe7ZXA+nMmwOnhLA5mseI4IemcbGlJ5MTIgsT2vezk+LDdokQU
6oUdxFnskRjfyJz99//Jk+LHmwEW0vqtAL794Q2qhGHE72d+QyYfihQdxOqTwZSlvsYYVdwuOkYD
MdzefkTZBecY07EvGMQuMKwM8OMhZDutyHUjBocDTSdSx9Iuyw4kVHB/3JT5hXOO/GzgNhFt/hY7
a3Rz97xSmkEi/VslbdcNL7ZIsQ/mN7PiwX6plI7BM/mUd0ThSpD9QotSZoRRDhjNQ1JGoxJGhSpt
Axf/x3gXXIz9BY0OPShNndQkggIuzH1t148SkNQABVeDxI8x9/MJn2iBk8X6aLY5jS1xgqXBdEnh
2MSLoxVOtO5HPjlfmGunEOU1JIQ8XbGCtbHl/HVWpbPHXEHKSivga6h9ZWyn38IqNBNK/8pepjln
h+xH75rPXG6us+Sdzn/YalroPgeqd5luyg7yJcJWupxrqdrXykpr0gP8k9ZMXhSJa8hzx6MQlc9P
ujwYSRvfDz+ytw+wnOwxeE0U3bo4iTRP5ZZA+NaBj7zOozj7O8u+cm7f2Kn12aP92iWErgIToYIr
Rvd0iVEyU/nlE/E9/aWG8WDuQBufWAE6BUAY6JflgDfyNxyBk/QB3OE1b9lGG81ggRtwwTyxdT2w
79rCkPBYT2u32c3A0/ApAmKCUVto6/72sWyk/BL4+kBE7644GUrDFD+byGS/h+KuQ6PA7V4n1KfS
OV/e63ghB645TLq0ZHlKXYplw/IkWMbz8bAM6JSGAviCKTC0T8u7c/MK0V5wMygbBVo6SgjN/qFJ
B99KQc7YtKkW6iRHSAxmXTYCpgeArcAnBglAXKqBMenKSrWBpjWprgSN2aMFVJjeNzIvGt1e8s+U
Tfe2KiMOknDOf58QRKYLUxqQ/YuKN4N3uLyW1E8GCA37MvWJMLwNbFL3d++0+I4w+BZeue4aBHSF
cxgJPpmU+hoFpWtzaH0BtruFufTsKsKD6L028fPznUEcr8q4C38NhzGCT1HSuTjib4LOPb+eLTUz
hkqT56HALeqw7Zedi1/V/+y/97Nvq4CE6T0AuY5G5DH3Z77kHknPvudRalxGIAT1VG+GJXMTOnV6
eI/PD1I+3l0dI3DPJv9bgZOf/GU4hX+lt8iYLQWCviIB0kOJ7TW0Pq9tzaMlT1cjKcPClz6kMkMm
7rQAdQqLkR6HsXh0xq33bdkNAPkacju0P/Yp04s7Uw4NP5Odfr4zTn8f2if8OJ98YWPMhqRMLv/y
KQTCSHpJs1748bUt0B3495r89EVgtLyyuGt332zl8JnEZX5YiJdJymd/3zomwMRPsa3wcXHadQtj
4NWs3V+YcSZxEFNOxFHGiG7lvaM8VJallG1a+QIcx49wOtfwuRozK3XMichQJS8dJoOfvZzYLPRi
VpgIBfeyfuC6Fv3TbkJxCxGaoZPlc7TYRwnLH6/tJTUAsD15SVO4zs9s1g6AQS7ZHFmVo4SECfOP
08D6bagqSjoQd/XroUSPioYcORSoLPDHIi43yq2qdwlXzreogLpxWndPRriLFsCBRnX/7GJlfRoC
ckh2v8QX9A+XB8I2WDOsqE/EJhTN0hAoGWu5IvbJwp/mrUYfJiXLnZWcJ2ihUk4UvNb8zWM8FNGo
frh2EkgLqyLjCq6TVNL3EhQ+CE23Ddod1QVBiS5EGqKjwTXNB0bTyqfg/cD9b4buhRiwpZZZgG1F
8oUzPSkBTGW5U+GlVUSNw+vwTJYgqhqtmMQZTdCbdKJVis7w1EaS1obeK8PQ52seG7FosLY+Bmj2
nrwtCVrXpnzh+lNVA8s5UdlmqYm2wVuEMTIFPygGSdxImkeaQrbD0OOdT875RZF74gJhkblu8nyn
7kIirbNz+GPF5bEO4ipmSONacgj9R5RaYDitys1xTta+cglJTtmm+L0LsCxHgnvjP+3JvfsBACf/
9gsC560Hs4VmedQcKbVWBiCKoCL4t1W6YC61eeRkO/+TcEpQVFZfu3lmATJPRs+j4R6SCInzKKPJ
NsANI587laLfNRewhWMKixG3YqEV/e6WbJREcDRxIxcdWu9xysofGJBafCgWg5sAF5n46kve9rOn
2ADpqKRmNmKK6JTrhkeJrqnT+SJVJUG+t4W9UPx5HkW+nu/vpRFUBUbN3icOHckhNSHcf/nTIZTP
Ozl4WP9pN3wD/hMUAL7wpFBhsGv9vvTktAtWIMVeEgdQqBQ311nbpT7MvEH1wHyQYg/pzpn5vzEV
pHt3WIgT8YaMPtzIrtouUJkjIHlbx7vjPqAPPHtl5vv2MNzAPNHDB+SnEhiBshe3SgfajWTO99UD
4XExVcPjA6NRhFIrRt/Fu4VkZHaMZCbiLXAbjHGbOSD1AY2l+lbI6uVLluhjrgoNflo6weoZI6v6
0o3ThPlBP+8A0zFti04I9elA6ETnOSzVcbcM+BeeO2jL2jN6jvUpjIpmG91sZC67wAAr7kZKSSkc
bKeA+Wfnv0pc3SImATzAiBicFtBmeLHxRYV0WjuRMjCzrrpxYjhYbmPYwBX8R6b0XHaGIG8e/0FQ
ZSJzyCsumjc2JSbMhRK/5MGXyu0VNS0ZBrntR7a3hLPZEW0VqiK3mugqdsWRX+40DmKAY3WR/5l6
XVQ73rZOb1YKuvSYGkow4F8M8GGFynCSqWepQkGYYckYWZQddbYLpnzgXDGy0Oe515rZygAibNUW
2Erp0Pnz5AQ37N+ll+ANJSFkZuaYrfcKscu5vj6kES7AWUSZBmIGC6GD7ll3mglM16NdyhyoHJjv
JxLz/m1+bbnbzGyYGW9+lcJuczfGiK5KQMACxbZ2LRwy/W52qowyeZPhiKVWdoqN/IYLJKwkybId
LKSujeWoNKDiI4FkWybCajKQJUh9x06HewYJNaPH0J7uthKk3bC8jww0NVru6f5/Oq9VaGHaYObz
V89o6WoyF3eypkMrv60ekBZ+imlLs+GAsFTM4NXUckf/2TFks2uatTllhrNicnxkn6ARcUoTEIiU
zRF3cHznU0pQ2QP7ILJvX3eSe8V/9eUUDnF7cU+2WwcRqpn0a2wsslGUthyidNj7bX1Ik/y7uzrH
sb8tVZ/RxGJNcy70FHJNskjCciOyBWdWiNTyRgFmmKFShYQbDNYOM4OIwhVqmOxWyBpA9yLk2jas
i6xwZPKwhxEf//q/vJ2Nl/lTb2AumOKsp2zRN9ApFZrte7iEHkaVBOv8PmOfrqK9dc21TQmJ4z/E
YeKKAshGKSTS0bQiTauaQ5gkx0UZwnvmBKnWYZOteuKOkiI1oR2WiegscrUZv48ikP8+ymLPkK/C
TX4s4s6c5g6kwT68d0yIIjAvNsotfBPBVA2EJW4LS7eXm194zh1P789pWl62JopOZ5LgUDNELnVg
vWmveESD7+j79RNJ9K+1HMhtfVUAepNN9idx2YHMnplnJ8SYPzeumVgMYZ35zfvo2aUA90dFFpjJ
0Wi6NCaWkUjdzM6+rx+f+VVHfpZSSa6wpno3p+cCNQ3RoNJSuU1Huie+V9f9128dFpsWBn36hTpe
zUjTUzknxgzd3C0VcNbsSO7rs7KoMxX+U8+7Yb/etnCZe5dWe7eOV8gTPNHJiSq97BAjbBgiwcMM
eiFNn8xcjMBGHyFxhtBpZyJ9LzsWRY/ZuTJtFjRGGiG0m1L6T0KYeS0dHkIOswKO+5X1fVVz/Rue
h9UYsriqOwJbCof7vGsJILcqr9CbmKJkZ0M1qN7gXvkzLmgPWG3q5ZzW1a07j20ok7+liW0Da9s+
ytnjAse2icQjtS/83kpZ+MED4PRTyQgv3KIYEtRFqo8dTaMLnJDeOAA2AiEsqfgx2mRn0tjFVfJx
80XDXz3BUtCqfYBhTyZbSG8nIxDVwyJqswg0uiPcp8PEgxWpvogzYd3aiGVzIqhCZ27IeEus3jMI
rP7Brb9wSxiI/XcVYzsoHfh5YhC1VhFzVsYsWKuyTjsAxMdk5ZqBM+bAyw3fokUyuR+QBZzHipJa
ktDGphZ2qey+Od6jTn/Uirz0+51nDCTDgTOZkvJSvKfqH95Uej/qa68IszJXUAyEywEfeiWnyL2o
qbYwlHJjS/ITOfKeMbNwvz2D/KACyN61vfqFpcKDEss0/rX+e3FrefPO3NeNuajaXBkmQWuR5/yg
ABm7SiFzL52DEAtn9gvHFYvdCS4VpnJPtK8iw3pJ8NRScNBp7gMGWqVHXRQL5HGot/eewzsnbegS
bVkV57HHBHC6HLCbfsQZgWIsapxq2iv/xiW2vwCp5jWnvh8od33mSNsNgtL1OMTcg/gFLDuws9Gu
53wobvbwYBjIfVv8g0IEGpraZZ5HouG4YkQ631ifjRjNu2+guUUTt0boiC4ctjKAIR5lqFhumXgz
F52nsZG8Cx19I/B6CSVlpUhCk1PYOi3D1nHko1IV6Xvsi54TF8a17eNuIhf4SyLqMWXJHT3NV6Op
y+T1hsGQGJG3ERYI6gWTJRTKYvFGKtmGY0TmtqFGxiu9ah/lV9wKy7yJAykEJ+zNGSc+z1ZpVjrU
C+YRc7JH3x9La6j25QxS5ZUe3BacBqPJUSDiHzc3FGUO2xTYqp+AjdWvrCSjtW4Jw/0fCTu8FCA8
51cHw6Oh6evKv2WNkianFh9ULAk9GHs21IWHXvFvj/njRedxLvtuwEQzAuaJrdLCyPMxEUy8ZCcN
e44ZzZUXetd0DZa9ve2l/LwPBr06nA/YwEaXPgviLxF13te4uL9zf3vdVsbdv9Gj0Zx0vSJOQSYD
/f+cwRMcR8MD814gqiGxtTPfUMCVU0R4U3oTajlB6e7VUM+YYQJ+0num0y37f5ALhnGRSJuQsh1x
GyhctR9Y43CB+S1iSPVfS146BCkhrh7hwQCtg1bAhh4HiAHb5o/J6iej/qKhdagR9pttksF/Xn2e
04trpougXq8l5US0vrbGPIed1TnR6tyE4F+EN3WkxUi99NQXqHfbOm4DJPy8pSBhzt7x2BNEdghn
mI79l8lF/4o1/hOWLHnPFArgDyPgaVcWx+aB+IMihNMeHfO6BIlDGRW6J44DDo1v145Yzv50WkrI
qGu7sxuXMXa1SXu/igWbOkpsYiGvWZEzZRJG2unMaLkAVzvy90sNf56FglUE59Ys7X9PNe2Itd+P
mvY1/8E/WXA3Qvl9X8TUUy/prxbtAmEoB8vePUZvUwMCpC2QOAJjN/qIzPsNhCqNmxcalV30jveb
5Xet6jrYHPHy6JpgRjTVhUKbP3i7bCbb23He3P+UYQ05a2soH0Pj/Q/QAs+ZbcPEwrUugXA2VZl5
iGq9JFW9gZz9FoqWsxAKC+ww0WvDuQpTNhyoGGQOG98es/Dt9kwK69HQGhlaWQzwPifRQGdyYNvR
l2Um1WUER59uSYNpiOWJcagN44Bon2pJ0qnF9dg1rvTJHYfGDQeiLYiqu8wHGVYn+d6IoUVNEK4L
yZSpSrvsKjrTLSH0mMH/uGFv5zlnzjEImkyyA7J0HFZxOX+vtlmvQWqjAiRI+ljaFhtW2g7Eui8L
YwVAUSNayQaU4/eZi2yXwpx2oOnvJNkCviVJ1agKDUCSKE4xtZneiBfb/Wd8dXl+SI3XZNxf6RZd
B+3MHwAB5BusV/CTc6bIqbQAMlOkZDQBUTox81ogt0aQCqVeRn5rokvRdfUfWDWBcnJBirghvPXG
d+01uW9yy/tDi81poy7sHAn81h7N5IB8+dQ7LuweuRpS+vAF2onYIghqUnbYGL90NPFLPUbCikmC
Yr1QAHIoq+ZGUuQXz6BCl2fckVDEO9R9NXL29fD4q4qP3WbPDQ2OrTb5EjJF4zCHVEw7CAg39PTr
t3bFO4Gu5SQ6g9S9VcI2rU6RhInLg8tX1MCblWkgfKarBvB7Gbn0pV4K5vGn0e1bsLQ//6MQdprD
DZ/allABO5EbU7vvJiWcIYWb4UNSbvZWFM2P/21MrPxLXWY/ZRtEeHMJqvXcS6S3Eli84scRa+fK
Bojvxgl7lVkWpf2QtD/OcI3RinpDTxlT9sVcKJ9x5Ij9Ht9k3ftoYeCQP6F6625u2bP2v8ZSGpRr
2rA7xZPFNFaOaHff9jPrP0ThTbWvXsC/1a78POaQVA8fR9JLDCU87LI0zjHhsrleZJrRx+YKVfe2
kmHDO/pbN3Pys3eqxZRCcFv7/xt7j/42B6M829Cd3QDK7sjQdrjHZYvwDTlxne3DvqPznuM4tYan
OugXxMeUM9f+QulCfg/AqyKhcrbzg0rnPozjbrSWaJfdlIuCZiW2mt1TbkHlfKyPBqko5ooivNWk
huuictYxGghqm0qHi6DXyU9OB5r5JF0/AcJhDalvkBl3mg5oALlQzrSmTYXdtegOiYkYfLlLT8wW
G57htOpUCOJM8J2Lgq+5U+BqSk4SrO2tvwDjefUUQ8ETTNTTiepwrgh8t1Bh44C9wAz/PUXWIMcF
YqZzHNf4qBDhyO73p39lG7kFrdYnU5Bvc5hnqf+XFxJkdRhlW8eP7Te5Pln3t6FOPM5XHaEImL8V
VCWRAdtosNFaaiOHlrvpCf54+2RFAnQik/OjsyOlglpZq6gdVvnh4bW7eOHnVLxZy9fyFYxZyd9X
PMcmWt56KjrnOyPJsrshcgyF7b3PRSTy4v9irg3yaIfmXVt16picKhgy5nr3ix8YiTseSMKDAxbO
pQdJFXLjxhXH8kXfJdDFBtd/0Jz3Nss+c8iMcZwFRrUosk2UQr5Tq1+RWyxYahv+WbMhNxwWNTci
WCadBfZ9GU1B6Hi68D2cls4K71FBU/IM06VHH4+/T2pNU5ovSO8xptBCIxAZ88LVywtAvsfrzc69
CFb8WCJXxmaWPTd1t6pQM9V3LiZkThjQzyGXcK4zKTk6gFdM+ziom9cnyj5RxVlxj6/MEHQzS/WN
tS/CCU7uzv4P+lsI+oHfzMNl5sYmCl8S4BjEh51Xe3AfssrvBbx4NdBxNZQsrX8DtTvPwF1/u/D7
zdYUq/XnPVNeMF8YNbEIYNERQGyBFYoKOojXTMB6MZ2MOkukHJhjebC7kmW4UdYc3XAsI9POB8ch
qs2PNL5s9Mps6QAnKJ558MuPi8UAyUkJqRyFKcCA0JH4ylnDBEm4zjTLbByoJccYQtletls4T2fh
QrCSUWg0/+MSElbH7AjScfJcNryyztXMGiMLMWmHBJk5RtMbIAIl3tcezGPZyDsPghiANjyjeltI
hQqikHCUh9WEbuIgOJ2m8K9/h006hRsbLrACkxzNF23K61o1knXRujnyR9b9AVlxLAvwGhjSq7Ko
XY8kpWrdJTnJGOlv+Q7uiJ0KUTXHuQ38UhRQ5Klxs8Q9kEnPh/9RfWR6Zx9+gZI6DtdhSZgJvfDy
N6bJ8ZlI3s0l7MG1Oh5i5TH7cizMYT2P5B2T/XWWXUv4cdL4n3e6mvLHm0thaWUytog+g5LosivM
OCRwEqGfiQUKlf86ds/o9FwAAJ5UnYHnlHu20i1fOhat0XUJKLhQ+jzMkQY/rqxiR4eG2CHKYeva
XObFCre1Rlm9NPUQUfwRoiC9obrov+CNyUfHAac0p7x2/N+JFvUVrIc+ZkEsU+pHWovq6YZllUQr
isyfkmziQPjBSpBxpiqehjONxTCOD7r785L04RdKVSMiU6AFheCo5tSWcUUCRtMKWepswyZxxsrl
Js97DA4Wo5fK0K+efjPPQ3CSiVHCElFDRoIvOBKh89EfM7V7eY57vN6SPYoEHW4AnypS2N+fShPx
KRTrxLqHZfPkcyeXjoaISQ3WbECj0ga6y4jSNSzneswO93Bdvi4tYQCt2GIfIoIKpmODRvwKLw0d
iPah9LPvqvpQ8Pl8IR52hfZqyzY1qLJdK0T2d+/N/GvRtJs6a9GLsUp5oXufja7t4ga5S4v0L31b
/PH89gnhbX21KK9tIpdm1X8PmEKj8KS80WlygzUXymxmxpOikfqxS1FDgZgkmpyX9y1N2sbvMcNC
llmu1tHzOBFmGGmLcvKNyVPUB5buLJWeNpDGD2JXEgB+MsCZxrMpWqkHx4tOdkLYuKOHH1y50GI3
24vVjcdGr3xfSqv/UcyZDSJzrrOcPfvb6ZFAXxWXx4yxX+A9n3YLeUytLVyhkTe6Mk57Ym1vG1bv
bekbb9sP/NZG1QNMbOYc2z3Ejxb/KnYbCrqokWnYMOli745VRbtHHVmVz1MdzrQZHBIQ+e3We8JE
VrxhXNC3P6snj1OckzGoxErepp7nKrJUTaIKxcKmihS//vLeEIO+wy5Y7umEIwvM1+ajl6bnLeTM
MZxn3ZCr61pH4KWA/W+PFSFnM1HqDzD0GG4ljb+3Y46FpEBDSM8dXAim9d+NstV3l6XU+USgr2pI
j9x/e7AAZmZn93eigC4BATY3Et8z52IPHz8gWCtyiSN3bYEW/vSy+NUJ5vEF8hYLGmtfFUJaB1NI
lucxBebFZ4SMCVxbM0qiKaSG+FtoY0qCldDfXfM45wV+GTLMmo0ImQy4zw+Puj4USKF6D5JYtWUu
fObTcOpLC68xYYVe6y6Q/rryEb2AryjQ6YmsIZoS7ANZ6loyeDojkwzLVoXLTT6/N5+BQmXd4o7w
OrMYGslu5qBiwt5vYlb0OmDmO0n+BeU0gN6zu3T/r6+cmb2G2RvjHVZZ4cXFzvcyyQr36wlCFJyo
n5nFoha1TUe+w4KnyjdABifSdsHPyiCUQL+QnJiS/V17HDdnALHju61v6B0+pI3i9HswUjr4ZUqp
4kQB6QriKGrxKkjf8yLe0mJGCW1VgN9LHqQz+A0bsBzJJpySue7gT9Pb7sZaHyWYeziuQuZVww64
UeZgDJ3LW6lMPIzyFNjc/e/dSYVsf+3dO5dsqQlW+SOMtSanW1r46Omkg5t6zfx0jqT1Xvv1PZu+
qoD1bNcmjvFz081TOHpwSch2IDbYp0x6rtNUeMLYuLjpIskXirOQgKKbRTG4qkWSDhh0SPBqNYDV
0G7Wnr95qHiHiZy7pD9IivfNnqoxgCs3kUNtfXNDoCgnu72gcQ3pp1p4jZjnJ6lgd5wXm7u8Vf6i
dZsAYhuacQ9RwhbdvKyP9xUW7fJ3OEuFAhBedNwoeBx2d+n0Rap+Ds+1oxBKne0btWbUkrcXlSqM
DieIZ6JhNLZ7TDiy14kF029U5SI7Fbt4R3YUiIaYubzPWfufCWFvUS92Hesn+YoxYHUs1PALiSDk
PdGvuZop3xcOpgP3YrJqo8brTmuxLUPeio235SGECR5gnxf7jGom/wXkFDxx4mWVlvg2N+0BlXpx
ulGvfHWUEyIodk+t3fOYykg9fy5G7xNU52kw5cOIHkP6JIIytOgmi/S5RuG3vCZgND7Jre1TsGQE
Mx9vcmajMg/MO82iTAn2l9M3bb0hGS2wTwRWxLZudLLg5aBVCz4RVEk5Ktz6sEOQcw/lBGl8tW7h
yTfKioMQhbb3GiKpNOh123/o9qVzCnG28wiUe9lLSt4PWfZblFnkGlB0gYnTwTZlLD585XtJ+Kh6
be6TcKAB3HPWg1Z4dco+XiV8JWCk4OHrr9cupf68CoRu2NNHtgsl6Wtfwx4DzrlA5vFP7FofdO4t
uNztnPr25IEFxlkfrAtict3hbe9GPDvU047T/AbY5B0faEGmd2rcCiSuBGQxvcNofibEoAebAIkq
8QSScV7tFC9sXxoWWYL7Yg6WeFm+CqziNyyqwnYKoNMQAIPkQQ4VSluuCFPuX5EpQnfvRTQVt5XS
q5Vh3DCdm47Z0P2/xBAWOtaoOFoBffCeDRixCnhO+E0Qhkc0pbOshS/UNZNNePfOYnUVpTbxiAz3
LUmyAbxyC2LZ3NgfdUU28MFjvCvGlMOVb9d1QMLsbDlRqAcPCt8W294vYFIXsppCDeyp5GWpaXur
jT+c3ZYryRUXDo2lJjICoV6zhXhkq/5GcDnb3Z9HZg8+HrF46Ql06O1t/ZibSWtvE67gO/1TpcLs
t5AxDaxt9+4y4tbFRd7wmzMST/BPLAyQkQV/0v8BIVBG0lmScva+zq+E1+TNDV5jymQ/VJgVA/Di
nHl/Kfvx/OqEhBvLMibEhek2XzmwqYQ3Wu/4Zbiu+8kbwojcXaCBV9GVayYZc0deBqIAQX4U0i6F
nSjsz56sVDikzzaFLBRD9H9tJpPzPmrU8wNZ222wTaE+5jQoxvhT/5jlxSz99kPlIqSzA8nhoGMz
RmgJFe++LAMerYr16FiA8zVnmpJvgii8zcqe6LSLPCLjjC64l9a2QiojZPr/hZv7C2Prfyw+7cNV
i/xYFatfIGqfiHw1fMrpZjq9mJXNpi1nMi1ryKTLld4zRJ1TlPLcu/UPB5OBt2Aw3h51fcq+Z/aj
mqP6fhuSHIfvDbAKuWuxdUbC2tobrw+qfm+rWrmn+BfX5XDLdx1tmyf+lVo6XcSPj4W9HpCidaAR
Hi6JYDnYviSTOtMz3YzPHSyFodPG/4AJHXbmyZxc2FkQ+7XxcfQFhoNGG1ORuF582+4tH3BYjlcy
i8Ce9RefEMkmyvvLSMlq5H2spmBWZ1MI5XEM3U9vVJeGzjw+YFkmh/m14Cxcyar7Fn5H8mDIEZtE
Jd0EdBmLbOVYDh2X1rK091P1ZJqfNv4vDCVOYuP9+G6y8UZ56c1tdCvKB2U5R96aqCGSIC0DddNA
jQrXheDijgdRiYdpFjENhB/+fin6NLGaex3CX3Zopq0Bxmqn4Jiw2Kw3l7WWfTRUywvNDTe12ni8
mt7sRUFThNg3qAXmcwBQzTx/4cDpHtrS5cv8J6zqvzAQMEOwRvOCMllstgqXXTiEA/WOztZnlYev
DI1GYPGEmMIUIEEdnR1KT+BMAbOEU58yt+4sa/NfJacKEzGAjGgyc5tt4cRMSCDrR7K8J99EQvCi
F4EtVCOEp0g9FjIZQSoQqbdrrGaIZO0wjurCf/DH8W2/TG4mKDnQtAbJeyYxKvFomnJ1iIxXL2Qa
gFbPi6yy/W2NRqMS+wmDfvQpPdSZyBJ9zr53St7ggXLSpknOfPDgiR6Uvaf2/8VgnFowzAVq4Ap/
+p4T6xtOw3GEzE+NS486nCRqrdJ6n1ElLzdtSEBskiJi5LsKl8ghkS4VB5rWkFdsP+ApA7bL4B72
/bmoIfkRpzYltJZseAYxAK0OK1mZDAPPiLLau6hhnDEMBKOAcOwLqu7kjd/ibk4qIqYdyRk1qaCg
F7lA0rOBOLXCpPDpvnCIEJAOczijC8dXrFiWFvLKH3ToFsEoYRe+k3Q2Pq0mN+zN8LI/9dd6tKhS
+KWBK7ZdCqqKHP/BhzIYu0JZi/Ux6XNexPr3ZUYS8lbnpLR5b00R96lBKIwaIYIR8NRSsnRNGVYr
9HN85R3C7bE44BYQlTvxftYpwvMREq+KV4qeRuXnwkv5ABuig+hhrY+5SqeqHyYFhXXcpxWNtw19
1T9vuJZ/PoMGw74smlEoN1JY6L5o9/r/Z2pVo5MhZ5QVvgy/MDCvnnRpkHbYOmoxYp32m0J9IKhu
fo/hxul/q+I1oY+5VC+jkBe+lPhWjHPp20Ddsodsa/Stggct0R+LtxqOZLxSpbL4gyChOeh51mnj
J4zOxgzXfz8n6xYCDpVttBGZrbr1vDQrQNi9/NqiTq8ABs3VEuc8zRQosRTANKE3JCBQUfvWDn+I
DwU2jzZjWYce+MMZ9d4vo9w6CRJoCDJTkEcN20Zw0JWfJ0SLSHReQ5+tQ0WCA7WJEqNOBCzekTu+
dxfbPORSsKl2+5+sPB+GS1JFfF3rbO/jl5hwR1FfGUEfk1eYVRGct1brO3esRuSHdtTPC3027979
HgMB9WJZ1fBao5QWSu2S+SLcACBAIlvIdZimo7/rJQV/h5q7EYu5RMLGxdV3Fxih/Can9cMcXyNk
xTibIZykGQCJfw7P0xtWGcEt7+JUxJcNQn/JpxF9jd5wLIhdrB/M84dzR/jqtyJJCGNkll8VUxCp
POwoaWZQ/JFX3C8vShmYUJsdOJjU/Ui9E118ZWE1qaDD8n0U+J6o0D4R6+QbsI7ypFuqmrN/8bQ8
vR2VlWuzk++wbpXkLbQif4gTEy0umw1WdW+B7VunXT2NqV3YrnR4xSuzwU110hULhk8zd8830gHi
L645FB+j0rDtS6QLBSNLF1PwdRlrRVKCLokB3T4JYQZ7cfOntjtRS/AmrJVPCx7W8dvTahxBcjWx
BVD2IXu4MME7frL0VS2UOfRzKZWyFoJ3wtj873O6VKnk2I23rf8xaRDcNTxukI4exgP4m1K0af4j
xbKXxmRNtfRgbILF8ii+gMODb7E0LC3IQRlvCFmlEhQaTLWcsj390gmrTArYxSb8O2Ba+U5zP+gY
19pqFKImvYkCMd+M0u/pWoGZDg3BmJPP7XXZ2XxbRyIYL2HPEbW12WYLCKhZ+IA97YmU5Wkh/70B
OgzyqyZD3pGeZuxHCWbd6xcIf7yhfQCpOziYGB3XCsa6uJjpZUcS51qQ2z0tEtbp+WMeiN64I0zY
9LH+pmltQlbZgCYstgX6+d+qJA+WtCDTsgJZoBt9wp9cuN6EQDKfOKAy2p0t3L6zIarkaELxT0JC
+jDdRajWgLQ42wwTXjUFd/0MWgPCWQZn9qCSOWJ4z96grFeSKsGWrM0JO0B470YpFaImy3wq/Fw6
09ST7SDTIrIAihiJx1et5eemZ+YYPX0mWh0dIc9NAN0RUN7X/ohBsHakKNzuvJiOoy4jbLO9pGBU
OnowDJUj00ccgOXeDjMkV+HXqWBXYtQB32iOuUUmpSNd3KxGH7MzorCWUBjb3Vp302hKRQJEgij4
Nf+BoOM75TM5wFcPbVtTKW95w1ekI25tG/Ckn6IFrcEKNzQopVbgdMP7QkL286yGBwPC432cY7bk
PvhquT7kq5SMaUNdZQS6OKAPc+xB+xZoduSqwDOydCR+VvaOjVJ4s2ddHrYbILbcKkUt6NiF25SR
cZKEq02GLSXxGCr7TLCPRCuFSEdhOE9uSMDxYRkitVFsPCPL413WcZYnldVPHGtTer1vBfGRdp3P
Q1qz/oJlif7mAWaurMKqwroOdSch3dmmDowGFFZNJzPx/K6GpFwToMuHN4Ds/5UOJmCarqKKriC0
zbTLYcJ7pZgx/a0YW9vTPNc7FXyGyVcfvgcPHcHq/9ez5fVK5cMUgG9GXWZX+dc3nISeF/BIckTA
PBXrE80GYx3mCPJEnIhIwk5RjBbJV/OT3zmGL21Okp8mijuuLi4I4/g0QeEWGN/gETf6hOVN/v4M
VawOzq4owUPgPbnq5X8UfTWlQ5nL7ZtCJtJwBHr5aBYrPgz+ew5tbnP89bF4k6jbgwUf34uqrclx
w3euLNo6O/N4BhBjJD1Mw8h6C4Sa3dYvBj8PUV4OAqBWK7zJGFIlHY0AqZwxLzFJVZIcbX2JrNdG
fW6RkOQZmYf5zI+DyNBvPm+s9Ba+/rGZytiy7IvY1TTtTRDE1/ri2WEpxEHxZDakNyoX8zIqrdpF
rgHFkIoDnyigXNGm+qzEwKRamu9B5cv33N/h1Vt81Qz9d1DfzHyKGN2H9qllZsYhlp50gHv/lVDM
P5vnePD0BBCEW+JXF99aQmLba0g45W3X28/yuK3451CSFuCARfIBPUSBOF6YJoeCUPCLDPMcBLe+
9XDOj/vFq5AejS+9+h+7u6OLd+m1YzDfzeK7T6fbxapxym4lG4ix79M6Gwn4+XDTMwPEWm2pl+/u
PPOM6Orh4Qd+f8VYMximEeaVWLJ+TJhOWafAZVq1V/CiPLTpWhMhPTDXt0R7DCZMJ32arIyzZBQ/
d416NREMF+ZSD0+g9gmn13oMC3+f/0CvumwjoCtnOliXaGVY7eub1tVdezVS+QJq8jpamfxUikPJ
12V2tnEFBWH5BuaJHMfR3qMi77O03EC2rFjm6aHOdNBpu8Ss58owlNPIYEOnWjBOMtxH1TDdilMI
T5c8h8Qk61G/zVf5WNcmX/9zCRhR0tnjEAnB36gm8SKIzW+zGUFQEGm/mS4LMReoT0t6jxmi+hmu
Aep2UbsXAq2pzU8TuRd4lXWGDzukpyaSzxBUzhUg9/NFmDDgyPvItKWzfi5mOJnjXsEroSR8dKMW
rrWZpCCTBsYxiC27lNyQ5g80Abj/zqjxgthCMA5eAUewEQFHXGcJQUGwy06pL1N4XlNUPxeh+S1o
ud/9hNgaxBvn7/VRcEnHmuLUdOq0/cM+N+JvqEf4mAUiV16Sdi7nCR2IC/nkuCcA4D69q97GSzZN
tUqx3dB2XZ3fVCpFEadSIHNKGlTaPBnV2cFHa3CLPdOCDoXeJCR+zO5wBCDkElotYHYPTOW+Rj0O
3Nan/IRtuG5fe99NdjMD5edhVSgCaGHXnOhD5+aA8JkSPXze0EDogGDHqc2yaWXHqh6DC6CDh6rr
TyAhsT+iS/s7LEJygixioea/0AJ6HWQhfu+CLsxgj5YjdFDRgDfFyVqvfuLl9uYi72Jjh2pNauYG
9gXFrE3JJBni5OmNYI0J7iKNG4EbVU+2KH7WKjbSd7MZZXtSRk1qkSLEs+eQLVyfAlIAd2nU0HLv
ED4/MvCAk/pCKzKbO3fQowLP3BSuztGgUjrMSVRMQRCR/wX3bzWb/40CYUGsEHGbCzSsEhVSuROR
l2fGbcZM33HhSuh8ay6DCzul/DByTvIigXG4ihOP3J6mYBNO++ORMX/elJN2yJBiApxXTG95UgiA
fEThS49dIPllRl2o6GzbfoqX3bxTvyfIWJwQwq8hkYovjwrJ/3rIzeP14QdooyuRShIft+L2YA+h
ldUUxucRTwXyF3Ioej3KNMrR+Q8SiYg0l+g/z9ryVS7fGtHJ4rrvpHs9CCZwB3SF4PlSwtNjLNtr
uLIPRTmb69z4rkoEHxR50sYNr+0fJm9OXYIk0V03d08ayaFkccOxnMXsPs4I7K1TMpbkfShhIdPu
eNzQYZg+RC9TQOO+cCKcKf0dZj7Cy1mf/Uxe/t2NsDHUz2ZbO336+u/DtimSucV2jBx5fG/Xthhq
SGqwApOPiEgzrDepagibaMXs4J9lklGVbU1TbR3PZT8COe3K6CqdVhMxdNpTdQvt7DDsR6kUaTwe
AjR5ByGi8cyJuqCuS9fGUjxIUB1Um33uzxfCMoNYcw8zbkTa9FRIRz6tmOLuXxmLhGJFiRsApbnE
wpexHLeqpuGe30S7jXDX57Iq5cri1m6Ys9BrwI5qiLwZgFxGvW3Gfnbg9FOTCGLXfp/lK9iFO4dI
aqRoLCUlEFxhkKSCyKaXaRVta/gElHMvbuBqhFsye/glCHB0tBJnPkRoe+MiiRLImOGuykEGgZBo
X05MKUcUbrycuxGLFUjbd1C9R2i7wh4HqujIoQsoOMHfkdfyq7SrSxRhoD39C1W1VJ/diT9cIepc
45VlYpj6JGSmUiRZRWjeReq3NjUEiyCBz/zGxV9PfJLSMEQe60RddNfwkYglHHLUEse+ukqHrPUb
/74WfC9sO0YjoVWRbY1p3n/j8nOwe6H611wnSqidKgqOnERDl+HXgrquwSBU909XzK7PONWXcFnT
sebvcYs/TB1X/pgB8ydyFajx/5Plk0TLYJZYIffgoOBk91dx4CAarz+bKfVroVSBG/dGMPa05WR3
hPdQ7GlDKxL2Uv4ihZX87FpG7dW4GB6vECaDCl4YU7o4FVl3HQrOEe4kUlZkfMOeu02KnI4WLrUU
HHv8kCi/jzM5AjeD7kDG7Byl7+eP8eIRMtHNeVINCLZtdZwhpTFCz8j4L8BOamuKj0aiZ842Xw+m
WE69TpENXA+vCDMuPoNG1KUAKOmsiV+Lcs8AiYU6E1UUxTix+SUNfD2pVBvrrDIVd3VifPQlu12f
1OpVPKgpLfLdOo8NzeNniTPkQUN6TSQi7NNFVcSuVHh0pzoIWZBSS4LeUNZx3VxxqAOF5WK1nTi+
tXMsK80aZcO97H6kq7lpfgtRMNcDF0VOx4VBhOKNqNtoGw6zZcLLR6Jf+hdNoFOMwXmtfeiIe/ty
N/G1tn5SCOWBXYgFvj85/aIuGPdtfg8imk8hFF7ZGDU51U7OHV3cCmmwqvL71kfJUeyPMt+J0k1G
7jzKJPSNeR3b2pu97MDKZKIIDnG8nfs2amaJ6XPOK3AsNYw4Nhob1/mwJ0lC+pQJsrBTl7z1lQyq
p6TbdA8rZH/LBZUv3xKzIF+FpZL9TbF95cfRDFyp8sZWJd/0RbbRtqsFp53yoH2zT/cIGpZm2bR1
V9nMY+lZ8FnV6/iBo4coEmxDFDN2mce01vuLkqp/2UmAk3ih6FfIBVb8xFYnA87IjsYpamM61XjC
HIqMwActfsr2/lZVbi0W1Upu+DfwtBP2oB8GCcyHf4VFUyoaKTtS10MbEBp1aX/3itGdO2+6J0KK
b/hQBmcaL6WGAOJit8b1idHtO2ZlatbdiWvowXkdrfio1xLXR8Cdn7x37G7Oh7D5zjsmcN+EVAFz
hGyix/jB3fYLOPEimVTREwZyaKPdTvE9BrJwvCNCvnhruEuLqn1buunDHXr8DbGb6vbD3tSbxk2G
hM+3UAX45jjAFSe+Qr/lQez4DYuICtfVyM3CAx9GHIkZnfOwi3YNxk1cIwYxeQw5l/g5Cap30ELd
KONzfItP5BtLRgI6Ff625iJ0EKHV9mTjLKPg0f/g+icLi7zuNDJrOhW9vX3TxOGyLgEvYoXgro81
ehpwAkYQkaiiybJng40E7vdFflxEWjpzie9+oNH99mfDrdn0m0SVl1YiJYF3z0OzdAJibh2DCFBg
NvmHQGRNlJd87Fc7/tFBisREMiUuC2Bo26lJl8bt9R00rMUI8VcUzBkwexV4S3Pmim7xl+XbF4DJ
Mq0UR14eWFrKYX0vnz9Nf0syUkTUIJRQHgV2HaP2ApaeYiDQadnEvs4VSlOJ9frMj4CTOk0fj3cL
CJXEnZ4Gs0S1FeV18ID3kuK34D+JKJ02pHZz+apcF+ltu4M+gQcGcCl83TSTVTwpQOex6tMH1keE
EBERdEflctv9QjHUT2HCOIcO0m9T1xfLd1EiV7vOg1Bai+DlFu/s/t9+CCHZO0k88sbjM0UvC68/
P29uqIPOyjWDke+dWJktYb1ruchtz8ic8jMzsyqwlPHnCDLaEYb0WxAVXyZsxUBzCoMRmoWY3vQ8
8L+v6HL6wWhQeIa5cpj014pbYaVJZ/qHFd9pga96hzg+6w65jxQmg/iSPGMUxlNN8lqRglkLfCwA
yeqQ+/v0sIK4QWROsbj9B1i44mMIy9V1IPoofNu/5gtBJB+3ipnxSf2/KsdYQJfR7TshdrDUzO+g
wd41EIQLPpy6nreCXd6V+9K8sGOc9DPGMdQcixzWEkfpoq6Twx6QC9RPutsv7zqYo5H8pRxzvRVW
CleOrBGc13Wj/AxLR1jRpVdLSqOi4CGJ9zRtCmjcfKX/899rI3TFTkKwKeIgRw6oNMlkRQ5GZjyy
qKYdmaBfXelsX9n3IPR4mK+g4QNKPirWVMchbuTdg+uHXPe4CNMVTYz8WXbFhHm14+0cjDZtxeF0
96BAYe6DUSqKaRnHcP8nlHx3btzHjjpARB+m4qu76T2r3SNVUeDK1k9iqtuwXyUYpgOIkSK3FDK5
L0JbR5qkDNrAhpYQOwkXE+fWNiI+nHHRB+JE0VYfOCi3NyofIbRgwZgMxQ5vCVY2E5HtCPItYvkG
Num7Oc0Irf97gBdKh8OqeDT1H/nNwbScYRMYeowNz9V2LfuInkrzBvPRyWX+1FTknkTLsGTZNdeY
MZ0g7NgQNz++N+QH2ZidT7+lDcNYvPbrAPeSV4j5rKNNJGTI5Z+QUGajMwn6X8nWPJXuKJjwzMvY
dzxPzT8w/kY2ogNLO9vAzcy1k/bhb3ERheTLWpwA4GtT2ALpxbEnukcWoMlfF1Tc6YN2gL6vUKMu
g2M9z2uP1NiPZ5KXjWyjliwD/GfICzkXj5Oe2lXYtPGSmI6QJSpgKROFtLacHLkA3f/1zKUko5eo
Zkff/+2r9d7qmCjJHqbw1uL0ZDs6Z9Ry0u/m/VL33klHnbhywbLHHvdZFz0g/x0dsg2JeoYsegbB
NTXxV+vbYxbItAJpho3dK2PU/UopnALanbCIeYh4iThj/loLCAhtEf8Hm0ozMHaG+n5wDHR2YU4C
HWiTyhMND9HXWZp37n9rWHwt5+BLCcWZjjLc3zZPYVIXpaL8TEVlQiZaiyFUKQwsTp/y9mXAFTwW
8NsrtAwi4ZdFtwexE4rIoy9OqpWEylveMd3i3jt5K7sDGCykGHGNDmHHphfVc7yjNHmTPLRPLlvC
K/9JF6cqr/bjJjrCx3dyzMFUf3HWsApAqNbG72sDKEoBNhOkHfClS8XmWvMJLcJOIKmfa2AUWHEC
GOEZHt7SJCIQ6CGlPjdtWJyqgA0uRnVv1Z2dLR9ZCVeKx7ISMxFM4OtfwuBQE2T/rtM6H3DFCJep
hTlLAUwxo5Rd6Po5ip/T8djorLVLEvQovd0Nfn8Td2Hte3hJz+w1GUXkrYfAVSKlsTeSJ0rPmFXU
6tXgyYXIecyshVUc8YTMHEgBInvkdbVjlaIDAtGUDNGKy9jvX886gq+w5ewLST2RrzoxETNWMAb5
Cc7hrt1qK3sYDPDYEsy5qeQuWqwTDGELJDbW9y6Q8zelAOurDewu9GwSvZzsH/swuRvPQLZ3lZL6
eh3SGwcPPoRIG8qgwVoxULTA75o3tNeYzzr9GbBzna0dSFVDTvSSJMDZGafU2+VPiyKejsTI/PUk
Hc9mmyrY9iSM3uvgYYwRM541UTA4XY28L21KD1iWOnlSJNJEmNphMtnUcH1PRBBD+RRJQh2Ek2bN
P56TRedxo/hXD/AWoQlQAB4akGNTV6UGtXrGKeK6mF/R0Qkrr+wLxnkcfbABNxQgBIEZM28uRRmS
QpoleG6gDgGq8YHpr2CEfU7Iojd+GyJYQItckGrO7DqqvHaD3UdsGrW/LflPPUNGjRMCxUCTpoqp
UUdLyo7nx6GdhhOQSiOVKuvGAmiIsmeAvWQt3txF+U5YtjJGxtYL2Rxh2Kg9wB3SbEzRkcdG5tnL
wVLuMk6/a1ajItaERmLROPoVYWWwWPHxCWpVuP9l5NmGD6Bh5sB6ULyTpN9UWPGoznMChIj8eNMw
3sVz6VhcUR3eMZIzQ6VVFtrCwJl1HPvFPS/2OHKLdarBSDaFI7YIe+WDyXQHx3/ZKvLWopeKjyzh
RgQp36bwTp6IIZFfVZYXl6ELKMFqO0P0VLvdd1BrLGRYCNUX/eGoiBR9Qm1ZPM6VLNAkqGYBXak1
bGCQoHYB4n8d4itdYLCf6WCZfYSMuROqYF7K/dB2LF+JzZnMJk6687Vdg1Ozp9IPUKghsKYekfNu
PWoDo1M+G1h9Zs06XwEq5bQlGfh1GqfdO2aUWMQj5HRHZRsouUCqh7HHD42wTN/AFYWgZMlnE57z
DgJMw+EewFBJtYa6Gyl68YRX0RM1fEAoNYlB/Xk+HdvoChaVTtHQu8sIB7/444nQsY9X91ZOoLnU
KK8U3zAX+pidoZlH1rodPHZHsXzrkQFNU6IzAt2NuCvlanR5IwerJ0RcAadJ1LeMpKBjUU63m/H6
7TMmhAr4bGAQaC2ZrkQuuFxSFwtnsjypKrakhcsVSpNlNasRW0aiiPUOf2h2maF6q91+hAVnst1C
vQg1su6HG/1F2LeYz5EI6+YV8bvax8J8zR3qUsjNij78nJQFsY+x7GFl4EaWyZT9dNpzDYQ+VL7K
mBOyP9szumTXyOq5saL2+T5ZuwrjIwYO4aiC6p1FFoYtTgrLoftkK+tAgM3bN5sLkxJb44/2xPxj
Pm3W8rUP0d5sSoSHtuscYIVaTicfrcl8fAUKbS7W/unKI8COWG1wIU4r051eZNH2BeDxG9QS3zrx
++bP7r1q6F5EQsJ6Ar59eVarg05hwKr3hkT6BnD1BTlXmztJk0P/tW3G5r6S8NBmzuXTbrHqrXVj
FCB2xsQeyMLpt086Y6BK011pkW8XbKqMaT3/HGA584cwWR3j5snU60KzLm96cPWe7Q0agBNGbGbl
Vg+CquCbHkKi+RQbPm701O+Vdi/ngoebQ6MiDo/6oxMpmpc9AWLLFyOFxO30rlx/liquawEn5KF2
isM6VdDWtpYZtrBULWHu01H1piqUEYYcIbjGe3eeHGz/YOBAKkl2oXGZ6bBpnVLi4yCMdPtpEaSy
k4LeK5fBPVBpm4LYaJosKDN1j257zLoJPc5iAWic0NTZjdVbeoYsarTWmpFDkv2Kza39F09a1tOr
gRi0RfV5DFHwTCL51f3zAx95MBIw5q91OY4pga8ZOM/y/ZU3A6w9ERk51ZAE2nEEl2d/TZrjaaUQ
EhxQsqs+wN/BVNqvgRnYhliAvgQgW1xbCuAnWYa16QoSovlY8ihYakZUOLXTBp5T8H3OVibfUY/X
2WuKf+Buh2jsFhlybuVG724J5sf5QdxpbHBhfgppahimKmkXsBiu1mS97o2Dd3gKH06X2AmAI+fC
WN6x/+0J6WkIJL/kcDyDgIxhf0LLy74NMOJ+tKm3PsMILF+Mqx3vA/kOuiRaAu/KhQMnbr+SAub1
+FSYWugkxYOItfrRQeuJY1ULg4LOSLi7GDQQeihpah0ChpEqNiLOHSfszNq9QA3SMEgXPAkzdCG2
dAVmVEvYSqg7jtIRRp18T1AcVIQDTicaUyX9b2McFqWzHjsoimmlNFcDAq2qIBL1R3Xe0ZoFbF0R
UDG6cilBuAu1PxgPu/DiE53cvjEa/nWbl5WdNF39YBnGwdUXuU2YVkCE3TUJoyY4HCfO1G2TtUsl
Q+2Qoso+lJayC2MGdXQl46AR4U4dYTREr7A3y7QXTo1nTJmz8QyfYBjmQHVBRF8WWskdC9jfNR9x
MKU7/gGYyFFdlmevMlVUPSuOURD/R2mEFlr0i5ogjADCfJiMyplBhf2oP1VmjoaYNkcYR9D4LNRd
bGhLij2zp0mA8JANalu6sXa2SukKjdgDwr8yhqF+buMfYuzbo8ZLGtCn/XAvybqZymV1Ozb6bsnm
267KJulk5mO8QqyV3fG9xaedN/1l9p2ZI7sIQodc4Jw+ncaGSQYSREUE5P1HNHmYoTysqgPX1ZDW
DRIA6QJfLh3YxSjLCaO3JA6zu7FVzhbsMmXQLUGbaBZ5cPRFceanxjmZ2pnqmXYFty95ineHh1vY
Pbb50iH1TW3AIG103pnk513FSqTpsEIVb6wehiBy+m8HmPV70AJl8hcR8PwN6+fWc9auEl3e2qF8
lZvl5d+IRg/3+a+UaOwmqUjJ1Jg92GoezQeXeRLHVDVEX2ueaDgKA2IS58NglarrooMO7VUmcRbQ
WWsToZramWkoN54Sih0Vmvh2FWRBOJWVuWueWP8cab0oQ82jewW6nxLtypBT34fdvG+joaWEbHsw
6K5h6K9vNrsTCptLmNxDyBBm7evvAOtqCHDe5/DlQMPIv635RENM/tIkmdqggSjbp9I1Hv/i7X2y
SlghbsuCxqqLLiIW2eUedPYutFWn7Tvru3lSiDH/l3mbuAMpOdhW8ska3C9LM4CRHhAs5EhiGOYx
57TQgKFn4IZmUCS0Hy6s+zTrU8LtGzHsMtt6tjfoCulzaOpOUL2mLf9rJ+At9MmiM3dKj8iB7/eF
qpjUVwPIJ7Mu+2yH+KHBK/A3EVKKI2j0Rh5IVTey3SIqPIRMyxf9XzatfxA6JuHd/ztOPC0Iohxn
Za3EDuWl8Ue8jw85/F7f7Gccyl5/+lxqHfYdm3/zAQFtYFFHjALK360w1fV5WhUxN8rU69icM4w5
8eYfH9ThIzVfcZXLy8hTiK0d9H/jt5agoqg8XauZJPQis0LJ0BF0oUAXEdmDCfyQ1jLvMnrUzhql
/5B5NXJSblihc+zrUDSRFe7zxapcnG3e2/GQt5lJIsgkr2Pp3WQ8zr+0XSgxFJLSLHusXNjSWuwe
2HZEw6MZQDLh3pPs5QemUIC+x1YMJUIlDEzdNCoWTq0Uv7xHTAqE8SlDBf2p0dW2dAZ77mw7ueZR
ILnyVsYp+DVCd+vhV+SZfrogxIGXF7jLg611vSnTCpMIPrrW3WuWpUF6wLOcskYwFnhUVhdSGQFV
edHwH2h3NAkse75xTeTgBX6idlr2isOCA/xNSoKrXyH/jpjX9fXkPkxNbF8j3cL5lU0DBPbBLOYY
mJR4NweN2glC1NUzTcoKZbjthsADqyFfm52iET/aE6x4xsvbjiZs3pd+Sh4sFhWTwjug+BfcZDi2
dbKwxZHxDsL3/jmUxtIMK1Gs2nAFzldS3UriL2l/+sxtkQvE2+xSSyLRFAbA4ZRV/ZVCG6RnZESn
R5XO+brkVIOJLA2cnbf7q0FbHxYl2DUmgP07R5l6xNxYmRMytMKQftym0kyvMTajne4x2Hr6oh5x
BC2udJ+PDGsQt3qiQKRR8n7E/QERUltF7vkd3sQ/32W3ib09kG9XGEQ2De0sKB6XKriU5bVSM3/1
7DYifcuqAMPtnFy+vML3yI1foAJA5MtDpMQ27lDaUu7OUq9zqAgKW4/7lzHRouK6joYY0qhfnzNH
YMXl+u0XdCj7HDwHtn9z0oK6gLguu0DtyRJ8USXlTLaFVxspSj/RRHOTCYB4UBtdSEHQrhRgZVYy
6LdQbOaGw7FLfzV/UWrP8le9QlAvQI/UP2VKXEB5/bDBWW2siGDKO+dejfrO/mbzOx9T38BIhWox
5pNvhCqoFUWqOCsNcUKPolr5hYe6VkW1bHY8kHWPY3nsvVdd6CiNYycu5Gm5cwBzZzS+9A3lo2PJ
MQXWikxCTClAv/PDOsCGxGVDBdenUVMIQK+yRkRgZzt8UY52TiitO7eiLf1JoO2DrbZvyig8n/xC
WYfimJBWAFdtiBYGJljg0WKMDXsk07X1L1uc04rK8CP2hH1LUZJcmsDs4kI4aICgLzIWBU5LUENe
Jo0QCXcdVCjE0kXRkC0DFwkxSTYoO+xzdPbSPpM0Is1yFxSA11UOcWgXnTyQRa9yt8v9wqmIUmp4
GkeMl2QDUSWmLOsQmCAj2DXeHaJGpX6VX8cLzQ/Unhr3cw6vggwrVcJteuxDDFIkPKkxal9N182R
xkfi+pKEBFauxWg9F4dTrRY+r1JtTHonMu2IN+sBzjzyvqDriZrk2QAhr7/Z5Gc+qUreLxdKGYuS
88XckX+gjIdpC/ThtsMSMbJkKlyxDWDikuEMTyljXQMW5Dd4Ih+MpSFVSOHgtWa8Ug3q/5ZNah18
bLmaA16B6XUkP4upEw/oSGS2GXPBiMCY+i4DJZSMAwuDtx8oRr9g5cXR0w2vf4V5IMuKwWW1gs6y
XdYmT7NKgg84Y/Cc0V7th4lhC5/tCHemm8gerGrjua0szuJPf7UIbRo/KOJJii2IbNjtjNh4OxAV
vHvkQ1Swj0UnaYkl7erUPgdu54j8eUkl6TqEbkFdaiL7Aez4gzz9RBwcT9L9vYR6AzuICGYtIlub
6Rdoi5lFjpe7uBIM9KzgPJ22FI1JiPzKpoRKGVNPXe07lCCRd0Gk0HrUzuj6OpV1sJVmVpXGFZfJ
hzRYrg8NWCaHov1CC2CpIK/odLLVoLLLV44bYpjZVhrXIBXhM+nOvvbQxSUEFvx6Egv3Fh7LX816
GSgFHIanVHKhCoejL3K2LqiMLKAQY2glRQU4L8Bw7DGY9U+UtsuwooeXo7oJQ/ZqYLGnSTmUq1J3
zKvCbQruOazdNfyGYr4lOzMtU1NrOfi+kEqsqPt8yeBI0K2fCA3/hPC9Dtnmun65zwblJsbnq2Oj
m+06JXqeq5Y4QBoSkYoCWpHlnDjVRR6DBn3etufypRUKmxlhdeEi3ZCLIbkeAGXumrRDSLESOtxU
WHbkPQ9aIjkZY9+G8CPu2kmnJN0YJGmO157KDXVz4kOEksLyDbEZWHdqiQy8hQzYvUA1q1mBbh/F
EDi94Os9jHYhsqSjkFujz0wC9KVFCwz7UfFYbI856GP5wTS6GclmVWDifVdeGHUFWzKADlYUIi2y
slECQ7dr0d22anXxfI9dWwk8Jfw/kstrgagmPTFUf3VMXAMSN786ohlwhLtkk3RpS79pFf8yW8zA
fYJkZ5i6o7sfWAEJPR1peZhcNdb3/1AQMDNNUHkjD2EIr4PYF0zO5bcUsJtlIhFxtUqK221mYxoR
w8Xo4v79TNZHxQNXVG6khlceAaHdyuKBkpntxZriTKeXbqKfmh5u777SYmlivy0A0MYkku3fDzqW
vZskz2xazBDIgsM8drSxmwExrvb3wBjB+NpMZ4pL4HiehZ2EWVrGFe0+lS04mnpfn/D2LX97rIf8
7WbnnxwF2Rsab87RFHn/t7hHBX9EHKbJq2R18ZQzzKYClUUiC/nlLKTERVmDDCqAxUFFVvHBp6np
ClW5eAbav7QY4dTgmWF2eb2FMMGF7oU7KG6t0iYiAcbngPyhgwhjehvjRw10aeCmN/5hNKNE4Fk3
/IFK4BQzBCUljvPluZJgNOcqCK3QJYnVLy5sZNSsJo3HLD3M72VAgSHc/S+bDe/QtxWYKaDkWkE6
Z9id8SU6Yb9Oel4aj3H91rfNyk/znW9nqTv5okiBfUiE414HAMI4BlQeRmss9hojDIqCMBGRrnO9
mBfjEcT+IAda9IiF2EffiP9ruZhgjRYD4MSZJUs+4dgv2wN/1mYvQYrsTSKfucBxRyi+eu7VOJc9
cBSY1az+UIFdlttj1s65f7SxtNB4JQt63P8UVBjgTdvSVHmYFSabgoSVJgApe2FDz2s3mDju47NT
PE3zsn1IZmMFZOwe6QI94c5n10SSG7UM0w/XJGQphNDozjKDBqOoBUpKy4Z4jRKAk/YQKia3aAk9
wtlj5cgEdSY4sftLt2sZQd9hCI+HBixvs10xEp8Zps76OBVhI5A0YESsuxSV3ootEmh35SSpNezc
oPwRbMKcWxERqA61H4PDlt2B44b1FvcEQeIwR24ncBguIOyLbhLvRCs1ycPoIg1tib0xMwwqD8CJ
nu4Rt0QvKfGOVcBBDB3/Dd9KwN7A9XN1CHe9mkAUZNOLm550wTakdQCc8egD2G3sX+MKt71ExVZT
UBx4V0PDNBelRRY2+iIJ2depFSsep1uwem/yXF4ovUJ6YS8w6h6KS7yIWIhbYcu5GSa9iYNsoL+v
DIvAZzs7GKj2WnKR+bNpOOXL+xOKInvYBHrmiyd5pGwzrMkvfIWJfGIzyXzNHUnXlh0fAXoDcFFQ
mwLaxrviyyOm6rmgF5SotXUmXbcvM/xaiXni+Knw72HW3osbSFROAuV8MFpNo9CRikVwhafHwblF
AcIYfzPOYz7XpSysyEwSy8LAXtVuCo32Gssfn76QXBQFzp9WNFzhQ+slja7dSvZx7q3p0h656Pxy
perik0UtZR3ebBwG5WCs1DL6JaWKuQ4VjWCYTTkjZjCV8UIf1ycNn3F+kXFulfnbBz5SovCwEORv
hdaPvuNZLq+X5PU3n+cFbCGP9kcO51rGfFMLUP+bo9/6f04CDtMnA68VEJpOulAoLwu3HWDRSA23
zjjHAyW4x6bgzYWlXmKHczyalG5PXDg314poeNQCScDtQBDSP8AlZ+YlBpViFe/hHNaRWROHz7HJ
ogpBQeUlxAOaBTpCZmkN4cZ8JpLGxkvz/vIyK5eLyTpGqWBvPH/u6Zy5g85TK5vYoLA3fPpJWHjf
YGJzDAtFHiO3LlBUhruTZxRd2Un79HFRazGPjj5NbzjaILuQo26Q3olQx29GfyrZ+xHGYVlKD9yn
FHxp9QX4hxOuS1ypZlZPW++K0TsbwdNUqBFYTNAmlPIipFAPHMg9uvl/b60U/WM6FFxULcY53vNr
VtmWPobbyJ8j+XN4sMLzyATZ8vdG6BXPDJAyBfT5utw1UKv6VV/jrwqfVCKg6bpgxyq3gUtSMkoq
6pPTP60c2Aibh4nwhs7rrBFDVbXx1xCLpG98gZugGIA3qQNVvCCclVFA4hagqgWTYnVWvFh7UqpT
oLcFRWccrfqmZUAqVh2EPKe7kGw5yxJsK+zh5irnvyGRIKpL1EQY196cJptgX5mvGkrFzA0g3V7i
NUkb57hv9/Mc9uxG01T3V1N/+tEJCNlJj48yVrL1HvkClFLBBj7ga0vMxqsKpqYaMxb2bxg83o1/
v7jljCIFwpjdBlaHKqds7Cu6KIiI15XjYSbN/ra9vDpilc4lS851fqM5VMKEg+TcPax4SzSklrOB
H3omLBH+6+t5f2BeI7ART0Zfe5FhCzQJ/0QEeCASwyh/L4Yf25O0GgOWf8SukkGLz688l2nV+D3l
nDMxKsibl0w2BN21elOXVR3cgqzgxs+x/ZGZNLHPEylf+nqdk3+NXFMR7K8NlsrYLCpFO+PwVGzL
+Lh59ppRkI7JD3lS7/lnha2uuoUD3TZGWgNlMi2nUyYcu3N5cRxMAPfZ4oH71Qsg3Zur05AWnKee
+kaESBd1YXVkljQWtIL/MWT4NCKxGA670nuWBFsu+xtOV42ZxCAk2aZ/9ectDIrKP1jcz2UaPFMH
Q52QjhTdzBs/1Ozu+OzAyfB12oNzy2hZdlUQSKrCK5ZnQWD4Xm2S6YY7VrIYjVaNIuwNXDo4/Dwt
vDfc3OcjkA2yG0Xo48XzS1n5EyP3Ag6d/Jewz/qwwGRDgFzal0dy9Bsv/8tVfdWUEBVYMRzkpXjP
NI/9rysm90sDEC4zk7Z2G3zuQeNUpq+vyKT5aGssxO0eXrkmFjemvLCyRfsRS0yBPmUNAvvlNsIc
Ra6sURM7hQgDMF+ylSqaCQTTAzEl4hnoN/KdfDh9np07DDKVeAw8C6ZeChKW/EYNcytkcvMt6vAc
JpIKplbnv3BfylSvvLia5pcxnnI0SStTwkp0rVYQqdcoLn4c5gDUl/bjXBCb4b87tfqENnFKQF0f
N58/CmFJ65WmMNyN5O4mQSGV1jVgE/bQpxXgR/UN/30tf/qz9kg84uehbawtjVu7Xh2OSjUYs+4i
jedBojWxEWaQRaq96LVBrRTZxL1LcGWUlGREpLrA99BklCnDqQyHmwxUo1uE8t6kvrAfb359CJKJ
AnOTuF6Td0wmm46gRLEWOncxsv5zRWXR5YyokOWaUR+rXEM/vV5zPQJWRtAPifWPafzjKAasFUqb
q2oYA1pYv62g1f8INOFwehMNCQVd1f/eRevwpA79xqzXQjrsAVXqPILHPP7zAK3kzG5FdJEv14Y5
W+le+htQ2aXNs9LGrDB8GHK2FQud5k6/Xyewj0IfnKx8QjlDAJmMs6goQHl7vrh5C6DDflydF9vf
t1Gd0NK+zUo53WDLR2Pk3R8QcoGdjVP2fCZRUY54whJ6lVhl/yzKvp4YQXpt+K89gZSbHGtivALh
/fjNe/TmNNWRVw18XxqT5NeA5h/IA1tES1/4njHQmnmcMBcD4+Ri3a6NX+sKBZkHJGeQ8ZuZrO4l
4Vkf64dku/HyTy+1hDjxdF1ddV9JUht80K1SR3t92JBsGU8GHuRkkeNLhNCWm2/6L7cAv1oHNSU7
E8shvBBjqL0RnLHPFU/FrCJBYujtuLRXtLmpKtm602txqliLmW81Q10i3GF7IFcwQEWiArRXzivf
46v/cKb2h6M4fbgmHQeI+3DoP02Lg9fzR5BvvtUcPgLg1riBRRksRxaVgAjBQ9/FmocSGLytGiNH
AEa6fvDdwHnldyMKRy9lmx+O+6+X2nPdlOmEcJDE8ww8jBc8xElg51QP4i4UdrZFzG/BLtqFNlh/
QTeBHDGnWLGDgvjbYUnVSS1WplT0FXLG27uH99I7VUGRWTUO5Pa64+E4lZosYYjTec0jEgZ2iTaI
sSSj4FzmRcZ7XRoAiwdVJoFAIbYa71M7Z1lt5yMh4HTTPiq5pMeVVwG4OckPVjjoeQ6RswZGqd1z
wLZt7IqSGNdARojkGHi3wINIOFVwz+vwiKovd3uSMZuKgdsYEYq5N0D/VF9mFE6Up2OcDGqQxhfW
q2LBA5PiAEemyLSWMhHacxPrvblFU47kVus2VCLDBhjuVHO9p5AKCamZCdnu0YjxF+YcdGo1BTPJ
bkpl+w581Ldv/3C8KjyLnM6RoTT+d6pMnbaweX+Vnf7PPwV8gtDcYTHgh6HbkPMSOOj7B7Zw2Ht2
4aD3/GSc6W1GXWvxp7Ks58fA60gaL3nehooW64REVwekWiYY4diojOJ7oubtUfKFpJSeKgPXGBx8
eYnMy2PFf/uESPhwhh+Zq1GTtYWEsLQdHVG9jSbfbcq6Hn+6s1clS7oeYp9DF5gg3W9Ek5p+x+q9
Hwkb/Og/r6x+R7pIU/1n5V9lJ1fXMIlAVDwyt6oMNnHp1/PWvljz0SV31JWfeVvxM/BRcr4ONADC
jMk34IIGkVepYzrc9uDf6LUgGVt0VCiSClWJLvGKg4ksCPDarWYTUeAw8zJQ3qayoGXZTWyIdKqw
eiTOfiigmoeMRIET4A2RuCxOQOqpoB6nGACpxUKwkFeraP63O+IBnyJ603AbF9erfVS28yMjVUH3
8gEVB8+CnXfLJyUz19r0Co/vxHKGXEsEEBMda9sOIP8ish4pJBEx/5xmaez6U9HugFt/mTiUgHhp
9ZKa8CbGRw7Wwlt9pTjJfI8mYaV/Zglphg0kkBHpsAeNtrNUV8Nj/Lot18U6A0avqS+bUZVxcRjN
wbFKvaJ1E7s64ANhljIsrjttO5F5Crc1z5hhPuX7Y/PrLq5lam+9l0oYANxo5RMHo3c9Yroj0WH6
bkz3/T1dOzL/0in4TWknC6UbpRaDP3vNEnfo4xpHQ911BfUGqyejc9b1EdJsZpFjf45/yOs45ngg
K2RxPw2uKWWSjXzBLpONc23yw8yD9BrZMlHNUHK1XXGL8MXHgcqtq8ioNY6B/kAogLLJvaCs0QaY
va2gPS6b0znRlBYxneVOev03VehnFEN0eH9PttVPpPmjeZyP1EUBtVKDUt025GLA9FI1YEItENc4
A0gde11dexkiQbGEOKhhj4ZdeWJfD4Fw3G64tjh77LBQgvL08Q7PYKb5PsRNcekEe8oLXYSTcvQv
Cp4sjOfGWb0TrURKsr4XlU0CGHPZRFmydPexog8qRQgfXxFJz1pS5Ts4jJUqEGxoogVJZUdl21Yc
xeBcQU0ewNinafVX8LZ9ytYWwLgwVkBysnyRWx+D9y3GrEPTPEdSriUwxtu+WELKRAnbNOiGBXv2
gVFv6uSGag/JoIuYV/hm1hYOWvaI+KuRzs8il7V+cvquwUF40T4ellwG0EkuyYPmsWVvsoOToH4T
PN7sEAmI0ZXs9Jq1Icpyew8mv9L6SRV3tjOIt/viJfyHR5hzJeLbxJecy93rmgb3c70yHSF6OvzB
2FJAQ9bEK5TKprF326FZGMLjHcDfdIHknV3PzsxPP50C+hOluvnaJ3yUWtlkf3J2GoOmZFA5WuLm
zGQGGURNUOuSQj3TRDz4oE6VHy/JLGfWdW/Kv4yRafxiwA3r2qvBbBIJdnb9fwmy2pRFl6ZRo4x6
Kb8QfXW07LxJr+Wwgbw/FEpOENHWXH2Dff0JFOQ2as9Ev9GmpPRa2jNkcSNZMRrCFvcnU/GlktCt
9RkzyQ3TU249nrUqEHigm9VV+hdcBKS6/cNBGMj7Q03f4vXvHBGLyV+fXUiAqEF782DT51tSCvBA
daShjrbIYkYiR/qEMIhzLD25trbHh8W2UnAPYkLxq44RPvadyRX/5dvmn+pZukel+IWBQevoXvHX
jEr7giaI9jhCXKZcFV2v11OqxmfQarU5YdnkNNvJbYY/+YWz1rNUiImMPlz6c8SexDM8eA+u9qNQ
EBn7BTlavSp8ZNZjFoDCln/Uz8tOFki9JMCkNhwAzNVlRHgQBLdqtgN7BwfA2TluzyBSTTghpRQH
r4K6qupfe+uN7sh5y3J+owqeJI8sdPQ+9yUm6KRwYHBqvnk32k90nmE0QTsi8eFVjjwlq2VAlnFT
EoYgCjknM1QgOVUzuhvpGrpslUkWpXLTjmqRO0NI17Eb/44kQaJDtHgabAf8UBvwNW1h7R4qLpHL
b69b+VRP+c8M2DUR6Lng8vO5bsBL/HrZWmvue30/qWLpHzgvUmHapd/kYZSvUXR4QlD/ASKYD9bq
HoJXzvKrGZeU+tJ8KRAFd9BaA4/HYL/k0KazPNkk0tDFXXNqOhYxbbzz9rvKS2FajqemlTRwmBhF
peGxJh8MnFt2eBqJu7/VHs1UQVSu63jlL6WKUcrGpsxGUm0qmI7pWiNh+zHPEe55zpWK6HZDY+Ea
9t9J12ihLjg1iwJiaCSIfCuYEYL/gcQVMYKCrF4c7vv2Bp7LFeIWyp2jvqe4G1TrNx/4m/YVx1+2
JHVu0MQyn9ttsa0HG5Qt4AwKQm9tw4f1zdlCm5EU+XVdSfOj9HkXazk0bj2UiqauRd2uW1dGRJ0R
hbPFaRUgaCBqmrDpySIBErg9/5KDjJVcyp8By1tHVc4+GdzLHA4Q4xDi/2rN3ulFj+eB/DnMJLB/
tw9RY09UDavUT/TEV6i6RYUpOgEVwFJk+wGRVtHLDgoQZdOh59zBSEl5JXdggFWpUfPLSTtqbK7q
3ws/dsxjbOsOsssIUauzQd1d3i5NC0g/p0IBL8mrIdMK+KxdjrbKXM0IXljGlOa/zAfNIEOR/oSl
CcgutaO9AD+KGGeO1bRkvc7ufG8r/ZcWQXYzn83N2xUFrwvDuXenDz/a2IGdb7PAA0QpZUHN7EQy
2iQntbp96K8s7LjFVbFn6KkLLUVycH3VywC5DSsbqR8nh/105s/vsyK7LnxJyEKtYrf/ALp6vEcT
YERaU4v2UWObyTMk2EueZDOyoeiGxFjtEyPs88qXR77Us2kVvRQqSUC11mE3OOCB5HwSYPFnW5TI
acko4KvXdS14OlTJufPfwQZ3IMH2BkFB2UhPAIHUIsU46/aB32Mv9kVi2oW4D0PahWZQgf2yLbjk
sCNyQ5E5SH2KTKHJliP+kWULyRzPzg1K0x05ZZTpA4t6TKpaWde/85XAxJzDKfY0Cx0NtrprTkcJ
BQsoXYZA/Igu1LH7O7GpjlWgnB1DLAhSrhusa4Eh8nyBqM4r+dz558ipAF81RFsXrKLI/ofkRYl2
8gVYpYr4qF1xyYbxIur3V+HqwOAwIaAiScSCf+eoYFeMxWkZuhZ3uimsLCsi+ssV+StpKm/IOLly
5xWs9XJ2ET6CkCpMtkXpTFFEYeKvv7CWvVdm7P3qFpvsQC9UlnElW//3jc4CPGg3WEGMWFzPMOSp
YgJg0LRt+rq6rzC9ZlDCJ2ud+Mz7W3efNjmfYYL6QZiCPJ70TPj3w1X9LTqSYJTiFQZrggok4/OH
RuwJ+o4mMJ3wLG45xchJXS8mrsuj5wc0/ffoPMyFdzj9073+PRoeQt4GzQ9j9t58VMHsKqNF8mrk
UnPpNektoIT1//TZe7wlhzxd5hgBnzvYt+RDP5uwzPE/HW7WAODuQDnS3SEzoVoyYNo/i5DtwgVb
6/lXyihz/O9gO+EYOJ8WEQLgD/sSaJi3JCh+XQIiONlBeUt8XewdPHlacM5BedAYYOyzjgPdL9JQ
4IY4cnkkk1WFlsxAtBDTM81Y70L8CF4yJ854rVsQVJjKGDhOmeHa8SgGUkrwhxrZ1OGfS4sA7JOw
uFU1IwhSUuMyOMTK/YyBnJPcXwA7k3lxuA7xORZa4UqeyruMUHY2PWsWz3kukWKwpAufmuf2kTsM
okVawpSrq0ScBloWrKhKHtnRC5oD6o0ib4z1HeaorbIaI4tbwf2VQ7baGLqRhwUdw7xLed0c+CBV
cfgmwV8s0pujSdN5k8IiVK7OUcYyRQH2QJ2+cYge0VNB0LiLTAm5yi9qX1LB/0UCMNa5JdUIfugk
dT8xeCDguQl+FMxEVdH/Mesueecz4gmkYWi88Ay7Mj0H0RicGb7G1Up6zB8FS3Pzw4eIO1rFVO7o
/eOdNzIkDZk6xuAkOycvYpBCmc61SHxGFux8qjLrWaMwmnFvHXRA4WwuhrQ0peor7V55Qo08m2XH
s2RVKtH/ZeeyzS/GkT3SueV1VHM4295GGparY+FbEN0Wx1gGvowHiLv8Uv91ZcZO6c2BK3zkg4oJ
g1BPEK2ygdS9tISrCZnTjeJu53FgKNNWKxILsPMjnPDPSLv3kjhRfbzsW3bWej2XUFNwHd1yPYWR
cv1qB4NUtvijPPocs8Ir6PW7xr4lqyOBviHI5fb/iZCEg9RvaDyK78QCTzcVaWTGLq4zrTnO19DO
5jY+ZXyFb/z3I6D3K3EoQ6bwGfzM9n08z2bfjmmFCv+2WJfTDhIYzrVB0wDWtUwchz44KaIo8mQw
qE9whn2gIunboiQY8+XGEA0Z24GC4OqHOtGbCwZZ1KTvMXlRcolnDL1bKmO+lgejVVxbOV9lgO3M
2gF9APthXnjfthA8QGNghco4uaXWJqrjIPyr/H0nYfu4CoZ5OkUr54B8IVKiRrSFqPMxZmvu5JOe
CDcqdFSt1e7dYQTOwOwQyqFojZBAHIv+Z9c00pSjGzFSrh2CrWYVURWNnAXhIetshNSXO7bvwRQz
xvZgNpefexOp1UykxlgZD2lUQn5pqGwOnZEa+UNINRDktPEnApg9kt/SlBCZJuxdGWoT7Q+6z7vv
bnA+t8uSvUx7WFCCbB60uaBRBNICSreqRo/9YRZFsc7XtRrzxnaVAC6KnMt2MUJhN1ywV7BAuNAj
00ZDr54X915NWQqZt7AicjBkhmVmlFjWBlDqkzB/kEIttcrGYzlhkVdi1SLDNGyxvd4/IzuOolhQ
E6QetSoHjE3L3J2xreScjA/CqAMyylRSsE22pOxWlXEaJgYS1+AngkMJyc/feY5r7VjO7gz2rxe3
Ts0gIHJDfZHXFuEMkvfy0O+qS4H6IOfl+H/HcBa2DMi1uJPKkSMNo+Fox7Rt0Ls6QZPudbu6VWKY
y7CwYZ3PODm/w2Y3JxAzjMV6ioPqsHtlhL8nvKkO4zQWrL7JdMKRsROkvC6tuMNntjsZHtPpLGer
kN0kBDfy9PkjSkUaSA20rmNVZHtIk/idA4J7VoaNCFpTCyMdo2RFgILAbFErkZiorRoZ+xmhjIVs
ga1EVvGfGe4E7Grwo67/YOqjM6P49JzCkMq8Ao5q8FaQ3r6bM6RpbxTMcZ8660kEuq6AgFmPppcK
dRY/y/AkWCfJMtNsXUl01LD9r4CCy/DfVFhRDLzIWQSCdaz8wgVvql35LdL7hULQKH2ZqGZgrUbP
FA4zJneIpLZrILAATKbRdYSeZSsAObGW9czJh0lAAiYvsEy3VG29ThKTN84hps2HnnlsGJ3jSGBL
eVJU46ngvRDBMZmodzKEJHTOGaUEn/WtAgX6yF8lIDGii2vrVUjhQSdsfsfSxPsLv9WV4GpHNptz
ae6KUsV6hNBDO1yGc5I4HPGf5hxf8xknG/8lN7c7GBAt5CyTuos3ax0MjbwsbLcM8a9wZ5om3udQ
bPN2sKbp6Ky8XfSqp8nr1XI6bzdlyPRMH1GB4DBc+8juWTKmnJjZ1YlpWAnL9lAS47dM6u6Saxiz
cpfJud+EpTyz5hyjfsl0Q6OEvMXu0dTuPV1hTwekwUuxc8hNvST0UIybWGf0LXCdfhzVJBKxAr3w
mKpA3lV9TmD5195inPFvvFq7ILQxjyeyfpJRPuM+35udQbmvf66DLds+F1iRBmHHWtpOMmEz4mKZ
bHjEU8xXGeKooA3WssQI3pHdRIyOYTpQ2O788CFhdSnODNz+sQbLjsoN9ALI16OfyU7dgUlY1mkH
CbUsBApFtwG8L2ofMJXqfc+4KWIi6bONObMGBZA9d4sT2EFoZaGFGE/y38dMXoh2C6J8b0SQRZyV
L+jX13EV1QEaF7h+RdJI9v21dziIwRIKzaJ1qPHb6/xekC++GDpsvr+QG/eThOiEHfJ4yLgPneXF
lUETt9PUcfdKYGtkWgG+RHViXGw8/zi950W9RDNspCvfNFS6SEYOwkk8vwl/iW2KjAWgqEJIlFL8
18HEawRSnbsbhhakzVDZJYwvSa2VEH1ovFsi3oqym1hqj2KeZ1X2j6GdsO+aHcNZI4dm8B5wcQvF
aSoM/z09uHuI7c0cYvb1nyBztz1C5TCzmecis4f+wW16mrSi/5adI7SDs1k3ttd2DG8fXiLR7E/V
DXhCVPsUD0NQL+AiUN6fCI84wrgOSrhdY4GR6eG7Bar8N+QFZllM2jkhTnHUJxAkAM48BZQBc2zz
bF8owrS180p7dDahqbr+1m+f8TZphvOawdYa4XiytQ7bY20tg9RUY64je+jCS4tpyITnfGq3iwFy
HQYRBf8cugK/6kQfytJvf3jS1Tvh4kIFCur2pqVBRKU3CNxMK37srhI/Y4VEVPB5J5lU3f3VDxx/
kpUcTBaHXh+oGvKKRpIVYUnea6TkYcip5WP6wg7IZbNaSFeNpLt6IIH7MgkSySsF+Fa4LB/BQehJ
6tauR2Tv6VKII/8pp6C0H31NcQnanjPYKp74v3flglW4etmxb+v7QKSN73eLKHRBI363zcyCpZ1+
LDW8mNy5mZjUHTBxievByM/J+Xhi5NaIGlPoV/MWSr3qUcDz+Kt9YxjSQQcs6gwhzCAwQJa3/7Uq
l7TfLtQkef940fSt+JVET+W/A4tBDx1hP5grG8HZ/a+JejgcxpkojaKFY29Ek3OQlP1R8whp5z4p
qvR9NImeKOWVQYBBK4Nt/eE1CQmB+cSx8OEd8vlfWzfpmGx/r2C9ohy63NMVihgQgvXdunFqYQHl
7hTk6RFNPd839YtYR5cEaZPDqCPNHRqzWWZwX0TPbMRPj4GyrdHFQcKR8+rmbFbSKCnz/MzuzcIX
sdDHutC4QLpvbHcEdlPdvAP67AIgHtktLlFJjkGmzxexhaDYNBmaiQw+MFjc7txYWBjONkOJvHeM
lgyuCgbi+8lRr9CX/jB6H/fVHrZ9OsSK75ViJfrL2zdW3UOpqkGy/IIYsQDhL6/ap0Ko+hvvdwBg
0KQEndbFqsCgHz/FIRkAwxf9AOS3LPVlCe83l+e9pQb9umj+QI9DnZ9l4y2koh4Hdphzlo83G8Oa
vj0bDR4PbSwxCM9UTbFKmhzxFJZ3FNiNgIqjcCxR98Mis60nF2z41wGamvJeDxAR9/2N6PgwdjvG
R8ML7QTVsCuGazgxyaI3SXitVaWJEEh7cirkcSFndpauWwSq0tCdBhYt9vb4cGDbb8ZhRoBoxvcV
RBmWovVLum8ivMbneHFAGcHpUhLQlUmN3KhCsPWNNwqwsme4lfMeA060GFqwlvwb3A+8L7fIiHeK
4S7bLnuWVxbJBkTDfQC4yGdG/Jic+Lk0dtdTHLE5cBeKnRjoAwoYvReKXAYEurDDYCQehGdb7rkJ
s1D06azLF2QJAUMBSfkDaL/E/f7CrjuL+53u7NEOPLMPoXf94md2/MPFaswyBwEOfeVpTVVnALJd
ECz/eFwU8LTAFyXhucPzI5RkeuRKLNXum4vnoDN+BtIaGwZLqgXIr/K6ECkHqafEANuMGpoeI/UY
VytelrUlxb1yUiVGkDVZUsBdZc/lywivFloFyFLw9K0nWRuA/MFwfEQfSq4W2dG005/mNROpL2qd
o8vh+tIdBlfScxZLcButfNvRvKM/mOdsEi1TT5lTEmDNL1qdxP4wKIORSWaBSHj2BdWAOnpBhbqn
kdie7VlLpwHw2gyVRXnwLN1vRFr5wGKFfJJXRiPRlfbSJ9Qtp4+3hEdgA4FyARu0D5cVqXDSIRJ4
pGu4L69mxSrnZvOmlHYGlGS2JOSKlWhJQeoukmKi83BO3/Bja/DjzW2ro+LBXcAFo6DhA5F4ppCF
/ETqU1a/6Gg1XoloaiZsf8uia8eT8SM/eKWCWXXRsgK4x6BQWn3QYK0s6LRRqUUmFfL3udD/Pm+J
M/ez1W7r7AtpUDSMdGGaX+ramc6ld03Lz2x5xHUSK9alPw2HXtPlvYuQxkIHxhu/zSfzLnR/Qy3P
W8IuNhReSes/kXECzu+12hSt4izFrU+kOeHnMPQFox2fFuHAEaFrL71SpvraNQA5fNT9SLJ2J7X6
NZ1/LXhnVWPjhdm6e0gMMxLTDoMCV2kt3wpweIwLgMJdQQf4+kI4z/15sMnWzTHJ8XnzneZZkV4w
S+cOT+1RE2G47CbSTAb5fwVcAKkEBYISUHjXF6cWscQqZfFzLrKEqgpS+NMrlrrc1gj1dtRIUfzK
vJmwv50Ci5HRlqjQddODZ/yUE1j0cE9qWZBNB2vjVuvK5wOwlynamhPN+8bwhJ0lHOUdjrS1JPOo
UCzjCjIUu8UE8DYPlz1PcqMTXTLM7Fh1tASoT0EWoFWBsDMIU6QqMunj10MPKpXDD1egiAfyiiBV
ZgvCivVTFMJr2sVWZbDLOvFdjxEEMhkuWT6H0sD2aCdPQFm+umx3NW+JC4Gk+JlGeHVsV32NwD8B
YpuAZURGtXagY7VDCU/vf9Vjf09ZFijIw4LSzKZeXsLN7gPVZDIanHHQoC+E8iC8TUjDtfHd/TXG
e13kvYYluwyLF3qr8UhIrxGcOVsbuiogHBVIvmn/t1SiqqkEYgiP1rvXreYnu6gAnfuV4yg01xfC
PiLZ1/sjHmbQzW7cyGbrFCEJ62IpqKr+8LcnPx+8o+qeF6MwdrLX0rjJ+u6nNGImuhLqPKUGPDr1
fbxy9llsTT0H/MfeyTNJQyKP+aeyZtaSZsQfqtIjk6zEmS4b0fBfTu/1CVGPCRoY6lna5tZ7CHs7
1ZRWklgA3uDOKC0Zm81W7rlJkrzqhVeYATMQdOwpzIpolVqspX8ufJaJV3jHv0VBYI0ajXX6a1qt
DiVH59IXBYVOIIxFs275C8UWEAMwoNbPKfyaV7TVcyH+su63wpCVPkBSAlBqAebl2BgOHKtqtu7B
UfGTJKwcD1mCEED5OA1MBeDjx4MaK6eIUUK4FtuWmgMfegrXtE2Jq8ENHcka87yYVmoR4sIOW8jX
qAJ9dzD7VaPZcO8BshLW29X0L3mt+vXjcobU9QUp6QR19nD15MMGlK/ePQLbne5R0TvEp2Vg+y0a
NCZMFiuRiTKZgZPh9j18fdenvadn9Y6YhK+EDXvXyE7/yKRVi/2XgM909YCebB14O8uYaCMttdOI
vCRuEAqzdH3w1O0fw83XuUZ327rx1XD66Zoc+nz69RVvO2cuFs7lIjFsXjJcwkfRiu9odh2COH1a
9jLhOqaLEP5rm4rZjuO4CCGNfMKFK7pawqCJ46pqWFXjsNWwAfhV0ghgkQqVorMmU125nLH6+mZ0
t3UhzNCEWuCC33mSyKf5QEg5z9pBeg339heaHuiJzR1Mvmhi0IqpCa22vo6oDaERZiQ0WvtQT1OJ
WlGz1pKIl5YpYnaOFqVJNDOop9G+1o9RK3vPu4pD7iRXzFd5vXU1P4rV2Q97TH7yBd9Q2yx2TorG
w9h4zvS/ydW2KSksy3VHy5PpnaRvcmE1gC4wxdtE2LtuOz2UCffkxmuWflU9GRnwPIP9FXNG/vPm
/n9tsSVBhOHFxxmByDlbPfYGS4PJSyCAzh+p2pASWW/QaAcmiSDYoUvO0kgcehWO6OG1fjFc2wYu
z7n0mxgJmuxwCMrGNv6ttc4FPzuY66049mejemAky36BijB0PhHnKzb8YqCLQv3NSCS71fiBD2TK
3S9aXyA8A4JcFYPaqxa32n3pS6l8cakCg22YmcPehCiQRvM+djfAS+wuxzEURofuDqyqzX3ZksCu
EGCj7PhjsYmyqWFowNxnrfCRz0VE46+lcpK0zqzF6Apsy1q7O366j65vQ8Bu1jotRXJ47uOR+p78
2j6HW9SdckIslQNU/s6GC/XQV6ek4Ab9vU1aExVoZ0+SUww0LDBRqBezC3ZupWLqbD5VU7Z1cnEm
GHPvTzsp13kEA99nwOEi8s+tCZRvjVt5UCtyFiSshQb1pMeWIhCBKwhBec/jaytAuW//f1lx/FIr
lN2t/uvezvDHvftPs7mZKvpa8XrXPY9y9N2urUVy6A6/fl1VocfjmdukeGFT4gnQQU5eBf7Ua47J
5Yv861nOSPZNs1w7FpMbsXrgeyY3Oc5OxjcjHWBsB00yitWrQ5N4be0+cgwkyuX8IL7t56zV7Ec+
EtsiT1l8uO0rFL6GV3ROSGGxwZZhPNCtEBcVXbeYuhc/ZfUqXIVI5l/wCjUEud/hbo/QSZ0LXnU3
UC+xnWPCTVAGLdunRh0DLG73Chk+Uy88BWBlOYR5uHFl3RbX/6vKCFfSthISIeJLS45MglbJrm9Z
jLoFmQZg40Gxr763BVosC46OZ9uIUd+C4g8cRItjXYULy6fsLt5yBtgWrLVWuBWwzJk8N83VsCjm
RywLNB8pqIUJ4YJe7Yfftmx/dPqNCcv7+eTdGvjzO3+UX1lZKj/c2NXJv7LN8x1RvXXfZThJ3C+v
XMTQusiQg5IUpBWvNZQlCq1khN4Gq7R/XYia9ypXIyne07tB7A9/qc/X6IYGixNGUmauspT4VD2t
b+RFxmLVFkODqPQaofzQEsTWsemeBseL3w3QoQNIIFfciCZbcCCMC6jBpRB2l0phZ0YS2urOEK+z
uPbHyz+juOzb/0+axl/Tkd/LBK8UxUXaxkSxgM8fHdxFQJBJbQkZkYefeFNDNdqhvC+R/e6R8SIw
tqpy7k6KmrKkccTgEpTer09oAw0baKewG+mtMJ63AnxNd+KvwOLl/DMNZ1Q/B/F5KSOWsj48vDT1
WS5XIYIa/fnnu3Vt+VkOam5Kk9296zDQ2svYq6eVpYBlSzAnaPdb5ZiiHK7I/f7EBecKfDuObext
+s8ngss2dgkXAy4XY7tTGNKXYXsJeG6l9E14K/3Z+caOMEFHbhYL9O3echCFNu4vSWNddfydgPBQ
D3l4njWu+c9I/G87cdYIVaQI3qmOOm9lS1njWA8kjrVq6io9XNPX6w3Q++D12kzCSxmvtMqtyjv+
jgJSO32mB25SFG12FwV9dW5Z4sW3RMQazMpjhoxeKOiuvYnfH/SLgiZ76P/X4L2eEeWpfPiwlVLm
4RzCy7+LMxx4e1U44PUtAx1crhqKAe/VrGK8mjQF+O/iW4QvRBkjkGzWuhfx0SHGhdl/SLzBOXQM
i11IUmbWe2rEKnuobgJd8HaEWCdxADrF8g3mWh4Xdh134YRl+cRLAjmFrDQsvUi6M4HTk7jaCkTd
7XQd36MIRhmASFpGhZ8l5B/Vuq5+ynJGIU+zEuKW7zDXaxa8Bw3KRYB7F1v616lKvOlL245yzPLd
Dv9UwKhBSOiiBypivNwiTSyuhWx79N/eQsvVzPzcYkGfe7XgGe4b/T8z8/MCm1X3WGzqdpAy5Pz9
WkMnIl1BI9+rr7Eb1kqbnsGLqwYCSiDADvuZmgnPWxb41iNTc+S0J+2OkEDh/zTxSh9I95y+0t3e
iav6o5BBCFj1xfyTMwHIRUzdYXgBwq2HN/LffcaG70YzExLoqJaySOongqBLz5wVLtbgtYD9aI83
+++3F2vlli3GyaarXN5z+A8TQu/ltWbLtX6sbC/EP7PkQ2+aNZ7PQD8gnKyVN/Mu0+W4ZGLIsase
ycM2ZxPW85Xb2MqK28XVfD7OLBTSqlxd1k69KoXl5dYI5iEGr30cbKuBUOQzK7lenasqkuAPyIkh
bPGQAi3y58fHN9qQqBB5HLLi98No4nEKxfnM9f1kziaXwVPxQrguxg/iVT4iwE5kMj5B2GxEbvP+
YAmuO5qiAAr+UhLb7+No30y7HZFdpWTZrHcspE+0gIz+/mCCjeXp9YvCm1xi2dM/tSF62B8+wzli
3SfOcW4NcaLMR37b/d6CSSKucd7kWnFwhU+xP/MnbjgVrPqnR+9PgnnY+ZyAW4S5/14ahbgHtl78
PwFkobQfRyfgGvHs4zatZ47er/tHsLvS6EorAYGclxAwMCEw9xiemRoE1nCbelavID735Z7pSQud
GKgeRtEHeJhj0j3r6GQn8TVFLrbYt0evfpBvlodEO5NKNiJ7IJYRvfwY+c+TyyKD8JZSQojlurg5
M86D0yVi+L/+h/VMUPXlYgCbun/7TM1V+Y5RgCjyF78iCscqcS7tub5i22lw+fe4VvbOfjgsCElD
NQ8FLobtQno2GvK/8Ao+C2L52hUVEyeJBbdcled5nsouL02l9tOkNm67AostCsbMTaFT+QgxPANa
HCmx2U9ip+og2EMA+3xedzNDDwQlIsloKgG6tzg6D/JYdPZmUO/bdExrNVycJU0MAXauLHqkpIae
ysgK7exRrlfzYABL/piErS29p/EkbwFqJC7JZuYpNMuqDI4TdjzhA5B2S/h7LrdFTfiYpdRsdAmg
fmA0IlavYLkGeK3BkXdYKChKas0vwXPnxXZCR2Vu2KrsBlKO1R6CMG1HqFPbEmAMIy1r6VRvN0N1
vIK58jrnpIPIED9DNksF8X9g4LjqDBZa7cgHSHQLLJYVuiOpw366UbAngzfi3tIBu5KvhKzjM7js
gvRYkD3EvqSo3OYnrYmJujcCHPzda6e8qG5wNZj9xaXo0mUlh/vwPRGAUuVC7MyEevdRxxkzV1rd
i4Fw3qGWIoEeqwnmT9ZsVluMBpS15vPju+4035DfsAu3/PMGCDkcePrNrfCvrisDtP/aJW62QnwC
tH8Z4IP4rLvGLj7YGY8WSpk8Yw2neyJ+W8oXu85irSfDP7O9OXAzchpRmInn9qDAFc7UmEYWPmcp
AhJDn1T1lmAnc43qtu2kqsYYQqIRhxHDdvhrzWtukFkHbrJ5kxeKSN8qkdYArjUCC9Rs3mixsv0Q
yHGRSku7Oi48fUVot3cl5zZK1chKBpi5PJB3SYt7VMYXfq2g7W92ZUFai6BArnwOq6+NjtRn543N
YK7fN2phCIULd7dty9l80iGpNfelqv4HBNjZxiqh524ey1X0QPZyO0Yy6hZwJq2waXRf/Rd9EumD
d9dCczee9qwGG6xtzk+XnmJx8zraXqrNiyIgocXenW7rrxZmf1L8Fpz+aVXtxXOWe+K1ZSQTHG/l
abE7yWR2jaivzJiiDQPS8UjLRjI+m2sBZhVmKP0ElnlHkUyfflDMOHP/pHTPtR4I+OCdcodKNHQc
34zg/62YUDrLR4NsWrGKMWlN6XIqYrT8jujBbQqPhF+8Fyj5IJXvcjXi6KgvlWeGSmdfeBgZb1DS
EjSB1oDVEdC9N7M0DJJm4Vz/4NO8JKtGN/+wjCbuAJ/kXx+xB1bor9OVUEdFu9s5DFhoBadd1/Gi
aN1YiGTm0DLnv5lls5XYIHYE4ST4p+kKwYH9SlQa/KBvKPH/QBvgvdMoGMZ9WSgw+mS6mpC0oBYB
X/KaYT1rwA0n1VvFJyAruma1Pa+CB7b43BFF1UFkoS1+N5mC6YM12+zMRiYObH6KgYH/9iEPEOof
jbHKFnHU/v9vu3+uGKyD8jZZJ4AH8696rjqGp9MmBI4e2tMmY0NBrnxDvdMIkKNUi2CJSbglcXt6
Of+Y6M2H5yYAFhio/N5cATHva8a4lWJNUvrMQ3Dj2XdMkTTKdMNKSztNIvTYogBkow6KKI9gFpRE
r7bRdTwqq9cXOLA9OrFWeVafma9SuJ5Lgb+zY4xZ7d6tGBGWC1+XWHrQoAgkVhaLcYGXVwwML+oI
WGzsPLR7YqXWxDUVdsonOc0W4exnCJu23m7dpASwZt9cJ0fbv56bykjvzmhtywDgo1YJuWJ8IWzJ
XBUJouM7ncO0jzUiL1A33iSYmp1bkzcGGnbsIhcLwLxF/ucmYIxUJ+ZI1zSWcDtxl2aZHHT8YA6o
5bGBHwGE0YlyYq2hKHmlLnwoMbXdC2ip0oG+xjzqq22Wg3YhROt5uKyTA6TAfVT64OCyp+DV/OLd
uo8h2+gC9uuKzM6FL/5Cr9RpGiaPLqBdFpaRmskvrGgdYmuqI3vnIwpx6tKS5TF1eoQLrrRbyp/1
NQdlW6rkZpxHN7Y8FZuUWYuN51wfzRLRsTkbZgOYMu9D+PfZrtZZZkoOeiihdg8kIXLQsgsAhEhd
q/0xqQ8MwkMGkti6g9fmp5LkzLQ9FM/79jEZO3gpbM08jBzwNeC71sH+7gUWdnuGOCEZQFiciOzl
M96dLEBdmIU6m3aIs3mH4SlmEP9NJXRP6yWeaXKcnQRDNLVF2WXvYmjrNT33xBA4QdkndUs3yD/R
d0wvNKRBWZ4J89q6hvw+rn0+hRMiqnt2wJ2a3MSP6I11kytcGE6ZSWULGO+muz2g5MDdlAMdaKgi
d+Gsai9eg/CYa1i2CDclBalkxb0OkArO+iqnic6WjFeHFRip6QtoqYrmJlzIiNSFIw7PC6Il2hb/
WmNHfQyZlGvI3239XAVgrIlWds//zrTxrVuK6Hzr7f2YltBMJHNFVyDVoOqReQlzmGwuaIjZTnra
vCotDKaLwNwV8FSewXtBJSSLVhaCgqYF3weIlThKFbL3j4RS00xYIZgPTTqmgPBLXRI+Un28+tDj
UNr11hdiFy050ATpsK6bzj1SWHTkKryQ2VxbZRmlrJuX743w5dRcWXqBEpzXwcdUiVy426dh4S4e
cPrbAgQRIB0B2emgIygAKnF3J4osMhIF1E884sOxZc0CylMMI2ROulLEtlo8anO8tlzJxQhswKZO
K2XOkIT84t320Tn991qON3n66tEAXpKYuQ0iXZRk0TxArG163I+6bSQA0ZSFvMywToB5sMdLZ2GX
B0dRfMJ7zYN9Bz/RBNtxKK2NKLKXgq1HP7Hd76MpDjLtGdbUg4EvJsxFRwG2y38eBGnBhybMA9Vp
GusBPzqjyV6tw1YptyOX5jMdS/9/VAVoj3W1VADkZFswLaJ+ZtW6mWryraeMw/v3Td+2NeNCzaFR
hxnifHxutpkEZVs0AQvCD1wvyFxVRAjCwiEFxrgQsswFhYN2M/PevoEo/d6lNi+x1YBWvYfONwys
KeNxSjwiue3CG8/98opxu5mz7ZvytJP6ISq0GVBlhc3RBoOfAu9NFmhETsTzGD9LaOzUY60OMe5R
Wt/yiY4W+TlysVgI9EoxRQQKrfHhErnXXDyU73UzE1b0jpA0D2DXeafs/PDht/ISDIDLkJrR3tpW
0RdmUT3N+TilMDivUv0Yi0OUjLvFCSPj4MsbWlXFpu+NuO1YFCKBzjow5WUVu8eEBhd5TCCVLNsp
9j62xR2ZmuKc32bEzpBnhReMVv3NUaDSV9vXBQVzvx4DeILbldBOQEkkwqbUjRe0AaS1QAGLohzE
ck5N/HdmqQjBIvPpT3BNb+jpQamYFFHxuaEfeNQy7R+dUvRPKj7pn8S6ZEUboZQs9i3yPUD+a5eW
p3prTG1iP1z48BnVSLkifb9uC5pg45G42BR0c2gqWKLL0kM1if88iJgV83tzp3Dvq+WuBFetvdqw
q0DABaDQTmSGD0hpA68flnEqq4BNSEdXbaXJSCTVrfpsct1VuTOscOSDFuWJHUd0/nh11ofmQLmD
sFwH1XMiZeXRQrZN7aYQFtcWx/USl5xsAlgcLoBPkBXZYnPmRnEQ39brgHvdrD2uUmQDtw1PBu97
AcM1URiPCfEU2FYYUoIk+u5TGSM629kZoi5CJ0qhPHh5bVgU/5o1qlW4hwX5k4DRYqkJ2geLVLQ3
ue74H852Bw6dhf5pVBtOiPIIK6mlv5PN+WEDEiWxdaYFpPNJ6/EHMLxShGPbQ8gySU9qeCSHm2/c
/r6yiRaGTFx49yqBQt8FS5ECTtLZuCQPaaE0TuWiRvMeVksuYn3GdwPtV1puMXmS2X0XY8j8blWQ
7xsg5bMoniP8zxD4UnvaZoEldwfePthcoJQE6ulOaPaBA9JWhM7tsnWEw+aL6RcNbv9d03aVB0wX
aB5bvStnLGAmrcR1q2zc6na2bXQx8UCjNU41lqcy3BGi9uc80be6n8d2XGxEIMi/gmStLW7+SUJJ
/IxfkGVPgXXRwF386bD8K8+EJFkt7UHST9Vk3miHmVKyhaVNTL91R83bxtz01pVkan8x4GLjy4Sm
Kv1IExCp0cfg9fHv+RTA0KLEAqmkU6mDlmFQcJOL3sXAawDsBuX+vec6u9FMliBQU5Cyljn+xjww
zybgsvmB4u+HhYScmR0G8BaeMGGPdeBRvI9K7KqwHf2aUCTS6mYMhiTDhqFXR/0eybY+R58SRW8M
XL9t0MN5yjSuurj2QeY386v+E8eibIcVUKX1WgSI/T7kL6ZlyHGRV+ZPtlJ+OTRkid9oiNkMkGzH
KLND8CmYoymw7wDG3CUysvOTNUaG499+5OW6xd7TfJ6zNSsG2UHraDuP1ZJ7R10rhxPcBTux3K/K
f+ciORPmxva/3AmU39anL4dm8V0q/O4iDrRFCNJ5+YR/v7NvfEynCgtmo1ch8qzkRWEuoHwOe+TB
Sdswi1dVL/NEzXDLTc2iqdH8Tq//hby9T3LtBA70R9xDIqbj+h6o6AR7UFNVugAl1VcKl/XCik+Q
HHEoTz0kIvBH9CzAdQn1AeI5w9Nt+pJj0EYBFYABwd3wBUn4tw/zpabcpzEkRU6v/lFwlSZmdvQI
Q6T605K3PeWa/SlxkxNcGp6p3xvU5kl8Qn7egaBhavkgA9UMP195b8xTaE954VRjPLtgRyGvjg3x
+eSIXHTs3NF7EBZ5/C/ScuMYgCTPtl5mHqBLjbZTfApKj3GIeZLibqu57Y/ipJJnZ5541jefKnav
mjZrLgoVdjCa68jyBuT0pR7YECUD2uWTn/0/CFKHy1gef2VfdDQZx+Ev0AVyhydac9k07rZYH7B7
vTEVL5oRV7SbB3qfuJK85HjIBjjdWwp9BGGnEo46pMPiMxILD2dqaDI1qladxATej4l0rZVTX50l
+lj6wWO7noNu++23cqSo1UgdYsLJVNVuKZbqsYboPn2USyi7Aq2uEhxZYsMrN344qkXs68qpjLuX
aVpmFaX3MK3e/dVaDY1xUMF+ZKGeE3gn9W4Z8jjuclOIV0RAc+eHW3hb4k9Gez2bm+N4TYmhOk9l
sTrxko18XlgYSDEqurVk/dq2tRU+/wUqnWt9o7HsQUFs2QCUSpX5XM4zZ3sZaGpJV/fD4okduRm5
oDl1ewikfABce8z//iupYBC/PRLE4bdShQu8cnI0t9GVQOkcaa2zemMmFL1hD5sz9egPWfBmpgbx
qIB9wo5RHOMiTK5/Nvz96dQvyZZ1F5a3izj7Br7J+d0NaKZ5AsPKhWF2m8xcFGYLoEtLOitqwQjg
JA574bnl6T1fQWtrqSErc5x0cP1y1QCTCcw7nY8MCZkWgN09drTuv2dh2lp/K0IP4wF5X71nQUfR
pA9aCthPRIfr8qM+XzgI7Ve3QPypJsSn1mo0vFvLrJv8v/gHq9dwnClSiQdDyER1Jzd8N94P3hKm
x+xp7O7bMMQH3vHI3gVBDSr6E8zG0t4YEN43YBOwsls826JjXkJScm2nWbbXwwItdGUsOmsKgS17
6OBJ26EfeBoOq2Q8jyDVAT/jJJ7lDIGKpUttA+GTbkfuKXX3XRfU8joVJM6dJ4gdtrzqdRh6PUIu
7oUEFa76qcekFUsTRSWc/bDvzRgPwH6gbI6HRwEJtR/1lHPiFKamKXl0zEljLUqisqanMXdmG5xb
seVDLNCMwpC9lI+nAVLyZDmEskW7zRw4oHOdq6wUBgj+bsW/CoXmfRdtlvLxCxkYVqlCkBSQoPzy
WRDwvUk00NJanJgHMmTjFnzLe/IiOnOGSvpDyN3VaaQVJk93u5SdmcNs3nUHIpq8UouRZV25a+vC
FrF/7pbbR4i7OHofwp38x/SLAtgx3dRJN1dK6E4Iudt+jmv+HEOMCaqYtq9fdmlWhA8fsGDJAfPN
yYChnzs/bEvw+YV/vQe+HnywHzK3bEeNEKecXoa3YMdCQvB5j6Hht2NQic1cJK7eDR96Cpf97iLD
59xQhJvUWbezOBd7BKadoEPHStSMhxy8Yr84zDazYtsyBXRAIWx5fDrfZQSM9KDto6ga/CQQ+Ver
mLy5NihgM0QAqAoKNzHkc9w4vpRXLl+iIKDmvZl6AsVjmbWw1aiO6LFRXHsAPYGsx5jUjZJQA6IO
aaOjT8iOBpvz+YYC5fFtoStHHeq6gNpZoyEWrW5Z0eVIRP7g1ThSRNHA95Z0rPdb62b2GQwVpHD8
7N6SNjtmNZU+RGX04L9Q4vcozFEYHi4iXEqGiAWKi2niynzSIt8+fEszcDa0DnfCGUYiL3gA8DAY
/0nYhcdr3AEqaPNHsT/7tF6DZG+NqWrdM/6qnwgcX+wqbMFfyC5trdVkbcwhbsl3ET2bRyo/KeTo
b7YwivCLSBOtN5Ihy6xpHBISNnFXmJSEuLOXwDzEq+l4T6PidxmKByjHtpJjZSkDsbku5TdnvQGD
HT3NGYw3gfb6ceHg+xKLdu59rTzpRckRfbYGlYKOFDC/uqMH4+OiiX/AdmSeJOVJvuvx5kXra5kz
TmWz705LMjUv07l6hEl/ggXmZs9S6GsJI8ndh8WhkZ6/OozF6G5/S+izjtuoqPVSk44hnQqbc9UC
YhSKq5aFRPqzfWoFNBnox1XwM4jC8xtaOpV4GqgHSW6evnrVmPi7Vs9FeH/fU2zg47GfvWoc66VS
R3DeBFUFAUP3Jzsu1PneJ7VBjLpdFGK67N2KXUevhQNBn7mCYSDyyIpawMjgAoku9QvvMBmsp6tA
Z8Uk7JbPo9rEDYADK5gFWpIPebB/6QKulsq0LOuR3GKeU5ZkvcO1V6T7LAPlNpqqZKqRccGWgc/0
Bl2JO+hqF/v35OxPcY/I6VxgV2DxWmdZjMJAltOAZUPJS3m4zaE6ivU2YvTjOraFezh26CzJ6qPw
uLyQoQz3Ucs5FNlm3jPBfa2u0ZT+Xq+uiK5PODTLGvrxLD6iKhc+VuAO+wHe+QFHg2QmnPt4M4q/
NmKkmufPGg0ZEK1PJrDNIkUCjzD0fDKXYRHqbmkUlHujP41/8qqj2zdBWpvagKkK10FwX+F7Wyv4
MdnyDuX/eRyI0DaZy/BLg6ez013AeC2wa2bjU8hXgGcAgLyzr8h0buuvUA3Vf1YVWktTLCC8TDPW
dWv3jaU7opbTmcoMRdXwWOioghnKye/k8yb+1y/Mw0KNk3tNBhMHX6PbrRbDc3xYGjU6/pEtaoY9
tdUTPTWLAHzkDaytuCQ7H5Xpm4ZA+Wdwfrfil74y95gRz/XhXtxU1Y0mOcJthrCMAQHhUc2lTYlz
aycIsU6vFOpMgi6kzyQe3BaX3lGpJYxOjyJuDvq5V0VSKxuOxCnFgYhZJQ2sZgudMNYPjvnSDWga
bqjOiFOvJ4JsOTnr4lUppNt4WPO/1wy4JhYdln+3crFAlCLh8USWTstehq56RYAF+slzosKfuQMF
BwYHKdJPjbRurWB6uB4pLM9+Q98AaOpNGpQeTuTfyNacg4wYPgpUuimJH2IepiAFU4AIBzC3UUUi
04KkekHGaZZoGK+BXKdGjHC6XkorSClB9UjFYUAYcWzNXNb8DowcWel610aCMtQiglPj8O623T8S
Dk/jsInGZodR2RQDgVXk0aZ6bru0bpsNhgsjVaY8rRzg0yu8yRvmQl3ulMrvTy9CT5y4KGCkesjf
38Tlhve8yFhCP9llD0wokZ5x4WlJTjdnxkTYi9nTR66KQynTKrDexgz8rLFvAZGZ4Q51WnLHWvvk
bL/XJPKSKLwoZlub63lhBKM4OoYc6/hMWk9Y5jeVNXuJUADx1GwM7lQaagmxhfl3aBH5OABL37IC
1hhDCQaI2LwjCxrnDPn+9oZt2UAx5KQ4kuNSO4nt4HY4XsZVEakMflahAvWrhhCpT1GbLoGfTBLY
dLvjk2MqqiThpS0fXWHOwq+EVSgkIaTDz07TVoQYitoFG4VAI2TY4luzXWfQeoKy6WCJESleqLM9
zO1i1JcEcc0+r/8XB42opw22LMqNRiS5MlOCLq/QymzIdCx5Ai/6sG8FCy75CnaAu4XJN+C+O6Wn
mxt9kilIzfFLA7M7DhDb8k4dCIGakExNx75a/Qk1UOeUyeLR0zjG3UMJXVdsswh5Eev2OzKBWbgS
JCs6JkV4m5kjnyNU9dtjNkITib+8QD2gceRplkpbZBMkVbzgUkc2MUZqL8YCHKwewAV+DccCX/pa
/V9k1nxSozO1van4Zb6EYZfyEruRH/qQrm40/Xo/VLGWFhtuEpZ0tGPC8ltIMdi3QxgVJQ1KtAzV
ENJ/V0AC1Ce2BiqeOJCNUx+0n5mmNqUOODFppb/9gy9cdj/EYzWDzdX7Sq8naa3CHisgvLsTg0zO
rnu+ce3Nef21Rkn0mmvAF4o2al3yj2oS+ldsTBpAFmDo1Jf/4hMUTihn12LaZuHuesMKCu7NpQBj
/nJs1GjZi85Nu8GOi3DJseGiaHV1Broyt3zVCo7GQOCBn+P5jOM6AKyLzfBrGRvWnA1XNQ2THVos
QTUsocjAHDQhs/+LKz201E/isSd0hseAuoM5/UPAMAvo2z74/zHbaJ7QUKFFJntbj8axsknZTK/v
Dt75beq9a9JuSbmVW29kBb8U8TkpKWDU+b0Y3I71gUEAhGf8fk5lqg1VCO0KaOFZkQcchJtBA8XY
HiNYA72lT/KAAb/kgkZpCxs4tjLquYhvrhUoZVlju1cp2YBoTBHJ2UKeQznJo8vpuVdr/O08HKDi
dWJyUvdddMjY2vJ5Rxjl99E3tdIlwLvz09lHRKGW6dcyE6V4JHjo4u4whCRcWuFf8rPnOAN02+7I
NItCsBLcbibNY1MB/E2s+26Tm54GL9dw+4fn3RR4cQUb9FjN6WYii6yCKc6UbGr6j4rgqwhc1wRT
tXPheciyGDiWEF4FOyjWzXDld72cc+y6mdupR/J5HdY0fnEcd4CjcnoiHaBJOC32U97YVqbCMtMK
DIqVkJheUkd3DuUXnY2ARkkqSmrYqKCPv2K0wqUB1NhqWugqaSwWL6GfAI7jjfwcXSx7noVb88y2
ifRZcit6pmVGtfWw+4IwQfFIVXGWEwyP0E2HQyfVXj4Aj8niKKPuj+aZc5H7PNvlol8jpjNpn38b
2mjSyIFMXiyLHftrDKt+1C9xwSuhLTOkagHo8B7rBbU70MsJNaavRHsqPuYTldWYuWjHmxanJvuQ
t6vquoMsSRiJCbcZy/kG1Dwv4V/li8QbhvyQkDKhLUAEZGg/xP/cNhHuAFxwN7I4TgfQMXwy62kG
VWgTPubtFNnVCat40SwueuvWeaaxV+GVxHBBAfn9hzyQTp/9sR4eMCzS+QC8tihYiAEaWajgp3u0
EINL6H9wtGadW3DLI2qN5c74Xt53YpOCIc+ilL5UUp8RJlHbKXfBiTJYwVxxYe6Tk1YDFBpJBWUz
c+Ta5o0M5ksPiUgd05Wm0D15bsRXf1TZ5Ji/SRzpj5YzbxZ6m8d7h92ZuBwiQE07ZIyOQE+5QtQO
oFdH4+nQ6K58VGfTxbwwGoT2zpp45NrPs66WPh/2EoRCom3KgtU6h/YPFjzqThunuso3s078/BSu
UCdZX5epMOf2BbaxCcgSDQiWuNJV1nKPHeHRM+Sk3e3fJ4PMWCMNkcq4yV9ykc5pOY9LwdF5aurm
rnb/TNBqnPZuYrDyb8vBNulXgmgQMl/MTW3nZCRh974tjYK+o4uQ09rLadaFA+pHF6bME1WH6izT
rcLk75AHHf4FvTAdzkcypzj9nyarRZM8EMQ4S0jMKEI/Q7PUxRSk/8Ji+rqB4xMtmUQ6MypJQw+6
1SP5ZSkkL5eMvnOxLFruJ7+f2UW90ovnOgV1akMvNSc17LwCyvG4gxMEL5tRm8oKayJFm/TUfQNo
q9+gcq93UO/ivygZdFw3OGIn/d1TDbJJj3+42FZzq87EHIaj4CxTDcWHl0LgkfbqxE5PKcDBmJLO
GEXbkFPqxMKr63gPvVIJnRzoHDr5SZrlP6pYvl9EcK7a3dSe12xBYOZXfagb7ERJI7OnQFGljsj6
9ljKtBoC2i4PTVYtGCXkxSBI/+ZC2xcO/WLTxpPlOGS0jeeVHhyL5ub9oKhsGR3q/VkykpmwlHMO
agRTjkoQGR6rhferEeF/OzFzicp59x37ueQq1Ppamy86XzdmnbKQxrL7x9fKidts3OBEqliS7GWN
QKJ+KjJNO1Wc9gJE3yI5/5pRQq35hQ1SytlfkI+Hw9DM7Plt8LkW7DeThRI79WHR0+1vFOh0YDlf
vMeZFrkFoffozUTT/AqWcf1bUHMy94wcHJyvBwAGpC/a50WFqxTOCzcjAJqewZW8J+wvch38Hhs2
5kPRLu2AH/08QKB6E7dYVoRSyAji/yLi2QjojiataTvmIHV4NNmuf05gtUNmW3upPu1rvOTTgBvY
lQ2lpLDqC8EnfDIMQLJrdM3hvEMbu9dVV4Fj8bZ3VJG9Sy1Ra8ZFhPJXDuSnEcWQiTnPWAcMGO7N
DgMj28erN7HzanteKzjNXOd9x57rdv7SWMtbCOFtL6WeVaP9BGVhAfZl4/APINvl3k+QPWF2MvB4
yH3iAm5242+PN3n2e2D/zI9Fxl8ZvFBQUrhtjeOcFTfTxReq1YdOp12iMebLkpWi6cHUrwxzE9Yz
ArfW17209lOlFFBlPQ1fA46toXm7XvCW0aoVgi22gUnMMiFfzHatmwbEvCaIeRvHUiFo3UNgkcWA
wocCE0FcEIQb0WRGYjkAKYwlQ3CeII5zZuOeEbzP6utRsK1dhgPzIhXq+g0nw6yuuUqehzMmfU6s
GetxGl9QTx3zfvvVh3giJEZ7zKhqCnheEOW0mY1W3gbpVxdx+zZQcRCKIvbi4IJgiT518RcQzb7f
gcaTAgfwOjaANDMrE56boUX2jvIW/+zmIDvGUj/dA5PO94W4fJPeaUcHd/hz+meiDUTrLtVPhZsV
yNamfHEnmzh/EH7WojzcJlR808tpe3nEGIpWFeOCAEA0PN/JRojLh8TPeUHaldrGfAcf/p/j4bwi
HVcPUBCorDxdGSvBzR9Misok7CIztj6jorxvwHiUTco4zqUtgqHE/Kg6RtFG8mu0PmGE0K1+LJL8
CqKgWyQUQkEP++ScQZN6r1JWoTdzFd0VnUP+6QS9E9s2+CzNGEnjtdDUf6unc5awVdWa4taNqGc9
alMwyVLQfUumgA99INmECaCQzGwPO095PU3aMEk7YtE93qmSha0mYzFKwyrhqwEB9mEBMRtWg92m
0o01Dv2ecVMpYznA4/HZv3nO5Wlqi2C3f75GkaaQ6YBHNajS1KoFdleUo+INrFxHjIKbm6jHlOlG
nUGGqhjouX9DsAjiTMj/LBlpNpnDzVGNs1UYIsvC0K5g751sZHMUACM9ihGMnAlzL9mpeT3ZS0Ih
u1xHiGcgT7cnkkq2zdwpUE1j4p9fEaLqgvIi9PX8g6R/4WI/vjFtIKqHiiBRCTUShnRd4bUUQWWP
sokQs1bOFtHS3kG5fuz+F+G2aStATt05YCK+Eb9BjdlW+cY5AtpRw1m1VsfSn0ygVX3X9EJEtVSs
eu5mWoYBypoJeOqdL5ekk4BwMfMbnE6cMtatyXto3GqN/VjJFsESmZCU9Yif7zkYahscWxVmNcnv
VBcX7VGW0nxg252zIeUmXYpeVyUKUH6pxFEq33GMheXAb0hvgaB32qE5J6EiIxOfeDe1u5JLs8H5
amJxzZjzfHMFpVtjpB5eabcHca5psXlMppMgej932bO7KIO9EXWUY7BNkUusHNsjcVnFN1gUg8np
PBmv/7/Nl8WSeZK2msuGxJwazeyXlukoAGVO2tzBnqGsk9Rewy7uktwsPlH5rANTZoDgiKQHbkkp
vdtmjd3xySqYHDlKnDW3tHjUPH4+agzvC6VNus2ndn9mcrHyHOixloRk1i2imQUz/0dZqRymtBpd
fDWupVX05fRhU6p2lrW0fvEOZC6KO3k0cOQZV3v5lmqTjUXZre3oYwCt8mXyGNvyZAyjl+tkVkqj
c3Nya2eOQ6QGQMRDHYpjOW2T1PtvTZoiUpSVGM9luunIeXsHZCajItGIMvxEkSjVJYpEuT2Ivvc2
pYGiDvcW19TNnQBBLu2etKr/CwkKoCCnIzC41wfGLLshFbR3X4GLMY3QwBkfH+LwsKbmgksrTxRM
ryUT+tALdUXfDnJv60UQd8iwb/tYDMw/p/OY22Hp0bnKhznICwB0Ufr4134DQiGejltBp2VT2sp0
qjixQHcwfyXw6ET2Hcv/9IDbBwJMUDbyMBnKGe4wjBp19pLCfh602gS4UPfwbEMOmL4DArmqI8Sz
QI8dOM+9BIQrJ0K5NGZcfJ3RpeOyXHV8/Dd2lKjuS1H6hHijGhO8Uu290Lj6FTwKYH9yEqxLnOnD
fDwuLKo20fKVZYi0eHDuELJZ2ocny1KAV0pSiBIajfzixAYJPVzJE8LjS3duKvqjJ3DOEVwXZIhd
EtuLzkPE/hxk4rMsBsun4vkJCDjKwxIylmphxjKZhB2H4kmaUDGRKX8BidwP5i4ysTAP/5o0B362
2aAG12DJ5Fne/gMoFiGMVjjkHRoFBFFoHjwXqfbJbNaVpnGSsnSqnlgfLMf12IprZpAZGp7EfXuP
29w6sTEi3DS9lWhKcQdMfAZc08f3MplP0K68YTokeZiqzJMGUh0pHCpaCqL52x5TxtgGurlLWOWY
AlKOSRU7qlqFdBLGuwwJUoLFpxzlg0fEbb+72oiUf81x25e2umAsQ82TrMA4SVLYkYUjXFg8jAMH
n/NuZHnBAlltzacIrjU9z+X3yjxEBpHZ4EuUj+awtVGliBwTx6mKd16//iBnTRwAINSjFo9Vz/Ko
hDn2BfDPT2zyfIEEZZudneLY7epHdGH0G9+6ohyO+aU+oM+By9FACq/gTMbvMviKVKINBu03eU/g
wn1eqmFxJjhGnSNB/vxukT966hh2+EWN6i9veYsf8Bya5UPCmkZHWoOk/qH/kAruLlc2WMOtvdvX
ed1+gRvumYfx+yKZERNNWu0+GlxMF/SdEMUbO6JPVN76V/Wix9vBKm0fVCgzv7DscRUPdhlycBPW
rXQ0pvBc/laBLEkEphEUYOTCfukJcDuy68QcmFQZi3NYTwkh/rEEwgqgMhzHDFt+E23Y2GyWIkjz
MYbL0ukeHN483v0vMHRifo+0HrHkJhU7enDlgD3m/JDUrFhamfplEPjUG7l04seBLkuxEePBir5X
Aqw9DEhDFzdKuZVA3t1i/T//+viaoJc5CdeGtDnbBa3Y67YJnzQO1r/u4hrVpd7jomzk/bhUKvUO
cLiq5UXEhBSpZYEqSNMR3Nx+6MNppJ/ZGedbQFjKHe19bWdnACLVIDNm6D35MTQE+j58RJdQIO6C
dzNcm0c3KunuAjqfLBa9HhxvROjPP6NJqevGKvNKNEk/2Zq58PCkssI+jhtWQQHaLrHZgb4pqFVr
cefWgNA3o8lmo0s30+W6mEooowtrKyTzqva0tnmsVq85+ZQqy/fzL+xSI7areGtWUBI8Jq1Fw6/6
fi0D1Y4wO+ECodIWqkjeP1IVCT3dyHUksBkykkhvZNdgvZyqNNe4cd8xKQw60rcyhGDf5MWGyP8v
l2do2vTV/fbvD8t01me1bn9zTNca278FEywWMnR2lt08mTrtPWL3QgO1b1Mec2rT5jL37gPfuDfE
ye7f3fsstEkE3rx0v1KtOh6kEfD97A/iotLijOwLzpCA3g5H+65BWESB0k0QgnUnupVHi0HxMZ5+
JrG60Ui530XndppmJG38nse+auSXhrIOlhQ5xwo8CZLi41nRcYujUDk4vVZZrxJRFgA4WtBqf++1
zlL0t1qD4ELHtU3yx5UemYuDekVWxjjokrt+4+/+L5lSd3OYah4FcuOLYNpTVLk9O3rUHOpr0l1N
hUj0jRrxwIlkTIFaq1Sm+0IAqALTozc7OFBEkcra+pVVyrCvSLswy1XQ7fq/mCe4Yvuf0CC11h32
hlCx2lI2vWi9IhJlVh1PGIlGfzPiOF+d7omaDRE8xkDUs6nGsRzqvSDNH4apDmTSl6Vs0n6lULkc
VT8rFYKzJ/q3+ZzPi5g0QW+cviHiEow1Hf1Cuxl88wDpMeC8pKKIn1WvjnsPceDjZyWt1KQOK1Fb
MdClfNoicj1WEBXPsv8A9etBnqD2yOiX3BK+ZO1QZSOdpujT8nLZnQwns2dyvyXFflDHM6AYCGcx
5l5pCzJdFtISeGLV7VFuP8leVpG19Q1oAakcxfbNWghS0h+1oBBU2ESF+nn3VWYwBZiDK1Q7Kmfl
DxSP/wLz6jjealAAskMc14QAPw9iXV6X5Gsslo6HdXJbUtUszDrph3NKKNHYGeO7HqUSZKn4Lx3e
uZ92dHxdhxnZZikk7Ekmk98xxw2OU0G7ngbUTpebKPOMpiZJdbsq/KP+vPo497oKdwdFVvQviWPU
8LoDtWPVv++liQPYcKj82/B6izuC0wW48kKnUocN6CCXJa0BSyc1p5OJvwi02c/TVyHglwkeddMK
ql/zw1JcbSzlv419QikZSg0wyWdM+HWWPDqOVxoKIzjhYP+pvxSgzK2/ppsiN/90rr5v4MS6r1ci
8Gt+03dt+AtZ/QkkhC4n2moMMPnCzpfUIvHJ5CxT7kWu5bIMSO1n8JuW3+aHcPvKebFdkeHdChR4
Yun5h9b+P3olO3HPV4KfTmOUZkY4wAOtYs74bMd/NNbma8wrIFoay2ObvYmBJGav/Lcq9mmVQblb
xpcGzDE/TDluqbyajKIQRSD98yS+UHvpC6wPTxre+ixlbKbgVP/5nyKlbdyBaIVVpJE4AwoJZQiw
4Zc3z5NEoHuH5GpbQZfZSPUu7JT7mc4ArWGe4c+RFQPiuE/rRw6xItCXu1o8F1qsp243aO2ln0sA
OVXL5CgoccLcNaRIx0GNIZ0s4GJO52iuWGvwhze83WxCqLuCZGOUBj1Z3C8HgNvGsGJKhKcc8Lj6
twfAEColyan9TORYKjVfhD9QyUwqWrybqeZ3/poLW8j8uCtSxcTXf84Eic3xaiYkc2tlI3TKojBi
g3S9GhP/jMf1x9rkDPr4/QRKAwBiiorbU0zQl3zIDdS2RC1W3I6rgXuu9YoFiItH6kzlGRe1pRLf
AWPGNFUJ9E3ypwlfNzumCRSwx52ON3cOcKviQuHGF/4i0wjU5cteSaEm8l4L/LT6IMQSkvFH7P6q
XHLXxq1lbOcCQ73ureEQ7z/hLFyqKEEnNs/dkCRQW+lNKcvaa2zD9ajbs7vbDa23r5bwBaXP28Kp
qetTbVUiUXZcvyqshUm4KRMjGvobD6hq4N6WRT5Cv/46SCnw/lx8G5en7Wi4tDaFqemrOpzKhdJp
GVIQ8+sqbY/gfWXaSOmcRG+8smm+CCIX5Y19mSziMjtolmtzI1bVgtpa2TmKnSxsiJRy2v/gRluY
QIO/Tai7Ck4jdjCFlEqZX8K+V/nK627r6QFkJ2+PDBbmY/VQu3SgNbpvBTOxzhnap6wHWfJqNo2R
EL9nG3szuIh2kH68EZQ6J9jgKasuDNgWJP8GxaO+BVa42Vl0UF5GDeiqlWx1gR9KTdiec80seO77
DXyaRKpllmd0SvJkfYml2izR5u5jSSy0wH1KtPgHsi1SDFGNdZy9igZj/P2IQsGsEu4O9moXRr7p
fOKmUkC3epjIYDvRcQFhLwurcGwuUTs/5/MvhYh8P4sSRC4bwV7J88Omaq1eR2wSQyQGK56KNC6p
z7/h/pVrxoi2SfKeOP397eajcvFfP/9q1sgkxtG9gjtl48T7o0eiOdSWwLt/bmSUDWB70x6j0UqW
f/ce6PqONCpaDxrADi61kow5SdQtrgzKdpXBOK7v25Btc+TjQFZcaNY3NgTyb4t3THwrDL0ksGfb
zJPSLPHkOF0hJTt2t3tGGggSfZqds50/9/5ZRvye9NxPz1I39Mg0IRS5wldh2Og1l8Z6qwpTTPQc
oWCsYa6sMvh1Zj5on8HvcOgtO5Qrc222gCInDzLDkV8D/uQXgZV1ThCD6G9dKEH4vGDxGCR8ZJA9
Gow9ReK0H/LjnGBt76IRstjU9rVrr5NVbLopB/15bO53aPyd7IEtafhXIoT6QaJmLfccDxs/AfDt
/whmhm6gz9GIUZG/ORCwrDwtFedMjVPGaKNR6aR90rq7RSQpabjmxgNDD05mmnZzWQc3gLBlDOlk
0sjR092zRKS42C8BqYW4KFr5P63A2tS9WJJ8VohN8ekmy/XS6RnukgiWaceB5W4Q5FN9iUZ9srrn
RtCPDayV8m2iuZ2K8Jw/3fRx3MyDp+DTjE/opu5PLD7Nj7fZjXpxrITAtKYeQ487N6zWywhWN1Cn
2ZlUGSxwW+Gjs02llgZ5Exo3hSLocLC/Lsl5GqA4a1uEu58n3BZso0+46CkTNM9ahxWJaCoD2yFf
Wh4bZ6t6h9N7LnIy1YlHtoPIGRh8A5MDKl4Q2uXt85U1hhbAXb+gEY8vSU1p/R87BIlVyixGzUc+
cJ+46TSC19Zb3VnEXG3krqaP4Mt0NOBj90Pwx3eUinzLnbj42oYp8BDe1FVGMrlWxi4Aj9OUIerQ
WHihB9cRsVSV1YU+hVJ3Yfz/kMoULJ947mE/HZskB6mo3SkOD9vS08RUXRoBMa9MbFuFc7WohI/3
Adn6cfGecDKiwFNHPKB2KfYFheCjd8yHd88b0Q5MVaMHj7dp1daapmtN4SjMrlZJLHACYXJYH4Ji
p0X8f7ZhC7wa9U/A5aGk9AUrUEwMMXCcnCBXEEuIDT+XQdUXFb8pPWJNLU8U1HsGCa7mzueda+IF
eijU/8w4yyP7hH/HZ+DYITCh/1Y62Fb3Ciqmf7waHH6owbOlKy+b1FY4GK9FQTQ2SqeFKknJyB2+
lRG+SdZN1cx9knlNNG/yLCzABr1TFsWE32MhanuHZ3NYXFjqfaR7DtH9Hu2K8DVoPKyTZIcfOH0T
IQNpGZJS5uk1alfwTkACrUSlWsG8elzYnzlAhzXWSKKwGmSGzoUgO8/qRfRKaUG3Gfomdc0+7H4D
3M5xhomsTLnAfdtpQ+JPCn7taWACjy6BBTGL6RQWZ1nqkH6ZQ+1kVb5XmjJQKjGsOBiTFoV+8OVZ
f7ZcsenlZsCka8QGx77VLM0rDJxtuY9YSgfXs1LPgd/F0IMXKx2bdFuTld8elc9w78WcXpA3c89o
PB2V/qO2N6f+bpb4yY464OoGhszlhZlzzmhndtaasWHjawH1f6ZydnAOZzx90NsPNQxsYXnNtJch
2J+KUVW6A6FixAI1ywtT+IsF6wNMUx+KUb63uSYzZ80Cdj/H2v+mHGCvtP+l9TNM3zD7w6PIGKis
NBh07H2m2uGjG0s1/EEaICbkzFS8RqPAP3OsbUakwJwOKQPADA8a+YKY8IFBQRzINZAGPC6S+3lZ
/mD83+o3MChTw9SyB0n4SsOjJdAlpzpRgybyUe7vHEastrXqZMD/TfKFSU6n5QsB0f+2688i4yPB
lyeQ5KB2SFHHPYvGnoal/RVgw+6TW4cQNvNwemWlNhLyLYcObs+liAh7ie3NX6sBR7EsjmoV2YEy
uchDerTIoXY3I/nQMri74lWnUEJVKYHA+zUQqE33htOfTakaWlbUnAyVHYrFIswp5FSZkUGDBgu+
ydMVGofxjZueu/QcF50ZavbzD6PZ4UxjQ5DGrwrFKCbMZNEBoJpKPyiJtt9xwwzN3mFSXXs4SVQQ
rABQcukah+fpYqG0ych7iXDvVODBoPTjSXIDBly+eCa4pbjYfhvv/Lw4Rj3UEttERUuBfuju+h5N
PriYPSaYvQQVz/tvmxENjpEkNnXL68QcDOLU+2XfQyXNfrshIwuIoNbVsxWZdBRn8LhvZLW4MrW6
QhfKLuM3g+wri3h6+689lZ4GT/8KqjErbhYFBq6mYdioFfYSYsTM+EVbb0TDSx0gqmUlfcDIIoVb
Ri7oztENQFE3gwLULHWmaLOJJSb2I1Wu0HSil1CKR7u0iopPd+zTnhwSFT2Oajwqh9AQiGphIiLN
7ekY8/I/L9EgofWGr2PLypIXEAcUJsi+qbI1bTBGRjXeCF1MAdkFj/CIBB3oHgrbCx2ypnbaHLvA
WII9IiggTOJdZc6zxyFoRddolx0wEIREdz017L6zOnUgE5ZBAHRFcRVPociTr8pioG4+07/PNoHj
Q0Aaxsr3KNMb7ooTT+vR9G5JVYgY6wn+kw5/t4uJWxTaSZPzJHVjrgj0t1AVfjiqUXHVw6JObzcP
JTa8Ky7l5VX9YXZQcXfrLEQEazPuRUttM4sdrn2zFvfjwMmhV7I3RU33vRmHcuzkwi9kLopc2CZQ
hWTD+QgJ+2F1t82cFVQvNxJ3AIpBsWIfqPezZca+jLPiSIQC6OuCNxkBOKjKq2GL1zTwhEgUR4tL
BlfzJKisLxBn5gFLs5OChsTf8GbkeviGbq8BuVMd9R442EEwXeEoZslvu03Mzf7oKE8CQ+Txvj+R
zYhA1lx6uXrrhe+gsug7xpVu6+vzvDn+kJzYWFLEsWGsqiT6YDga6+iwQBoZT5dUmEHkIlN//u4n
2y9YuapNhvRsLEHmL7ryDBomvI/ij4BGUOnm1i0DPl+wyfx4GJlvwxsW0lvd4jyfx8WbJK7yNUJ4
XdHhlOyP4ZIOW2tXKa5iet88HwCErwJSDIxLv64G1TJNHnzsXZstgo84uRN1zJthR182WouiZhR/
Nn0P7juvL8Zz4qY8Tw4vKNSs36CopDGFkd2b/LBRXFsbe5ewjScTC37+z0SLCIxJH7kSc9UV6XcR
HZVxMaKy6T5grtMfGlHM3FdWbknlVS+6lOQpRvfgrSvVmRp/PonFTqxDgpSDhmYuqXLprpLcocKe
xc9SKea1b9t+J/Humtrin7YmL6hmTwtHFDWtBsNoo2z2TzocWnp81zFWUf1OFov4Xh7pnj8i/3P1
7pOsPvdHo5LsmjSQL0Qy/iJtdrP+6PZuDI2QTG35s8NauHihs2ukc5CHBb5/Q3CqZ//1e7COjvoA
FnNQGm3UhYHKAg8nMnoU8hgaqXwtxqHLSuc5LjqghwDwOGgixItVeVdFYaJkIsU81nR9owL4OMiX
UdUBQmjNjFrI2sYzkhLvfGCinlmg4gtkckFon/hC0R3a5qfvqAOJhw66JrZcekYty9l6yruHEw6h
YXGm3oe3e/fR8BfMftVOuX8So9MVYmJu4WPXFsBoqtnOQ4muTcgywcr0yJbsHn/B0t4aBTeiFzOJ
h7JpQyPnUs3yOEtuWYZuZCQRAbMLFhCQdEc3O7p971RQbQlr5mohL/ZjlUQwYNNdVXEnyyPSzVDP
aFj5bZrKMduqBufdeZyUo93KZ1AWqmhf24n2swgO6YgJfgsRD5iAHTHyhRC91iXwn7Xu6oLTgrS/
a4WIflyUdB/w+C8/r3XHiqBAkHODvXzLNo/WHJkN6G38D7y65A+TAUpzOs21I7bT+N8S3lnLWxHq
lltAKmr1AcPu26XEvJs/xQFUu0lNW2dAvtuVlzPeqq/oK/d/KvOujOtIqP1WqvLts6TpX9GW7aBH
cdMHKzRHv7KgyOuAc0uPllWfqdlXYprYTw4tce1Tqc/b2svPKUB/XAxAZL7UMeA51g5TdmKNDUjz
MHakst7tBhak730z3sk1MK3U8TCQhTmISvIi1VcpBW2yXUcPxuhJFpYxo0A+Kgm0P9kd3bhxDeVJ
nqeJwp6oRNyfH+vJHAwwktF7rZ9l95bxWAW0lZDT7VpYZmxEblrOQeQpZaAnZwqNzmUO90zhoff+
clKZj84nqNLmpCyA5hmo2Itl3YPz5sDcM97zYFIB4XUZw1O69e1xh4g35pzkTdaboHFXGVACk2Bk
c3yE1LJTM+c4ccIeveKAfCLUOvX7hwzk7IVZz0BurFjsKQ87PJYSPYiY1XntbxmKiiBPnVc2iA7+
5WTzKtznCjz4o/F2UVTcIp2Pa+CxvwcfYtL1Cdb23Wvq0EbhSA6berHwjFugbKJd2NCw3H3i+UPr
CFRsrcjJV7BLN8qEz327YQ+1xZuy9ls/CNmlCVpKu/DK9I9OWN2+EzvgEDaNSFIzh42wEL4gvxGZ
pb6MOS2MbK8bOXNeL0zXBAUY71952inAl/0x5XaQ1nudhVHw8B/JzOQbs+R82dqJRB7XobovrCNr
WfThOhkNnwGlcxcxXkdJQgmCF3P67PU/7WCwEpy2aHITpI9vD/mtJEtAfkIK9eNDoB7u3E+DEsWa
lxrUf9KkaknFJWdmkEgIKBVLOuQXuxHjpeHHzipVjAivuOmfUDGZSwLQF1Rh3WJGxMZE2+8BD8ek
0b7MQo84WLlmu98a1aFuL0HYLikAd+25Bz86WHGa846ZKtt/LhqgstAiwHn+6N1MNFmhr07c4pVP
PdCoy+yUiCzYtMEyi39Me8C0QlbqCwPLzITJZi6gm38Uz0s3x1doWtuQQc4fJ2Okb/TTJov1gWSe
tj0Sf3DO0vOqJRyDL1XTZP2nhBWvOV5LLER8TXBDk67baeDFTKhXMwYUOHL1DW7hp0QCxG4I7qTp
ByMmefu2LkLS3/EOvSuKacZMunnJxzB/hgy6r/A0SfYUAuETtEshQ7L5J45431Jf4XWalw/BV+8e
wx6lz+pL7WlRQze8BVuyPkyeI5l1KsWnkeIl7IPuXFyk8u67ZwqyMk1CZ+7zlbMsRpXkSyXNDCrb
7sMbHnqKXph10hxDFdeQLz6mk3hzW+zoF0UfDHHs9uA6NupeO+Q9CBrp07kL9v/sMhy/40lkVnW6
XV0sIlgRYd93qYbuH4uRmSBAyXCkqc1UW3OtZd0iqQWwqzlYy+aMaRbwl/R3q3IHxe4IpTOW/t47
YDhii4bLCMpIXWQtCj5gV+lhOidxt0ihMu43UFNAP+9JZZFaE8kUKGyZjy3HNtfCUc7Tdo/rXimJ
BoKmAwEL6Xc8ZWr4UUFieGwKtot2hznIojTwiG4qZEWv0uAyd9hSTNt3OFqWmNrE/Gwvtuxmlr9l
FhxRcTimty8O3H2sLQTm+UBr5UbRyc8tx7Grvf6XdDggzhwvaRfEgiA97jlk3gnfXqlTQ+AmzjTL
mFefckVsBnlPsKgvkxo5yw75ekRWpcTmwXeJf04BJh0+H8MAWArdm1yCgIh8MsaJRBAjr0+lJPFM
Kkp2ljPw7EtTaOn8LGa5tosRUTD7WDoJh7D5KWpBh/I6XihKHdiTtiOone68p6byq5vblgIY4QH7
oFwdO7GytyslBmaGLraiX4ouFwCrR6QSIUL7UfvS6lgG8iHAaTTkXOLZ1HdfVpUNZIwxW+scSs4x
E3ocLLE26lZqXtOEsnHyObkYMsuzm2mrz2+W4iAcmksljBE/PuANh9j1ZLYN/wVmY5jTdo3FatD1
b63G+akg3TcVUon939hO2KDxeVyw6VvP+mQH87mHN6zCNWmqRFHa7ESJ6fB1v586noL0qYkkH+Z/
Poozk76xBmeglwQ1zAygl+8BSvmUfaFsOMpwlITqdlnkDjoGgHWls2waMc9GisdyNHmzscWjybGr
ct3uEB34uHV1jpTduS1LQIA083EKvHIcAHPiIcBZ46HFG6OSuy0xZGGfa73Sw8+j+Y90SdPIrFYu
xfr7wHWP9B/NcJB0IcQuTMdKgp/bJjdY6Ka+foPmukPmFfhk4+BX10jNDLmsc3mlKHtf5s8lonkH
8OhYw+WQiCi4XjC9sV4eJJo6qQzmbaHrjeNYY5quAEseT9dhNEEDBo5qTenjvqh3FXzaFpjWiJhx
ajnd/4udbOM8Q2AAyEh2eSZstZJkKLWfyDjIw4JggLawNp+ewkyOTITivHAnazq9BofzxBjCnfEz
KNwPrLx+x+eE4qCpynbzxqsDOC0ovbWD0ON5Mai7wB7rTxr9vgwA3SyPcfRSCU8U3DyQtsnB1WI2
4KM7fqeSeL7i7t9oV5rqSEz4C4sgVGSVEfUKMMS2J5NdQvLf7XFxkkUqgixzpbwtcrKSyIIor1uz
aWURLQ6kk+336vnUuMFVa0MC4OYRIavxsZUYsFJoXHuyAyMkILVKfbp0BRE1yLoRvz2+eTJ5lmQV
Vp3e9BAIri/34GOH9yODuK8DgBHO5LSgw1PCH7SxlxgvICfGSXXk3Zntqe93hY910WLOkZz984Wz
7LR6ZWvw/2EVvr3br03oQ64oOpKIh/znhCBjv5/4IVWiCzPrA3idXQ6Lh88tHWb4NtHXX5ZdjoTH
N3aCcDEdquRxUUXm89LjfXgVo5T8BJzavtXuIHOqKP7SI6x2oP+NYo4DSnFo8tgouJ9cIY6G1hps
i1D9raMo3y3QYYu7YolkfM3bwCRi6EwSA7u41tWI8fJp0qsOpwE9lxFZeUZSNbfuwIu3C95oPU1A
P8SBgrBgCCqF0YLIC88f9MwS6wMg5jE6+t/WebUTHYqOe5Xa4daO84UZO/fYcmweVMnlG11nxzXQ
bWK/GbohgYpEpU5VKBNijfihaLh8yNWC8E3M5gmV/3Bvh4woqtk+Nfxo4V09dpEGg0LiASJaynYh
XLwHRfzbT04i2P+pwxmih3ybOaO94iFo54kL4g+k1FienvgCTT22D1SQqlTlXYgCpQasEUrLpOpb
p3+KxRRcp2E6BB5VhJ2a7MULj0iRyK8naCm0EOUYoyaOxWkZPQcJBOGRnjVT6d1yL1gai8EmBflp
dsWvdjMSYag5JSXpdwNnXRs4m4IxuHjz1tc32Ds5FZO7rr3EJPgVAqKVMBtS3LBnfoaYliVJkexs
Bqc9KRYDqvyr7pC4i/KaXAKteKM9qjBZLP40QZwac+3LvFdU0cgekFVY8N73LuuANWaGVNAnoCZP
ZygiKsehZFB9fsJNToRNoD2c1txBKOwN1g369oF5ocxCTJCrPEpwUZ6WOjWsasRKohN5B4Vg7Ob4
zlJBUPg75zZsTvac/rMxsBOsUumhWhap3VUX5LDf+iNwnTSVziehZmSJiGtLqluEF1ks8QKYOCqB
10WAkprnrNg6gIhBwNCbGJfF0nDvrNFvguHk+kQFC0XLgeQyqaoDJ3+lRoqb0FLOB3ZKVNifgXQs
MP82abfaDgVQiLhkZqazKuSuqJAV/iPKrQ28VsaNjE3SlfQr79A1JkZZZLezam19NfT6c/WQFoQI
Ugpz8HBMGLb/qySUAsG5nHdNrXrwjDOnFjA36C+gUKEZrUykrD1pyHWbzK4yEdQ6fvqYO+0XAKdw
h5zhSDn5PxZTY+BTGy/PrSbNcXYIXY4san7bCYEiQ78pz93aAiHPQqtwGT/1hLhk6+lsGLY9+7Wu
rHPnmgGdlEghMcy6ai7F9bRfk1yFurDWaI3gCu5hPSNqfloOOoIbH1R5fFvMBbq8e8WAMi5pvnGr
KN1iKcqnKgDsBAWVYLvXQUFZbD+NODy53JTfrYsZ1/FwaKzWUaIuqMv2RyZeif97orSS4MY3Sbbp
y6lPx9tlCGyB7uHjqW1NaYdabCZbv3nwc+jUnBct00DiMyg0/CK1Khi+jgcb3cFVYI9FwjrmcEOC
+HpG/uMaGf+sIdSwDHsYAA9R3emM13uEAG2UIhZpzMACKece7bnMT+negg4HXnpIg+XK/XreMOzg
wenRMUsYkHIfSZSzVh7WtpkyARUr+goAGa8LlckBQBLt99Gv+gdE+A3cpWplHTnBXTs1wgOEmOTV
f7W98N0I7NoPE4BOfiRxJZJCRAbUS5th86kN10jFSoKOrkKwT3CshFSWRIKHNKf99zWpHm7qZkXu
bFFTHG8iuJ5dsaps5xdQL3lnIx0HoDgKptR2uOFoHSnOSwRsMog+3xQL0oQS/4N+c/M07jVXjfZ8
SsHlq+axSsZ63WuO5XOLFmJlj6mZLt23qG7ANS3CZkR3nsiWh8n2jOGBTr29uUWoqTTZ+/yYFQYL
cwYbMjZCql+Sa0ssi39UVOvrqKxK3sk94nLhHD+wmHXOCuSdWP4tuQrjZEzrRHtIi4mAdt1DFU6X
eaW039lX/wjrzHmimqPuQErtBqBj/wW0kcx4NKXdFGhAlLrXIIOGWwJXUZ3U23O96GoiGNIPNbl1
ZwbXoodCCOjP9wtWa9X79gcWPvXxYy01z0zmOk5vhNZcoZ7ZYb/96cejRSw45Ufj+E+v2GcViyMY
I594H9eaty6uIG4UyTIxGe8WpKZganfpoZZK3HXCfikjAX44rEPpVvnqrQTmZ57oP0/NGBbKNbcW
Rj2vMZHOUcSN1eWOwHTwMURVJvF2sOwxXHa40WE6NvkHSifNMAPvFZOqMfuhGELDoDPvCeuENhtH
9VEv4qEqXUYy8i4QG4HqfPIdmLVK6dP0JsxsUU+yw7T/4O5J0TaX1TRG6DhTePUIGc57LmaNNvdU
v69hDgVC0LB5NttnKQYaprbr26hnxLw1ZZ5kVWkK2EFT4dfghdD5F3kD6GsO0ilEUwnW8CzfFhlx
UNHC8qjQoSvC5XglJn29OMgHC3xAB33/o/M2M75omaWOfp506XdfqzwGgS1Ytb1FAl98ripgWhvo
J8Uc0ZMrSB2En6X46Ly2+ZKQsbaRbxmlyqzCv007RWNj4FNuw9MoocF59OX4IJfif8BFo1vHVXLd
VkjZbv9ePhdXQiE+aXiiZT7JzPtmDQOvSi2ARCZvXw7uMhflgpfj49mnTGVbfrpnJazvdwP9kWno
dcTjGgEqudyx4V9nxmzU7wVavhvwZhBN51VpWjwrrIvS3ysE6dcWp8eoEhFRuMfBg6vfzKPwJWdU
wbgspVqIB6y+0P0ml+HwaSPtgbEu7BfIk15HRxU5J/hlHkFeQfxQznEkoN6l53dfumhdhlPOdgEm
DCWExKGmKmuKL/tRW15m4uhE4pt8UOWyHP9JPyQs/hfXE3sfCm6UNPBT/zftcslhgyKpzMXIFyU1
+jHT0mawKPePmb+H7qzXYWKTNPRkUQVocS+XuLsbUjMYwEs/Oy2VmreyqPfy8FNXe88HUw7mQBbg
ZYGyQNNwUvLsiFWqHG0+DOkgbdOSQksmOKER3JY1Tm+rI+oZltUfIIl/dkPAObCdQw2Qqo10gC7I
e9AeTFuCb21Ptj4nagO8tFjgx5ZyhPoYGVbdExI/N5QorDLBol/BLMSMNtdYuGbgqkuaJc/uT0Jf
8LgEzs2GI5E7jpVAaoxuAmLen9gGD2YlDFnnvhbyInswrA4JIYpnIoWtRKohub+q+niRHQSZWP/0
NNcP42jcyueEy9R52OhNtan40Y7PeqvVLAQZ0vECBFTdldfoPqKZXFkCyoa7PfiWt3EtlMTT/wit
WbxCUwbJ/j0F2wgAITAmot2eF9rF+ZmkwIAGpJKhOTSayWB0xxnjLzODTHw9uRA4g4oZvD6rr+pf
UsSxPR/ecNVzGMeT//pD1iBCFKasuTPIBbHQh4O2CHK8+Phpi51X/Ao7jLX0EUnWCcXzHtSoCXks
sJMvZNTp9UtnaBNzbZhQBXmhBySJ5DBJJzoh7p3S8HdwIkMe9HFknSU19D5wJV1GwDas5B0vzis6
UjfmedueWiMs7oiwI9sd237h8pM2OkCcrkCqsOYSAJuA+qKnMlozSraAn/1OT20pYuTh94Ptmx5T
gfJq7qC6QSeBNcf1iLCKZvSO6fHzARDCmXDlNELdj0JcgssjDfxHLIQxJUPGB/1ixeUMeBeMQyDK
Rq+a7hPl9aRoyHbkDOf7lsyXL/mJeCH3fP2ujKqrWobPnJujcxPAhRNOb+/n2CTUestevQlucJ8+
eshBffUqOXGDIV8foWLb0kQJAPPu3q2DruklIjfUGeq/AirvWtt/qU3pgxCDHTk00h03HnMKUVzC
CzG0PAxrdpeszNslT/qdb5bDVsmoJgK8D1clcgtkFlYBoC5hhsdRV2P2QMx8ziyQ58i5AGYXEg6D
CqARUFEBRYtVo+wHaiR+WHVKEK/HJEeaOLJcXyUH2QJTKG5Dv4umwqbbdYMYdko/RLDsJNGFcQgR
ACbUuJtYjkg3TNmWDq2YRp2H94fyASQh+BhxdoqzSDFdwt3lGY3UoG0vC7Cn4qpPkEDOqsMzcbHR
+lj3S1sFH4FgodLpt9BQFJv11thRjP9p/3odmJPJiuI82RTIz4xHBymKGyUVAhwBBezMS2zCQYa7
QcrQA/WzTZ/1HXRpyugbpdo2FTtRHfCdw8Vfl2/CHLrg0X6fgnTCmYvFt292PTJuc+KQUmmyXMAE
XLXz0gEDQe95FhzUVnT8asDZczPU6P/X0hqW/8xiyN72UQUKwPPGfbKefK2PJF0zBeqEdfdtbWpz
ANsvtP+kfgSPTvVPQip5XoUjUALZehSwd7oP1PW5oVHcCpBgaJUVRQsaB9sI/zUbIXASiMFlB769
efYHirRdyNfNtpCNl0zca35Pker9o825OwCzUiBum/zHIEbIeolOikSfib+Vz3zad0DNvOU4cBU+
MRrwgUALNB4fNY3oFGRbJtOGEiEgIY+5XD9uniV/qf9UDrz/Fj+1PE8OkU6fj46kNTheItNFvdk5
oWP+cxeGItgrwv2DN5/7oqV91g8CncxPM7HGHvH2AcWFXQlHouZbTPKLgjJZJs2n9ogxOU1mnWOf
w8iPiKTgVqVHJNNTC/jCr4bXKLFRucWiWNHNN/19rDklCZwUeOTckBRvEJqjYmhEnWNey9vJgAJ5
a/XRFJyBShqRMujjuxY3HrpM/l/stU19ozdxy1/p0n9tv8iSXYJoQBCdxeNWW0FEIQlux8w9VDda
fGmsknuo7+F2lywV1/aecxAn9OdtR5pBXJOPUTRnKhRDHp5AYmLBVVIrMHfYJy3dlcwqeh9L5fdz
RnH9ls4snuAVlN4jKiC9LOwm2PGgiJg3zTvR7ZHv3cvkTgHX0+Zrbb7mYEnzJa/kSv04W3Pqi7c9
ukth9Z5r0icQubNbkU1G5qiRlKCHc/X7BEedSL7kyO+Wfc/PY4ZChvpG5i7ET6yfdbV7c1IARZK8
7QDG39SKwujvyl8DgWi86npjUgq+O4zPBhroR2g3imo2GHGdy6WEoKJ92iyMS54UmPpMRk8T9Q+O
9U3p+w0fW1kqxDNOmks7nk8AfybYoFwAcymnmbZ7AbGeUvxTnKCPgZ65g+jtC5a0967JryRJrZFy
xjovknEChk2jpS5CQhb3jM4bcM140lvBKRkbDzsEjBiqd6HYswmPAcwmUvG5y3q2ezDPqYuU4kJf
7J0wzKQMH+TlBMlnwEWNqtjPOsR8xrKTrT/MprvBYIXrgE38sUGpUW50XHZD7/Wdx94MVW0yTp27
DlYZKq8Nx/Ii6UxwWuG6JI/yTythhZTerJLIMX1VSScRhvpVHun5bagNxybEbJMoRvf29S6Ug9fV
ZNlCy3dtBkojeUoHhzkXo4646QsWzioKKbAgXIp8GZDG5h9C/qocxS7zSdHj6Quj/+cWY3QIs+iS
egqNWQfY7KELN8zom+kBZm0KVNXfXRu0DTEuifP6x8r2y6iXqRLv47wfbxorWDByBXAEEC26xyBS
cPXVdtdWgnHdBcKvVUAUxZZO9GfWTm8vT0TLGzgDxdDtONjoHunCJXgDTT+cKnBhIutLJQrDNu3r
xpCic2n0ZYYtcR5eK6mDNtn/XmQ1P6Az+R8pykuudwd6k1P+jlv7UBHzySHJjZptYmXxMbtSaoKt
sZdTlH30JSKleV/s57a4qTMCdfaYA0/gbrHnjEt95l7nyGlzayl5SFhMfAvSR4WLech9P4B84r3H
vH5PFrI+ZK8M/1sW6Jj53fw4CGD2Br8SioAnCM52FGnJjho4mPMdJ3OPuLTKezOZwoEQLATZaXWN
17jC+1kDq/SZIsezAIbXzwjvqN9+lIkSNux7XWm/wIwsjrtiTD5RIzF4nPFFgyuATJyO0kwwvvcH
Qo+lAMrmkNo/VRGynqYPgVk7rwjXBEtofk4DwoYVTWYHhJTqc4WEqw7D+b45dHE7cdJH00Suek6w
9Sc2cWhwz2mB+hOldg7NoBp68K1IpIWRO81Kv61GmXv7qkHgWyjdxiuH6yzRqe34b1awiZ6s/KhH
irksJqXKOcZjTp1k0jGEL3N1II8rAie2OXR7uqwMwcpGgiwYkkhDcTKXY+APiFAL+ARGSBnqwtIC
uEdn83tzV6h6R2WzVXLuw61aetgAbqaW1FHwJi58OKSkNwGd7SHtj9seLB1MTinxiC4VrstaCIDd
NjuVUynMH4g/FJdwEIAqgmljH38+9GjqQ8WKBk/o2G4SrQOMFzzQtJ9tzCTsHWoVpLaJYLpUFpjo
Q+OpnKZYfpNHeu4BQUK2wIvuzOmOYwudP4eePVa8zdFxzBexXNh/NpppKTHU9V6YqK6RKttciohM
v36nRvagl+XbbBXBw6TFnWYGKZFHFLgww9o0nYwWs5cOcfwYdXblsNDru8VUuMgD3YB9eOx1u05r
03Pww7JWjzhmkwErO/wAqYXs5NZ+tH42KIW/bZjDbt2Aq4jpOUZY4zZrDluqFX1i6qsuxbURwgKc
lo8Opmk4byX16EP0xYnEhZjWYs6Ny84na6aHldXbvpin/mlB4oB6eGGv3DvXWhEuMPowVRlrZPNg
s1NiYVvcKqmsNMpeh4vEDsrf/pRGwJFpdvsUtVM8FAsHEuPVgp70Nbe1fqJxq91E56D1NcnaGclS
7YKIxxXkPrRPK4E6j1LpTRT/38jYaj3+WyfsswhulkMUXbBa5s/LagKo2VltCHwnLGSLRwtjjgWp
SqlopRhJl9Z1CWfXsJaujR6J3FjwJbRgIf3Q/Bsm/ATNVbmxCPnRT4nDyf+QWPycx5HPVTzWaich
Ft12VhvH5E8nbRShdmkWymqUd/8J/W4AhHQFTFIF0WwuFd9/tPDsAYgaCjmNQ418+nYWiU4oX2Hq
qSKol01/biE2TwyfEAC+thBp+x8o7GF6rQdtt+ZMHEHvxg6n+JJDMvz0MzP/pIzZvPA8B7f5IJXQ
i6yq/KJja3JoUqZkYML62rKdi0MDcQjiT3tLME6Z9p+DUwmlWHoqfop62OjMLeAtg1lxArcrfScY
HGiTm9kWH81sPEUFxQfLd5YO/eIqpHRpOpEn9QYJtRYF+aTdaPVkba3n+ORp6McOjRMT63mZIgyg
TdGwNM4ME361lX0hRoy5M6kO33fEvNFErglfcBPn+sOp7j7vhDX/Ra8VXSEpIXPgvbOZmPiyMkV3
+SvC6dflrdm1YKLbkY96nXX5E0+/TOhLsVHTcNtwJV0TCwQsnOXelahEJNp5vo407VLLMDq/cbHA
Jilv91tChQdsheZT4MhT2kxqc94aWCfskKyZJxTj9cLIj7B34tYDB2UEdlbbiJTvfrSq74ke1wPn
L7yl1YCyR4PIa7DN8DD1B3kb5s6aGf6IEE4rl87prnRJEEc/RHdaGuRG2InADqOEuKPdnylwi2FL
u0JICWNuXVxDdDVgSRQxPXnhBthioifAUoASjg4HoT4TJDCpcVTMplfsyhI/IjALYDs43E0A2M9t
x96txKfZThMMm1SDxRWw9LDsWCQHOdTOpUCp7Jocx1c1Ui5P/S3fmh0/dwI48+sLEQtVDCyyUppL
dBEIhCJkfTOtg2KZoXc+ySZEVwqc65ZDGqA55bSvfaj5pKVU/1ZNk/VF+xETBzv8b/za5Kx120zU
NX293ayIcrLtgOmzRiPhrRVvB2zjg7n8Du5GEIHmd5+uQjDvo7lVLtA9wzaG/v+58YKkvNPoJ7ME
sy9gtSrnlgB2bagGCKd0rszletu9STtY6E07K6v+U+j0DDbQ7xAR0L51X8WdLeMF9PxpKjY/RIm2
3TCGa6r1Ci+cWVy+gGCm5WSLy4jdPaaEZnME27zuUp3ME3T2xakQpAEMcGUWcuRKn73ga4maphOF
1alC6Rbd1cCmT2nukjAas70DBefd8MYPuS+cysMQQNSL7MI+KyRW0wWHniqs8rsRh5Tibo/LyCYp
gYFKXPLEt37MSJusct1bepkhskkPaf9FTeOuqq7WqqjqXmncRm4dNX64mvgM6OOjDvnrYoqAadw0
ITYPZ15y70wD9PilJa0LZyj5helMCOh0ITUoEwMVuf4+2I4iQhBHSQjJjKSRnj9JmvE4sV9nHm3f
JvD1ZAMLM53lfjCVnKtfL7d6dSYVLaxYaOsXgpsJHJMWVKJyrNA65A6zDunkgLrUDbiINQaZGIq4
XpnhDJZnBt/T8pnKbwC2bHKUbYlTCzqtHXqnsG8l7RMqqrC2MN3f7klimshs6S5jfdE7SFe8m+Z1
PiCvhoiZPEujWhHj1ly2sHf7w81Qb48Dl5DOEDITWPLE9jt+ITGynEigxJ8B0A4j+LPWIHSUkBbb
e1HF1/9McHMfviE2nwIuloehRfUah7OpHEYiRJnTs/12aHQeAv5rKRuF7e0eEFCCXB2SS66jaZrv
b78h2TuLbCvdM3vT4QaYBn+i0Kxd0d2GATeCDQSgN5mbiOEK7dL9HVvU/KAcuFx6eBnYy+XJEz5T
zCFWSDgWxpkWjVx1C+OuihmHoFBNhGyp+ZkZnPCaBZSjqodZiJBtmQWNMh7cGqSKG8GO5p1GkRpg
UD6VQNguw2Fy0HPRydLOFkxefXnJ0gKUIIpRJ8YiTnPRahYrOFk9FTYq7F9GifHM2F9c4/vxknbp
pH7FJLXHFsEYYEXh6lj3uBgN2BwRgwHVrviLR274wBo8S41uWbJk4/vkb4Fb8OwthMQIOUrYYHyi
IwzC0kB2hpLM19MM+ImSrWz8nO4WRyQ7gW+tStY6HctF01t/ZSGgCHhpVO9v5vhFQCPY3g4ue+ye
G3mKlhovYCcyDqzNL+fhkA5yb+QLneYgNMYEDmpUOGlzM7U2CmZnWs52rR+Gl6bD9XqrfHCm+GHa
aMSd3c3pw0mRFhEMXeq7wF/QOKYovQyxAnnGPPb9jYkdyo8KFUYxDuXqgZd1HmuYy57adY9zCic0
4ZoNN8IizuNkLfm2bQ9vqLLxIIchhizrVSJ0ZDiri7PthuB5yDspLSxzQlvk1A+AC1wzHNYFC75Y
dkPZdCReYrVUZdZ8QoA1lWNifSlmtNKYQW7qWnkOajnwleorE2qhlPs9Dsx/p0fWKgJgvKBVXU+W
zWrmdD8kOlkbHK5MaKC5TXgXm1LN+ythHkPXSJvn+8IY1eTeDI/QnYl8L7VQsUahwN2bepJFwylg
eA5BYIdxZBtB8xNGMssQvt4ZoT8eJP38rvWgaVxMOG0yP88FLztGWPbRg63bLnY9idrsegZx6ItB
KuVXC9FrosjrxERUMOl6oACjmW7xS0x2dxcVbNfPr7EsqziDQ0YfJq+SfmR9fioAbCVJsD1wgVRo
Zpx2VM5k/X4ImyE3snESYT2RVLZh1q888Pi2mTWtlEs0wmfHaKSWACyJvVbauqJRY1qojgRjzUk7
9TL3GjiyEQQ/E3zSL77gpnvNwgr/cJ4RlDlcIvGzwuh6CIdmvgkjCSb0WDp/XKxd1h5DtslrIdIC
RkAIP5jXLQABwtTQ3Ln9+WLfrp/SffBthiSBYal6uPEoBX2JAFHulpaIImhEhrkq6DYjQxuxeXPs
k8fmTYhiOTChYPMf2SJnRhDh0+3ex09SbQAmaySi9x5hGz4QUW3qylTmCQ4/bfqgT/szaiDNnYCS
08EAEK4SXkbjBVKUPJblKnHTWPuXKHyRByMkCTVLWqBPwcOKu7hfHpESau4JSBTuUq2eNcM5t7Xj
NGFpPPCHfMMtScZ8q2+4QFd3/xM9jRILQXO4LNTLlVo5pdlQ5MTxJA3GmU3QWM2whp7I1Q7RbByU
RvjiYezoS/NN+cIST/D/Idtxen42QIarnd8V+Zyw0Hl9ayyDdNa6rirKjA18NHKKtHfmfPzABPjg
Vr98KhwfoEbW2XklcKbxCaKQgfFmmZi87OxMDvdp/jCKvB/A7ChZn0Mjrqw8jF2zJV+uBi81YDpf
afOO5Tx0+dMy7FDOGKQWVec+POCLJ/4MXd6paMgqPLd6kuBlvag6zKl29poQaGe4fdLpiYuyibi3
oAKFBPrfv+jRlBLDW85GnY2AtcnN19aI5yn8Sp7Ly9GaKJiVO1L0yJ3ppSq/cM0RTKLgBSoCIbKX
uUn24MDibcegKyJY1FP/giy2EVKOdqHYxgkqksIKESo5EwHPqL2XgnrJv71CBhuHLvzsiLyGON6S
RtlhWY/pre72d1pVgYDFji74tnEqLbo8kS3ObzW6jI3cXZukgZyO+JC5L7kg0Vm/12PuPj361X3R
J1P6QZTVzm5oIPJ8RTAID5x0+mNTdqiX7iS2ib4Bu7V+iZ0S7bi1vvLUoCJ8d9Hy5cCqe0u0X6+C
uaFxAXTvPfJ4sV3p7VYOrLd4IQn8bfxoRmb08i+ntOjIq7FtOCSUUWqqy40aHlFZlWo7p3zGy1Gj
j7Qjct1xoNKn4MZMBIRAZqsaxQovQQgPxSdh/BN2OxvbisQFGUzTGcnvUIWHicrMl9e/VfL3ZoOh
Ws3TVARnWA54/5wmyZyVCSlzHk3NaTSoDglQW+vvdUUqeUq+O6L8eFHO4cHkjXOwcW7s/xTCXXvx
9UHdpB0JVq2Dyl+muLPf8Wh3xF+MJ615H8pAXJatDlZHxCbXewLJlHs0EMYZ5s+vRwcLErjRI21q
jMWOCnaB0LUeBCc1Ca82AFtTb7eLC+VyAEfbpYY5yfiMGk6AboIJwmfYrMTriP+Zi6g4P10zX3hN
Y7sJVQ3c2Rsjin4HmSHxzsgXsgtLJSKkxRYtk2AMoxMCGFVjOL+6IaQlSrKmCzNahzuuiRBa9Xef
K7g437xus50xRKtoyAUfEoQD1sM+H72qLBiU0SPQnJS2WGdMM6/Q9P4qgaSBY1gCJPKDvEfMpHai
LULZP/p8KlknVWBkwy+EijvcLSGYvLySIMAwaMaTexd9mT9cc8hYU+QDFPxYb7xtrQAfXBMd627Z
6XotOeNkzUh7XcIjkSC1sfMdmM7ePyFVdTIfm6Iz89EjR5vyuZeyfK8LPLVE0ZTooEG4yMAeqZMM
B3eW/9Q9aznwE+ARxFiQa7M2iEhSA2TTXBMBz5Zuw9CRlj1dFu7K7oc0sN5PsonO2P4KKb15iASP
86g/h57AGD+8FHS6lHUl7UwQClvmEipGfp7Kya4ju6nB9V1NfgnETWbJiIsvhH3GIry1H/kTmw2E
5E1wHKISagtJ2KHop+uFAOlNya4c3LSHR8FE9lgNbWvE36ap3YjAf8zCEVEDGRpxhpICAEsfMMX6
MiQKaB2v8hfY0AGbb+U7MUt8DIcwxbIeeKKjzntTyWoJxp6BwrLgLc2wjhvu1NTbugrbJAmwzF1u
TxnXXut+L4RN/MHq0hy/QN3FbxBEHvUctRP6ubCwRUIm4o/s+metxmnua0ZWjqqivSJC8dN44R6k
ZOo4ntRKkKhLPL65T6Fs7AapeWfjr5u+q79mVtbQ5vatRxpATjXBIDGhGjxGpbUsfJp/GnShAnH4
1DvGKMYBSbHjkBcH3LwwhxMm7yXwCicIqdkfiJtB6BRCUc9yywcEolygeVvd2TTZ5zduKAGbfsFZ
kejdmmC5Fr7FQySafzTOMxak++cqk+dVN5QBLZALj1ZEnlWYkr9xIuBK24/noU75Z/x7f1OJ6G24
NQ4fqqQyWSmj1WHy/GQZb4yPTiRpj5R+eokCVF2TZKnmFeSARwZeLdxyFvXNsOs6RaSsFCY0RZwF
PdSNxe6rFdNuOdBJqdiBthO2E+W53AMTv0riGWTRVZmdtnSiMJaXABNCfApEb5tZHfubfLGwRp1o
91bYLz68xSCZgzOhMM4ErTI9+gZX+YScgUX5LNeQvuaqT6qJYxM9rzC0iDI2XuVWo833kS0HPKf+
0+6rP8g5YZZWoUKYFBCY+WjOzqOsOGUMPaY9W3FGIoZhoOEVzChPkJqQIHyDYGjF0Dyhq9ZEiFhU
umqWTILugkOoc+beb+0vCzcvXrLrlHM/h5GBMsq4mAMRJzQ6FilAyjw9h6gtoj+IV+HpONhG0pIX
p2m2kfzGyNpHveb3h/Qqgg15RP0Dve2wdAlk00CLdKUVxnYvenxgR89d/lwNUzoVPrybHq3TYw7A
KhfeW0WTS8MWuPDBgSjj0OpGBSYB8n6r+piK+gK/oqXmoGP5NEEGPyCYN525s1VCNs2VVaWgk6ZV
3SGeDcMEIwp5oLYUyrPL34EPgw+8c6MRLGBsNqmTPE6XwWzy6UfWotE5fHCA9X7UGB5qcJSL4AgX
j2I9c/nF0V60cg4t/7zSrfWBWP3usjrf3vpebMs/kvS4O0ikxRJ+55uzzVoAeQpv/90lmDLS+CB7
+1T3TX2SAQK+NxWwLROI5kOQVzqKEbMgQ9qtf4xhsVLkxVA2nvjft3EJEctc+tgfJcaAiZjleYu7
7wVCKJuBJNjGC/zIN3mdQ4xWyHmAL2yO+z28bD4kSgkiyELmXhZNDcAwhOmvBt4debmUTPsqBJuB
7IMURXkL0sL328RA+vU299NOCjqgDX/NsrLfnqUAnhyDdx1XVlsKeLjiGVx1mmf33JJp8XdANPf8
tc9FjQNI/2PvS2yf4qXcGnYcg3ofjsGW2q6g6sG4usvDxFdS2Sq/mtQ7CBN7nCWqlEaytXgICIWP
/9gRYxH91Ipwu+ZpwkXWQ7tWYG4OXpJqmhR8E+Mh7kwZHZ9dRFRMzvHb2Fbl/m5Cq/JZ+CarZ5lD
RW6mHIo06ZxzJj7WRB3QVZr2cBw2EFWQmGkmQ2IjuAZ7mTsY11zpUOFudTGV/o8rWTk9lMEN8sAG
/rKF1J7nm3OiqQ8u2gHlvA83spEOLqWOdXXiEMh32+QN3U0ZQa/lD408TW54k9XgnOkO1N28OhFi
09ihGvVt1EollnEsTfI2n7YE+NJgxoj+6/3TuzLnNvCJltOuySwOq/KxMN1k6Xs79moMhxEBdvSq
i3qhxwkYVXnXHAO6uAUJmp6/SWcKSbn57gsGcIQZknh7wlE4aI9atUdFGEfBMjDDhLdmZTNSDQza
ld0k40kQZJI0GBuJ3CGW9LasQFD6OBpu7xnE4ss+8Yynxiax/tT+gvJOE+mZvah7E0THFmomwIe8
rHQYm40OZaMe//WuNXU58A1QUnZCHvOlPbz1Jh9vCDp//W5rhaFsHnKwA41Uu+ZzX51ouEofpuH5
jOD7+1H9G5hISfeIgksVSPqwAocoOktwQNDWLhv2C9zsgrPBWBnXF1M4hbJPrjfCyCln3Coorsh/
hUDnURX0cdPBZvAfSjfeo4oaPWvHIQhI/uftRhAccZQd2m+qB7iZqcKWhGpl86WD9oYnvdZnIdJ7
8uJcKJ5Fz3Xcsa3pBySrr8BukJaP4XRjJHTG5jxNRSBiQA1dGihgsFnsqhWHhbe+EtMD8Cuf5fU9
u36ir3e0LXlPGOK3dTQe628591BR0SD328pkEJF+Op9VpGLPkQgCl5URab4nav26DudVgaSN1SZk
3fVyVXmWrxJPtGVxbqhLnOYnaz7cbXW0udMN2SXY5euCtmjseHUseSp6qO155zvyVBrrl9dIWXfQ
rknleZf9GYdEQmkTlDw7WTvZ0W8gay8c10RM6r7u9TDovVMMdb28nJ2ZJgjSDpzCbjmehXE1zNe6
tEZW22R5dn09AAKy6Xh39CiRylgmAx2o3DM7Edd3e2V8+cDM/cJkoIksMAZMuOozTVa6CwDAjBGC
4Qna3gUgmCBBDHDbeZ+mY0wSd0OfnRmQkRTjGp1cSlGV9kCmrh5Q/+mfTLtOIWn1u5OngLXL57Gc
ENevQpKEL5bXxvAPixUwolJTcRYFbwoH0vgOwem0hiSxC+SVfmosOgiwTiyqXVPxVkGVE/m1aYUF
H7IJfLPM0ZA9RyD4BE99MWNx9y9l/XvvpshRGNblGwEWvITI3KotbozdRO06S0htEvdH8ahrBY1g
VswMCRq5d0BnXCLjkIP2KLIHs9zgTIsmS0L84oxvm5dQ/qmMgO2Z0qSSNJGtHm0h70yqVpDElGmm
MDIeiFBM4q7qroDEEKy5QOMI8Eoh/uKAoP+Q9puJQSeyxaj+tail2LLPrJqOvn8L8pqZZtxkvEvV
kWFNa82OvFCJlFd9k8rAq8DX6qxYXJxEyfXXVuikZU5Kn8GrKnEbAIp8yUg35dl9WWxsLKk7hHHE
N8OxK7umocNX7tzEtpbHQ8S9o0Ashap3hNo2ZFGH4UprPGSQqQhgpTTXSGM861NB8zG/p6GFmUjp
+vfGfDT8Wgz/HinTxxY1S1rpzltjzhfZYnYlnRPPjlQpbr/Nj0Bvz3ogvUVR6CtPMx79tX+ARzNK
zBlKq8nKSEB+02+8sFnEZxsKApIdILtBDMl9buFacl+i2cFNAv0GodZyAL82hJH1gqYoUNBzBZ4Z
BZuYSCFrM26vCLgqHNkAmLgac23bvWSvz+hKVU9n9VdIZKuv6eb742ng2V7RgjXx+Pc0gJyvIKZc
h/GNPAxjqE+wVx8RQF8imufpyEpz7pBplnVOu9O+qC50TYCjSUIPTSKzSboLeruCJQixxtxNEjgF
RD6G3xS9bRbaf8RDbdxs7Peej4OQikMuiUTxoiGvnhy829gLifhRMydxpy+npTPDtROEVZC3FEHv
fiXzG8+64dsiag4Vf7ewgzbvgtxRxQzXbRzdz6maleY0t+YfFwqdYA5S0jQ43Bk2cKCb6Jwn7IbE
F54/rNBAE7YEfAijgwvzA3M81AnkS2HjGPl72HJei4yAJMyFv5yXHiEPpv2emROBs0jg/MplkqiZ
91Q/6JhEha/mfLx4sF0K0pKW1p5sVjPse20xQX+M8JedVAFc48rRWiItYG4FE/dOKkFaSuMuKNFr
OCIsOOsYulxC9Z9EOY+6y1b65lnjJinxfVMTOhi7BzsqIp8i3NglV1kyqR3lq1QTrqbBOo7oIMmw
mL6oHFmtjHJTjkDF9apfFfdAQ5LcuhZUVroJs0883V8PjiZf3dF9VTE0gMLZACoWCE1VcUSaEM5m
o2TlhI4rOApk7eQD4cneO1NEN+E431vgx7MtgaROdIuyfHOPLZmym/QEZUdadcFxW8Gi5b59wSqU
b7SqBSb64kaMlnuldC/SFRUZvNApJpcMkMCMHqhJPmvNlHQ7t8lGW1X09X1JuEtzX5u3WrpDgw6/
MKxSBZGAbjg+dpjqWwKcQl0WN6dYbxGuG99oFs+nGn6yAJzgbfzp0Yo3wDEGwyx22rlRfSZfFBK4
66ltItIRjhRvjyN5KQkgPCm7ejQfR1vnsLbI08mOkIuv4m6LzN5YgIVXcIa1u5gwUCYa6Mw1n30N
QD4AA4uhX7NZPaxGAnkf6RLr43+I3GGWekCvM8mbHhUfM/OzfqMiNrCjRYCs5rEzI2aOC23+60oF
Q/HgwUXpHM21CqMCMyQ3fbIdUX39tLwAzmdF3N0UnouVNLe+v8IaEwrM75gJWo9U7RFjoUr95Vi2
hQNPrVXUfkQA3a7zx5kRUeo4iAOrk2e7xA+ZFlB0lJTP/TtA9YH+nEE6rsac0fLFRquUtMHYNVYR
q/+XpGrdcjPbbrJyWwoK0/4ov99kOwsAs01354fCXs0Q7nADF3Iysb4AdsZsO063wQIlWtaKZKMj
OiOktYeRhYMlHq1g/kbVzuiDnBu/xT49XUZwY6miP6JTsqY50IEYAUHqGr4N/kPzPFyGIYSL7uN8
Lj+vCmisblBs0pKbyVsArxVqb0rwpaQeXXQXXajn0ofmbcqCPv7NBlRNS+Rg8+Sy+UF+2OA2Ddbj
H/fCo592Uf2/OxU6pKKwkVF7Y1apNmDHJYbsIQFBc+qbU6Y1fwyl61ph6o9sXIwIt2SHM6Y/IB0P
p0yuoqPfhb/44JDU9pubzsGcPKrE0I9ZF58t6aobLb/D+mui7ZuK8MRqNj/G73zgw7QYONUYmBOy
YeRHMrITwC96s2H0CqjRlUpVZT6jk27CSRLg+O9XiHi334jWnhQpGetkGP30LWEKqgxQaYDdElvf
BV0Sq6QAJBa0gbBP21igVcv/cEda1pcp5hx84FkwdKvzbTyqTd9x4T1MRy0OV7wmlC1k+gqYfI7z
KMHbfe7LcocLOrK/pnCSZtSsBEAmpuAjyHhCQhf+li7szlLanORfwZn42AJ+kPVp2DQhZgQEVhKP
VZw1Pt3bzTT7BvoaY2pRwmFi5x1NJ6gORxW7VIaY1aOUt80LCaws2ppnsy4LTHwdITwycM5Jbdqp
c/u9kvbiG7el/+TULuXdIKPEfvh7raeFBB10zy6Z/RKcF/PbON24x/CNTwMOkyZsK/z/YtU7Oa5W
GiPBmIDM7PO/psnFPpmT09UNr87TE1gTz5BPZDVMbV93ECHcmAmzz8AZjxkK5JH+KDf8KEjrnTlr
cNsd3lwGY/4/a1/6XLsTxdGwTk9JbXDyRv5TpreBFKhR9pFspnIpAKV2w4KCMTYxOGppTPdZ87e8
/9bDisoDLClIeioukD6T06Y3agTIlKugfYwqhiQuxELNmfOfk2UfmsVG9YGW5+9TQZv+X/iAOX1z
gK9IwfIXGJUzAWGzh9lir0a9S51y/HSLa+xulO9lP5JIIHlWcKzB7mkwxtdlBRmnxU7bbd8b5UDh
mQSn7FrxHJT26QFJIrwdABc9MRZTQSzvIEqVWPpTpd1AqtKGbDBYtPECiAhDpPBiewFbZ9+88pZx
YCUjXIwG/hlGvSjhKXXWKn8zs/fbPxrvNrtLcKjQOEPvQliY9tVb1u0OGFPC4WSViFJ2Q1AJ0VWZ
HlLj8l3MmJxPIu7rBojRil59+HptCdDBnhRbW4y6rRo7NknomxxfxivWN+oXR0msLpqWEIj8dxcd
RXu8Rhsh1f5lbTO/xGkGaDkGvt1EUKhb6xTvGrF5BZPUzRUeEIQapQDBBte3x+VBNtObHRpwVJ54
J38LZyw3XY+pfRPgadWJBSkjUHHP9rf1vjav/j47n6WdWtfXougb1H0pszR6KFW3IW4tFgNW7X7q
vYySlrWHGXIX7UcMrcGgarcSMIN/R/sZn1+cRWs0a7d9j3EX4SZTMenQaiCm8gsZFQzIj+F4XTzU
0bpYtY8cYCUG45EEegrty1xRjC5Z16JFTT/rqSIMbeOaiXPdzUgk4Xt48ECKrcULhv1lvGKaizCK
PBo2v3zqgKyRwuIj2mZpoqKU6LTf0p7VLpE0JR0I4jmx6PW2zIi9vcFMVI5UZ3qf32e2szu8VOKN
NXYRzf0b/caKa/YdUGPlKqwsvNl3/cl8QfDImG5P5wrAXuIrZke2E6wFg5JCCxMMkJa9QYBtvkPO
s/uQxasYIHhVNAVHnqKkgzf4OA7Y4dLxxnDlonwzLf1i2dmQKU7K1kJiqnkfVtSDUJhN+SDmHun2
1UeHBi9kVk7zC44zX/KSbWlCdZdY7E/cifhVGkk4lcBHPZDvMIwDX8sbPCsjuUjYsdGjlqpFZzeB
860QR7G3TUKQVt1iyOV47x6pXGvuYCnhuHhh5pxjznRSMKr5TOnfVvySoooPBTrejSPpdg5iLblf
WMD6UgWfLIjoTGPbz/SgMG6H60MEGB0EaG0Y5CFX4iL7IwW7gzB7/T/LxRIKuLsvBuM69+MljpC2
NonEg/jhB3sBN1biiSRC5k/oDOK7Fb+trBGxtmoz3f6Q2EQNzBwCAs7qZ4YZhDaw+yAd8hpVLsEy
Ogep+fEIwW7K7PujBP5X1pMXgnJhtOXhjL59qqKj3xpoY/IC7Utzh3q8rfRpbRyLV5R4/YZ285CL
IOJoqZqXtBORujB5VNmb8rffZWB3uYs2qjw2DB37hC6jsZnuqwUCexaGV9zUCc1BxaEZ7z4/Cmgk
JIxTriMzIEYbwmmYYFxKnK0qV22jQD10h8LKHWSJ20z/h/UcqEpp/lCzqhC2+qnQTyNmnJOsbdw3
DfSh8mpmwf/a//ycwfeNLll5jkhGQvkkMUErhOykDO7OPI04rifIbk0hotMHbScvGYUemLjMlsQ7
XtsuzbISIla5z9jQBNi69awjSESolgALvccUBbNJ7zrmH+bgB+dTgg1MnRQIO2nGtt/EA+cdKFG2
Y5jdZOv1bymRIFGuIVsKPGlyRt3AigIxzinkkn7Mqe+yWoQxSG8+p+C2CzSLnbO0x0zQYErScj+q
TjJ5y8FgDlInQqyHRUr1XoN4oafikJmu4HkLuUTGe2jUv999IHI18nY1tDrEZwzLkXrDrOYvC9Hp
X8beBukX3cXQmxl9JHW0wRvHIEeaS9PNDxAuHpKGlMEDPMskeJ6LOI4Vjk7tMAlQ/VkatgxbJc+8
AJaS3BJEuy94lENklhHUsjTOeoaV7Rb7tGPLIp4q7DWoBVQkkXyOhg3Tonhi9x/HpcR1MY6lsh3M
F40CZaud+3FMQZwr0IdzB//bF8YQnj82CkzvNT17cs6BDnBuuxxcRpN+wxBR7RU1sa/6xEqqFRF8
TiF6bTLcWOl8xj9gbVyO1brY/IHRZODmEpCa07va0PJIYa3x8oANVMbJD4e5f4EhYAjxanckE6Zu
gPIAtIgw1/FqYV2xRdGx75Rxl4mqqIuxmXp+z3vVk/FmzBI7os1yJWSeKx9OqDqVMrb/u7+qWtCT
Tak0ODlYks7AdVIanABGn0o+lVJZSk692sZfI68Hqdn0RxqM1c847V8+K+ehMgrmj9sZE37ApSts
kkGbb23N+L8u9PH4yVfgspRbEtmfLFj83Sqkz9wX60XLfQI5Ukxxd4MLFsqo9dKP3jwX7scSiZo3
vOHQn0s6DLR/rqr6bX5HMsUq/k53LIuQ5k9Pv6KSsyyBdru73SzCJTBpegd37uXVUa+Us2RoMr2f
fq92V6GUgp3tTRLoLLZazukGYqx5PcSf2/T1n/BVEmW+nZn0+/ztuf0kteqP2h90g8+vgmIPxPG5
8L+oJyaDz1nUqJpPLF5rR0yVaLjUuuU3zgWxgGZNIvFzccUlUBBX4Io2pcAbo5NmMHXgcKcrNQLb
/FK+UzpMmu6d1u4VU3lqSkiEMUSt7PS7dqz5KQgp+U6Ai7r0+5GI4z3MeW2jE68Q0T1z6DXTgX2b
VEOWYhEX8oRfVpqQKhpForlUYn/igaFUg/YxgCzuNdvHxrE742PaXK/K+Yz5U5oNvjI6DZl7B6IX
kCslqkTtjRZyWO7qMp/+onk2jgEGoCb+9YiBrldG2KzPol+1YwTGLb4P9UJD0bs2X05/CyH3SUOh
OlDKy/3yO1MJjllUeRHzdMIHYGEcI80OdhWh7o7niilQm4n3Y5gY6hsuFO5h9rx8OfRQsBuTyhDx
hKjIDUUrDCxiX8Pw+GNlsb5vd62lzNf9Xs1Bk8R2o5+4jkaJnZnxyh990pZvYyBqc+NOpAXyNkF+
HjRWJoSopDW5asNmHW4hL5MnKyD4F/OQJHL1snDoaubXNiEG8dPVhUu1qylVkn6HBM+6jFNR8cX0
CA5+dbq0clRQRfidsQhV5H2GGnWXneQbYRXFGRG7AyQhLr/wjkq3BcRO9hpgnERTobw/fMmSxdyA
otGn1kc1S/pccK7tmQpuOH0xWPPO4xPUThdjHnya+mQsx0jwTiBDbxyICSJnlwV76hHDY9upCS+i
VX9AltrFz2FpcllmjXVYRFt3GtCppBbCr8IbdKoO1TsINP2W6X4IfMOWLxnx+Oxje5pWGvdNurI7
PJankJN2KHKlw20Nke8MNzi0NPo3Pb00iXQYBsp0RefgMUMJ600HdSuoT01qBLgv7g+Nk5LYm59F
T7/FTds+6LiyPOeVaemTBJs5EpyMjGihgL4OOq6PGZF8MJuoUmSg5v0Xnijz4TUSvB9eBlzyyg5D
/bRF8AkfoCjbm5DrejJkDNOjPIeXfBLbj2tXmdT4eEcHQUc8uonI3tpJGaOwpcSIKDQZIgdJtjGa
9PWf1IQ2jgxI6BNyHXGdJobfhzVOT4LShFacops0mRrYrjtGr3r+sggI/xEusbF1oClcUVJaRiyV
ZnEltVG9zLk3MvURnNbH/BvhQPYbxWptm2sd3LNakprCEntB/xipRaZ9vi110kaR0EVUIIGxOHcF
JxajwaDu+FGfKv0x6m4zpcBdxntbjHxYF2CHHhu1jbplefnc6vMnG6e6tqZwiX28ItT8wxvbWrUx
GLSBB02Vs2TUT7SZAPmWTurh1ca3Ki6F+RU6bD/D140PcewQ18C86CGNSQ4J4OZdU6mPuEq100nU
nF9AOHJLlk//zobugI3QIgqz517zKCmV4ZT7cKnpVaWtK01TO+yyLciiPvLOIA3j//Tm2FpNacJ0
fmxvWNNym9XP6Y2fz6J/fDjifl3fbLWNt9RDu1bqsQt3X7V/rOxB8dcP7YkbWcq6S2jm22yZGqCI
kM1avSt/lQgNWTmNwY+nrSWRfoUS9i5KodtwbCZUO7jJDXfOFLOC2fsAboRAcKQLdmeiqo4xuwmp
yo6OT7r87m9RXeHe6zjLA/7R7jpExz43r6fpTOK8mK1lgOnj7Kv8TZRwn0bSSYYdIqBpgs2pybR/
r/oiQknbtB6ROH1O2SmgZkkeG2n8Z5Z0UmjeN1suOUBlnKUo+uv/a9FNwfP00HlDiTzM1VlsTUzb
ViOnGx9ogTV6ymmpzXKq45TXfBYFj3PpAdmhCze3h2rshCwnndennuUMPE5HkeV076kMojkQHBtM
1YxXne6G+GtHnAwQ84Wh8z4TXT+3eAmtJvvobNFhQcOXgcuwmBTcUiVi/tdC7LFJeylBZsoTRjFl
n18u4Q3yqimkdef6T4Jfck+fz3TehBl2ddfluNUflUywv2TpoAl2WwffAqF6lQwBRgAQaKHcyxaV
lMbezO2tAceCnanuHvtd4axYjda/1nTWElBzw+6OAmnfIVLkSTyL+IQEKga/5D3zisU+5dxAzECj
mgAGhYfxxUgl8RocJrnyzL5xh1w78K6M1Gct7Xyt465czXNpenpHHIJGZs/GNb3W61A5BD6IMrYP
LUeYOjcTHL/X8YY9QkO+pThnfOEb/dsazFYcXDNl2scu9+2X10RvFfVYBtARMwMUqwLf9t2dirtC
GN+uLnt27RtzseXBcWEBovovX0Ghz7nf2yTl8IDPg7LWeSc2dyIBc8RlTiC+gPbrdGKmpQCNHFCJ
aUzkDqKreS3lYZ3j/OmmtWtQOXMWgymY6QL8yUr/0BTATz9peZzR2mtiS+e6qie6y6Om2Gng0pbB
UnWqTe6vhHPwZ+IBKU+sDtBIVvxPKHv7NjGr5MCSA4U8WaPYL+mQim8haEBgXrlciGymBJ6smI9D
NwJl/KXWNJ163NKaftkQtGqhHVaJxGSUB3oBmZ6tuo2gTKIKhvfrS8z8Eo5khqAyfuTgHJL6a3ur
q4MYP/BDlnjGQp25nyqEHgOesReWcFiNByH7JVB8++i2DyR9yXpxYxu8Qm5WpaqanyjBP31RERFh
sNwZdfANEnbYHbjKHS9GEHUWJ4vL7zd3lQpOfWUvt4/MvJ8yUrUjn9fGf6Mv5W2eTNFgIAHXnHN/
TjKVTvVGjctKv2CH8Zwiv2OT7fE49XbPDWEszLfZ6nbfNS8+d8HVUA1Db8LE3TcmuOHwSyxExtG7
vwxY/UBxAZRjFdMT6WDaQGHUizeOEZmPgAa+WB4wQHZPjW+GKcup+DNdnyyXkjc7sL6SpiPFwe2Z
IZAF6/EMfK7YA0W7x6SOg/cC+xVXMO9UrFUSbqMyAApV8eNXQiCwE1GUk25a2eTBttPBouqzv212
hLOaSovxHyuWq4uK8SngmOoSgg4xVdTOWevKirqep421gzUojd1V4J2ey/il5npbN881nFKLcSmv
c0/4mypcmSHz8USJVmo3b/Gt+PjrXQJ0FCXdZ1f9CUrzg34AXafi2WJbs3XjyfrsDi30KiGgXgnA
cZLDdiSoIwrE4a77imrzktd57dJgj6yljwjWJ4B1vxEK2Z8OaI6Aut0mQdemIaFoENpCjVHchk/6
mQwOAslTlzarC4lq1fVe5mmsJTbpIJiTtR7QNc4hwQvh6HgvT6WGEEXA7j7seApT7IWcL4/aF44i
aECTJjrybx7Q+WoPJuG0ogWQ8ZpM6kF5sKITEK0WhBTLaI3v3wH8mjfOuzP/4t7VGNxtWWQzC3P2
fc9iGfO5QIdHgf+oCF50weJftMwmG2o6I8whv+GGn1ogUrwiF+R3nLmAUiehfpaDINi+EhV59mhZ
uj7RJTlma53xxBBZhqVVIE7D3P3f4GIUyw+0sKfh9Dwhk8AYJ4caXgwRRSIC6gCGFLVobw4glfdM
fOi+0xUQ04W+4dntQFzS8/TpnfFBHQ85/jNH5RGKsNixapy3c3ZA5w242uM/4hPPEYOMFc3RABsi
FkQQikaCVCaQIIxzCatuvalnKVN5j+WeavuDY4zKHbVLItDnrKRvDprK4muM9AP3AO+bNod+NpIV
3el5KBtubE0lf+gdUthl+T3Jq7KjDTPTl/3Akudj/33vSfNyOYJNHs+op7IfbvgqUouyK2jlN65d
6co1pn6DaOuqgYk3G8jK8EWq1wBzVHyUTYoC3Cq+N1pAzvGxSQxW41sBhj5cnEN4YNQyP5LW2hL5
mz5YVUqD4vCSp4AxYQElQj3RzMY6zrdJCDVS2gNgivbULdz+8VZs1sWAGESnCP+GMTau7w8d2n/R
lL4bQ/sVNuLuAcLedyUpPCMWnJ6NUMTxSk1/tBGMR7IopQ1EzxURofdkq9hjp4HaTObcSai7w2Yu
CnnHO3Oh7G9aL3ofn9y+K9lVNMALUjS0NsQPafnNyoWgq+1SDILXd/z0+RWAljsg9xe+3TQOMSsu
+qlBe1lZOipe07Slijc2EhLmA0iEiuF+2UO50wWUFCid532A729UBxV5DeIEmoAMVUSwTG1Radbq
VyqWHhfmM7UPW9zxTPP3+vbUEeLj+EBuPj4Qu7D2wA9PoM3cdLTTQQUMdgz72dwaV73w2puADWnh
obhlIx29W91KjemDD/iVMHwXCjmXDn5Fam7DQ4RUqF9ztYE1m55IujUSZ5EM7Lqx9yfmc7/q/4XU
nQVh1eniI0/2W5+chXsqYhD5YKdyn4bdGZN5IAcirnT5sppvK0m6jWCqY+HU9Dre1CyHjb6YwBV5
yOVdTfOHvA7XfPUvarIW5RpHzlwpOdq1qVrwfABd1IH/StmHXBS11qWY44bKHkdhf7FeF26DgMlG
3OiLIrc/A1sxvtkTSfofZCzUe9w48gG/Vz11mzqhs1ew+n6fXaILnfBQrspu1SZZGlXwdtSCQmU9
YRyGIjcDP5bGEGHH1PJ3efDglm+M58CIDStfpQxZejVA2ME6+kbCyHPdq3GxLfmg3OwTZRgcP5Am
5IvpNPiLsYRINdnRb42Vzf7h3V/RZFKyRBctnFiNjobpJr4yr3fC10wMTfY6GCcruwNisS9Jl0Gd
eD2Ne8OLqSJYah30GFn5ANnTHT750P9sTZQPavLPm8ODOlBaS77Zu3I9grtn4XTpFQsp8jPbpfRP
N8dJ1XR+BR4X9cCqda8rhWOeAxDKyYtjVlRrIIG+G+PbR2P8IQhzdYUrYjPBJJx8GTC8qkaAF8Fs
ukKzKEbqDoclmY/ys/AeyhBrtOCCp0ladtBeRBrQjgQrx+7WOazVG/5e+vKpIVKNWQS2NRmNnVFm
MTgriU2Pwl20Vux/7IPL69BgirlLdrFaFPs+gZ+Jtl/RPQFGmM9g2m8uF1K3E6whIX4gcG3Pt0ab
8ZTGGVRw356tdzxr+2cgBVNTrzBRZf0qy+ta6cQ5VZJFtKucQn+4e5XFnVv3Hh6ehn1HwGSk70oN
3ltHY35bCvGr5ZI+162n6oCyZ2RQLTz77yCcuBukuqwEePt4UWeONcg784+sJkaZqeSKxLsjKMZv
UHLSZXXupdD9rdQ4KfIo+Ku0UlwvdMehzCskI30Av9TwF6kmL5OlWB0q27CpNXERK7YfK+eUJXyt
oQn4h6CRvJrjzD3KCQ+Rj7/EaEnsewCYgPA4orFqPt2klKokY2kBXntd+R47ShVQIPhpeeLMSi2r
pdaYxLbKZqmBrUsVKX/XVDgjBdXq+tK83SqX+Y9dryEtmfDN1A60638f4xc5JuHCpEqIiZ8OLKIT
PamYHFkLmT81/Kvbwj9ieq8gpzVZm6CDSe74p8gc1w7ySQaBAYPLHwQ0JqOsZjKbD+iZ2qyk7cLT
BgX+m7EKePFxUyhuDuYjIVe2Diz1pg2gbd/G+zLZxLsPBFQ4tc52vABp4hgCHkyfskHwKIrA+mB4
8Cu8a8uToQ0SNNiIC7D3L4UpR1RTlfMqtCkNbqQE/DWeErwS3fsu0YBoY4stJsiFdyz62vdkzsXd
+nRsOJ7CGPxFJ8uh4s/cAARnoRp/vzo4+oqeR9N1n7pflK/ad41nft2UhurESrN/lmqcbGy1wbHT
jQRQA8ZfVG6jLzo1IPjkla9UsEtq81lZkWYSUP94eofM1MUjH9jFag5FRkZV07aT4CmoPcy5N/NN
skOYFKa/hS9wiyHxdqgE6h4EaYBIFxerdWUumdOLG9psPeAUUKHNojoOrl5iUX6TVWCqLQMbpVHW
ehsWOOJS4Mxi/kT8L2UuraNpzU7NGXMU8RLgIfYkp9u74oHyX25LeY0xMo6uZ463TN55Jg5dXoZ3
X4PhBCsmDdWix8Ak3oABiFn8P9KeKFirQ9Pb2zKIb8+7n5SNEF10KW7Nxqi+mlynVqtIr+iAgpfm
nDIuAOqg4UvZxBQS4dUrElR7D/978HkW6JmfqAmUNmKaMCYRpxAiHy/hHRXnUg+youQhv+idhXxa
NKYpaMbAoof6CFINC1M8tCyUbCt6csPCD64X7xiaqRaFnuC0HeFoatNvmAtQcZ/yhuJzbEsrs3lr
Eo9+7HnLDwPs1/OcTZGtkG/iyZAdiQM+cQhn03U6qo6AcjXxTpuooXJEG9Kz1PTW+uR+zOUIhWsi
/OIYeYfnVoPXWQSW7OMChGw+i9ZiFkUSRWcWFu2O+QxF9B71CoaVBrOncD5m8vBKOQtp5A6+Kq3/
wxiSIqchSynOhQHMwMIKRC13X6ja45TSJ9bCzdk2n2rQBH8xU5FJKiT2SQ1/2L5OK8IUSLDLQ7Xx
Oldw5bhnfdgMLLNMfYHjwbdiqlUSrMtC9PzsBLxH82M3/k9rEnNyrl+1tlpu6Izm2tQNl/nxdmLE
zpzeRnUz5ck8xbaykjpzcNEWmQ8EefZRhE4FLDcXQx5tIZosTaFGDiIWD+R+ji7PbpYn2tAM0bBn
oYN0bnBhSUML7PbolSeBC7sZKcxeqejtaX68L90IpRmagdzkdG3VqzJ/A6akNegd0MMXaiTFRfRN
CpiNjwmP4k+nce7vlVIVc2dIe46ocMmOtG4COByxHUFlNUodfbw06EoYybQCW8WtI9YWTp26UvC3
y+OArna5smmR9hHSPgRZFnZoKJP8NKrtXvAHaQR31tHjkV4+q2I8+AkzuqSi5GDaW4Cck+raM/7J
EzoB1DJj+Uoh4NBPlm2RMl07imrUFVN+w5QYJXNfVqnI/VmZtFlIJAxZF/ehwroseg2LdSF8gAyg
9c111apjN5j8SYKl3lbfNPtPpo2bXllBZ3BNbTucieLL+ejhW94MYLiDC/2zp77EYnturmVliT5K
zMatWyk5+GWWqKu/m9PLEfwIN1XO97yz4sjI75yLjpibv1nzS17Fg7BdXdtffE5XSg7kgtrC1X/M
YR9yiSkhBq/UCs1nw0rO/Ud+75qArMoMPODxNWTl5xKbwbiPTkpfXllIuDNUkhKioIAPeVzWo0tn
ldF9iOJ60IYOnhJ3W5Tbricfjs6/UwsgeVtzNrYTkPmzaixHGXVPKXM8sjFp5xx9iHhOOY3oCdbx
ScT+Vw7Vyr7nfcxRCOz0wWpG1rpZHeyuGZno0VibAR8McdgvJ+eu0BrnaqCnkwwv5rR/9JUQHJPn
YBm9yliqL6ERQlShak6hbB2UQQph3bg8Kn7QvimsLQsDbrQD19XxEIij8FM5Sbe9gM80hfQKY9OV
SeZzYkM+/r++MTvRB4O+/Y/3Hv2u27LnmPgEq93eBWZrt+lLpUxuYySJeHez2CeslgnvKA32mI5G
WrM9e5DQpGsz4SFWIciYt3ETg9WqQq4U1yOA1h5vDbL4ZWW71uQGraKOZFV7p0lnxDV2y9kBtSw8
sf6B89yUYTmO2sGkXKS/RAymSHGfX3X6GD64oOTES0WqNdmJHtdlwatRYIw6qlAPFIAMb0HqL7Kw
eBUnkh7yDSF3QAHLUrOkJesIWgKAyPK4v49TNztJBnG6uYkgfcI94m42LRbLmG8H46yiWhPshEsr
o6KlUOrE//kNCBqlDRF1mPiSot5dWqvqa86lxDsTUs/8WSDN2A6V7LL3Aas+p6TxwkgbV2o1wc0W
21qKTC5EKi6+XKPrOjg6kMd5LsabcLYz4PyHoVQNzIls9dFl5CDlmij59bTh23q2mMIxwt0boBnd
QzLU6RC5jj76xM13vYR8WRlzNxVi4FM1TJubpEiLGyNQLUT2dbz/bGkYSqKbocUjRENFjxPdBDtr
ixymG0CqrrlKP4XxQLwiGOEQcPmFNpGYbtp/mD6PJIgoA9hp9zps5ewEVDAYQc2G/P/uHub5p9h4
gN405NGSlp5Ji72AMqCIocs2yA1HrznLMvy18IZxrRZq3KiMexipFMGU0VFy07Cm9WD2TKuk1PGF
b8fdo5qVXpa6wIY4eDqmFHp/tWTWryLpsZusf8igzI5BlnpsqV6dvYb7A32a9x4AhYc4Eq5rULwh
yP2LjroF0W60JuaKU+6DHUdthU9Anpuwd/95qeY/taeH8F+++BdUe4Sn5/BVttnN5Qjk+3Ypvfw8
CPog2kLzMcOBONcXogCRmBL22mSmgaTUUK33vIMCbkyR5zhmgfQgPutqdNbOHGa3n7UvWFvspVkV
CHQy5551FOlw6elV6Wytp+T45DMRhhMVpn+v64CaZrWVnxhg+fTIsuI/pdDbYAuPuvWkd4fbNzsx
l9ROyE4opS8CW7rMAbIqedVm1NHcpajIne5JY7iPghe3BbF+YRkvXQXlckh8qk7WDSgvfdROFu11
WGf7BYK+HtK6bTQ3JIMH/kjn+09OTAuqi/syte5oTZnpi/S4NsT+b0YmxhNB736nK0m2rylveb1a
w/uUIt0Eo1EY428/XGbrQDCAz+XlUWmbPWscGYETMNBrx7nUT1nAug/fpXv0zHifafLMB3C6gxaH
0/9Jio8VeQTGhpRr3IRaVmpVnp+BOEHL1cSYhMPm9J9v4F6xFCVxOacjvmsZb+41oyHEOPn3T2rd
AJzdQLGYT3H3HefcnlU6rwrgcrIFnLxZCoz7a/FvNx/X4Fe7pkJ79AqcRSWO+3Beq3W5cTaHWO/X
SmtzDL+GOwRGxsGI7vNOnJwH1qfLagQAGrK/AMwAvL7aVva7cWV7XEAtDQJI7PtOtrOL34hKLyGN
tcSVmsuoGUnE7gow2EaYVGuJLkR3nsqHvMwSUMXXDPDtEGcnMf51IwCB4qZ7SkrTelI9Nm0NfX5a
zhbolv+P9LmfAMLvCD4bGUmuA1djlKFfAMISrMABOTkRCgTt0nl7RYmTk5xPl/KmD0tmU59DFWJ/
AzUf8jEL2BWhbaZR7Swi6oMQjjIj4apLf//f6t968raRD11swKmvW4+Oi6CYYNO3Loj+Z0x2jUyy
NGUJcXE5p5W15PMc+MAxhjnxNNqOJPg18opb2cwqOzra/vx7RJEKJi1kuDNyCu7MqviYCCfK4Ci3
pPsodZih+SvAMPA9cY0lb2xm0A9IRPsvU67EvJ+PO3+EKBqHF8gh8k857jNw2IVz2rA7pFHWbgKn
ujyVBM2GgWduOY0UAXxcFvcK3CXQF1o7UmvV04RxTvvIhY8NBPg3qRS9R3Lu6yqVxrVaFjm/tzoF
D0jCxbFUNi4siCFl3lr3B9VcunZQZMpqx0qnWbp5W9dwJ1aMX4djIjBMHgY2PHlXFpBgpt5ZTfrq
6JHXXNd5YtkHOIoHFD8NWGu8UcpKnyBV6XdfuTPUW1+0p1hRERTKeUzmYeDaW8XHnr/nwMIl/ZPQ
SfMPg716Ac6zOHzH7nKda0XMhukvuPqAiRjwu8tP94+J6L2OQb8/WjPwyxMvKt5yOdPgasCYb7Gy
94tRNsP/ltyHlx0nzxFKuv5bew0VAh+F1ZnCYp6PgmZ9Ud1v1AkbtsKQB13MtKhwEWJsTVCLVBma
InFi3hQTeCY6PXufdYS0la/zEEcHrXtqWsXkXYqsq46kvik2YnfEODYu2RvPFfjlpAcy5T9d6p5t
6AJNN8OvNcXSLVSbRGDRmMsAmfAQN3Udx5I0N9qe7EsR4G7JLBN8RU83N8g8uiEs+RGWcGk7tzfe
q1dr2L277M3Jm+Gk1F2Uo1eK3H5oC4SSSebpj2+18+DYFoFNY/wnxUxV7NZp9voHUZfl82v3XEfU
wagiZHElCI7WOwXZsGQgJQKXuo7HcDS1OcWvAZrBjBC6ZrqX31e4QTlif8ALuSh6K+2ci2xNQbYy
tLkbPxZO53xeJ2+2BMh4rL1XCMt8QSt8XHWWq+hgoS4GVaWvzjYvu+l6bgSoI5/9fa+8zc1pHgks
dA8DI+z+6FcAQ7BtTZEw1yiDKrdnxgbjEgmVzSnLvlTz0q+b3YT4+stnye0s9WPOZEeQQUbI5VF7
WBDeCQvW8rwOXERfaNxcOdA8v20j/iLjL7Tl2pLVBO2DWrk6v28jpgVK6y2rWQoTjISNs+67wyGV
aj0xwHcayjwox+CqBbD74Bzl3Uf1xMZ5+zn1s9FoCuVZaqugZTJuZ0Wrj5fSV9Ci+wfLBhN3xuf0
SiLOkVe3jeQohex5lwV1uz0fcsQeFcNUTI0iJxvIP6Fr68goQO85I799M7KiRE1+Hk0GM2lUW5aZ
5xVvnZKqJ4Sdw0zn3S+z0gAo8Ur4Lp2h/QqjmRVceK32JkGs07MDNPcQjBSVHUyIIm8DKNG6s9bp
paVSQ15fWFJ0Uz4jHgncvquJbuIn0N9fMf6m4VxAt63KS7CloBulDZLx3+gyw8ZHN9ioIqTJ/69z
6WzPccXEGPq6vAkLIaknW4RcTkw0HyLDB6LikHAQYjv3D4EAxRTIHaJDIiZlEg2U2OAWgM1+lITA
P7g6eshz3O3+nvQ2QbzozOdW0CdLgyEjMW8dw+W3PuF40YARoeh2WHq1/1+DQGXlj8T1s7F9RJai
fuEJcPllU9SXqJKj2O8XHCsZ9dyjPImbxP4WKz6nAGBYLJos6n4VIy4qfGY34FSDwUjg+eNEb3Kr
E7jkxu4h9AtHaZq6Ol30JxuA2rdv2QG7EuEcv7dIUVoZQKN5T2CJQADEMP7DF0MY9RZns9jv2dsF
dOo60pn5qS9ttaIovF3ADlTRn4IVdPPEFNerHTl60aMHhHMWX76W4fhdCEts84XaIjoNatv3Ei+h
pnoGGxwe07hAcY0kr7M9cQ+6w8dvlBJQS/q29cmMt461TvYumxun8/Gz5IxeRcV2LbM8aJmrvjNC
blrLtztBuw0f38wMuO1xw/nXom3ypv7vOrnz3SE3KAebfOnNlCg68qu/ORcebdEvu3+tvCVHoAkE
nv8eWeo+CMsq8ikz3PZk4X8FXN3exFvoXnr4RuEuAJmOnsLHoUEbAXXG4KUEhuwLDAVO0+A8Q4Qs
WcSomi/Y+/rQctgz5Bygr9gTEcrVPoGJBp5kgAzatNl4ZIx3e/sH/9uMLChRi0JjDS7EhYZ9hg/s
M7+uOAYbYPZA9jSDyB6NzlXBEi80UQRRWRkCNF4G1iXYuEbYpqcrYkXxWEe7TPsBDMPuESS5MeLq
fboTL8ptRj2LUhvUjfNSDCNworyEOSjQ7nelQmiDHjEvK+6RVuZOk3Sp4gQ069g56FW9otG5uac6
U5BoRH1suD+r+gIh2JN1Q9+y7rfBkakQbeiONtU/33KKFOUIOjeVuuP42ifBtMq/1I+MHfBSV27T
lE0qw7KsUcik1iHVlPgBaYW9Rigdzb2VD13f6CKxSRO16F+cVLVjyc4/OM4LR+y3fIzmLi1W1I1p
rChdYBgLmW0sih6NkHxzIj8LjNMl80dTAnOEwtWaaG/tSsrzxNplbiTlA+sRVq3cOHah32yTr3T2
g8zav6iYSwKEvk+TGbezYRavzZh4FXS9uXRkW/AZ8MvTHAf3QWG+JZcSgbj+OyqPvbwCUQn8frqr
+f0gGWiQ2pmdzZrnumdV0QrXhZGU2oprE+eorNUFKBKNJXtr8ZEPBw62CzH390dNJd17x/240s20
9gf6gH+AOGwEEVSot52Uk1mEYKo4qvvH/xcpK/kAbcvuTgzcQSIuIYiz0jSvXDmbs7picc1ayBeg
vKhaPDpoUQ51rINc99YQSLe2WvvHnaHKcEV8A5gCo3cMe5s1MWhD1+JIvIoD5FY8geYtletYQzF1
Cqu9yLMVsD2eHF8gfjUv0qSX4sZqp8pYmbIJ1r/aOl4aSWTX56RlXSHeZorL5F9Krd7yPNYFLJ4p
WwLbSFG/Oi0q+2pp6KvrpxvW3kKGu8emXcPpAYgn/U8CT1LwZLgExVmG3c5Ew+a98jD8LHNFDNG7
xIw3wPaM0RN6nPVjqWDqOQHjozImqa3IGNwZ1DS304naKxmYdfn+8oamR8g36FuJejpNuaK8a4Fv
ZVlrTBUFcGhHrh6infm/DiMIIPJoLtJCU+nYJxcFZcA3mGjZGGxYX7AU5JqmG21pS6QHrBv0NJS4
srXtQ4AzH6UCDY/ACri2OTO+mT2hNDW2tE8mgYnJSmZdlcUmY4QRJes5A+E8Ddiy4S45XHKg7U2k
bnhPA4xCHPQ2l80PK8UOGQbYP5MzE9EccrH5hj+jlgoL/qeh1XNzZXQ3YLLnnZkvdp6VPYSEJ4X+
jZRZ5NDfz3/j3hUbsnbWPeG2MT3NhmWFkS0qDOjrNARLMDECOiRTnDR7CrAA5fkRVVu+f5igZ/23
GCw5oLg0cfL2LFXvoy84olzHDeU/Ez86R498/KaaYhn/UkFcy7NYkDKR9xzUdxmyF1G+kSqxaSFT
NwH1SbtRApZFe4L+GbIoZojkn3hZEinGzCSlVM9VoSDuLlnXuhQ7T8VmLiWBMrN1llnldyrjglBK
BUnHWe7W7dFT6GvarPhOvgdONYsCsLiVmlQTp+2S3lDs+ZY5+MG+kV5cyB5Llv3fObGxNx9kwa6/
3ywPSsx5nglk5b6J6DV31+k9ft7NTy/8WXhy0UTyRORPo5CqECACyYt71bF/awL452LmPig8ZI9d
0TaedUCe1F5JBaQWPomfkE1rhD4KZRxo5r7z8Y9iz6WvVY2HoS1cXUxiOfi+adreyvvjCeZNlGl1
16ub7XRc61bWLtaI7+S66X/+yR6vtfl35Q06+3i6J7il6nIKfcvkhA5aVxQxcADa1nkXBHdRJk+/
x99oOTCh+S1n1rbnl0BNehzQjoIzB1zDBOGLN8sjUGP4W+haG0ubDxAFhOql35QikdTh0/UXWV3g
EQMpN1JcAKGEz0WpdivA/JJRu5dQJvQOedYxJ6JqbmcYkPg7l2U4iqMMoLkBL1geXjPeirLVCI6e
1aoPhBBfDOgTzc2jDufFNItiOrW60Cw1WSMDpNjSSNzfsRMczjRTRdVaKs6rekduVe7U0wDq2R91
M6qwcIgsPEaR4F2byY7JW/sXZPaSlNSYWJvWpIGEl1XQcFchDl8FtABvol7+C7c7tQRGFCMIK1fJ
QOrieGabluAYYYGJJKl0LAvjtkaAWyFjgUPz4kAfjM23IpE0ck2apCNIxIdh0ovPwdAtDIQtzevY
UzbnxHKEil5Qffrh+ml53MW0U5omuKLE3g/mzinw8FuS8YfxmFj9DpiVncabRyXVhOI1t/TMHY3E
EtYSUzd3LEScGPpHVYGel349JiyqJAuzfWZZdiyxQpr6UNw8oYps15UFaKrWYj8LHy90qTwtaSai
uvz+s9eIKV9tv6lw5C2AoViOIwgy4gdUV+TmMuf/w4h2V+qRIRRkFNgEpMKnDYm7M1jXb7S+n0cj
PCWW3yWp92x6hWO5NOsQxLr6Ir+L6/er6DDuJGlnIujHUixNaeh+wHA+FLNwaLJ5Oq4IT8RTRbhG
TCYGkXzVOrPF0muuX83kNDwkGurCEGzqxm0xRIPrvlc/mEj8+uKcm4wnfwRm+0daWUq3lwQnP0cQ
3DbZbL0IXegWSsodb9Y7Avbqb7b6/H+HBxeu3XN5iDOqwx/hiZIS7q0MzF81XfQz1xwm7nymQtFa
f+NaCBfj+wriRlk8knQoIoLPpuRFET2dLMFD2iMZkwEh5MeX0MqU8xC8mf8zfiCfuGyC90Dtb+sx
nEvHvvYjugmdUP8Eqc4Ho5ELriE0OYWWCi+DBgr0JLZPHKTEcqIs+pp87EnvUFDWmCELJ4FqzmNf
8m2YvY/pPWNGNzt/j7r3vA5kEwkfLs/Qr1dVfBAQPhl5K4dYej5xB26nSV6W3lRcTzYlFyaUtBeK
ACwFDY+Ibuyn/NonLKscXDs0ezj3m6onZVjRHSlcU1zHWbrCrpGlQMJ36acovwI1qD60BgqXWtlQ
iu7LuBOa/q8VRrnaSPjIlyaZxITSr4nwZo3My+Zqo+rzJm0O/unOVZ7Bk8wS9iu+b2447DCq0IfJ
m++2NdZqPBq90DaDsEWrQYYOus3bovXh+edZOlsNL2oKAgxaOHqE7THWEA/QG4myNSo+C5Nl1Uzd
QeRD2SrHX4wJbDBuFyGKK0+XG5+IJWCahq1AM49c0kr+gCHxf3Jw1fNQUwHNSZcc9lLgUYDjsV3Y
S99dH1O2G9UBtV2vP232h3vZ3txlkUESRMK460v5wslR5tuGFy6AeN86D/VmNhepQy85QPeZefJ4
yqgzmiCN2Iu6sMzFcMVGaluh86U1PGJs2g2tBZnBWhBB7ruCmWCqHTg8xS/D6akPvsIEtAyrYScz
muGa1KvSCaEfs0JErpDl9OlqjGGjHm1BNR+HIcL2mQemorgMpLE75g70w3go8fqSwbjaKPSiktnX
Y2dZ6NTu8dVB8eE9q0FRfiaomtptGD6dM6iB3/DjV6tyaEw5wJPCEG5P0dNzE7oC3ioR1bSpCJUi
GntXkw5sN0TLf+A3tU7dmlb4UUacYqdB+c7otJXeh/sUNBqLLGHIeRuKHL6rVIbbFEPamAq0RmED
pElMs+jX/aorFsg6UtUdolJP+sglyHdhFgaQLRyqI0VMeXLV8PgPkdMSSWrkx6YYMa4loCeRGG2c
RwynteM8SJXn6xmJxzU6E1kt/zwv4UMzt1vn+uvlz/5LBorKN8Uf5w3e7XPngHyHC/G8jJeeeVXV
+uNIruiGHhlpiOInH5ufBWDE1zlcHeG6KrEAfNUi/pIxhrr5b+wx9jXZ5zLk4bERwWXJ4SNjIvY5
dV7I7tJ6F2xIy/vqHgGt7i/29fCE9fhqFrnaq+/kdPKoB+1kZnWhpLOUWziBcxRDWWtRnkydS5AL
N54BNqYzpfBM5/6sdUoHdb9hle8kZjHiS06HGGmXbFCLhW1EZSslq35vZXO0W5SuaHzrUFXl0kYM
OtV2Wsay7av3qwgkrJho0v6KGUoHvWT4p1aV67yYbE48wgf/p64iv4YfSXDdFlqD1F8om2q3bECR
M9iQy3NKA4kvK6jNQ9AnBlXbg3F6crb5l+3sGGwKphvMnUbeYcNhOkApANgLUTDp8pylbOycKcfL
VYcPtI+4VrCR6lMLhNrozdXYqMkdlxPx9LzQJAi1sUt5b3J/q/JlW9wX6Cs3/RtOeGpunIYdnSLA
BrwtVyEuzT/4bQp9WpC1K+6Ka+0QlMVTGh7CJIq3JVeZMuI9s+4wswAF9vCU3Nh1gqihwZqULMjO
fOoo7nr9xSo27AKjTx74dqaJc/PlzH3TpkAhLRzjAKIm+2t6l8P02YP1mIkkiuMho8kkNJo3m3Gs
Mj7hSYG+xXmTHw/3zPeFkPSb3wF/+7FWjDnM2wIPKT42wBxG8s/58+rIPH6cEc6/PspOC9llEy6r
L+ZTXYifjkHX4+dnucxxvRr9dBkzBAFYJFRHrBJipCtdZk8uLr+n3/FWD8aVWb/DJsm0QiFmi6wo
XHvk+nlSSA3IVxKqKy9IQq4S6NRsRUYw799DiDj7cI5140rpI/GGKt6whQi9JoHPvpr0veHdsMbw
ni5AwlU27r4sGP0TRWShJ2XZBrbZm80oVFkkTTlnNXVK/ZwWpMxcjZGMXXGL5LH34gFeeISl/CBy
kr6gA2GvZT1+c7KllqMdwjlnhez43d/wa6KfKGc7fxmqRIgX5EXoBhzwH0NwJFyoUC+x6Buc8nwc
kQR9bpAU5gUOk3linsP3+bw3/HsFVcmgTvRmgC2L/2HDXEJfZaw5iGphfN9fdBeRYLxX7fLAanmr
HPsdrlVt0ixiac9r8IsDYK9BHyQ86vi3rM+vs2ypFT7mnqqUDImfCp4BXb2SRdSH+5eCKUTPbaKy
pml5VyF9pZ7PD1ObnOqqkQMh6GqLZNuG4jH0aSYh6ekMAfCF9w+9h8TAUSFK/AntJqxfAvw/n/UR
vnbv1iwkIxTMxWr2BgJ4reEUt/C3VE/69O8VIDuau7bA7yzZlX60Da/tMRUlN4LZyQpqGHWnMUnY
fyRfnKc7fONFY0fE9MnGLR0TqxEgJgPmUQ5NVk8HdxZsrTcUXaq/62pXRNBRXzufshWz+UcruZfy
ls8807zaYcf5jmJDx/0h3yONvUAtKKr9rvI6hDRqMc2ZQHWgHg5k65CpHVytu0pJFy3mpT96I84y
Ts55j0YGSB/2wF+RONBfbp3P78POJTMjlYVfU+kQ+kiRZ+e/H21AZbmROPUxQDAUUPjECN2SFuZK
GEKPtzd1awAI0y+zcRqaOXvjysQ3UwfkEv5yvpQxmUOqePnvz+Za7AgCGa8kvIVgVwRUSUZe55LN
Nk/r33qFLXkj13O6ppXs1acF48lV4n+nWSJhbvZ/5PunWTZFJBWqsVhRwxDRMpsMAP5z3GowZyGV
tmiSaWKL5oXbt9KDdbcUTTMdL5WqA0sQZZgDbUrEbAq9h7VOCX9btNuoTKaijSfipQjzwhPpQvBz
xrhLPhAV0on8HINZcbwbeZZhiH8cbQELVafPUD8K+IMvfYmDYo3fHhCpLu9UHq0woGfPhIFOraeo
3tUMKBsEEQN3UJOqw25MgE6E7uNetjdsFS3RIUTK37hwV23I1SJxVJ/OAafQyF9KcTmjEy0ZAFSf
HCpGVp9FpWnLj7c4i8gKF3ZAbT/yNPT3G0Vvdh8k7HZkCIWI28p7IzZoQNFIDYi3nj6i/7x6zaea
2x7EDSumMzql9jC9HMX9euRnBTVt8NUOKESLr/4QNxTUaHI6SH4o2DJ2Ilh23T4BvZQb/fmdna/v
aIQFQhdhmWPNm5NZntAc4+3bfH1UEqnGgkTdd8uYapET1JPsDvy+q3QHiNM9xIv+mCSOQuoBbqBL
s2I1OM0MvCAdQ3HFObLcwUXJNVYRWQ17brFbUyeGOot9vVxPLis1WoV+mnzTPtaY6ZlHm2rlYMb8
ZpmeFKBuIIO4zjx8228/deyBTF7kzXUa3s4P1HDOFXMB4BjfcoG0HD+qC1vvQySAzQS6qm6Bzy99
VYqmU4tl5x7ric6PkPfkUH7EgFVFdNc1fqbhAK7BDpe70iglIVHpsW+OEU4YSQfao3SIPLlXaOU8
gvJwwDxZx4qmfqog/cxe2eN9nP6AvFUGO11kNi6uHmljeTeHy54nWCoRFaC0GsX6/oaFc0Vzq/r8
wlyz17FHDV2HCSNZnaKSLB9UQ34l/UcyEXN2JUMcZq68E822Jw+d/oIG0NpTOnXCJZIs482AB9Wt
NSMPo5UXl5WVlfB+VJzsmXnNXis9T6E+3jKqltNA+4qr2ZHUMt1paTU/uEV0Qf1UMF79rxFIXTzL
RtVIwaPNV0jKLHhdPAA5yYQINfFLBAc11ffheU+XXao2Cl3TJbH8goNcyfnetNLlVtwHD/3H+I+R
3FSV2EgOaKYIEhozEJqeO4xkbwKyQEq52cnBgoO91J6Ps4vokMgW37aOQyqgbuEPubCTwOKhEBlj
x2IH07pZPUO9FvF2vY/h+8P6NXMTQFWdvNGgHuzZRUaCxmjH8BN+Ujr5CUsz63T2I+zjNBfQRTRu
JUd53C3Wsz60PEKQk4fh5MP9SfCb7jEuxEM62d7iikA5m3UgIxNIStkqngXbKCtlUqHbwxGEKFoL
K9zACYeh7t8k65aqgsWfOhqKOA5FAc9w0mnQf0AbhVjFuga0CL4c+NosDXzOWKQLn4L/84xwzQlU
wNSKHGKHI2YM3PvXTU1LRUuTs01GZUVFYVHriGlKrPzKNPd+PQG9VPG7hbKSyEYPdnWyFNf7Mcpo
u+MDZPCYM0R0gH2pBb9Fat1Z6YdgxkHtpzZATckDbaOuxWOE8ug0TBCd6kqHTmll/ZqqRvG8LnkE
Gk5WUfce3FXQGMlS+9z3iCTlkjkRY44vlui7YjEjW4JbzKycQlEvXuhjyLBDZDiHzu3AE7oX9b2o
uXEjKcN+qflmnLa/pG6CCipB0rPHkM9Nmi0X2ETSR+U4fhhmp6LjxPKoLGBHXqsxWQBEz8Z38uxn
wiImz4ts3tS9d3VHhAcj/GMtS3hj5RU+JwIfpQNg2p5Smh3hX48w8BX4EHBjcdlbn6W0D/WZJLRW
LYhgVuik+HW2UvMcYJh8lIGy2S5EtxIdCnssO9Se5syvmM1XNRAZ267HMWtNbpQleYZdSubF7pI5
AWrBV+9DBpOTtICmK5HGB8JXCn6RoXZXpt69OvZuyQlrIers8BGPzmogFZK2xtuTvOs1rRiWtLXs
UATAdzbsgf617AdwzqB/bHCZR/8I3kKUOnD0FncysX9FYc4TOpR0z9D8JpUrYF9yb0kj76Z0R2LV
TdnvQRaWleldCODiJ7UPJZp5Y3pWZ7s0vsZ1FSUDOZ0HwNb6P01z18jhd69eCfVwHAybbQNB4+5K
oYM4gyapoIxn+3YdZiKz8ZWUNYJ9qL0p9jo97j9RF5GvqaseCDacjypCqKHqo7HMmdV1P72Aw0oy
dRYpH9d2rU2TyIUfXXDmnc1GxIxF8PQ0yhCU40RwHVAiyWwzcTj8J6vtsSIPunqm6OlHvizbMYBv
WRBWG6Yeogvu7N6At1FvQqPu2ARH/a3by0rxW0PNELKGKQcyh3Iec2dIxUTDqYtztB//R7pMPcKo
+XUY6kH67Rg928uyrun7XGzS6WzjWDi6Qp+0iTTAms+Zj9gIbWDB85eldaMx842MyML8gxy4oQEN
M6mkXrWqaUN5cacuj2bN6vp8dTeK4WwKYwYg3ZGIBuHN12kj41gG1KTXpfmIIetsze9StU+KcmTD
7sAba3U+lLjVoUfI4JixaIN8WFh6meDlSEOk9V+UdiYg2ms7DmrKjI/sZzXxyASEvPmJyFoU3f4y
znvtrKDpszlC1Eeb80+hfnVS9IV+ozwJ9r1mrUkPiganTq99i+wNxI6VmT+fqUB3SFzomg3j6pAw
pTDKJO934+otAZNgvsHXzx+sny2J/FxGHXQ6ifTY+LyBwTeL+3F7YeAHSHFZRoajagQKM6ct3ac5
h3lIsKmx3qy1L6S0SkdMFVMST4MMq7k7CTW6OqIhzZgMIj/UfFgOhOzR8UF8AQDT2KZ/f91GAC1N
9Ev6kSKoA5ldys/VNcV66rCfz9OJ2gKYQHdhMi7WuJWIsPuN12deyVLvvXxf69xZVaCfLqIvCg0t
Y55+12HZ8yHYhJdFlWaq7S7tywQ++E436oNZOmWBFZ27lgS2vIYwiKGzgjMJxMdRIxzzSDR9Vy+0
fEmUL+Z1oF4LoGtdki0FsMgGK14o4RBILotNdforrydD3H4YVtXl38LKcRfLQ1xG86p9kKDedfzL
SIBS/5AyiVzNSeWdnke8n+xEaAZ8HnozUesH0NoOwd8WJAQGnjYB9bFCALB+WST4lHhxshXltB7V
pTcCnbEhcAeLdVlgWVMHuaCjIICkEOP+LnxrGbTOt9dAOCuTx3JMtO/FybblakxU3vXr3W+xo/rU
mg92ZsNMxKcJvF0Nj40VKcjrSe+Biks5L/YX+ow53c1ROryP7XOxii6i5NTnm5L4wirmRtqGYLZ1
QOUJR6NaKSfIrB1k3r+v7MvFlW47LdgnFR/Te+2bgyfbPOO07eTUz1QvsyhLoddPJv77dSBNE+lR
mhjiJf8orAf5Sz8SMsAJ5viFhhoZH8iT20l3OFS8SjekXZv3+Jn+8IB3YgCW2AwPz8JBm0D9Uf+1
xlwkjX5mEIZZNzEXiix16l92cHH51eWX3cGt8YDyzNOnF+SHgraA4tu15jzrhLeueZ/r04hqSmFH
5xm84nAoXk6kb3/zYZEgp5wN39rw4SgjJ0B//ut3jXk/iAWzf9tr8T4wrZGgSnEu33dvQMZstPR0
RcE+JCkoOVzMOMSJkLMVau/r5v9Y9Bu459wPzNRmjJK7PdG3EK3spFeDOk25/oJqgiRz4ncw8A2u
uj8KVzeklU5Q9FSFciDLOFmRqnkKdn/pgRxOJERyGcdOUmWv4rqQSb/KBW494UYGj1tmtKAJz7dd
5OkRJhmmHR+qIjFvbxnj4QRw/LC8q8gkA9KdoeEL6ZiP3wu3couEoF49ncn5EXi0NH2UkUs5sz29
0/mtftFfH/lrB+7BjYcnmgw/3GDkrWCTS6IiISSxEp+oS2HG879yGVl+8j/xIjLZHTxY8ijt1Ivh
PNsjAoFZ8gycEfBh+4HlWRDEJAUsN4dohQJP3bA2pdjpbhK8/zsGVk9BYoARX33C/SLfYjXSkAIp
lNSYxw3beJeWCr8C5543IfEDrbh+z8lY4Mtv6gTQvwFNLnu45nUa3Ywh1bUwgvf2hSgX4nSY1hfs
Sc5ceVi2GMxODRnEH1ungKQQrbbpZs604oJjcpn068BI/cbFC62Z1LQ9X/vMNlksNT8F/BlG1Aa1
59qDaAZUZ5CLfyqY+n410GsJAgSdmv/6Zj8+lg8B3hg9nrT1RWW0+IGic9I/Ny3y/RQc+rqC2l2L
ybKrs6ZlCThvGnfzr2EaNJOEPmx2+qMjY4UUIUOWhJyiMRXcG/Jrtu2lcMS/Sg68wqE0rEXjdebm
ETz7REpxPxTx0XzivvrEH+SAN2VnTj7KICBfo1HmWWC3TDaDTXszUjRboPx2YW28p5BRa2gMESG1
Fp+D60+oi5/K8J+dY96JzIALZBRn+l6vrGezHKcNvFLV6c/et6Mg8Ll3Jv5gFuMNPbEAvWVJy38E
n58lAm0bO7YeTQyAP4Nzln+womoyAI/57Y/9RPZNX7j8zGfgpr9DRiNr1FHfJfFeROJD+rstn1lW
XLB5fWW6v+KROlahTU3fq2FW7mv2rw4kIIn4Fw+x4vOsVE/UwOWHnRCxadyWL8OLUxFX6YSp7/No
sNg5+OaS/sE4QCr1L/tGTRQCHZnYfVqdGro+0k2GrskEkZQ33NtOwyyKbbes6h13wu7+JObqQf1F
AYvks/QhtHjJRKKrQ0XiOo7AUj5QEzdB6CeP0z/ogej7wHPwLHJ6+kMeTD7r8Bp7WPBPq2oqrzdK
iQoTjnr8ef/VFGTe54d58ckK+PfU1itMK+rDy2i24Ph25+w98vJ0pvb6Qq1BQHiCWgTzej3RPR5Z
TMYdfO89EgaEA1510vd2mwzu72s+Kp8rFRovUKQMDndFBrSpecXsbbAJubbwlZbz6skFRSWFMr/P
LAU5MdLxvyfbex/OzKtewTaHi2yoluVSgjvdRofDm/l34X/TXHXQxCYiktRhIDQXg2zn0HSYIF9l
RMVu/EHqUDDwn7L7ELSzURc3sCSgZMoYbreofoTZYEgNm7Gsubliw9/idLvJu/a8hDG7Ib90NFl1
jMWohc/2kaBgvda2rdhcwJuwsbVYrSCTdOChIt47hK6KIB1xzxd5fBX1m7G9JQVKY6NtvXv9H+Ck
0hdXuinjYeDhZskoySEB9wmlMdvI9W5ifMiWJ3OqzgUaojJWsGj2ua+ekucVrjz5GZSoJQj3djaO
IKWpQgB7qn62LzqwRKevWsUGBCCTyn8vB+uFFweb2SupM3QjFUywCOccYqPRN+VpdDeqSk3AJZ6d
l8V1UQcvQziPzh9nDDlsBvKyxOeKVJkWtikPNHOSI9W5Oe7gndH5bvA/Ew3lP5C98wJzSe7KT1He
F+rELL9ujbHSD/Dky/LykVhS2DG7aSfN3nFdAEViJ0Hio64GczhHJ+o2bfSZqVRXySZ0H9PwWM97
1ELFF0Mp17GQx3HWVljnXOwM4YUkF4VcjKAfVRqh4V4byjL/Da6ENemvl0DqIRa3hQHkYkiFnxk9
omab01WdIR6TmYuvpr3T73L2wCM2o9ChM3Kt0C1+yALhjbfbD4qvqE7HSV3lU3YujOxEyXvQyS9V
pUG3ipzZXsao0sAVoohDdP1bczpJbfPr1UvMZoLDnJ9vbuymot6D9Xq8Oq08Mklff9EplbSplSS5
xsMkDdmX0fv0S7gX5OvMoK0WMFI72/yDlIwaWjrMa2UA/dn4nNj0IQ5jSdgabS+uvzXY3qRlw/LJ
btVa9DkdEiBvBOPCFr/31Nc/ZiPagLJxnUGw+RtE7lxEDSlc6GdgjwI8nh/VhhX+4YwGAJPdnB93
BiatHZ0PvIkZrY0Bz0U74Tpkwu5CRzM6wayfskX/fY/5oq+MuY9SZngHKiJGvdxqb3BDSF575Ve3
NArebIWjq4m7yufwhA72Pk896q4pI7sY3TcV8lnazTRrE/mrmSAlAKaZfuTcvu0foZ28u4gV9Ev6
Zt5a37Ql6MQX0BkWfksX3X81XrDVys6m6O7MCOElSDSSJRZ+WleXDC8T12p8kmwIo+i0lautyBeP
Urbvjlzs2MzMe5hKuo9E89GSnB7NPGb6FWGSuhvkliFHp4iXK3b+DW+0J4GdGmRoiMN/4xuRcR/f
noQQTpFQxGgG+faZN2DWScdkyJ282S4LHYQc6OP7JXPqP0SnaDiLdQyiOufht6Nz5GfnmKUpjx8g
CEqbO/63LaWl2j7a0DYIBNnxbhfa24JhLypQ3t87MN4kNEzEtzfKWd2Z8A5YftE3cLU6L5+L7U46
I9Q9WL396xDSh9zs50zfsVo93pbJHao2Hk1z2Us/Mj48Ui2VlPXi9+cmSgcpv43EtzzCzXsJNmb0
PL7HKM92BA/OIeNAdAGE5JaNsTrEGVd5k0FKU11zAmuXkNpq/rMcJRKw8X/GKEZsgKswdyRwCO6T
mKzYmUacPMst7YNtEDkoimJ5lPbRaH6bL+13BenyuoKdUpSSyKCtYtpg/G9BStHcJwcyrbdpA9Ox
VJ0adcDN1kkn8tROeVvqR71vEpkeMovrKmHsDBkkDxOzblL0IYV3rIyDC6ThPsSzNraN5DNGUIXg
Z/rac23tiWw5bmTe3UAjpKTOkiqCWS8oFfYhs0o3Yyso4UEMT7AZ452D7K8gnADBpyr8gVSH9RPu
fkijv1K4ldhe0Tz16jyi4tr4ppcv03NCZfOteH1oOZLZdpJwEsRRfcCMwlOM86TFrzXq3x72TcMF
r/QXEQoUrgnMKoG/j882+GxArUY8IxVkh8H/odK1cELifODhjJVYLf/2NXoAmIPTvG3THBTUXUqZ
+dvqprc3ZlENCsAhg65N+t0TJ/tRI1DNsxaZIhJQ58dGTpmWbBbt1+gJcpLpszRm2QexeavQJC7T
qn+88k8ZCyPfSD+69bXhiNDJdsaqBNsdmjyR4PyXgQTwDpqVqi/aEDyjg1tZ1sqmPFHLaQ9LDAc5
I89jTV4G9MT0RC4rmR4Bg4Dzkrzx2LRfv2nQO2Bb3pQnnOmcSqnbFjjqbjU7jj4Qf6owMe4dS/O0
XEvvAWsMRvuUJvTCNKtDwtHpJ51O9QSqnOXVJxMJLx5cGnZl+97mcI7vLfWzEIJ6fUAqzvQ4K3Ic
XvDwO2aoCYD4iWyDs/R8xqR14PBnRpU1uWAVTBghVGRaDjaIZB+5Etj+MVOjpfPrJIsHB5sQPNIJ
sTnFBvPajlxqtDkYWjTzO2vb9pTswGZu2RfsuKIN4KQaY96ovToBBNtDoXwWExCtjSrL3CgN0GKG
fv8gww5NKz/ZQcunGlfqZIDWA3wPa1vMbpZusj1fAs/kMCi5MiyWpazR5yM9glcvvigFbtLAvB3z
U9lcJ1R346sJoljoHvXr9xx5IRymnVUE31xEOocFQr1HogRzHDOLfjzYoVyePr5IyqeV1gi6UR9z
nBPij0qeVaiVNdtdmG3t18b9GgX9cW8Erxbxgfu1oY6M7FkKmU70eHV6gBZt4YgkpcSJiEz9NVZV
3nWFOxeYIrzBHiGorckj+vwHjJNjphbcOgYWcS8V+ybuJt8XC5eMzWFBZgVm4rtg6TzClOzABtB+
XMNKD3d+UZlvT+KYHDz9DSMVBOKNMfvEWw48xvUtr6ykOtS6Ikyu1bZPkC82d5j09/ieIvZotj4p
LEy+EaNgimYKUeyo6pDw3Mxd9cczAuw1bSWss5Nz4aEhuww7tQsCX6NGOMjXLQ3wzrBObyP/gWYl
2/lYMlKY9fFjJ3oeat2m1lXI388fDbxW8HKQQDgXr7wGQVhucD9iZjAS8w4n/mo4pec5Ow+YIT64
5ghtnBYap/zxD8uwjkqr3lIiie20csXhFTyC6UHbibFIfdhQyKH78+1cLUUqI7W/ewmIEZhC6j2c
AwbwMtLN8WgVTv1c+QVfa0H6NqOy2yXguhpImblX8fvwC1ChNLn8MxYRhQc+4ZmRy2bTw87xFA/V
gS5rCGFV7ZwdTQj1DblQLEJNPj+KaTeIhtPcp0nPEv1ASJmt7jUSsZJtHKwKpFu2EcfdfIZYrprI
Tco0o20p9yHe5xRZumUug3ir1ThIOKmoRNHt9LNKyKdoZjRj5SS73WfHZm2uhRPLKOoCNbZADXYM
+whH6DwQmFgRHS8xUiL4dlJhjVLf3GcEcWGLnL8yrQf5EtMW/SSigSCqSU94KHzQjw1raARDebBB
KaZBcRcPDq9qD4g2T8PG/tdxKj+NAjgM2SI9u8fSVPeCMn4PutKOZo1cFf69CQS7LKgZ/k9MLMIZ
vb7mFZAlXuTmRk+3gCbuBefyDGuBbGxmZ60A4JxxPRvmxLCqOPj29G/p2aCVAW6UsF6Ai+pz9jde
mM6Rge64eMJ5C6XXMEBmlxYkAnkX9aJsUtJuchc44qrA8l9Ci3vHpICXwP9ZstJD0h0BAMDIMDdA
3jyPv0ZVlEJwUjTj7/KePRldWLq5DjklOoTDwqgGxrfSwjfO+Ty92tnyE4hYjrjlg0sqZwc5uxIG
gYyuq4V7f7i73gNLEwJkL+9AjM6oKAKexq5UFrNnD0DDH2r2HzkGfVxU8CMjUYZ6DdpscFxXa+n/
2TGzF+AwDs1OqC1Icrvs+DJlJDN1AS5suTSY1Nkg/3VYQADPMvBbrX6/0fy7/1zrKIF4aMZeTZX0
vw3ZdrUJtzG33wehqfWVj8bIin2dQqdsrulI9fefn2dtSasoEzVdnpulX/36/LjzEZtBsnCAYJ3T
9QvI+trRH5RzgqJEMti4ofmU07xfkcVeCTmn/g38rCpqS6gm3fdrABYhnInXVoqU7TFFp7SslW8J
ezBTMXs6vhriZXc2UjzYowZ2WTtH2Zo2mQdoSyl8NicC7g+xSC/8x8PD8/QT9DkMiijggqSUU9bH
wizPoms/iHJ3Y+qr3VWbSKpcOSr0ctdbP97ZdmJLHaYWiHu1W5lGo0fDD1eNlk2KShAsh2dS+Sjh
SZhWWHZpYl7gOsKDR+APW7yvuqfMdMZObra2PzDlp3Oq+liOvDThE9Bg3aMxESqvm7dlRRTlYVdC
z5HBK/C5KXQ13p+39fmT5I2ICpnrQNnGLgDcFTStNIYhSgH01PpUexZZIgBYC2eoeKz1qWoxZA1z
a8yc2TP020PduLtTOvXpJNUIUsbIEx4Jn8cPDEp562+zUjg/a6MeknVRwNblx/8tVLkH3CU0f+hj
SXhd6cpuuY7dBgdABIP78BQ7w2PMfhXPQE+32vpBRZaL04yGIUu973rO0vbdHF2fgeFBWm93lzSZ
ruJUmxj4v/HK/3ze+SZvh7J2c+6/jqW5ckIv4iW312owwM2NCTl0yMshD/6j4lWnHCa9hFiKg3/Q
uMIeyRUSSrXJHrnDzJVNjbbvdgUV3yREfVCL3JLkRwRK49s/xgVJbkzUkCEAdOe9XjbY2dtvJtcv
djx8UrUYS6KmkeytHCLQ3iWREgKkg7N3XCk6xaLQZV/US84xEVYXHiq0IAEHOxufDijDWtw5dS9E
4yx4FP3rWhlAa6t3zwyNbZrJN7Tx3QB0EuU5TQybrUeu9UC2qDaQAGKiUyrROqgoWaneWNZJGgxD
wTiNK+MzKDN0SXR5BYSa44qAQjCzQ0U0/L4SSczjPu1XERu1Mqw6ucbUwBdKZ3K1Ts6PEh+Iyyaa
dlRY8NChSLh8BW6K/ua4KmbVKEuhTdDc2lqgdKsn8s6RNdPY7OowKjWlkSOXB/+FK8t6Uzfk2Nml
BuwWPDGaRf2gjAJ09le98IBOwj7m8ZNsDjwuWwGTmvv4L3zRNlFv+vuCuVYtQ7aZJkBntYH8O2iV
BHxPFq84MaxDRj0P+Bc/6ZQ0nuPHwE+9+cIyavYuEs1v9ZNUcBMFxiIRIZsZcVob5a+4u+55nYoP
ugh1HC6xBRxxyuo9/g8d1qbjAvKIiw9ntr4DcBCYTD/57lRFXlB+5L3AfUJe1p2nXIcdYVZQYBgY
wK7Squj1HcgRf2S1Tlk4zE5BLXlD/sMXPZSFo02MrlnQ//EI8GxloC6TDYPi/ZpYqJVhYGRwxqv1
iVhtjSpd5fLv3FFLN2ruB/gLqQW6RKHCsslD7D84zyNPSpfYvpTbOWKnIgifC5ELBs9pQPRHICjM
mn2L9TnseEpZHy9bkZ2RNyND6QTk6fyiYDrQX/krwnBS1C8Xuh88MKMvOEv27BLN+/ofymHkTXbb
uB7f+Fc33rO0gBvAVb+b+kbWJy7bYtEY4qCylNEZ3xUF48UG/wstUz4cVtJd/v+Crwude8jGUOOD
m4HH93myIVtu2oNjNztO+REFijKcwBtuuf7Sehd9lydizxzKXYFUOJ5PmH8ft2jKRXHibCRKHntQ
V7Td9bhi084V/tM+UWGd9HF/HT8dPdEyCzM3MzJQDvYJEpQGvk7QI5svoePSt1RC/r1TVh7u6QJ5
54yRJBn/toboWe8uyyoXhjIKhjpe/qSqjjBMNl6P4irKdWaPkNOunqcjpzen60siCsVBPH7kYZ54
opZe7QD6EvJrGedNq72O9JzeKCOAfWKwUTAPC+FYwOZA/Zz92lgZdBPLrtnDz/ebnL8VAGwqndM4
4o2wZQbYzvLyeLXPWQsmrWLUYnYe0lWj5lx76YGIxpV6Lyq7ENin88dSyOMd1zSOVmQId+Hy9Hbs
Ifsa5Rl/Han8QikJXKQh1tlUhNvrfpMt8g4y4jz2nZp45Uh/WUUcp+LlSoeY5taiFQHusFIKaTj9
0U8poa5NWoUnVXGlUCyO6uq0w3AJSlSlMVUwWlE834hvDusKXNVZaCBK4J+RWfqukxdxq27QWq3/
6OM8XElv2cZFIQRFksXEYbpYGRygxjK5xpMX7Wt9LrEJt/NKvnGLTG44NeYKYviKcbK7rQMGowoO
Fc+h65s6M6w7nUyrQN5Z0VXiikgP2+ay1L66+/58qwKMW6gO1xvQKj67RnLCOVT8426M01rYgGrK
KxsstvY3A4lhVoX+CzPgEAhVO4ooNiT2J4N9Do2M6skoeX/Pq/vlDDdlmgtJev6XlUZaXpdjZDb5
kduAsr1pkJ4avwJXM1Q5gSZKAko8tDuStoomJMFZw6kCMmvzk0FKo3o08GmAAiqJj1U5HtDXDm1n
1dj61ziYVxrOIS7TAUFhBjVDcHXiXyH99AgyPj5EgcGhYjElo+XG9S3wn9Wd/n6cvE2+7Zoa81GV
w2DGRE31l2UFvckH9Tgtp76ljQS0tDOS6GVlq/lTHumJF6kWmeKOkqTu44JhqtzU4liStj3PEAjM
1K/x2djalPA9rTVsmWTLccqvNlQnCeAa1oLc8Iq6c+AkXejqWqlQBbO2ewjXMvqlzitVrsaHzmqi
1tJf3eefAkyc9xsgM3XyQeM2FXaJTut7bhZEUrFrszinRLGDRo6C4Z/Y5j3L/MuhmDIIxLe5BEGe
w6qfMb7K1SlNTkjgM997COOMSDWCk4V+verfoJ7+2QDVJ9Ny0Stg+PHluaU2Ecgkjsa5Lnw1bb+f
FfwgkS17fICddOl7x2QeNdY9NTafDTtK8WpBNabg4t1ldZTy/ZyHyu5nb4byKKstKMsMPIJAk3C5
aT+uWpEWitWQp0DRfM3o0oIMWYWNDSJdkgyp9NRlE/PSJbxzdNLWTSl3mkEE+bqqyl27sxSdgLsG
YO9XCYgbBvn2XeGf7yTFq73LaOLHA6qvQ/frloRG+FlaNS+T9DIWw0rJAEfZUnSTTtESLEk+mD8X
OVZyuKsyDczWX9OyXK3ERa7L3G0mmav5D1kbWsrI4jGn7NcxZVSu1KL0SanjcD/hbYwY4hvTPC4d
4Ebryb8+oOtRsJ8AN74MV1HpPvSfC9uZnGe4I7dXrG30PC1cv4CptYF/XwkWtXBSv2AczkaCt3xf
Py6orG2e22P/1bFTGXpDbc3hJY49nr6t2m39XAZa9cwb5cvk+nerbCAjsXtgzcvnK4bsMfuZVkvw
nn57RAjFmoX7FdcArIk8ahyuluipL25it4Y3KQ6CVM8n0u1cf+oQ5nG9fVuD18JlVJeeDutBQQQ+
yQOWw+qNh5T+yd84YlM98g+gCuPdjcdxV3LA4cRK+aRr82gnVnKv5uQA6XDsTMVM7nItvJoLTpNd
hm2sumpCb3Ho/7r0yPyNDlu8MsAGnMHazWo9fmadXoulQcfJPDNqznjWm1c0JqKeH8jOOJVZImlq
TFFTdc8nOf+iymPRUyrWeOXhSF0rWus/1cCqr8ckG+l/srmRgZuufdQZfq7HXBIESGleCpyATeOn
zY27cRpP0UTkBS7Kqr8E9WLw7GCegRhCfDfEyNCr73YMKpvtA6zdEIvUzQv9qqMJgEAhqMsN7ORe
yayVXbKFHt2d6vwioLY8xmYpbOefVsfxnZt7CTz9LFBFIwG5SPXLyFtBgzVk9YueR7M2BIs1d4Jx
bIJ0RP9W3cCPGJYm0cr9dm+MUa60BaJ1yjfGNoLA/IsvFHPNjKupk29S9FaKcyZ6Co4EwZRovbDh
HiHEik3Fc6iO6ZAkCk4sLNlS++naCN6nxOmniSdS6e4/QgPp8khnLiriIPRHkkpj3EZ46iwmGFhP
ZvbDKf0IWzl0VHB+xXGVQM3EpbKHhhOzPMVftCngbQE4z0pGMkX1PwcdlEofoZGaDOkJM87Ou2QX
fj+L0OVUbqUQbwJZbeF8WvoXOyB89qTu/wDZsi+ePerYXnA/YGBSsVwy4+/fXsqKhHxgwyG+g1Ci
rHDAnJ1VNq9SdRY6oSJcHVBRRahPeQ1GmKMC+85AWGeebV7jbbAB8vRk3gY3hAkeFlofijMe/yLa
Z7XcsVsHLJjowK19EKgNwn8qiLITc7A4PCR1XUM+RMHtOHZomkKYk3zO1zrFnjWTXgnLAzkgbUyE
1ShPmORwJxU2a2JIxvNlTgRGLjMVpXKMd/GzIaUbrJAEER+JhEieYciuYI/ia0+RAaODh9WGJxSV
xF00+nvxONVlpH7505vWmCK4yDEWdbGLWjUazWxhFAqNyYGKeTfKjGyAkhD4ahxzY3KWAiFUoSaw
gsSGVHDKv4Q8lmOkLAmCeqAtwttfQbL2YFskaqPHQULp5BvQoWWFce1Tq23m2TWFxj4ZIkhpXjC4
syt53e2gSTuV4CAmTbM2fW6HSlAeZIR6mDMzkUssWWR+eRWU5nn/Ifg+ZoW4gF6UTLnBbeR90B4z
jUuJmGHTB+sOHdCK2S5A2sRfU7Fv0OLUXbQS09XNM1hVzDTkCi9l1X2RMX8PYT0w2G1y9GyofXRh
0lSOHx18s8DlA7NT/FuSy4SDDkrDOsge/IsDgo+4Fel9VuhYFYzUY9wzcEMRY7ZHDm22qknE+P0v
IsecmS3X1T+3jIG2s3eLJNddFeZOQptCL3FiuGw5nPQyQsduGPGhnm9kViE2n1viv30SMQNSRzJO
JVLvZoCwvOC+8W2Ehi5LZJI7gPUR9ZHa3hvgrKbGaQhwz7Zt36DbnCsXMt1a184v2YtFEV9I75o4
Ybe/4WVSYqj3/8VtP7EGWVYe5xZ5h9GspHdvScAK2sa+nD3FG1VNcq71uagW+R+KIHO6WoF5b8yn
Q88sYGyDUdd23Y10oP1kyd+lo7lrqdXjtAXUjXU1LJFgP5cgB7dE1BGrXre1WU2wmH2ZaRI4/1/g
glVoHWoNiYVdRrUQOl5nZE2EhozmzYkGsHweRRGkD13KCp+chm1/LUpHK+kdYX25KKXWFGOosTg7
rUG6XE7/JEJu2hyoSjH3xkpK+wY/ykshgCTSU1XK7NgeDlqrQrYH11SZXGnOuQFePS8m6m/alAKh
EOadBruP6s6Qss7d+MlQBA5IdBvZwYhRmvVU+sICc0oE03P1k53QzTrf2/7uLkVe7jO3Go4uXkkV
NZz0r+KTcO8bkUBfGpVqSNS/c/bh9TSZbXjV1952d9FezzCGEDvAuQoFkiJamieC6DZs6z4hdOOI
c4STSEk+fYL6QY72+oI/oKb5wGLfqL+D2jvoNNuLT8Xe1QXDOS/a+sdt159w3KyVUYcYmxeccUH2
533pLw0/+XRAZe0x4PIO9h4PgXaByLIji5BB/e1UlFIM6P5pL0nlOh6Jgp4YWNnm2IHNthYezJTX
xyJqyA/eA6TCpeB50r8mnoJg0402coPErMer/cV6rHL3HykVcj+DDM/cnoVkrI2uc2DFX66TBmwI
4XYIN6VeXBLgCT9ROwa8QygP+srn5802diRPU4+zGUEfP6f+TogBzGIogVLgu6XhmBhBKU2gVPxt
m3ipFipH39r0qgr+InrtF+H47otWkhNV0YMyQDHHvUHf+w3RNWbIHAWEmRlw6ye5KxtB02hh0B8G
D2ky3k44VYNOQN8znq4sKE5a6erX3rlYycLS3cTOCQlpMtqg8WeJmJ0MsZfew28IK1VPZ234SsAF
982Q+JE490V3PSdNaK+Z+7ngA0LCUDwjd4K98hdQnroAHdJcgJ9G6NFOgajh3/Z8HBE5GuFncMxj
oGV1zAlXyNQ0Px8g723tqLFLzKY2DTQCFvJl0nYlXyxEJffnxeDiHIiGrvcbt2uJMWQtQhlw2duP
sC3BXaRyR9keK2A67cJH5Pnw0DSiVfr4cEeV4KcfmNmBZOCZ+QOYihnAJk1ywR1Xlma/31/Mfjzc
QPgXI9nBfvNA5L3FRvLo2xok7H2utWKxly1yClf61aGU+ez/YFTJhUm7kS5H+WqxYtKKyxgymSvZ
agH+f1l4/yjAEqgTFzkrxrkIn/QXph2sdROkAOtpVUyzXb8+5tNwFsade9IfgOPCHOgi7Yr8xt2h
OdccHNsrg7ZN4XNW0GQKSwPUnOILrwBVg/hKDVWDKdW05WZko1AlkfSpZ7hnzR2kmFx7jYznWqGh
+0aSeBCU8qQX+IZi9cYZ+2RX4RmxWzPZ886HLxPSLu8Kk7MsB6OTGdAZRq0z+mSZCyAK8JQNx/t8
grsVvNnZD+GbnPwEst9u8/z9qGwlrA5cYlZDxERxp148Jg1e8ihBZCr7ZrO3H3YvNz/8rFprFWy3
zuTgaQ3bbEhsdS7S0OswsVXC6Q81vLMzDgblp2txHlJ/Dtiq8N9swPgl+wVvMTdv6MEaurrgR0tN
03KZTP6YDvHgNqJMXLHVF0B2qKhEd/AqNKForHiDDUGYw0ViXXPlVqbQ8YeunLuYXLgWVTDYboV9
SHSS/Eb8mWpvZTOV9Dl2EODr7AFSNYCk0QjEmuTvy8Ujvz+M7ChAma6elSqP4B5+002fGm9eI2jj
HDu2D6ZgxIxH2Oy1ZFmqvRbDGGAVQLfXCtcE1dcz7pyyYYCOF03a+24i7G5VGIkP4KLghm5FWjnY
KxIZwBqRCKcF/carmXg5Evv2OyXNlgq9fZgJYn0OGEb5HO1VFMger+SSdhlgx9zTewusdWBXS+Rm
UXMNwhL4+UIaD2drrxu6u06jkE3j5pINIvoW63II5Go3PQIaZeuXb/Ov90Exa1bkzSublT81x0dg
ofxR2n69eq2yi66RUuTYOd/eofjJK4v5WWEgLN6c3r3q+YNwdqmjguBUzki8Sf1SCq/ZzHPOwVp3
KaTnYHfwQHeTuDZ9mVqZGvAgfG7MQYH087Ek/RbDNDtQo1gdgxcZfwMhRrMm9Sowcpu15bAMpzBH
UP0f90tQ33G4Bc6LxwjJFt1/ivzU/5A76By3Awe1xKnUb6H+kzg2b7EC9l9WuRwZliB8EDZyQNXo
B0isoNsAFLX8fiTbhx4KJ+m4Y0DPe83qrm1pCoVA3jNeoRik0ZqlIeq/T5z0HVo/Ai5MbdJvZ5fB
4yhNLZV0dN9WQs0EFpiohItAgmfXBQSfHVXh6682P+j0zkI5xy7oe6Y3Efx+kaj05SeeTsBMZ7Ik
Br+7VIByqTmGJMZtMb1lpgZD+DyrOc3/dckKe7E36s0JLwYsTteAAHMRunIxNkWz+mf4OcLC1jrt
7ey4GhCKO5PloHLN1M78lphz3U9+FyDxFRipbTPG+QYVPCOYttfjx5ssfU4JbYk5rzaNnVX5+cgn
MYdms4fo5AfhikbRS/TlnoJy2gabKRYi1Ky38f568dBQGfb6YXttzE5AwDvwGf6QxV5xggAzjrun
XKb/dPvqktUMIMz4E4Byra56khMDBMpr19bcyst+DCjR6ezE8chLjk3PWzk8OddFUm84nID7fJgs
JJ1jMk1QKqkXXp1/UDcJBsq08k5K+IpiMzL02YoQlFMgb4Ruj2qmvtQQ36tCLf99rLEMlnua9xxP
BjIJ6C8CSV3IA1b5GjspZ/myodtukcODgShr7yRuFIbWSjWbDu34j8O8g3b6KDZRmeozqQnykziF
hwxO4G7EtG3YojE6khZRlKl+pq8wn8Im2WT757rbwCjYz21DdH9pASBbvaCNdDedRBwX3aCKY6ia
/Qr5am9FpOA/PKdZ7VXgUA8oFevmrMljyj83uETP2q7d5QLzrfHHWEzvY/vv7/fcfGtANqei4h/6
8CQzuIfYg8xiGpNAJDNLHpU4swLMWu3LB1bgZLmbHpQ0qVxjrlb5GgqaG3+ZpFZPYSm6w7iq9OqI
ImkuM9WeLtDrM7l0KROb5jKLsxY4I3mcb86En3I/9sLogT6uE5nLnZEf7pzLDV/qg82acm1HH9P2
QOiBhGqdVpYRONnyVjxU++aQeHn/NNJSP+S/XDxg7oWAgSmmXjnmZ/dNb8xVOl4i/AL5o6l1H/Md
B7GCAsVjMtgSyQMcS+2xLqFP35GSq/6qZK9q5kLkCA21456n50l3HskOXLvXZaQ/Gkt3Kr/8LqfW
gww9DAr0GpWMGyr85DP01FQsrJSPp/X3ATKceJ+bw61vc6948wI0TbSL58ht8frzVoNFdjOgsfQw
0bzQ9LcB5pNDcqFoeMjgguJ56R9QPe41nN4xXeZ1arM21Vk4zt4ELhDV27vTVRA02fUB/znXTkgm
k83iKZXevAvK/FIL0T8OHkPnmEf+nBhuL7ZLhTiWo/YfSydlY7L/Oa64vEABa4/Aqbb+IIjUKKa6
9ShOvtOxaTh0jm9KItT5kiLWIJnHWbM3ibxp3ZoGZPFCi38cw3vCV8aNT79UdarBguPLrD97ZzY4
o+K7REi7s/9B2BJtw58L92gWMaNRhdTQxOtJ7soe8VCC5IKtNJ4ZAjSUe1bF+v+6icuDaK1Zwuo8
g2Bcw+wy3ElZ8tWO6w4GYJ/HUWpS/h8zdX8ZcMuJmlW7RnwKCeq3JNMTz5U5PJDmGxv2vowAl33G
fY3B6lpvvzoeAN8XSx/3A+CvPQuU+5qsGz8yrsowhW18tdr+A9yV5s7AaNt4a3cUoVSKtTERAOXS
bXEj+XtHrwDpotlYyfYLRTg6bjLOHO47vNyya4Va2KyEUh5vJlsNa/pUoCAjKF3VFwwfOZH+WHaC
Vu1GhBvFMnbJDup7xmDqFhYB20YSNWBPRfDEqDBAq54Kbhd7tx96MSHAJXV0kA/3NQUogxygMDpC
TGUAOQvk7N7aakOUihjnuDzuKkDEkPSWypPBD96Y3kYGwsKMCMsJMuI9mLICZB89ee/8gz2s9wd9
uvV3bzjkViRFF5ZyAhAz/iIcZeAkyaAqFM3ZcyZNtE/KE4y0IawRummYufwk8en49sXlc551rHzY
oBa4XLrdqEIuv+ewkfQVPqck1Xc5X2k8xnd93Nxc645F5YDJkX77qE8M8pFv2jB6OKhDWOcIti2d
ltww4KZEvAqJgRcVlPnlVJTMtF1yOGv4iFFuFqio/N0VH35EHWdvYDWdTPKwnyKdwunKDjdQ1nBv
2csWGhXVeVk23zbYcRusSKCJGwj/Z0iGixTELZeRGeNWm3Bb4fOCDYBlc8YUvli0Rqfo/E9Fr7Yj
dVVPLpiGr0xTfCw16J8iDL8zAndodTgGOvpkvSIgtzSZU88A6iBy1SsYXQLKsP59WVGlvCKDYmBD
5Fs9+TOcwwg8YPoGB6HzQ/KAtHOYIRcc76NPrk6b0u6fZpxgv8fTUTjF1Z6JmVFpYJMXciYkuWkT
ATYhwxQtooP2lLzVdWiefPxJN4PFDiZnp3N3s6MXLki5J32c4Up6LNfjYUjjgiJKY9rKFyFZmPKo
1B0u9vD5PEDJ6d3CVqGsBUPlyHbBrALj1Ae4Gvwwe2JN8NInupFgMUxudeENXGShfuONdGxoc/kn
spZi5rO3qWhBXmgKOm4HN0miCdI7oHibpFTms4FGk/LIv9keqc6kIRlUcd3H85HIv1420S/SBvZ5
1Q0lRHMNMLM15k5Gqwg0qN7BlYh0DuSZDxou+2bKqAu+msFb0hh3o/PWLgSJgGlHDDMNP70jSoa3
VD/IhaKCbkvtsXYvjhjf18IPm14cIucTEIjN+do2K5AoP2NYH2Y3/XvOTyX5U8UHH2OKULDdFFAZ
gWOh6VNBWRwBFG6x3Y+xZN4RHJ9AbDcUe8HGQCOo9KVrbaqoGpdDdn4OV2sYYNFj7WP4SrAxzVOv
hQFLJvMOSTJsAwHAIQthU310G1ZP8j91iHHPb2+mqy6MrCnWRURoyUg4fsHXkO/tt1D6rar8747f
Jmyib0dTebxrqk42J7Fcowq95zWExEfoIXvVzH8miXsoKnQo3rzm6emMQYmzfKlHcz3wx0CNjMBZ
NNGs1VX17Zj9azaL33VJKKUZ35rYNLb6CMHN1me8o9HExPTZv7Y+2313DkdMPMeAQ3U8O526d8sK
sCfWZsggESLXKbseXDTI+4hzc3GgDtgHsJNIztYGCEcagijoGaY0VDz4ZD3KKhb4f5fpC7E0aKYm
rxwukCK5omWMSMFqCRBHV6aXS3OCa5HGw5ZCf2LgjG7Aj6/lRu+tyUv1MUMf4ddcK5+fxG2B1wfo
LJqoCJ6jOAPg/k0OhaC3q+tpzUmYd+kz4s1rcpNyahoCNG1jSdZiu2WKjK85jj+ZTHIgL0r6klCV
uov5+yBRSh38bkxOwKbptrvQ1SMJ8qIRmwgVsT3ZZhpKm+uXmt18/Mx1cIQJc1Resuy1xo24dgtX
i2LdjB1HR1EvmeTrleiLdNV3TPzpcSRAosros9dbslyI3WBgW21Verw3zSqfCDzSZ/6xR8D9+VHG
aNVuRUmqg9etKa663VkiB2jU88N2lV8wgHTvoNKYCsQ7neCC/h313jvsIWvDzRpq1JXW6eIuH3o3
gYNWu+WSqMTaxcUy2sHm05UJwsc1CM6xRi7gcHZGuUHiFuzQ7Y8POpzT7OcSn/oaAE0wZneEMsmA
kSh56gfWINcAHTj3dsqasokcRdRC6xQNRba5WvycNE/0xmW2lJwC1RC5O994OYNnW6x+1CUP0H//
a+pdgLHWjo0cEnFYrwvEpztxwr2NKf7E2jsqgtguAFoCUvuORcztf6Qw+e71LP/cSvNRIdmpFgAv
MihFyjf57n0/p2zSW1wUzhdBQMzNdGyI5L0lQ2HXuzZL27eR0pHo0/ITQkwcijc2+N5PVBylSDAi
i2M5Grzzewmsf822w08MeThy5rpzagJiX0eXtzvTBroExh36fnLAEtPZt3rM0zs6drBMB8qk98YO
al1pMwwZ9RDNR0+bu4kv/A8J0Mev946LtpNYWy0iRqaCriUPA8gutJeujp1gMDrTdMZLnx8jt7+m
4UQEKA30ojGR6rXNOXRx1/14E0p/USXWcHqDAsQzaf1rd4Ai0VST6pZnmObY1KiOLf2Zo8ZvcTfH
Z17XEmu5De0iNQ6I8FwY9rd/PMHhrPylXRc1ZRqokaXeA/+9iYs06zhFdfN5Gi+J8SkGQDFTOjmj
C+yBwsiZl/6T09D3W5Nwj7Ak3oBUNbA51JmtjEIvXrbljHeja+2oE0LRalgNjSJcS5yJlymK6Nuy
jbia0gk4i6qaJcHasgmym3w0TUbruHAT++E88jpJ3bMnmtDljKzPSo+knOvf3pDeWp09VdbHzW3z
gwbJqGiCFSzauZpl4SVwox7tY4QvoHrlIXLdwEuewu+96od+f1Vti/2L7RqKnHRRT5PDqnhM9/TH
+EIak06za3X8kLUPB9h3lIklZimC9/9ntyIVdblIMO63VGK1yhjULIs9wKFSw+5vEUpE2I7VtPwy
Pjk7DV93wdxuUYU9BvFLuDmHM7c2LQT+XzPREadba5YsD4OGe/tXsdd6zmwHelYc+lqhTBNPUr1q
Bk9+eN2dmv8kayAiitwGoV1qN1o6IbOzSfEEJYBNRJTYWY2eaaCdpKiLCcOZclB9oq+Tb2S9/n1M
ACf95ShVGpMdh+1ysPwMDm2qfcXgww1ADBAKfCM0pgd6PAFyr8QdMhuNjez1PAgnddFIW2Tz5+6j
AG5HXH65kr2d6jjQSKv0gh3BXqNBec8rJxYpo/HZfzbzyA9pJCxwGHGbUZvGW+wxY0teAiHJ/fvH
eQdyg97/9uR9TTjJujsRM91iv7wQ0CuUV1OWfVDiGpZtwlMUQ7swNMoYX9Z4oFiPHCetkNT3ryKb
cxALVtc1rCEE8WjWISv2rfXe+7Hq+6cueDprc7lHkXfccMRgY1CBE05/igaWzUW5OK9PbFTxtmYh
b0D9pbdAbkQ2BeocaxCD05gR+kSJOJkavcGoqJTEdeObXz/n0T+/HO3p1vVQvlNZ/O/+0xFS25qI
mTOaBU3+uTfr12v2KEIRyuHEj6J2rjJSpZTRvU66wQy6Y9IHAvRwkXzjQADayVaZsv48RKSeFCJh
XAqqvXsxlw7kVuDce7jzHuy8dOpjCS4pyOgpYdnenBtj3DeY2QAoifKrbP6dqKXXiL9b2DygP7Sj
QJA51NjgeIxdnwsZMz3rhcI097DYXuBlE4ENjiaPyWof3WEKwZYdWxgNQ4/DIOJr9HaJTZ1+atb1
OJMkv3i1c2rQjBNhVx2cYQsK8/mXZlAveadAw0e0S5yF9bzpusW/aRiarS6LlWbbwzQwHCLvpJX8
6RRlDfKCdtS+YPY28rr4JTQxB5mlweUVqH8ptmxF7Yal6b6srzlfbwI55AeOGrb3UBD73B/gRqoq
CXF/O8MREF6bIeOBm0LTKV/vnK4a/wWo/0oF/Fm5zVkuWHBj+uT5q0WT6SDN5PIeAuGhHAn+caoJ
auSBnD8Q8a3kX1bu3rCE5XdH3SO0Qgb94zfA1y3IluBJ69J9XXTQ1urec0zMtUkHm3OgY3AHs1yj
rSHX8B3tGlBpTKWInjNRsp/GEQJc5RMgkS6aJqBcHeILRMeKvxcbphh8+WxA+oPHwy7QKeI2lyEr
8JGQ8wRB+ZcTfOP+eTt9teWhNarSLIqP59vwqymE6Y7iJKrcJEOJMmDCN8KAzTDYxQPIErIeCI4B
vklV8MQkj+TIhgs+IOuxv+9ycOYzUaZ+wkEcClOQAz9dOTgISU/P1cIe1Q4WB7VhRIhre7mtft5O
OI0EJY5vTEhj+TtNqIOJEWijNpbEyt9Wqqa7ycy65Bo2BVZEs5dyZsYQRyeXRHxD8UBbkLErZkAk
5ZBoO3YUvGitFF7szz/se2PSa3bhzXbiXmQIxVp7EEPfG70409KlqTThNUe710szASkEMvaeaR99
BM4ixxSETzSIAQPs4a9yNNxTpG80+wzCgAMSBd/mqAhGyEo+0xtt5zqGfIo2gHygf39oMfyiTfv2
az6mbgidUzQZybmOXPcPcpR6OMiywa0FSh6p1v/CldUQ/8vnnebaKBWEhXfR2lFtzEs89vJwDhYR
zBpK1v91U+Cp07sb3jmelJYGzOwHIHFuXs9atHnaietZRbyJs/fm4tdCIrmgZR8hQnolFx+injht
OmWLvO4WgnZUkiT1N3hGlJYjnoafhZyV97b/TQ01GJQiG59J+5LKNAEIFU8WmPfP5c5GHxK1AZCA
JRM5o26t6zhAOvfb9hl2DSgL4ohNIcG6uOECGJ3OfztLl1d+uM3X1uolkgkJcA9Sdq4YBYYRFKEU
zxqhSF3ipS/XxgH4jwsouKYIIjfu7PrN+873BZcT9EmEUj8ako6miSjMZ4LJ4UhTpSMZRhPgngIs
pjepGy6NnKBdRIfE2p1dgBbSS9DOO9sRmMHzJ3eqNsiGpMhGj8OzIX3XdfLl4yfvKWXWYOA6xMYY
4D3VB65JStGikacDuR7C1wjt+v56You2XERQ+Bozy8RFKnPswSfyniPNKs142d2S1dVWAY5wWs6h
KuXfFtmdb797qjAmUcqCkmRoyIo/+CGTVGigXSW1LLyfaT7nPa0+kDCtDowjJSi6lEXRSevT4c+n
UPiLLoyVxWkj+S/Y/2ODgmd+0GQRZb5BrfMxql0PXFlOJnpXstdYbNeUW0Z9tEbZNswI/j4cuuhe
lYiGsXWnKdAfobrVd6OZ8i9e6GYNn31B5Pfj0ffjhyg4UTwJjRTFuAaoXF4okoWIj48t2++Bom4+
COWEN0on8nD0ZRXIrJWaTIqtGjrvxJyF7KyHWNQP9VwKBoTqU59CIuDHXNXguFRQWi9q5CcPSXMf
jzzKv8dwf5ZyIHkOr36P73VxkOcNg7crkwsuZYFU7D3EPODT5GUqemcdBo59/hnjmN1LLdqFxgYe
fYxeUlyuYS6a4om8WpK1CO08ET1gaDtwoaojxGt6/UthQEt7aQ+3reuVPTGb0oyJ1yHUqcMjOWQY
2TYuC+C8CBC5ENwfz++jFUnEtVHLSlyITRjTwmhB/TZz/95KnT7PDLq8mLnZIPJRILaKRP1DCKxq
6F6F//IT0uK6/fDaNqf9cJUBaMK4MKUljzOxcWBjUhPyyyzyzsweQxzwrjUHxo8X06dxR9Mqfd7C
UmQXS32vVQFwe8V7tATkUShFomUJasFNrprno15GODW9um6MGz/JjVdr0CHsEBzoBUzsLkMp403f
ibhzrIsuVdDEeY790gR6KUflqRZpZ+p7ljpeHrXynz2aw8iXsSL90NJKc3sDcG3W3ROqfHuk77+p
pNf8TALZ7bP4ete6J9wKlckMgEG+CHM7zOxHsvIMo4G3UwKeD94RebqeSPKFJ05yFPeXuzwmeb9c
5xCapMQq8Lyx3BzlOf7I0+hFIhhWzztil5GQKfbh+SfzFkeOWOMTjZECYi6ihExaxYPSjWMyBbbE
hGGFKpzdSv7PectCycILjSLixllie3dJV9VVGx3P0Ulfe+QD3RaYlQDU7Z2I0tdxt2eV/VKsk1j3
+RL2aFfJMJ2kuaSjbr8BQHYC2mQPUeh7vtOMoECznurjIWsAPjldw0wkh02XDJLEAJWUL4WPC9s+
wjG3p86P/27+hTXARW5/gbTZNZlHUj/fs/TcHijY5tjE137QZeoiKTl1gD79Gs4jsW2M75DdmbHl
UrTU+vk2u7W/O7nuam4DSgYXHri9S+/eiplCn0RWweLg+oFzSArkACkdSYG6S2Ebvi+100bGls1P
GBVF74JdC//ECrFp3OFzY/xvUP3qvoG7Hf98/ukiP0WW8HBWf11EJluASpJhmJdkFJ8zM82J3B9L
tFmDtKwxGzwpkrJU3siUPHM/4f5XhOnSIaA6Ee8ortSSLUZAlq9+XVqMFeY1wm++ruMXMpgKaWyJ
tgWkFQRyd9ChEexWWZtwB6LM9ydVBhq8CmIiRjsTty9JVluZTN0jLKDHwim7Qyd/AkiaLDPATfSb
Bx3muuO+Ll+6tQJH1WmVyXkONI8onr6gCg138kX6qpIChQtR0zeDJnymhyZ0LuWFB/RTF07vwwoV
xshT+pXOE9AxFjU0Osz02DzMUj0SUFOzfmQrCP4lrgphHHcKQNN6EoK+7t/27/VoslFIYPm1zQuJ
TSX0aujwY0pusWLUd9z+W4Ornw5k9wqbjWjDGBsE32IqYgiNLw31NZFa548CeezE4pGt4ODkKOV5
36o+bXJ+Qi82xxGBNGdNKDR5W5lFX0YTMp7sDMCxEx//hTIWrqe+R53KIGXuwwV0PeLeOVREnf+m
VyohNbN5GGYQTP2qF0I5JAStlo9zKObIuHM/stSfAd5HM0WITEoB4UPv7BzArLTcLiI/gVlgi7ZE
nGsOgpUASMOYNiT4MASuojUXyu5547+K1ag8cKNk6MPw1b/PAs8BD42q/mu6g9U+3OuhvGG7R5QA
zbmarZxOFp5456aOleBn9PjHuLAwbN9h3pfOfHMBFqv9R0XwsH44uZPCs7YBXiLdr6LILuKdTRd+
RKjnxj6FaTxevPORIFlWG3HVxIK6OCt2ucpgjZvBSwlyoAbw7m84c3BwXXvGJzCAgQdyWXyvgQNH
hGdHzZ+Sjqs3Mw2oRQeFulH8JMZpqhwV6+8k3fJfcZYrRdbY+M+IQjy2dL2jUjJu6KgLIvrdJ3+5
tnKdWYb5uBCEspbg3hiMmDEE1co6c7bLvIKN8d5f+Qd7QYn+tlXz5TnAG+imxGF4uCGH05m0Etaa
4IRxavp1GD51wvCDUeYcy/t/4SprcmOFVz55VdcKEMCF42wL1l6hym9iOjQXlGjL01tXNhdq5hT6
+RzevmlcL1ur0sn1Dhe4dFA1jP4tfPvHNzp9JdyrVip7cC1z42p6Zn+UThA2l/D95QjiH4/iM4WT
wZJQ6VTr3rerRvcdyvHwqBoHffcBOh7Y7pzxtZBBi3278eLvw6rIvXNwWcsAf7RarRWDLPmWcMMC
NZ7XCDw4Z/juWDMft3jSNXaAH5XQ/5ldfxDBJAadh61ouI29hMBHCNAAshotWXNUVy7MEEwFRuIu
wbJlOA+fXLMsWg/qfTwDZ/BJIi55uANE36PD3QYfn2gxDBBIhD6ZkiVxhTr8NqcSE5gTgKB0K7nU
dMEyxzi5a3sKPjzJpvm8h4y36Wl9N73KSxbb1ib/6GghYxpdLcKgsTj2roTFxGTyvtQ4A/nGtUxX
2XA8BPUNRnUFMduG+7dVWpmXYADoGCPWFKxxcRVw0Y5sONh5K6jo3uYiwIrWgyNt4THthZ7CGhNc
y72CoqCdbk3+jzWwPd/6GOkD03G7FW/JRPpAW0Ot8gY2vQqlAQixL+tEu5iMyAxOLQQmTR0tEDph
bDoabnlvVAMSm7TllWPqPp70u6zB0ItJYk78zD4fldUnlzFICVD6NIbm6+arr6e9gZgjzwL1H+2l
3KApwNMD2/x9V+nf4WEH8KG+piZDs6mliDuNhlJRI5Sa53rmu8y76ez4e6bMeY7j8LlU11xnZhCo
Vez3lduD29Nin218LifbCNoh7XzU98EadTQz4INpKrq7TalM993aVGhktIag9+IwK983VeB5CpjC
X27YVqzWKpGoDy7lsgXzBGhy0iloaXi+UYVzQJOoWHTLz/zeJe1GeZN2OmvWYAVFHCOjnS7pSKfj
wqJ64jt4JxeIDZOIf2Jqb8Q2U2mBV5vpqd4RF2/38GbJvBAjSigOS8mySCbu1NjsUCc39m658zeS
43jhBT1Er7rxHu91z7UHjbKzxhL4qHWPsoJR+fcj2fo+3wFnRdaxzHEKOBv93mPL3bwC2iNiUub5
70EkLvcVoorTsL2W8PEBFVG/lT91gG9NOR+0wgfTlZvnyYAdJ8PmoeGAu3DoTNqHo3/S8jugpyLs
iQAlaFP16Tf/cyMxBpmQclkQV97ABW2URnvAAsRkGT0fSHT7XGuN/vIsCjATFu9J+aQJimceR8dL
WTKnSUhklAH23axy28qm1Jzi87H/FMFlcSMzy3W6qKFr9DO1+6I8LFyhtytw8GcC/C/cnDifnYpw
GnrGT58N9W8DLz6CA5EZBlFm76JdX1r5NBxCqYdW47gQ3UajCTYrQ/87/yRB2n7j6QpgzJ29fAhU
XvwxIS1tDRwQPCqk5V2rtuy4AFDGgmiCIeJxLHqrRzOPOIB3Iiq6q8n5pOlMDBgRR9Q9EYk0yPvF
neqbOHy9gXdw3EaYDIoU6x20FVZ8rAZIps60j+O4U0QwB3oUuBYzyh48FMrZjCk95HyxNG7fviTv
UdrlCxKnKHddjp2Z7cpCzzK6QMjP/dwu1Cd7ZQlN8lUIbu0BJZNb2PeJZcsv3NXSjG1bqQkf5j03
mtbTu8iuNXAcyTqNwaa6tMZUyUIqhitj2tLwl49OO1N1wdOKRWcOULTbhh0A6XIjzDQOrM6wg5EX
/em7V5/S1ycMgL8H9QqXjo0kqlJ1wqEn6KUF13tlZpKV1IzJTCmp5+JV2JEpfQVgFDi9mB1DZfXI
SfF9cG4cwyAL0C2kwRL99V0RDlsuJqWp0nrpXIv3SV6ghiVXQ/yHlXy/5m7Zs0uesmdzM+aoA8Cs
F97XeEsS4LIvhp91VpBiSdODGdv985tvIZcns8DL8ADDQNodPbHH7F/qwIt3wsxeFrdk1ejvj2Im
Br/WdjOH1Y/feH9v1FqNX5IMw4RbKy+gU+neTETXKlKaLCiLwThzKagmU5jly8bf6lWAP7acG3dr
ZYGNaiiDw74VEtH4NHaEOpYJDNwuiMZ8gOF7DtXwK0AJipwHdY0NNpoKMCgdyynb1lFPz3wWOQ6d
u7gQ27AQD08A8851DjMReNIP22v2To76cuGtj6qx8XNebg1uPDOwK5e6zJP8lruDbU+yc4i/uwmV
gJoAQfeR3uH2M6nO8dbULTDfYqTTYLIefgBe2HHPuSxfClTRF7wv6higxPtrFMOYWF7aWjRQCJhf
ShD6cxufzLTR/a4Ewi03zprYe5QUe6ejuPpuZRdoc26Qr0AwVMGYU00Z9F+2tJPpG4o0qNWmg8FQ
2LQo73wUEecALj8M6noMqVWK5C8nJI0paf53SjPyIx2YVYKcd4hHvKEBRvqZAU4b7k5gUFis+6n8
FU5kjYPaHnUUHqjspeNdapBeGeqmkfbuxj96sCgF5pb8amT4qP/Rai/nbcEHOLH564EdJn0pCVzB
wRZjjMHJnS6hQ7iKNEK2PeeuRDlEwUXG8KyjxsHm+aqrmHZ7emLQofj6EM9s4+80viWi4r8JWJxu
j8v9yudyy6l8tJbxMGjc5xakE2ufLObThnmN9ps8Z6qmSZOajQyGJk4cuww7pJHt2lWsjXXCFBmz
X/9jKnq5l5ozw5dQqUCY0NITtbFClSSH++eQU+X2sRIbjyNSorzdJ7+LGBxZb9FQPeTChTaNnUzy
qXUCkGYxUwED3CZOtEp8iY07J4/5UEVzKRZdR7XBepOm+7SCZi57lg0h8lKX6ao1QQRqWBSIN6dt
34cL3iik5+6YY6TbWDINrhYqv4A9zzAMtXvOLQBWOLrhez152TqrJP/ddc5qJ4Zh9Ntbpox05wYi
2pi+otwICslqXDhJU0Co71/nfwFVg8aAAI05gpfMwKl1DidFg163vUlMRZsynzeuZX+YqmP4Pv9J
adDqGdDsY7u+Fi5arCNPWHvs1J6rsxs0n99tpIXZzqtzP4Yqz5y8wUrSd+c1efd70+UsumqhOFNz
lHuqVzvddGBnVqoV2P0M8KgtRuyVZViqijkXSTAYAG4K2PfoavUku8SYtyoERkhxCqq/tGpR36PL
8NDNS3t3hKVGrwFw/7z1nmAAmoXlRQgNahg3l9DRqE/R9Y+nLP+ZZIeyuBUl7A8q91vALglEb1qU
Z+4SxW1A2kcuU8rjspSE+4Rp1OwAdm2SEnQZCTjEmXFWd0czaR5tw5vmRcmXt6zFzwjA6JEM4g0i
WvuVaxKMNJhqJtILQ8/DnvS3i5hd4D6nlBRBAIhmKEAW6xhicCRRZqyOC0paDKVHB9no19tg7ybD
9e+Ta9O4ZTu0DgHRuv13KzvCij70V+k/vKWwrXN/ZX8lBcIM/MxS2zRNRckTX3WeuVc/ObZnrM2N
QJ0iWTWooCSf/pLmgSLgfWdloFcKMzBPVOWAhsFTfGsnJ7ma4JA4qDbGI7cbrEC2WVPYiERKwVSK
oCyoloJBLlT4+lxw9jE1mShNYcAmpzwk1MlF2lr6VRpCp4+5uydIQWmcDwohEjJR/cFfSWVscPRI
nNUrcdGpUNiQXBLZFkqWXoBWpSgfLASGnJEDCD01iWoGRpsMiXZZKN3SqliJMdHstUoN2CFYbzck
CQC4AOPYhi3kLwYE+XaK4/m/czuUnSqDHdxQq6X1+6P5n8Ijc/rFg/WgLdTvQzo72vn+ZeFVkv/D
Eu0q9IsM4LAgNk6dnuk6Dre1vuNzM7y/ynmNeOlNnO5yWC0jWoRwlJ8Xzb6B6W2x3FJvBsCLydE/
l1EHeA8jBr8Q5+I8wMk7p1pem9HlDQQ0+uxWNF1HBgV2wC2DOiSneMAoIP5VwOReXSQecYTm5QW+
xEZ5DRkxmv7EJPmAzYBfPtRemc7e4c3FXHptgW4t9rz19CAGfKvMCZc3TGbTxDGpc5eh6gePK7fn
7YakCFZZsFlOAP8YEJzUvVP5YhHKQSYhMaoRrcOVcq8hgzOQ7qLLdLcc7B0hvGQuApZRwLMQ3Ch1
+qX0qkL/94P8M9pJJqC7Tw5dBwqfsfY1xZfcHvnux3PIdUFdSl/oPBNZpKKoXLmBIFfhHi5DHf93
dN1Ed3LQzNeedN25aE2JPHe8q0iCKIsJXtgsUKckv4GyJ5YhFMYTE4AnQ72JPJBnEoztqJI9MhWa
4bsVdGS//BPmtPDSiNDWYpb3ZTsYXc+7N327micZpXCHtKipcNUnaKJEQuFPE0Ra4/ccmB0GtV2k
80Qgoz5p01HT+nMBnLKImUho1yqRk9LhRSl+I7WPj8MjRm54GmWIBL4KsnZXph4SpcS+AfKaA3Ai
kIz4NNmZFNvbIzFE6FG2HPQvwmuek0wSO0rYhAeBMNjfdSTT2VXNzp5yUxFnjkxvK9KO2Pl2eNrK
Sj0Htu2KqHbN8My5O0xIOxmG0ndnLVK3iKe+HIiqXffzqC+5cQed6JyZ/uxyQF6Tr5o5uRd+Rhkg
FnA0dd50/qmCBxQz7Zwugsw1ZkyYFPM3tcKcufelvU3f4dtBzroGnKVKzPB1HeGrHsLUR2KMIh0n
5QUvoVnps011cjhD3d2pRgpbCNAt5phNr4xk5LFiN2LOPYgLajJBBPnhG1rrkLtG4rlJuLbnocX1
YJjEqSOnsJ384fk87fFwFNe6X4gVkm0c3Z67zhCMn4hevY+jx+MJY7xskA7tZrWf7BF6x2g83MHf
zGK6vXMltvphdo4t6mn/SG9pUtk7n0r74fp/idsEi4ZPn3qsOcFV8KrId/1Akr1nTJ3eEySmRPn4
3xku1Kja91oQq90Hjqr/yfC4EYFDGVLNDIkKkf2gV92whpebkfgM0uCecDDiCJXeHt5456JaJnTW
pRUQZjHg+Gew21qsAu3w+/tbAevqlTVg8PTfmC6dGLyA2KfXM8xpj/+u4SYUTUYDeVj0T6SfH5yE
vlFmLOKOFBUEqJCeQq+S55qdAQpZfRywpvSRZ/1t0cTNyMQ7L77RVtklnxkQz3h9gCVnvvhI0wS3
enwisNk5Qbf+wMX4JcyOcV+nEQ1FP5D/Nvkch0BYo/08ufBZWAxiRU4gv5dI8tNRvFUvf8X9yFRp
WMWYaFKw++YXNKRfHJPBeHuEJjrd3OBs/dmWxdQd8qX/ZF5NThlHRbULR0nauUBonmXnEYm8i9wC
dsNwMfQ6d0iMacbSMsTRKMwuDMykrPJlMiPq32JhYIraWn8SD1hZpMfvDbbLbeVEN0rF2kSe3pzf
svgVj6I4RVDW/8xKQNuTYLpCdNBZpTgPpS/1WwZUTlMBkBo14ObKU0o+H1PO0hk7N4ydAiEjF8eu
2yPi3pFRne/OOZaiPbRq1gczG91H5vyjlFZ0wE0B6rOEDoqDTF9mTD9pTLUtvs4rIKfxGBSfMHpD
PUdstGEYROKrOtmmdTZaSlw5suX/440YC0I92TirCS+yymm9nt6Q4Et3f0gXkeYJCXYW5luS5/wM
c+wmiHZx4dHM1bHjcB37TSeh+bqju2Js6AdKXDO9br4jjmmOcKrwmQg4E5WC+5KcuMo+2+DGpnlO
/Ps5TAEtSVbqGrh77c3mHzzEsAeRRJx5zxCxcb8EHo99iPVK5zAS/06+IViiMPnMRdhN7XRBU4eT
u786sHCL1E7lqnE1m81oovUkmbOPXd69yQyJGLKPPSHNhJnMQ8XdSgl9bU60lq/CHF+vDATDaDGe
gCXl0nDaE88jt4PCapYtacNhuHjG+x9B7ZYwRQeE2jOAtFV7kKx6KWNicI4wNAiBp9Yy3p18XqHQ
80o3T/kxZR/MdqGiO+tmu4dsp77LoKBQiL8USkspq9sbBULQ7HT/VHR2Qtt4n4IPRPPFkpcLLKPt
EE8GuvTB1S08bZl2q+7AJeobN/m7Q84sg5BeosieqHprHA1eKlLiaTV8dkE45Xx/hROOmYq70jWG
GfvEQVwEbVpu+SJQaEmF5eIuaQ75MpoXv8pkWu8AFoggUh3N02hEVQmPDxwTBbiNzSN/4cjNxGMP
HzxANHwvalbe9Ktvuqxi8+quaRdE+b86K8Iwk0gLgngDndKOCUuJ5PozXZ2MkXWjDPpQ/pK2VTbJ
IvECiN8Hz4XpAu4pakQtpkB5TmKBgMmqX2vaoPnLU1sFt+rC93n41bIhb2sFcIeK7Dae3+c6Z8D4
Lxg/ARDrEbhfHN+9uMsqQd2bREAOH0X1uJoXJn/n8JY1hmVm5rMLbixhuj45i5Ad7JOfCzAyuHF1
92sw2wmrizMXgYJ+Z5/3WA89PYzsjqD9ZRahzBwKqHHtg4RIYRVh28XeBZ/yNelYQJEEsN+tjRV7
+TPIZKpQFmdu1irpk+GoKOg954wYoCXok3u3nXcxGIfFYehk1k/LgxhBD8Xb/0yUj3oOiwBlnLEh
VJWltlinXAqDYuJWLl97drTxjA3nK5BBu9APzIPt5n8SzgzelTE1wCcyrXGQzRO7hm/M4huZd3f2
oyQrG+OZLqh1AFo+oRCzcCD9CHD8ZLpi9SbvaLoXnXbLMkr0IYxb75uwkSSwyVH2UIgnyKZImm41
cGVmcpWJcC27AR5xNBKyS/U9L3HpigByuB0b4M0EsyWM6gvukscBWs0ca4DoQo7ZHtzltX8IiNeo
X8xyYrCNexBHYJAyH5oI+hC1glszNMMxY7XnoXASOqhsQPQ5aMZ9+ar9eeHyAgXeI41tNiMaOlG+
+VwSj+emjTCSGBpExgfY7Q2vlfWO+go/DUQ9aYZgybwVdNLgLbRcOdGCr76Ic3UUSnOZ8QKJnN8s
bqBY8dEhMgpwvawL2NAnukXcBQn+lZYdNzAVQMRXCuMlzOacdNav9vkzq1q1Ta/CgxI+crwNhiGY
oxWZFNNZ5iIXB4nIyfu/WkjZuiJO2+24V5qt0P146c6DAIZaSj8z6JhRbH0A+3q2zWTeri+3x3RM
jPmVqkgHkdcwBPsOYIUFg6zVbfYunfpK+UVq0H0RtE/VGCNDvOIHPHhUZIBhWRMB4JrWIR82pJtC
zcS24bkyav92zRKeaXFJ9vcnIggyOh2sePstSmHP652i4zkwXsshIThYs+eehURYSsKwdVHZ3zVg
6pjZv3y/WlevdQ87U2GQwGDIkjb1IvZoj0ZEJOESrULi+qR+mrUcYPlTPqQa7vSNdW3jCmuCLuYN
qTAytQBo1cUp5lUHetzqR/qf/NkuxLEJ7hNfmRoB4Z46ebb+GRkNN+s9gCgfv6+w/zAwVrtlIbbW
pL5rmazW3O5jDlXPWlLNJEo5Zxa6iWtIyEXJgPiXe2lrnMFrsl4ZROYN1ftAznp2DtRPES9XpFsO
vWzytSzg8HivG8YQli0H+b06IMdIL20M2LPQz0aQe5uVk2GAnPlr4Q6WtAN/mB3U2/TGvNJSKWUG
bTLkxGxs2Yhoeydnmbd3h7qdlT9aTS736pgJDP5Jt5DRSuD0D0eqSK9YixhhX6KU2n0sdMILtZ3y
k69NCdT7BitxAExxPFNsuYBxoq7PcW8palrbEoRQ8qQaH10LUG9kIkK7psbQ4u4WHqTd4dSutdg2
kN+BE4KSgLwg2lDdkAEDnMocIx9hdNeFjkKPw+1t0POQBDQf/UzMGq01nabsJZm1LVh20PDER9hR
msu1JtgX4KjwSjYo4+HgQJO9RugUw1KIQElLqi3dGKf5iGUdtlUbu7Sl0o0m0dru/rwqEcO+lNun
59JaVWbOu9gUoYby76l8XbD7tM+DOJA5m5j0S6BQ8lwwE82xrlNAtnANvFA5pSmdrqbam2jNwYm3
FCEbvBW6Yl9BsvwpHZQ0dScqzaQ068BBb3bF3L81xMzyBCaB39m9OdeE77P0jH2X1/aLwrIodZyw
WalnweS1CDDSkVq50wYTYa4IQL60PkHx2qrH7wtjFLbN7jBTgmEtQsCQ5fCI/IciOLwivMAX8fhA
RNZvhw8wnAWmij5KmJ1MFz54E2bUJ9flI/86P2Kw6fyBc2y1ZrlT5xwrUgD4luFLM5I3yGpihoK5
s+SB7DVbMb1r3eWs1CgXaFLxb+2MTbIH6r897mT2zBAOg/Som5McWiGWVwjZ4V/YJNybiBG9XuJB
l8OskoyZfWFu/+SFtlBA7Zrbeiep39V0xOETw/JQ9l8zkf6e3p9m9TjBQcR4Vs6peb52ey3UveJ7
waIYco1Gk9JAD/b9L98ohUXSLWTuVO2Oia16mte+6kps9Ax+0fAWe9lXtPQ9hYIMlbUrNgnOFVHt
7VbV369TZnP16W33969UFHQzNICCGUT9Nssz5mcV3bB52vSVSPBOmtRsKAen0hMXaJRJal9tK0Fe
hcNpGe89uzSGsx/XDp916SSoLP7D+cwBkVHg2JoKZA/BfXQaDSPIAVuxrycaTivdnbDuhB7eqzD6
kn4Cs8wr1GZSeUn8g2eeIQ2Vkmsx5AOeDWT2HT5iWMpBjQ+d6FTRpYDX1p2oUp6EAmMxbynkqoDh
PqGkwER8YtVVX39fptJpKYFQP1VqYoklzNgpqflszANS+ek+Zq1+NoTy9nOR9VWjlr+41pZHRcLK
+FXyWjXXj1kZ265E6ThAXkPWGYKK0VKAfZ4znQjbsUx5G42dcJvQuLjkQxQ4aPnduk61L1m5jnVG
Yc8IGB8ZbCE6I5Q5MDRUX5UUZEo3zbYmWCLMM51t9NPZ1YUxApkF7t3YbrWjGHUgmd1BIRFNeTpu
0F/SPYY8uganfII2diHP8sANd5kgXEKTHK0fEbUTVaSwwP5TKecz/5Ato/aYF5905YFumvDRxUZl
QFFJ/2rei9N/c9GcN5amJschnc1sYPnE8Kj5MoDzBONIFF9fpJe7Y5GZ7U/B97BIyak0Pm1dKBCF
PHf6jucBL524fx9u6ZdSKT9DpsjfY6AYUAN5AsCWXPWKWVyRqpBE6b++BD5NFXB5fz301pxfmA76
a3a0CdFQqpAMNOEkeNEUdn59MmOQJQEImAlshFYn6FomfDwykdZJQMbklFqi4ZZArNu84B8Dlakf
OIEguSfzESbFJeo8ivqr04+LB31f4rQIwCSwCGT/G3AuAkIr4yPejMnMv08syjYWTyR/qeqD4azY
GMCiWRC4Jc1YD86zt2/7GaqygRCUyGybdPhkfi2bv8pyfsEmMQRXxMOd7PX4cCr+E4oum3Ezb4s4
Bik+7/a892qnHvA7Aa0eegY0NbuyhiYay/Mj6J1cLgPPKTicgBwMLw8HydFWKVTMlbkV9Hu6XEVw
KmBz13olTgARkz6jjvU2LXpfD+T5eRKcbJCeB/DKq+2pXrXozCvxsbgHkia+o/YxWR1kLDVZjEvR
cRnjGQuLtZci0AIj3uahOFS89uUkrldnhx/fFTmIjiSjzRERdHBjI6PfJ3eurahVbxvuShWyLbKn
/4xviJwgs6Ah+2pqyg4e6khJZD4axKqy9yiQ9BlgmO4VOVUI8r0etS4dQ55cAUemouWd55b13S4V
6kfhIQC0b3z0BncSCMpnk2bwtnPf4AkwU6JwkX0YQSF24M8ruQyfYFxjPaZ9OsQdbC3u0cNLzwym
auK7Fbl95zpitWfTEHrb8NOSO07ph/TmNONK4pB6tO9/hQLhvPBZUhc8qw8tPKh9iVFJi9NpnxCv
5ZwBOFbjBh8GmoHoslDV6oiQ7orni8JiIrtABLEI5cVA8VrATrRFOoy1i2WZfh2LBRK8gHcvjyOr
pM+mAr6z99FC1i+t6SXwOZ2P6Zvw+J27oBeAk8bHQXY9JuIhYV466WKipM2NWIeklD6mQO90gGZH
0Cgn9cI+ohNcPn1DgajHrLvh9yEyBSS0MqIu7sIoWcv8EP9+yYYQ3krVQ/k/fFzZKclPuPQeAYa6
dctgiCeb7iL4j9kcUX5hvTJxSleb9WBUt60mSrpEZKOEg4/7aia249c9rQBqhRb/iFZx0Q19Fxa1
nc4hSiIC91+TrJk0wnmVG6b+j1q2XQffmwk1mq/tPznYV5OH/gGSB0/8OB2eF0wi0u/v3XZ8jBhi
mXPhfabDbj5BBAvPijBSFX7aOHJuvJKNnBa7RFbK2haVHX6kC162ooActqY8QkbJpyf4jOyztU40
9jYx0gnf5xQ6y0+Wn7wAD8ARnbQQZNqTPwZUYD3Svv5xEptWBxksph3+FTw7CBiZ9QnrrNcho36R
Ldhx2qaNBYnUaX9GKQ+D/S+T8Anz6l1IYYH0mbT4ttQc1INJsXrLoKz1EKBKEjWrvjQeK8ql3A7M
OXSZjweq574S0vpXXUXZh4KqfZ7rT57cUjR8W2OQWA4gcEi8ES5lnrhiLbQOJUKjPOV+T2XIBWyr
lxkHVsi9p6rdhbPcRqVdr31BHUO46soAIQRj7pHm78bszuH9yZk4eZ0OiN0VIHUWOkOagpDG/bKk
hy0kvn8x8VU//cdU6tQMjzINV0PwJ00peCwSbiWx+wBHd50dH2j9x+pHmR571imK6c1NvWix9sh/
bEQefA/oPkYmLfWYR/gsAAUMQSIvgoRVdzDs43Q+Hzi04C+JD1dG0qTlElPPNLPgiHCFXk3XYR8m
b56SER2vn0/tabXa4U2WY7hPI7WZdIkq/i5VtVOKgMd9XgOM39toiHOXdTX44GQkhfGgMrdKj78T
pBKEHNeAssr05UQAGPlXB0l/ItC5fwgpaTCBqNgh6010k75ENrJaZWhmUwOPwjreb6z+nVoZ9Tf9
GQrOSxr0473rMLG38A/6OtNnkPG7E5WYWPBrA7O8Lpazbhx1JyP5yD/5hFCc0ujW1YYd3L1q43Ou
+wNsPkkWghj24gt3bDu0Xa7kBRs2e15noC/lV/0VGKqM+8IsMCHDTpR0TTibDWT/peWq6nA0wkll
jg2dLbNRyqoy6GEN7zKkyKRAAspgoDQPJwzEG39+ROp+TQDz3NZ60ijqRGVd721NzZJl4GfV6e3r
Hmwn+gelQDTH+Xc2RsLQndwky31qOHOnqYIqILj25F4ksYA2YAXhfFkge1f3BQj1GEyQ0VoPIcQ5
oy2U2KOJMhTHjRQCZd1ZTZp44x6zVxbEaU2Z9sGv8C3wsjvoypm6JXmBtD6TF8fgZJCVaMTnKxJa
wBI1Ipf8Dpv5nm5kHGtpc13Oal60e97D2Qb3Qow3yqSPfkluDmsmSN7REx/NklYqNryWiKTrc71K
1OUM5BYLXkkvk8W4WC59LEx7hrKdGfJizsxSKxEcytpxlFBXyTJMgs8u+peXoZzt5DL1xe+fkTlI
4PqW4rTm1aT0tc20X3mPp8AiFAsSfYWQ9+vD78iOUylCrxzxlDPNi/fJTfs/Pup7M8HfwUJzFhYY
zKdlfu/IhPJlrd5Kz9MIPFomsbF1bX6mrZvmIy0LOpPD51tP9u/Xcp08VNcd0jNavzkCfmqiE4aR
zFRJ56vT3S+oh5zJ70y82Sr/nUsehTQSCpxeMgO2rpsjsipYJ+54LSOyliJ8UaqlTMJ3ITvhWhBU
jr/piDRDySWlaIKhxXUBTRYMew0Ms8PwtyN1/J2wZDQKvxcQpLFZcvLF6lEUsPRqDEyL/qBU/xbN
vfs+EkVKdoi3Xf9Zo5MtXxBtGQE3P2pS6SuPQZZy/secCOnBG+rv6kkXlB20m1w2r4m6G/yyICQ4
5EMbT1v7Bow4He49Hm8FZkwSve/4T4/964t01K4UTRCoNFdJ2yvMisgPPKG/gs/9RHYSvKwTbs7+
TFc/Ory4kU2SNlidG3Fwln4tRxhgpTmtkLUilBsqv3dG7Lpz954a9GXHbAMxlU8clgzFjX+SdFzF
2WY3s9N4Qd4d3kA/H/PMVhOG4OJ5C0F6769B/0DwFo596H/O6V3ufdJiqk1CStpcww15h3K0Ard6
qKHvtKgX1xi35iuuIlgob/XA7baLBPheq0JXOK+TU7pMY2ecWmdWI+GCjzCGxKBhAfWiWe5rdlIg
fJ6aBsmm5rV3li6n0Gul+KsZnKGO8dLZZx6EImtXfBcYKArNJ9zBvC/3FUrDRPCFD5ThIfkUrAq9
rbKF10Z1iYEdo4QsAoHExcFMECmYOchr1sNJGXtr8oNqxPzowqUbxn4CdfiReB1+2apcifI+QcF8
zo9Mmcl2psjEwqdSFBwqY0vM8uy3LFeVgtvOSxD8dSp+E0M7SkUnWEjkpZCr5OXYL6ULsdE1TQU4
MAZC+wGAJLeJRHuY55zk6XdzU83ZTvUqScdpLAI63BaEuKAvIT6copSP8inDvpeFg4I+v9p7t8ak
i2GekXoHRD1LR9849vj5Nun2VO60zKkzewwrv3NHYv9mJ0jagkYyf9Fv9wAuIX/w+LN6eRu4fKXo
m2nmVROyglK8qlcWNa83VRjAO0NHlJLbTEq6OxQUu1zICnFjVyZpOxFL06S79Nr12P5KWxSgc8qR
CeZQzCoppdfPEX6Y1le6+npNRuQY2HXbJSOLlrnOBzeD+HiUkYaSuUS5mhBzYdHy+FXWMJA4vcI8
nvkgujGI/etESz0RMVQASLTk3/TgpXdj1i3Sj1GJHSabvYxAJbL7Gstxfj5jUxO/bcnScvGXAJAh
iIdFKQvfU8nUw4KJE+6+9Ws9eQ50lUR1PGBEw695T8aCoVDYvfnBQuV6DY5XFQvLRf8VCMcRS2gb
1n9rGqniDFQ1B+YWYWcPPhqpzUYuLDuG4UITpptg4IkNaoq8vxXVcs2gp/KUKYaXtTSnZnxHuam9
FOEodQlhsIGPbd+7c/65ENWa59YwL6EmcG8VHg72xi4smeSEcMvcCtbD3HqS7zjnFEEsR8QrNreS
7mD4R7qEmntUMTYQkvGVeQnTAEDvt3xhvUv2knhLMhXsJ2eA9llisfkzZuOn81P9jTn5bQFe0jt4
8I7cC0jNd62h8iktV8vsrUIy+56PCWFPXdFC5Os5/7sQGBGK+qus32kswi+uM2emRpfG23N98G25
fG/kdsrMYYNfurOjfRrBdwmURLx9LDVyDtAQHLDD2EbO32oQX9gz3fUspMKnEzNBFwsvd7ahMmLn
LumJ2x6nzpw7W7Ltz3gAIy/3ERaQTlRYQ4dsE7r5KySQ4QMITmCsIfhWRbyOVrtT71YBUiS5bu/z
DSQxkR9x/3GLGPeTVAm8dtyKd9n+iQD6XIjRN90+w3q4So8RdQK0jAA5uqg254772dGap59fa9nf
+a6HSyPk/P7WDZfTxFkCTPNsc0rb0ev/G7BbLqkk9eqJa5TudfoMj/uZ/whPU8EIOD/QWiMwj58D
VQo/QoVwOKyuCt+FErfcv78SWRItBRl8GAv6prwN+Z6D7F23mlv44ydwuBIPPNALJkFodbx6QYPg
F8uehK0NE/clo/R5isYGLU9PsoRv7GWON1vh/nmrBa1Hg4SF5uXiTO9Y+7B5WaRXYsTSeRjl6xW9
4h8BD3EPqUrCziSYf2V1666Byr/82C/AvrFzvMywAsROyMqykYjsPPI6ou9gICt+18YOI7R9WLtb
5DttwXMREfoK956v89FNjZzZgpgi7RYAQm35Xk5TsHHzvODPfSS/2qVHbYRN5AdUPEJawR1thE3m
IYpQB0GAgnW0wCd4JKfMa+tkND2wBPApg5gUjz8GgXyHDqv1wXKBC5dhrPg2F/2r44NOX+nEu5SX
aI2MBc3lOCTNHP7hhT64fKCDT2hlvM+/oS1le6sEs5x0cxfes2/cRTlgDWaCvs9PaqYgsqeHC1aM
yOuHM+5mI07Aj2obJbPR3l74DvunEC9gXEEfyFx2FhR4MC+C5ugBPQn9elCx/oTyWFuyRDtJCScz
V5/yy7oh7iFqJmT3TbQFmse+tJiko2EBgZPzKlCuekg/KTEnlNfmmPbkvaZJIOO5a2SmAuMmaWDR
Lpyf78NTN4f3BBI2YF7chzB4YmacLQIMkMqYxXib0WyADrP4iGJAnq4Yok20KcnQJ/x8YxVIMtfV
hxsdFsd6ImHMBR0TbBRFLPt2lQYw+UnNIYQRdvgmX4kX0d3RIU/zEzWIZO34PDPsTMRpwzHYYvWW
ipGEIYp3OQih05rN3PJz2eu5XT0pyFKd3IxHofVwf9l3jNjKLbbIjFR33JzrKa/7IS99pRMnvBbX
Es6LyXL/YpFFRBeRRuT8BxpGI2mQliLqOq3h3UC9tIVUkGXcZ/2B+pDKuvOQc7Fe9YtRFgmEcvsQ
xyMruzXJR4YCOuIS/4b4Zd0RsNOwxmULa4JcDGf8dvV+iOfRWC9mGmiY7gXgzuOW20LVkaASSPFK
vpP7KVo4nAD4erVOKLOPPnHhPjl6M0Yda0zyz+yk1G/W8QK3n/FBebaj0FTqtgz2fnsT8NheRm9+
s72d5FIdQ9AXEfuuNnw3SmJa0PtZwXcC41MQaaukDZsqno27jJ1goc8sugGRAP0FKHNLwLMZdlMD
vHcemlX8HZHFF5/3dFRBJi85SkK4F8DSwQDxK6/67/YMWmjHCjuvI+SKKQrJphLme4S7D6tdJRyU
1S98fF8+ZdK6WPcX68ay4SBf900YDOwARHfQr+TII0sfvQKJJ8TC8vRW3ndIlHl0yhfRqGD42LWJ
UbngoWF94Z7DSdMfWc+2vtAwnMMs9QTgnBrg/8wtgAWVGsDYLkMi4PUPMBW0neKCgamEesUQktWe
aRZkZjQQ2ZZ9p6BsxDVRcka7S150ufiK3G+9HBmri/GGQebG0+YwKRzSVvyjsdD1XZxU9qvG7DZv
VWWU5HddCZYxnzrvdx/agHkwjPA6Pr0FQDMH2fIQvyaoKTL2JdAv3nEHui2moBpO4tQKwY4Bq5Qd
ikLHcQ3DDTMJsXSXfIc1nbsdfpjxMss1viYNbyHSBHXHrM5PMc2KoB3gLClUuQGg5OmmX2mTN8om
Zd34SZ5F9x0CQmWFTl33EdkDXXbdSgTfFzv7JZYNVvKnPQwtRHqS3eI3FBQVCYLBJznik0bUGdh+
vX9eZBz6/uR+g7Wjm98rnCJZUTwItxfPdqQvz/dpe5o3l0Q9F12IFROa7nK/GnxDLq6QLxmxKHzA
scwsUgLEmkIM7Sor0IMPcbxcBIDQStK/g/smReBL7S4F2TtF+dtBRT4RqAbu5s1Ljl7noQLbFQGh
PGkc7A8W8X9tRqpIKkOBEzObuqdWJJnLxuNrFktMQ5j8vC3uuoJl1FzH1fHFJQOKEE8y4JuE42Id
QJj+M0snpVVu5jwYcwEP3RdNCLLIlYaFD8/tk1jGBqDf8ebi5lgE0X/5X/pjGU083Sfis4PhdFD+
hZ5/iCgl/bEwl2hnkfbg/71DE0073mRyzZw7gmDPd/694XZhE6sCDQvTYwYiFgXAWdlai3vKvoXg
a+NfPV0VDhBUD7sqxSS1CU0o9ydey7C+5r+O4magIl0nv5lAvktzNO98kFaLFOF2hmfxk0QDmbLQ
ro5Tx5q4m7t5HlbZYaYFUaKM5xK787uOm/Yv283rjJsv5IDNAv2xgkfCPMjxC5wWseON2GWrAsvL
J1+sTMlNZbdACGXFg/ERPjuGwPNUFqSTbn9Lc+vo8lDg7FUuA3AGUU7hQdoXwlGkHRQfnP+NcZ+e
BUb8ni+VMw5vdkHwwnZ9osGA9RQVtpAxkSazLXKewsl76bx346WocCDYw2clE4xnrUdRSO5ZCY2z
U+2zBFoYi6QQKQyfM2iaAu2JWovZLuJzvyBYIZvQd2RsJenOL+seDXdePl3/P5eVmazOVb5uwKq8
CVv8n1GteqpVXrK4lm2u6GLm3HyPHoJkR+dvzO8edJM+TLDIv8Q1aIceDqSKUNnabzlVJufs1SyM
GebPKdDNAzXVZ3vvEskajJ66vCjWPFpwXc6K+gN4ikrCVGqMlC1/lSQj0iQZ1KhLeog9XqFo2Khn
+/QJHmWGxcvXzF4foir10Suy+2UoWZhGvmPJIzjhhAVgoU/HRxeLRwYftkukITXfFkGdl/mOUnaP
clfPl6vx38h/IAJ95hl3bkVAlTNr6JB6urP+ilnSb+p+sXiLQOle4EvInt7DRqqn+VjAZRH0A9iF
otFjJnx1JPi3MXXdTc7UlgIC60cRpscSfB7BNGfOQhxc7F76gzM+k9/qcIDvU3zl/of+oZcda2EL
7veAvUaB/BwbmRdnOFdl8C7lzgwvEzLAZVFtrNe3b18Oow/wJTMpDV63EndWXzDi+QhfMo0kAN5G
frFZRPwgLtE4nQL+g75i5R/7nKz+JuJh+2jA3ILqwniC0ahSDErf8NZoKv5ujn/FiXJb9+SFXdxK
uWv3xh870bTDNiW6ULp5lDdAsqp5ttOGeg8+RDHaiIPr3gcSRRB4vm0X5Z+4UAf15UjxelKsj3Zo
IA4kGwTL70wyJFLNxGjx9DwQrH/FcnevjlVm/j1ffYOsObPZYYCUVbVyojr3r1TQKnVGxWJzNkjq
5CSRIiE0AJTAtDEV9xJZF35m8W+3zdIMIkizpqx3YTRDsypHMu/FTgo8v7KyfdGUkQQWorWNz3h5
FPW0DcbaIZW36r8ze/r08mzeajgJyZIXhJkmcueV5kda2s1smiTkaYtsY+3e2BIp/VOJuu3pfCzF
2s6D3wu+Gractb76fPhK0zeECsw9nvhBVUREXIhs8IxtdmF3kollnjqV+mJVv5JFHZ10xuj2eb2i
NbWhuylun3vj4kMttPQVL0b5SysfNqs/R7GPe4/c3/VgS6KvKxY3nflbMC3SOOe9dfWeBPVFLilz
LSKIAu/3v6dSwnunqEcVmrMdP1LGN8VpI/jAoS5/sW85HPDpPLoMe/6QPvpGio0iOsRzWqHf03nH
RLCw/ix8PEX7G4OH+m+RKhzt6hb15SfJA21k1LnOUSrgKwWoOdikxTUcruibgwNpwpHKrmXwO+Jp
x6cO1B9qJ740wBBTCa3Tn1idK16lV0kJoQyJSuJQdSPyiU9ttSRxbnvIO5DfjQwF+RvVikwbbCwz
mvTi55NQDmFA/lvKkYA5FpVWrJSG/AY76xUHcQFCxIQ/sF9KKbvVFNcHjjEBsSrNKXKLwf6dl1eB
EhnxeGB+GV5ZMpb0I/8RfM0iWfs+NybFJILm43hQvKcAaXscIPyrAOgfcDzJ2nrBRCowPnKkIem7
2tU+sXmXsUGrBzJGGXb7b10cBHsmWRy68kHflvlyZT/0k33cTK+LCd7gXRrJ6f7gxoLuq4by2dxu
DwzbLAqwz69qUjk9QkoiIHjQgxAAcJooF5zf2FG/S3d9+bivNOxN/vSeqwJWBpBa1yhsLilG4Xjh
0TKVy8X1ldZQGi9HJJ989iEwBnCx1LU3QQ3SrMiwj+iaTaPZblGwMGhDLPU38cUNbMKkDiehFnqc
Fsz5rBa5RwSOB1JyvqOJL8waRtN+Vxhh4QxVPvDugAojyNya91DKPbtym6bR0fm/1Oi6URXqZtIK
oO95cIRvfnJs9x7ZSZ269EFT7Dr4fGHD00Ok4bHbA1Ap3OXcS+pMCLn2vK2mnWxp3XbMxDpoHoRt
8JeEXPnK2s22xjbOP/+8lz5qOt9+E7NkWUzZeRG724TezFYLPFEy/mZ7sSnjUNiOpJGxIr/FfjrI
gRbA/oUwnVRGIlPC9I9ibiCiawAj6jLxzpSKbPSfedrvcgxWqSvCMsCz0ymJWyQUBVe1+pY3nZsN
VzB/Aeei0un+Nx00fe1UHZnYQRQXZ53HOpiaD5Zk3JMvAbROFkBqxHHdi+D9sfEYxY9k3PawzgC4
43D1Ku3lmQlch+xu27lSkD+Z8VinPuDDn/9xMSaRKhq1nSPrNVZzs8Rz9T4w3w+vCxw+h86GmGtS
5zXvThieR6W8Q/5X+aSyDCIuFceEtChg2SglErPtWShWIeViwOWMmkmwAOO++RSIvcgZiRx1F2RA
9ycKp3ji89Jmcho/W4DCSlohf9IpdJXLPfqqypWjo9EJb+Lwb+wiXS4tgWZ/nlLwXsZHeaaDau+p
YbbtjaacjIm+jSxiCuhQcw8Bx5Dl2bgylvOqXMhK3WnlNuXCHVOBoF5e5f8L7q/Bkn3wrWBi6p0V
ZgxA/h77O6VztBRyq27lpvWlzHgrI4DWxlyuLScsAHF0iWG165mNSB1j4LyMsYWGg1515IgjABrR
LNk4wp3Vk2yFRJ87sBoPCED5OWPIIcv8WB9Eb41chzVrrSWzBEgIc22M9HEfzWNc6d6ZZjPgnD9x
rn5rGo+YwTWibpM1u5A+iiXLug293Nx0eMGACy6C5Nt1TwtSYTCxlERSVB7uYk0r5BqGRpdUkXQZ
tvZMlMTv2k2MYxqSQ5mlAgDrcWF+fMbP7Yd3ErCEDjAXvyQTPLMxZEoN2cMKu06yMEl1KFyQLHHn
Ok+AOPgAaIqUCa/9r3/c0WHbz6LZsPrJ91CLx2/H9yxn7h9fn53XQpbp+zNVT4Lu6UT5LWWQ4TP+
fRco5ct9IdlKTldF1zhzHNto+rjAr9vOGBRT8Q99R0IcJmCU13h5UWAIOn1QjiCWRLsb/XRf86x1
IIAhhvUat1O6hB3lEsxAkt4CAUOwARbskXjbER/yGuM4mHdamgJ68bXQMNvCtaUDcMy5Xl5VQrSz
HAOOIB3U4Uc+OBm6EjLQps8neRz627NM2YnDISGwTevIlxrCUVywahxPlS/puPWHVFjK+HjKF1GX
NaQGQjkPOtZPYHiLT3wXVqfcdvv62q7yXRbrOHulage7ctZuKBsE08DshMTVJKlgYwML0sC+HC3Z
k88bYhxS/4+OBuxDsfr9SSidi+7E+PpJfp06UcZjwq3Fjq/WLm6FxfTYk7PJ8V/lVyF48wLalt4E
UV+cSW/L2aPmCDY0h91/PE3zLPxCEZWXK72ROvkU6qMnld+PwcA2qh8GQmt7C2ZwtFXtCOTR1ZZQ
vJGbP5QaUPH/7n3N9TOKE3Fxc56YrPc/katgAhsUb0eaH7M6TBBb3Y5/vb+QyACm+UAVEMquzVO/
dUOEkzJLUJnOCHurjkIK0qTgWMspYIbrz/zahXPPAlLqCl+j6A9zktLiTNSDl8/AVGdEc2S6Cqd9
0RWrWWm5GYd6kJUo0DupdGl42VU0eWIrA66eEGyHblBBDf2wNEFqV9cE3TQyis0BWXcbPSImFWNb
WQk0G8G7aP3yJ4zBJnH38+nW/kBo/fGV6uRCigdOvDe4+9com+o4FgSn6TgJ0Ek/ujhZ78JwHlhb
iqp5s6nOhfHV3c18Ne6M+1P0O2zqPehtqZXB1qs9thHh510AzeY2SLf+trZPMhFFsWRAwjDXEnri
yheLVtNSXuZvuIGRCYCuatoSoEkNAzqnGGyLRhihQZbWfap7qWhFNgFx/BrKkGxih+ueRgv0lQub
9kllVRAy8cCO46vE5yRDxNXybhMMD29LpzXdSNhwlAOPzEHRpter999M6nAUwEqMziIcdZ5HB0oe
ou7in8aJ6GS20F1I8MpFRYq0FwdOVStvDyzypjCo1zrdoXs4kr4+shKBrz/5pbLTs2XmnGhkfDSp
XStR6Vo3k/2dXZLLE69GqMxYAMErKCzrhBS/MMMJEBAYmyGkquzPCYpv7FUe10uiHXXflfuM+1+Y
FwGq/IysrcZlHBJIHn9N4iuReaFoazCjFhiNzpCH5tofmKX7Yr5imOOYfUET3ZvO6fK7G2zWpSx9
6vQRchbKOj/g0gk5UEarkIcFHL13TH18LZKE6hFFXIK8DQgA9egPLk8D/RzoBI0UTTEzWcZSZdZD
y1nKYYFjPKP1i5t+MB23MJYkKXqx/ai+FCTyUoh+aQwJsFKyjLcgXCgBtUd31l6HRVaCAdvDRJF4
nX3j5urEh6+Jt479HNRhTUaXQPCGbemAMf+Jfur1wGvdRkMu2l8W34yS8I10kZYCrhYtDDaZFqJk
0Q+fxDGpBOPsAlDcx59LTf/sSQcbNCQ/JO3Lp/I8UYvihEFF82XDod8Z+CLWb6mZIAfjVQlO3H8/
eildLVmeTn3DwvkG18VSG+EFwYtrDposnAndJUVe7S9Ub1CzYd/lKKnfzA7xq9wP/HBzrAviHWPJ
lMTYeJAoyQoSZHHnyxnOU91eV+ENyVFDzwamNUa8kAOXKvhnhE/V7HM/BJjitmuGw3bWtI8JqvNz
geOzipRm9StB2Eo1d+K2G3zrIzlAqldYsvaiMwmLs81ZgD6lWAYpzpK/MaEgDJq8JbOu9mKUIrcz
a61M1QmYXTYZXlw2Y3GHbupZlGAlLGGXAqpVjLftuAopRQXmfLWgM85/HxN5XKQQPHZNFRsibd3L
0G0zTnR1dcB4WGs2zdwQnNqaFYoiBO85EVUrdVOGLlV2xQp99wl5Bn7gKATo/dYQdnIYnxLfWKHw
dbjiq9rrCLFSbd/t+gDUCjnoCJ0IXtlc1o+n7ZxaYx74H6bzEkNfzEI5EcmZhI1KLayE8tV407go
Ust+JG+vXAR5EQze1iwG7VZQ9yD1ER+kvpOoUei5IpJ/MzAXcI8W3oblF/IfRcdzBhPTpeoIK1pr
ygSOHv9uiZiazDSdl/CZRqWjYENNAPHeVXjQvTwc2PrHjbXAIieJ6dxpeg/YNr4+jswWWnf37baf
DRj8NNxQOUsN8Q3ADK+qn+zLuvySy0yMBJqkkUSwz1G0qtjp998DoxB8q9qQLKTdB1pR2uUgOuoC
yIxLuDcVz7N5hT+4Rm75zRBfu6QxnA9r9WmVtDuX6ENA8HhAb62soLt0wJKDm4605A40UrSAUuTJ
+MWR7DxoYzpNTrjEMYy5oelXOz24vxno4VR7TOtDfS8Ychj70HvrGzl4litxCxN+VO0lgokWN8B7
42f1J/WwUNzSs02IbZYapB879VwBsNHQzrS6mPqbXvGPcnZQ8k1JxQgC7mpj1SFMQll1fLWgDpew
unPbhtOg4eul0YaYZtPHm2wniHfnjN/f3qu0OVBjloeyvU5SQSw50+isYeRHehClCeTJqYWC+0Mt
jT43pOBngb7xtRcUW+/WOlD7o+ukJCSZa5LpQgbSe+JG/TKHH42x+n3aQjbhoCZnAe7sbjYAl8sd
M6hxQRVuaLI6hfBeEY7ezSnFxkVOkJ/WqAR8tkB0MX1ppS6qRI8chWi3oJ3jYr17L7jibQowQZnv
Ho99L0rjnZB/3DVsQbLuYMml+FfaGJsGKevLQzAIuZUzRPgy0WbZUkZL+MvA2lrfdpWLh2zHcRi2
/FFKuqSOeTeGHk0Ggcyyt901RTnBYqQ77uVs3e+r9Y72i4ibxOY2XSYnwLCmhG6mi0RZb7P2Z/xP
aR/14i2oRQ7zBtfGCJy0dqnr+D2WGqilis0kME/QapLSuI/efA1cInHYSRuRD1yugr6G3PDj6798
xzNzSHRI9s7UUbhXZUJt0WtnAKln8LgcW1cpqt9h0Jvap01Xr4Z2r0dPPeFw/UnnS8YRfO96ZpCC
s+fVWUx+fRogRNOl33zeG/hKmzbaLrOZxrDhKvAVR+j7W2Zi6jZ4rtVdoIHuPq6fSkdVSOqIgU+X
2o9PDemNUZtMEdtlbbru+ItZyD2g9PI7xfaobF5ZaOgkpMGmVXqWR4XIcwiF3J3tu0FntHRyxDF4
KWv0TD2eT25C+h9DBFEyPZ+TueTnyXaUtUShP2TUWX3ozb9LmlLWEjChNuNEbrdTMuZRy0C2zTxa
9UhNpXZ246MYJTYBv9ew711CXoOoOjocYZ2A8tTZALrwYU+nTpay8kfsIhDcVYaxw+ELoHC+kjmM
Mf09jINlUEecGm3tIj9EUKuZbM11su3B1iIri9tB1i3UkleKJtkageUnoU/M5OG4uopkrJTuFfES
n5R6foFNU68dYfdp2mO9VTLNN/MdmQrTFBdb4HMY6QtNCkNfYeo4HvIyPFDUJMBMA0kMtyxrKrlm
+au3xlhNTDEUf0aTx8Usd5nVvq1pcKPcMcBB9GxXAblNBAMcRPcNEfx1mOSVScHOeveGKHfv6Wea
8wln+UawO+X0pTSBfeNzilelj9grYDxgMsLN2iZDhEI83Ww2grRkz4p5h2kkpT3osHRw6vr0+Myk
Hj97AzkLWMwbm7cgq/GfqkLmayEULekK2cAROrXSfLswxgpDdSbDEMfabJEXTWviD/vQlQyMQczL
hMTfRhhfL8sqvdURr2S6EZWV4Jsr+Xh6hQsAGCSdT+NuDkusgpsgRbN123hY1NVw0Cwe0uIQ4cMU
TC36XzyINXcxeGDuk9f/EdHkcJ1Qf8H2j8VDMUTRdyurzqCyTCf2reb+6/iUdoQm0BDx1ZT4fsuV
BCn4NWFCYjPO+Alh2S5aMOBG/ZuFTIzsUJakV2GL1FpBC0c9UQUlqy1XGkyiR3J5OnYxD5vvfXMm
xzIDHetyfZpbTwicS+NrmWFldHohZGUJfC+GkbP7YNZG6BECW0eNuuKuMbpjJWOCT/uHKemA/Y7G
8ngd5gIlIx7cmDdNSjN6nEOtpjzM1nZvwF6SXqpvCLrH+PjjXnBsKV8tVMyHdqGBxM/+CTRJtJJm
yP2xiBCLIVtcUgyKSbDhsPTp/4ozqoTgGW0e67E4QwROPjdZakDqoI1fbjaTTZvCLM0+Evu0PEn0
YWxVZCRSBEDVxrSXw5HhHO7b3GOBfQ0i/aaolo/Bgm6N8IqyKoKZ9ej+Hu/rlIu2kmaBXMjjhNWM
ZzC2KsGzoXIpOv5JFHS7UTpsQ2j7LB6dBYFHADRj1mEnsY10XU50Stt6WNVJrrVUd5WbqvlnC1/E
YoufyhdsjMuq6xBoc1oDm+n0nWtA0t0Az7xPZCoiy8yYF5bPVMk+f1dFRrU4Y66YsZj2CkTGNA9b
lLELviF0d9n0g6rYeakvaOwYLpv/CIARbcZzW80sqV1ApuQ/KtI3CZhrYYHsFXz4d88CG9JY7/uE
yJviMv3NEsUBD//URCDTEvKw9P9ZW6famVGmaXX1lmGy99/I69Sk4MijWV8ow8QxBPYpYxKql7Dq
0fJGmEupAny2OTYpe98qrXp20rm4NhB3Icn1Rg9Br2rk88PbmmOCkrskW7HCTzuizcBpS9t0mh1u
ofGNzOr8jC6GvVJu74c0WM8QSI/2CdN/qwZN2+Xv93l94Hg0AsBwRHJTHjO5qfEyGcnJ//Hhv2Yz
kxX3kfnB3hZRHvdIoWZDthR8P9HQFDRkfnuUYeOxUkJNMbkdrZiMGLK7Q7PPlAExgKPpUyiP4RP2
v2yXs9PlNjHgh/tpmRF84koOPNt/yzno6mo3s6dnvxPKpl5PtDlggJfwkCaiIgUceLAtZHwhshWf
bYsSAQkPUAHpyRa3+02XGWGJ5ajfReByD/kQGH8xyhv15L/fdj+yLJlY7LolXX5wuHSq+Wm9SDAB
9ZYa13HmNzSycxlslTeUNmCWefZKnIYTyYAgEI/hHHXFINSjk8kdXUDe3Dt19Z0t100PUaoiNI0h
ZFHCpxzT8AVTZVN9bOwYJ5cxFx80STmFsQRU87AnZLkoVKQ3iJGNqWQrM5tGJ7ZkRyqUDQp/Biwq
EJqeIWwJH77P4d37BibaF9RcVxAdPlA1Ib2VIoDwj1cXGjyIbC2UBfKyt1vpzxuvui06+k/l6sln
B7zUKDuETnAr2zs49GUtkTRTt+7uPkuaqIz1pVkdg8g5i0rVjEfbWQnd30Z6TyA4e/m96VH4GkF4
msKPZLPuj1qXOsh8Nb845GxGTwRkXaKKqfiaCdXZV4d37oLAkBBHapBHCNWPfQNtHilwAWUFiqzm
C3lsz/sDK18cJMAXR7tStrGHax17p7HmJ+Q1y7hAxrANTuG18d6Gnq4hmYOJpV+dVZPSMHkfIV63
+JDrbgj4dF4ZeKOFBjyuxK9O7O5Xi7gmFW41msh5UxGqABw3gdiLA20+sNGH9B0nlhueseZ3nyQc
TO7CPwMI9aGJT489UKJEo4mNRV/v2onQScS+syprIXHD+DzqWA0uND5QZy96JZc9FkO9x94a/1Z+
ISgm2b+hrGHPmYHhzJub6VBHtZZkX9dorEbr2hBSvbPrMdRwHIolugIW4lC1gz8QL6I9AXuD35vr
xMe0BbNV3Ow+StIYRmtzPBakSV9l/vLDwo+mic/repWP1e6Mftlr1Zf4UrfY9jhwi4dDtMxRnJOY
P7wte1Km1iGwhjsJEzlq4On5bzJ7Gjmc723IjX+Yvd37Jc8vC6zJMCrwRnYewRvBSTvdpWiE/FpJ
eA5EWomv64jp7Iya9uzyqAUJEhpNagSvYML0zSxB3v7RZPSL+fYQSnJ2Fojg11s0nfnih9sc2Ytl
/CnAOrsYAeoe1Bn/7IraogaylG6cX9OML/19gocKj7eaquCyRkEshdCAh5mkxWI40wagufLxh8uT
vvC8WzQCyn0l/CHPkMvrzNFsu1YlnCjdzr7zCcvUqnMbVE69Az+4NOsxR2YDOUWVxTDEQ4Zbt+AO
+nGrmFTDLsGScn3ahQkl7VCdqFWIeVzRU8blu4+y+ZhxCd1fTYxUUkiCSXdEpvU+pVNNEsyXXS9l
LnrM+9DRzzC5gf2Erd9+FGY1FrPmDUt3ZN1LJVrqKqVNqYy/KHTdghHMrjcEcs4CUAJQvnpH31UG
MbiU3P295b5+GSq6+ri9c8xVj0bnFm65K5oTpCJzcOrxRCY0acmyr67974uJIksoHOXofWXwuFJ4
XG99yeuN8+zuHpPkRrfuBdXWFlLhHx+gVlwo/FfUpN2EV7i5qzpv/ZigBZ99udGjd2hfaBd7z+ht
0FdPRNADLKsaevPxeWnm3GWqLSupM8yQgwPEdq0U7EdWJ0KRdUAa1P4kSR1tWKfgkR6NnNZ/ZWPm
r8ZHRk3xMcKBUJ5Opj9Lfkp3ktSWazRhKAM5WVA6xFKvEKAyBNbiI1axbpD/U9ZwdKUzUjFbtZ9w
s8pIo9AiYGkEHX9nMK6wT44oDztwaj9tmqH1xeN0+e8zlBFLK/IcngT4gGRn0cmMGkpUP/xBcEjc
kqh5w3g/nhkBOG9S5hvRthPQvl05JmrxBLQH7oNpQLoT+J4Xv9fjk2bdpqZ6QALanjNqTOzUQ66G
zdEK2zTzPYZF3ZZs7KglLHrelNKtYK1V1I1/D1kE9ZVA9EU1I7fySNxQpmD+pi0U2j3rngA4LyNv
Ir3rfLZYonoOqxkB5MLharFA5uyz49kUsza2o4ZfqtPZ3IQNLl9Om9Nj5MfKXNyeySuvsGH5rv+u
TUYsYiCRPQV2De3v/HVaQibr0NiPBm8H04FA+ZzetSUBWdGWuAr1IXEUBSavYvzT4x/LqRI2pA7k
zSbrWaiI4Ggmt5JpxGhCpGJp6jbbNcujCBZeuWrKwoCk6Xh52cMVCy11mDcl0NxVo3RXtrtIZBQ0
mTlpLHpyqnWTWAVse9FcgDKgz54A/LO08IStxA+dM7jf7V/UhsP+wpInDkrsrxICeRJv/f4PQT/9
T+uMyxuTk9MLoOq5EZCmzq4XN4P4j8ueunRwSYf38c7kv/1ATDm8k5FYoOVXztDyvZIL7asc9LJf
93E4IPNGbEJxkssbCsfN+NJGCAm57G9ifL3QiaLOygJ6ysJYLYuu2R90BH7DKH1pH5zOS9t5+rpj
YoNzd5iBhrQzrQb4WB+OXSrnNogO5vAdWOH1f8y1AmwaMmek3nfd0JMsLNNsVElOEyvYByEwbDYU
CLUuKeti6qGqd/sNyaIbh28aWl+yCs+dZ2/mBKf2RZJvsPUN+hK1bs/KRdYvhiLKHCF3anDY81Bu
QSOXfYgFjTeans4VgaTl9y8Ufdj09TpyXooqZsYHKCUhhg4KAHE9fhtjR+I/w55a44HR5RxR+OYk
+hFQKBmSPjFFeMbxJvQWf8L3+eVP5HGKb6sUQYj5Q7Xbfx8YnVlOWLkZn3obB+gPPXJwPYLD+XMN
8w+WOO3surWM+8UfeAxWZp1RjgQzTaW8zBN1S9ylO4p5viUeJP5JcSXZkc98UkspWDg+98dyx4NV
/utGsYY0fXFycQEBRVgkXJHsGTJCAHwT5KqDP/EJZwbJBHNNKwWiVixijZsV7yPVDKJL24xcs4vt
zYXaVquRbzF3U/JYRoPXz15yw6LEilqe74ypm4w6YxpWxNWFBZk0KfqGwZ7sFJumm0Mkv1hkoVvv
hN63gmSRfibBDFmxT0C7EcUkkjOApfc7Fk1DotdOZP1SX0hQkDNPQqEGJedh3pVH+wZFvIX54xEU
DM5ZkgN/pG/DuWVbS9RM7ecQeW3dvQFBsFd+IHXfmNv8H+dkolP9OZLAJhvmWGxx9FPT7VQ/NvA+
IGYkMgD8BOegRzYKkoSnXOZBBjYm+VkgnnhJJBoR13VM/TY6iHKisrqX+Zh6u7EpBouUx6YI10Eo
FPn1OXYL9A7vMAd6wAXDNiYi4O/ikGzyY+jPKFgqZF5uuvC84qDgUsDP7aWP1NTxR203u8MJwxSw
WruOD8EhsBLRcm3JXD1qui6xbVneLzkteZ0grhJ1y6KV0RPv07Wgk9nGF2i8fZ4Vp0Et3sXRS9I7
AA+elQVVTbbP1LF5UQqzHuKoNURRB/KE6/2XFm484Tj3XwWDTsPMkGBKkUWQbe+EDZPIzj4Hky/p
HXzU64x39V0YL3lhYIw1B/wI3ERtAoJn8qNQ7fKYW1uVICWUsL/wC3ueiUnc+Fnob57BmnHH+d22
bALKtz9YI5lDMFruMUNnCB2dS9oH/KXCeNykUYiF38+R06yE+qeg+Pk7FxKHMUNJtAjMGaJ+fCGC
DfMiFKU0UqL6xAT4oAghHUxQitKzHYtjyDm9OPQPNJSB92u6Gb07z93Vg+uKSnehb6CFaWc3H0Uh
Fda1ypcWaKxJ4JEPDYdcy3NWuSB0g0qNPNfpejoKlgTD27yL5t9wFXsazEwMG/Y2kIAvLdySmWDI
ARg4/1SiJmSeUXgcPdiId+KpKPSd1W3vqAuf3Gtg3SZCwjy9/YUfJZ1i5ggUlP4IqdWh3+moSLmW
dln5E2kl1WOYEmHuoikwmrIEqYuklUw3ekyGfGoIlWJlCLyG1D0Z+CO4vkEpYM51nHvrVR61pS8c
5Tc9lYAGOdttKq2j9b+EWRj5qkzfzcXd8o5wZgdynOnrJ1wK9QJ8YhjwE4bazU6S4XALkU3GmRSS
OK8wI56hhOzQFIy1l4eJpVdC+cf8rowHS5tdyR5AQyjoKk9eDchB+3fsr39ExrpERAIiETQTosIa
rsjFdpTjSKPIya95EVOv5cTETWU02gJWdIZ2S7MCCpWZPF8TkvQzcdiALLJm222mqhA38Gxcxmem
aprgRBaiV6hb2u26IR7qO1tgU+34fpGfyRKXMRjd6x13jzwyY1VzxufDO7/Bfgc/O9wi36R/MbeD
sRQD+y3VtfDtcvIRALPEuL2DBhWMw5Lltahz1Q7/t8fr2ezeA6x3XV1HT3JArAP79EzAPab79e/4
BStKIpKtX9fjnM/E2/jk5/8hO+XvEIG55+eJvzhGjW/MkEa/38R/JUOdOdb91EQDKckoUOQeCrG0
M/Ev/Ck4S7R+WiYVafg2/dCAD3JltrcIO5BlqSCf56ZZitz5oXEViBYU6yvr3zjrvLHzsl5XkpfK
WC899syd21A0LU9TeWrsXKMPeCrhT2uhfZxpEJ47QZfU7Nd2tQKZkf6t1hZosdKKuzMolQV0UAdT
2zjXNcsigK20HA0/3zd7javtSgHRaHzpRKQDduwRI7sknqXkU8Xh9VWip4v2nAAE4+ugwu8oD9UD
ZOk1llfAqIlul7gou2uTZ+nWcyrE7iRFfBRhf8EHhpwXCE74Hxd7Uu6obTT12z5dEEwKdRGEdsWn
IAsP5gVTSMT2MV1jhw+akwy8wVqGsJ+vJ+AfE6frat1y/JOYoGks+JuUtYs+lKVmaJtBw0GM6eZk
TF4ZVdZrT1eTE/xYeBaa7GMEqedEX3cY6SorkuyXXJNxREYbumHEk3cNffZivyYRhA1BpKRGvQaU
T+/wuNTgfjZUuuc0Ute7JKAUKO3T/0WucRKwO1lVWux5bwkJC/TScePcWfSOivejN2jX+quR6zfy
wyT6Wy9Cv/R0qGpVGrQwpf6NtGVP1obV1LTQTzQkACkKV/+MHFpstrX+qUaKPb5vLTJ/Ke5YlH4S
bzC2CO56JR90CQ3pDHpd9d0nRV67waiqDU9UnkJXBAiwU7RhTdx4i+s6lQ+/l3zC0wWirAuJ7mIz
NAnmtN7BeHkhFL9KXwUWk6fs9Sxp/35mPapj8hozmdrIDyA01b4DdNxWKWP79DqaAEUdsk9fUv5u
NV8EETty6bOsazDgqGugOjOAGweTZiSMxH91KGp4aiOdLDEYPEa9uLvMZtpDQFkVnp/q/uAsTYF2
/0z1HJU8DJqBBqUSGkgkIMrCg2dCurLt1ZOKReY0lYd0KzGbk5x/SGnYmkNgSVV3miQsPa+Z0tOe
4/BC0n2ODyl7ffqh4nNuMIgM+RqBjFX1fIfsqN31/L0NDG4SYWHJAuKpcB1Du70qr3OfaV5VS4Bk
uBD3DhUHMbI5+3ydtrTI+e1kHC+VxVBOkgkFvSNX0BS17wLx1WEf5yX91CCinz+N1vvhhuILAvAl
7C5LwaAy4zYnvUh+EwyPdIpgUgO0w8+CUVDAvjYHhs2yhyQn6DiRy0/SGULBV2uLe9LU/G4N0HXx
bSgPMPhtu1lFDCSu0VStEHIb3O2tgjSiVwNbrB3DUTqU5ehrIeCDP+mABZIuHEGoyImmXS1aZypc
vwIes7IFbFIqEMcc8iYqulJCsRM5mVFDOB3+tTKMARcfL6fIIgert1p9qxV6CrvI1ohxA/S5BtWK
pZnT8opIPLNDUhTPVg1nsB6Hzurt1eTB8J6z+O6+9Xs9fyMUj7s/6sSgGtwyZxKD/PRllW3yVmk1
iYGGzV5dPt5xfqA7z8VghyVy8RZk825IZ8nUzcr4FtVY+eexz/3AoGRM4lk7up1K//+p8ZBnxOT0
ftAcfdzXB+m76EegpcuMa9joKeCbmO/sETUZBSMu9u5rWf14v09gAOlwEYCE7+uN7tzJFJDDrVFm
KUQcHTBG0c3QelI80LD011KuV4tGxWov5uI0AO+VxLBSwmHinAFI3vePJ2Npxa7zdq5NTVN2EoWn
0d0+sexQsPKN9bJZ2VA/rQFKPl128PhR14hw9pgyEy4nBB+AdEyGucc39d+OOHGBSTvgQs7tNVZT
VbB9dnlYIOucbCg2OQYKbXhXP6lw60zFok1Fc14vDKTPxFbKh9Te12Yc2JTdikU47HDtoQV08Oq6
Q1WZx9OBkw/A6OGrXd/SkvQD8nAnQGhPrEZxotyDP7TCA4dyHHZYMP5TA9qY8/Sl4Ylawout6N+q
FTthvXIpNaBbu0cRcY6WFEYq3SeZtsCWA6PGGwUo5ZtpVjU+t7ns1jaVQqig9yuvm6vIiXfZPlAp
oIJz6tj1MIIJ9MtxSnQONmazQ/8g7Jo2RYzG/OagJL8wtMNdNG7FZJyQiplWLcEytdKpdnvKmOsn
jCjpqoqm1TSCjqvMyQey/9CHimS+7sn7jGgxOt4BWzl2e4NYpMWHQ47p9q0il7KxVlXvChd7V7dB
84c+J67pGjznmpQuMh25+D3nDQxgb9H2iOAPzUolDQFD+z3IrJWE29XcEEFvWoUdIFULrKw/vfCf
cuAYJtJDZ/d7mucEC0/zhYcf44tZ0Pw56J7Cpo+0W+IVUMhXCedG6A1Qp7XoLTlkq1pAhoNLmQQA
zbiFa0OdYAvp0f0Mhy2BrluBF0WdfcZwyXcrKMj/xxR01nP9gHbPXsJ3F2tAL2RQhnU/esZzNr44
b47gJPk6FKczGbxl0DtTDJuv9+YwfM4/Mp3BdupKacCUkcS1Vz+6n8PglTUJC5ZURoU8/DQZeSMt
dfQiA0OgpthLMiqA9wYiebZ7wUJ4XfXe5qWAd5dvtME4otfWPZ+R6nqnPrO5sRABaIyD9XGVFega
e0LFy9BMfShsnHjb8wYkyusIUzyU0Jx/WTYWlC5jrItB0RU+RbRPevkeLSmCxvETMa2NB4giygPB
7gtwt3FQXNThSQl4sJSnsv0H9wMjYq7VOAyca1pK0oIW8WIauE+EzZ3Mq5WyE7rZJrWzFJODMGIM
6omSTOwVOeb55TO4gpzSLJA2jtI4UU9a8q18kqZyRuaGmBoWM/Ora5wdy9C9Fo3le69cEok4tQBi
ij9DxZzayth8BePG+kQl9qrAt89uGTMgsgh2SOP8G9l9hoF7v52KJJxN3B09uhRRhJ/ePrxb5qig
InkRD9gSue23t7o3UBW6KqV3pL8ZkMVKMVTRYtD810VSiKX3jZXqLpmSBU3EBTEK3Q0MpSaNLwPU
JgDSHphfCbLv31661kBkeQrQKJLR8aX79Z9p9DQcfZ4WC4s4sR4nxBmKA5AlHROXAxplPQdmVyL6
3/0bde8TBZ/ErQIAwch1LQu3asnjHf7cX+U4ywGKoZkUzlXppk2GUv4Ca1MD7Qb7AY4esyubyHDO
5k3ygU0Esq75V3jPR1Du1iNiUN4ld5oljgaWBSRKaCN0roh9HpMUgMDTxR9/KlRKNhOnDBKiDLvT
X7bG3qaaV8uUxrpMX8BeChBTrKzoY8okWZEUiQHW3bKmeodEGUBz/NBzh3Dk+K7roVDngXwv3r2a
K6rEE+271bifOBpSAKb+MFwvfZ/7JepMpL7RoY2fqWDBrzvR1fiwJ7k/RgJFJx5btY4qXvY8RBxk
POyW4CqD7aPpNUoz65r62PR/GerHQlP7oq1Ab6qO5xvRGsRAHBxQ82ioDDb83MFafRkbd1JzaTDC
YYA9gcymRNJtpNy5VaMeau9UHM2uvEbvT5r9r+3q5+3dJugK7Ah0lpXLnIy/VAU8dkBYVYQYjXbG
T5W+8gdeeJcCb3gAl+xPXods1xy3XasreEw2Q1O0VJfMm9hUL9fdxCOkrEPf3xbp5Inyvgox9hOW
++4ED697ZXmifZSbJHp5pEMOvwZ79/kBJ2Jil6h9Pe2/uog+MAb8g38CjDiR1WAMA/Wz3TqFimRQ
4EKsnPT+XGt4wCJ0PYmpA3N6jPsAND3GcYvNQy5aZuZ9QHvHASJ4zostNt5IkhfPJFGLmOqJqpm6
V+ypulNrT6uYURBY9uDg3xp9AU8sgMCh/vB82X/eCiCQ6Rn9fiWIzQ/Tyqye/RNxlJiM7GZ6GPgo
a7GTTPDELyVrUcGjHA6smZNlpzYAKTJB3/CI7dmIqkRagbcZH7mIMJhwcFLLKPMIkkqXbXtgxwys
sZY4GLG3HJwh/8Lz2iA1adL6C/gyBS6a7Qp2RC+6rSt/95ceE+d2dDduDsSLlTSSpjFFnyrYqKuh
mAmMDSJTTkU9cR39/bcIq8YlmJDiZcSoJPhN1RpioMHVQ3cYEh9Ytan9TIt/1toiUy8aDwFOwu0k
bFhSjgK7AmtWm0NIEonckNSZrYV8UPRBRqH0zsnsL2e+01SBAKbm6WY70nFPQfuKNx0aCxLQUQi2
GluGC6pxc257SATHBltH58Ocqis05x6H+PCamxxZfryW/t8cHjHM2vnodsp51orPH0SLcujo1HzF
pWn9vt/caOOmjpa0rmQFksiBslggLKiBal/w98O8aAK2dRSCbQaJ0sb5G7vWMcCyeVA2hY0092+y
IM9P3IdmG15cI5kKtG7Y5ko3lxZITx7avm6lQGjJmffBAsQRMvi4riyOik03OZwtwUBjFds8+xyz
kE+SRuvpaZw7WwWfOgMWRSkmt8H232Y2Fxy/I+tUvRak2buzBNO9RpXyQQCenorjKWGsLlqJAwsg
ICHi7qCVWkxqk/k7+6QmsVEgVR0zW+RDgrUI+9x0HKc6g3F2balRlX0PeBIji+pkE1GzUQCjUqT+
zZTgLhAwLEvWTL5tZOM5gdpob/5M++TMX9lLhXCLLnRJy0GY8Odi8VJWnCwTKm+EKl8LXaWjnrVn
5mylJeky/m/p3lWUEInzyyeX4/7GCDxrJ/9dv0HE58E0K91cIqlkeZj61BOj0Bvln6Kr5YezzhiP
Bl64mU4EtfxRDdJ6La52TKacLmmSG8Ta1mRfegHIARNYPFlONxwszIpn+9bg8nY3eQt8NYApWrNC
Xy91yKN5jMtGkCk4dFL/MOKgl9TWVDqZkgy1uv2H9i/ycCJ56JXcYkczLoVWtDnmlcMkOHzSh8I6
H1hU5qYw5egGZFLOpaeQl1in6a8p1JJyzPhQt8hvna4UoUlcf94RM2gYWhRP8mdzUcvyN7SPyvk0
8AF/bNUwegI0cDvgjqunuQwqx7ZWsoBIEAS81qzOkqiuwj0QO6KfvXLIzdkOMJvGqk70eekIPBoY
mQmMEHh+zmXBp7Lai6bZ3g9FM3Fx4Hw+eIKh+H85Ixp1ciJMCq7fzHJ47WE4ve50lfOcyvRp2dZx
9I8oCuPm70bkSA5ws+rNa6R5qohAiC+gw93kVnhXGsUSp7I0l8f+5h/U1raEx1QDelqnN96v7V0a
RGBiDfbhwWnGOQ4y8BsrFJnjV/Y4arQVcBVio4fAoHRdNrTQS74g5DC5EbTXhPx1HWj51rkuPjE2
0MvL6eMGATEJWR9kgTyH3nsYwb+r1gmMFXY3P4vM0ULUgvTO3Ip5gTzvDJbiZMCb1j1fAMtI9a33
+ZYUb0HCYPnOTk3oaH/Ty+JDCrQUCeA/HkT2NDBPokGQWoye8ds9SqwM/ByYjAdsdsaP48J38KAX
doj8ly4I0G+908BclojaKtxCdjzbVphG2mnp8eFJM9Fr4ZyUFo7ePrgjlvUbPKMItRELzYCSQK0R
Igos5R+eJ5+echkv59yW3t0jmmh5UbXjb6Czu3WA71UmXbpmy4xobUyBEL2IaDEOttKNuLLLgPoQ
xCgd/64qqfsN22+eEwjkOVHGuJj4MfdVg08wtbNGM7b2LcL+Ksxn1WCyRiRkEW59TIsZic8EIAXu
kuzkehFInU80jh2MJmtn9lxiG9nntBUA/jAtCcgcGtPUaOBsJukYEk14F74U5bPeQdyk6/rpRBxT
e1+kY0QQZAMx/FE1mAbc8v9l/P2sHKPog2UTrhjpCABnhBQMfM5YQzK/S7VvVs/I/YFIZS/dSxFi
ueIOANHrMiM1PGmFbg9W3V05d/BN+Rq0pjgFrRfO7VxvAMpdndTQSSVCpIWneZ0T+B3LZeLuQuWa
drZh9DUMfc3aS1Q8salc+GWng714Tswv/VRXp5DAZJ5XbjmIP+ajiQEodOHbUPg9MDSrURo6DE1O
PuoOeteMxTcArNCdD8zhSPMbS6WgOrxLpMx9m54AzBDJh/M9OB6DM9FdDCcRKEhxEBkAqyyKtCef
KCqlT9crWi1Wy5wtGtiQgDfm92QxDalbxEDK0sZnDxN8W+EuRypha6Iw9ykqEOMMNlDJRRhhmu42
Ke0S6k9DsA8CPqW+8YQkInqh+x8ULrFO+nwD6ViGAvPiunIO4oOf3LVz1XTQkMLWxuo1eHVmBKnE
hFZGYSK+RQT2CuunB4nPGnQgnCbQ0KHEeeflkACRN9oI7/xdXr3aPgcLhIA5afyPhnK+5lahJPKP
z0FH7+Df6NgTtVCXRphudZXow4klMIcHTx/KT3HNh4rkceQntd4Q5022rLQ7Gwxhw06H4MHpjER+
oQA7C3lYhow/bzjuxWkFhxOy4BtyT3ZiThHmAZrSs2/0l8ypoETfX5wy+W1megctpfct/Y9nWpdX
BiGwWEjtR5lCiXxrwIWfzGQYZaf8M3jz/KBSOthEbhzm5iv4QeZDNxJ4s3Ha7oLOslMQJewj2OLB
PbUJeXe7QybebE/JmmrP+dLx4Q7eaJ3qI0/Z9waAx4e7+5FhQx1Rdu4qq8T/7dz5quwI5y94vWNB
5MUQnrJrv4SAUloM/9Itwxma0dN2lg/Vr2u3v8Oxpc4ZmGFt3GstfLqvzCBM1Aa+YXxVDIslrQ8Q
CPvlIFLbsedKW7xf/5+L3+gRsEdj63Anh86pEubk8GDtq5UttjOgQV4OKBbsp4KePDdcq/ynm9lR
dOtK+5LGWDxiff9i/Zm7GNOsvWpgSpm4OSo5s592bqxPDHE6+PCSje4rLvPVLxSaK1BALx9LSVYy
HFfmoxzXPFhlj+vsvK8Myijdv+6XE6IR08myr95W72WwHGGKkHEYX610Ewh60092fb8xUbUiP+Tg
FaENFldRE31pM748LPpDh5PKSyGuDFzfMXp7k6eNZhjpNmTql4fxjeohlxwwyYwzN25iTQZnqAbJ
EtR3OsNqgL107f/Wa1l1pjiybKLViUhMawyEs6WYdZw5LsF4YDH64bwF06w7fKs+m3NS3M54dvD1
Yyg2NcVv1xp8MkztirlDPNm5eSxg2vGuv+o+usXMT1I9OBjyI64Ucc+QDPHii/dZ7uIHxdXecMze
9I6zFZFTCHAdzrH5zKH3wlKwUV4n3gXi59UXsW4+27JPuNOXIDoEmT7f3VOR957CHClg/qRXpCS4
bPr8gYDhkdPtZgYyw306KoP7Gpw1VZkGWRl9LDCjGKpNJqD9VunWdc2Xu2I/ZIlYy69JwKtCfai3
nfXNT6VQ1NICGP9ZLp8jnks7SMbiC/svDk58c05VU9dxQNg/GDlIh2GT0f3I5pLRi/9JfXRFh3+G
ciWagSD6nh/4NRtHEN4dMx3sOwh2/6J7lmwAEPuUzHoZdYeQ5vx/Ekg0R3DRhkSQFVeiK5a/N5wo
5qTmh0szehOnS/lE9crUHO5Y7gmY1yWOYPOzD0SUuMtSed5oGU+HhgWihahuK80yxsLGwuL6BVvY
OJNUYK+djTMg7My2+aurBQFNG1SrsjB8i07yyvauyKefgScnZBYPROl+JXrovI5I8KF85sHh6lRV
LM+q1FP2ZCuxQ8rmE/8EeXjX+2Lib0sAh0X/pqB+KVPUeqluKg2QRZdMHjmSJNjvWnvepkeUm+c1
1n1f+cyCuiZ28gG4HtCVaaHzIomVz2O7jp+WSMAfw4pnI9/fuq7hqrsmE49DfHXdXY5HaJC1L+hG
/8/Pv8CvVcd7o99zhcE3jstx5FQ4cclB/gP7qQbwGRtODjRvNW0YIqkunM/Jj9No0/7tt2YCC0Av
fbiDLto0huJYHX1FL6TaIdcpzIAPNpT0n93dDkUKzt4eWaM7kUTTVORiWBnBU913HMn+ofIdUZqi
l86R6hhNp/0px6o5tb/NM9q1M3aZo/OSWLjkB4ZG0Q0Wwu2yAsoUCL0pAzDgo+vxZdukF+M4qbQc
1ApphxjtiWAJNWwFwuf9VM2H9IM2qmb2Df4efQZD88lcOi31gKS+mAxMFTne7qPqj1QhiLnUV5ha
eaDRnX0BimUeok4GyzAhzG+QmnMSuTHRFft4q4rP/k4KMgVAnBK2e+SQEVvGLoBpZxgncMm4q/AK
RcnekOpTwtBn4DcWfMnweZnBLQ/aL/9NFQAZHfLNQkqYZz9GIawK316Swot4CCVqPc96sMppBY9I
+aT2kMOWHYecUUpLenqnq0bGvg4blnaT6WJwjkAfMcRPU8Vv+u064KHi64vp9xbFO9EZVzziLqZk
WDITqA2NOW8FLcIpQPYjeC99VRD02hW/2kvcxB+5prg7X4bGQe8yJix8VV9nLJy7K9K5GEXtfWUl
2zV7dd4avGgdjqY07eqIcKj8R2ZkP56ATkwtAuXkmoUDd1xWktuap0DxratKJcT0Ok6dtAj+Rznr
EMELk3tujvXVGocnV7CK+hi7MRbxJ5LeckxWWGRoaDSWapxhKFJVO5CVblEK8oR4VH6QhnK+vuMv
8Zy6190RwsURg6Q9t3rccnS/fAalxq/8ZZ5DCLpEpRsXSvd+UuPN67dOs8fy3Ee2faQm6T4gYowr
DQQaTMv3A2Z7Lz/BCnpYJ31ULODiLQlAGKR+9c19diN62M5ijSjo96Eh7zUbhmGdGzCjERTkYM01
RahhK6kSuvyH47X/Ra9GDGA4IRu4DB3V0QZPIo7y6cfe2UQCstqgR5P3uNwxsGIiVxlbKc9/ws1A
hrM7ScJY6NIXDrSb4QnOSGeJXRQs7e4Rb9DS4Y+6pRHXWICbP2eNpGJznCtGRNmxDRGKiui2Tei7
OUzfIBYUWcJ8QaZU8UaMknlJ860yqGdpJRrXihXlv0HkfTG4x5bffqiTPods4a0TPZw9LT0SeWOe
gNZcd8SrwNYXuC9Be5Sj35U4ffA7PGVxYc2NnJD9uF5Em8MkrSevQUerloGoqxULN771zPnXN/Tc
iv2dZK5+mBPwy5pZweFUwiHeTNId0d2UtaPyN24gYDOAWr/dccUYqbB88OgA4Y+MM+0KWLcJDDA+
PCdr38lH1aBu4VY5MG3XvvdA99DZdNpTP9wXTvRR+EFwctkSFbUXFpRH4eK2TfHTMoMub01dTX7u
5z9uBVeSYiFzsS66uB6zNok6BtGezrkzmotxZDMPOAZmHILPkbyJae9/HX/kc+oLjO2VSkT2REql
4hJi9urKdt/8UIeg22eehP5LlN+vxe+Q1/LwkWyFiDVYFmVHHZQD3N7a4oMLQTTj1H2ZWujDZr/J
BlhMNniryfQ6/JpUfRTq032CExg565NtgfBEJFm63j47bBVMLlNgNdFWUbR9ZI31GOPSy+599ule
WrMD/WJOnZndtqrSWUjMA7M4edRpGk0y/uZ8u9pjABUXPfZnsePerBJ6RwgUpvxtii9WW00M+Q+n
01tvNw+fG3cW+yae/XXwt8+EN4DqJTiDKA2kmSHW0X+FlHOUoMaAgEsYXCAIRhUgYqfnMTv39SvR
qBtujms14eqlh9J+hSMsUK0Z0OEs7xeGSrKYGi43k1q0H/vJ6p/P/51pVkK1WDQhK7EhmV0b34IK
oJYb6smqGH47chEPvPowpie9KJiL0D/ftzWjEpzG9U2AtntvmoFr4CBw9PKSG3aYPDVVJx0AN4qh
XxMfzmN7nffO2ttxOKJqB/bk+OLAxYuM5ref42TajmLdWEWmPcZChf024VfpvXXpQnDFeVYSg1Lh
nONGTqM/mXkvzEDPVVhOQlvDRTO9zWhPYJ7uMyOer9ZR/dzhode/uF2lWCbOSeq6MEMXQf/6zsBu
MBimKqfadXtYD0psUNXI6NyJX6x8bKJkx4rBWBbcJ4ILYjdpTsJ4IcSZtI2HIgmRHhuZ5QC/+759
xlyVxqP28RJub6VvstCfYW73XDW1XewGsEuS0SeJvh7pr5WbOKxbDFkTUlJj7quCNfaJEwx2ZV00
cNh2dnBsm8nkySU/KtP928K4OKQ26C5n+1WwGR6+OCRYUMyGYH1lFhEEqbVVaAUGkzp6ZuP1jO7E
w+e6XHtdiQIAS1M+zvQIjEfOMFKgPrS7hu/YOqzlEeobP3rUeQh51e2zs+JpiB24wmVxug5UuDdo
DBnKwTKOoMgYHu3ZQLt8A5oTIaT8ZVq53lIXoto8TDUt4ZYQCwvLHUXDcM53GmPKQmac93cdsabp
oNbhtyuSUAniingfAfLsfEMlSUMB1YZYsn7tuIwdULsL6YXyQlHHophPmzmihOo7jjLlG6Jh39gk
aFMGhjDNCN5DOYvh05ZJ8fWGq/68iCi3AxiNzO2doodc0TOwJXnm1jw1cbClQuVdlQA3hUjHn1+z
6DVuysGssctfyNulWr0UhxBEZFQoMbh32SZadyhlVt0QAJlqsr9uPyEum8mPPvRVleiEaAXWyQun
h6y73M5IjtNIAVzirx4QN4YI6SuMqzwB0Aq2L795UGhWNigG6CpYVAcZtRF1UxGeACXZNddNmMbs
eOdhFJTx9+SJkDIrbEa6ZqHz1r8NbL/wee3esBk2OGorfOG1rnfkAA7gkXiP2ZEb1dLcwlm8dVl/
haGm+nltgnC5btY4ZR7iDjGObdxxAb+JHK84e78XNfQJ8bhYjSxGNZHpK/fkGL+1GOASy3esfe+7
zoVPZXVm9Oe3LCdzQw/9ltFC7grd5z0ZIm2vN5ThJE/lamP710ZN4jmHlL/fz7AXwIKMV58BdIT3
5y2CcvifLMoMfn/KaYpWFObn26R1OSA9oncJ/0WoD4eh0HOM4dkqO8UaErTWgtzA8QafRExItR1M
DMUVnmKrrUNEVy5/jDqjmP14zh+aAvtmRz0GBFkSlbR5i7eECz7FUwdHobIrhFVaTwCym8G9yXP4
OhEk3HgzdWgsc3xww9ZEl2yNrMYIv88RFttRVsIfA2xHT163mksfordCc3Jvv6gxOS24CKtOO9TY
CgTAouC8LO/eDHbWtN1Uk+Ay4S88SoF77utEQHEN+alwVElLMhJ0/LCt6s6Rj5lr3eWISemV40c2
o82WVzJm2tP8PYpy+iH+QLlKXFiym69gnLXZRejKpaCzbKXqBtB+iN1rWvJlkcCFpVZ5dEgPny3L
DedObKvad7M7SEyz7FXbW/p2+x8i8CRoobZQhZOqxSq7mCZ9JQpatvgQyZMxMrGT9UCpah+XCJeF
oig8u3/a4re65cBH7YzvrUK9twSb7aultHy9D/UaIebQx3/7l5l6T2LgYLhuUs5RUzvLvjHGJeaz
TCVSOwaGr1jPTtusNv3M+i6uCLqpRifCxPNQaIiQAT09bXkt2Y6YVSvTkoFHk4kXpjVsqCQ0f6au
7rDHC2/ZkhyQrA+SZg6XRf9MRM382FhqXV1WBbCi9cpXBRKXvIlD4B67Q74+cUh0cTpLJqstPbEU
MYGgu3z5rY6R1NCNAhFtjb12whq+aZYC7UYEIn4af4Skcd8YNa3kA3vo+MUpiwN2ql2fZ4RjBRcY
L9zUFT1K3KlEBC/gdXPGFw/jC6T+bnfypWjl8QsrNNvmLoJK5yCfTob9baHnPwYG7EbZdWisrzrS
P6IEznT4q6lXalpIs74ntnE5foJdaAEjUcEnBvaIsJVLBQqxrnbTZVPhX1fWORl7Kgt/HztxZ4Zc
Y2eX9DjhQlaZBaFLt7ysy57zM/CIdSJ5Ov4x6/oQnjVg2KKhmYJJBJgxVLITWvT5NjkVR2FUzLF8
3snYSsvp32OoU58+m657dSRrzWE/I/Bj1h3+mQwuuBwdP50kW2I0Ywiu501zsldrQaRlr96KI1Tn
VCgK0WaBdFkQjkR3S7+lQcg6UuIvUU6XA48uldg6/hiEvuyRF5opZsEqqkESiBGU4NzS6T35Kthg
Nfr59DAwt2U6sddjDGv3mkpYICqTpk3bCBZdZRKXWeHRuNKAFwBLOvehkmQucKgik5btVnntx75R
qahtCGbCqFVLwaFR35lpWk/X5XQXuiIK+5bY6qzi7WJR+SExCxeEj/1ylDMOP01B819KqXAlAQPM
KpcxTUF1kRwQEqMOzxe5pOccp6o6+oK5xyi7pHRFNmLLWYToQbS9W70ZlzmsCIqHLNqa1/yZBF3O
M1q2Zk8KiNumksTP9CFo7o0qFHy6eLv8WM1LB081fctlXRBhNuepjIAYEJ2jI7rfeJADEs3BqNVz
Wt+FPtCebtczEHFueHGp9skIaMdt5VLPZARY/zpzo1ap6QWMC7P3Z56cO5NavVLth2KjR8ZveDnJ
lB89FLj1R8wbioOgi4utvdORU8sbFbtjcriEcRF/ZtcDTZo8+OINQyN9AMYa7j+mapaJbgi2CBCA
yI/NFOtN966BWtmJWTsq+B1S0BgCTHscE95wnr6Q7zY3bnQf6W9uoyj4SZSt9Qn/eLl7HuCEH8Wi
BXibeWh4SVSw+nt7ZPCx06up8OIZsx9BOdIZ/AU4jywpVtw9R6pqR3Fmnin3ghY28PXnyAi8c2fw
zSJbZ9u892hMQXXerOCgCV4Bvs5t8X0SE0Y/UipZjf/Tlh9JCU1md8SRSX7Ai7mvAfyxGkw1YHWT
OZYj8j+naA8qEoCxlEamTvhfDH58OT2a1NE3uvXZh9NNS62xRbXs6PJlZ8RqL0QcRsTp/IrqJNgQ
pl82Soq8JTXlV1GQ9mBsCDexViVUf/4J5QRk+WckYnfPB4ZRI841x4OlLLGgphaen5LR/wz9uff3
Z4YdlgzdBmLcus0O2vcyO3kNJq9iXAhHLLW8Bv+YDYlesrZBwU8zSwq3LFPriDoCpt2KrMtlmo9f
5EXjVFZUVtV/79+ZYb3ZsEiAnJfok/FROI8xg+cFoLDYX4Y5LbUb31+KQ1Th7X5zQduXznw2Ypo8
/XlB3duH0MlQt/zdwLO7XlJ3nRPV683XX/yZobHCZPJFLU8NkkQxzLFPNMdrC2UUYxWGi/+/l5OL
HbtXJRMHtCZUmxp6DxDm4Zmltwm+g5KbZfCnhSEzpHo8/3AhfiG0GA33d3T7WMW7QAVYTiUhPUVo
jST2IJP1b78wctVctgycbbH+opJlPw3CvYR68Q3mJWFg3W6iYWsV0ftCnKjz1TgOYVtzAJgVEtuR
EVnDIjpG9EcRT3u05UTHm5rcaRtpdvkdxayNp0laPhQyS/tyEwYkQVqTQNghUcusBG3WWL2o4+xw
xNTE9OeIz5BTna4+WzAjUz1cfTY/7hNPLatSTlLGE5Nk70YrcJiwrfqkeEEsIGAnD+cZ1jeCht3E
+xiteHec41GDmTcOWnxhBh30tjiYo1Vv+OirvFkPh/yJzh8T2zW5rX4kQRh1BJfgrIJREFHGloe9
0rzmbOvXBgSUUZpupjYz+Ld7oyAbwYuYFppr61MoqpMRi34mwXfv0K+FTl/DA0mHsWIpmYOqWIpx
t5mbIqpXXYG499jJRnpAZXAKaHYY1j9RRiKgWqvQWTFrEO4cTbloP3SpjyVQG0BBkTHfQVqnB+S3
A7oZNB3I4AIGChL2ffs5Q26dAiJrkAmHzXZNMj0u+Vmsq6ETNDpefNdG/OnU/cQ2E/Zhc9JuEASg
Hk6/0+nHRwv1fY4IsQMbuHY0qLxnjnsKONGL/mTVtGdpZKIy8W0faXuCEaXrHnJkRAi4yygdEgb8
h42T/WmywcqTPqROC1xqUId5Xale8ZzOaA++BOek6mntKzR0ABXwJ8E2thBhdLAxRx4iEeSsYIkp
pEO1JhS3oRB0sb6Up7vmWcDSoyU1h4djp+Ds8gELbJnAxfbwDM9VTtCXDVKm13RYJxvCyLjL8S2K
dv85rQVbn42GorzdipPX1IFryl1bB7GBjfEFyiR6Pq13kNaBdKIq8/CS7p8De2r9ZavQG0rhHRBh
j1g4+lKDwBtEifGRvPZw/d8+n1+VEpeR/X4P40YGSiWGk0EqUDvr6jhkkhc5nNthUOZxpEVXGnVX
X0MAmlrvVungL9h80IKi3VU1RAPnJ9xbsCYR7+O9+SuTT8wFjDRc9xzgPR+9xIe4FHZUHuVL2Tsx
ledU27N9vKQnUqWkouPxvuU1xSutamJ9gOEH5ML06CWU4F8GwONItY5ggapuGOPRpL6jk08GaZIQ
W/4kiYv8OxItJOIhe24V0sCBOfO9N/lsc/j/2yWBAUpPsONAvTyl2QBeCigAk6TQ1L4U18oHid8q
mEptAIJl/4QPcfVeFdXtrMCbP3UZUqLS1jzIYNWdzTmf40eG9bUe0QoxsY1FuBqnwquczCobmp1j
tmFEGmSqX/6tvPlOiOYL0s+Zc89fkgBS0cEzNd3AMduTjIk5WT2P3vFjaLCGQ7gHx9DlXn0tNDf1
rwUYVD8DF89TFxEsLIXhhYsg8M5E5CvknkhKZuhQawoUL6jdfZuEsV+AkpX3x/fI3rKw78+ajnUm
zGKDARbllPrQjUmDN6irYNwIxxJoIOYx7gWI5+OWqtPNM3pAmMoLza+TwY0AqwChYiRwCKddNlS4
VUfcvuN2IebfXa4G6sBPPnL2P2pj8ZT4ZuRjYMNFoLnDyWZPA95hXOuSGp7GTFEulYtb3cxboPSr
F1T1yQA/hqaa31bK0qlqxdwl4Pg6fS+G+/X+ZGOkjesRPwllZulY4Q35ybwznsTxo0k2d6DM54Zl
quGqiehYBynBa6Lz6Z+i5aPLb3pBo1oXzUbEhyh2AWM5iPEke7W19VgEupU0y//ihBbKYlK9a4Xn
yoIeBn4bo/z47W1SzVYGs9u0hvGNZUPK4ke0JkMXu3qwMBDxnTie+eeixrtNcnZkJNAiXg4L2R+7
UCZ+lMwEJ74UG3hyCs3dIFOiE8eBf5mitqqWACP7Dar7C4/NkySyhN4/1JZnLoi9HgNI9kXLG3R6
JT5Z18pOE/JdGWq/0uNjcZ5mx8hWtOxUlJV0Fj+S80r7CtbMgKL0ypsW/4uq8AX+2Z6B45FCIDkX
BMGREf6ogo+6tX8OvHt23ROGXGKByCgK7uIKyfslUTuy7F4K8nKRM20Bmc+vaxH/bHlIQnlhgTep
AgfVnDjCkQaUKMbqhG13A5UlboW5leyyvN3c0F7KinbNiWdYUl1pF6X/FLf5hT/DBqnDzyovrkmh
DIYF4ax+HqZfbFVZa+MRWi7FK6zuEy3Er3nK+2tqXIojsgp7iQrZU6RsxgNDN5zAFV7wFiSKcyP6
2nNqDtgd0xPKUoq9kb0IzyjU/zyHcUthRf97XtePjOmnUtmXOS8MropbgTC6X/AZ8VXLf6rfVmSy
CMCN4kHY+fs89qDb4P20evzDEDhJoUuO/BJZvcDLdjfFyyLnwDxD/NPu6h1nVAxLLjLYEnI4jvpd
WQYw8yHyfQizAsoiTa20laaI7VtN3BW4mnE8BGHhEPtZRSONCCSgDtvuxdHsy2kqQgXGurl4ORxI
YV2XOJQVyO11TJqvnYqTNc/OlUnVEh7EgryblgnizwPFC/iiSqCWavIOE/iyjKat3c4Zz0qyydwk
BNRk/R61ZhQAHHG/5eMPjkB9v3qdt30I2BlT1sOhTSU66KRGAdqAPd4TY6bF3amx6OnS8Cg2RCUs
YBhmn/TsamMWqzd4198q+Tm+aDHe+VVk7np0BU/6ZkJxo+BTuAAUBR7a6yTbVgFbXKYNTxfmDoTw
YLPRA4tU1nms+AC/oSAs457pauK20rem3nD+nVZOXXFKCab+CSxRiDFmBahWTD30su7VU8ElOAT7
0UpL3pExleEmJirPGrdHTSRWoYw1D+AGU66vlI84U/zmywMCPPbAbaUlx3Le0Jyw0cLqsv757wHA
hXVGLG7zek0Ny5ZEprtP1X4LHCbViT/MV+ujjrgl2solWPGWYPBdXPj8GykLbSAg/5i9V29BprnC
neO2Nbx0knL3m3TGwlUIL18N/ur96UJ6D8rMHJZOusZaI6frbV004mMqxXqO3Ywxg82QDbM28DuC
kr5bHdl/wRZ6j6TYORFYi/YDDQg/+29AjL4+pxlG4TGm01j3PND7IMaKyjMwM4YYckqEkkN5/HoJ
/zJoh05nMvCztgnI7Vi/lm7/dYDghSGcseUp0lMQh0Jwtlmi9tEo8FBtpnIpS4oGYa1ZQP3hwloy
ut/XsCNiZMmkv7KHDkmwumnNr45fhiBKQuAqHlC2MwrK7mf8uFbvzPrXMa0kkHrObc5mZnvdEk/A
QBqHCbplFwWnvwmOdsaclIuEDu3aQPMg90du/YZxrjxmGQcpAANYs9kHrc7b/RXkqmA5LqZadAEz
MiDRC6Y942IpkgfGke/P6xsh9DRBQkp/u0hyynH8+mDPnFApv6+15tt474tY1TuJKD8eWN8mbme5
vG+lr/Rh2J/fwJ9VFCy03h+laeQu8MrZu0Qzz+FYYk42fqsn77TyEyVXNxhX6Yn8sNO8mzAkuIel
izxmzypdXaMACtVfzDjHAHDbSg/+GJBKdj7I1rlDe9kJPmFop5ZtY+jDjl6ek/G803+azd7Zm03T
bTcFQcUVXKMoLysC2CLRLvigI4yiiTC2SAEwxNkjjwOKDhFflWHk3vmChApCLsn884Zpn/i+N2ZZ
EMnNsrbydoZ2BNHlDIF54CNcvoD8RjXmdsGzXeifOKlkBGS5XOplasFMPD6XKHvxcavKncDQ7Di0
ew5kIE+YtRZLeFlWi51KZHBWx0qIl/FmeU3ACIcYgauEULB+db16c6TV9FYqCJpYLE/TcrfiDO63
vd82h6lRaABuSO3qEQbcMGR0tkASOi2m9Byu/N7nJ2EsRoFYcroi+RpSYSBx76iN8KyffT4uF6uF
qLaiubGw+U2+d/DZMjv4YjOBX/1j7vmbHepFkJQIKWS9geP9B9HUcQ5Q8+VLfw1xzumayFJ6GMAp
5h8tYFPaefXop2jDklTGwk1hz1eR6qV8TazNLYiwY7F5BngU61DObynvmwkyk/MGVXy1SQSCUW0M
A46W+dP6YE4h71g9SAHwHMekbPLZ+FEA+iJMA6SAEdxIhBTAqkp/zKPhfVtYYR37C7qxD9BHKDYN
sp/MpPaeJQoEISP/hahV3UhOhF+aNmLDHkXVnqIHLcL3ia1NoyCu6W3bwPlUPF4sDkXtQ3TDUhXF
8/J+sLD/QGEK8+Ti3EZ+yY2b1p2x2J54o18LG2wWuf4f2UNQMT9s1N3aSfKOy5Y2ctuBIxUlrWez
0u/tfDf1GpGuCtmANf3I0WiUgHUfmt3ClUdxCOHU6SuNhvpjEnbqlJVxJXky0zkONeZDmEy/QV8h
aTCqDY8ruamIKZMJWlAG9pU0sqA7nm3FjbtZm0eCmAybkBtgsNl+7mQP9UElBqnev/DlBdd63hR+
GdXv9NUFgsxcFPVnA8mJA1HKqxP2VfsZZwgHvMaPLsT9AY9fJ+XQQlqWZFGZtahC1opuCD1bey3H
w4GGmdENfrHw13Gos5HgOkNttZ971HNVZi9zgzBiQtJBFCtHYH2mRW0K7gnCt5cOonnzhttjirL0
+uEzB7v1hl09bZYXVyQkPyt0kz740WhbsomZBuUZe52SsFQxUyitG4vnfxSjJOVrgIUIJ5v7asSJ
kff/kfQH42dHkZ+Q1aE2mBeOfy1J8tbrHtXeRCJzu+ynPuMC2g3xYDlMDZ6yE/LJAmHa1GJkXUHw
BVWdnOdQjoFpujlJykUIV3oWaIwr9qd7aftss99PYiDgGST7Zl8t15s9PSPTHk3T3FxkmVk4QW2j
S+rSTbb6bH2piv17bAChlXe63K4Xtvdj+B85wbLHZNZ/5RD9PBm2nZapKFDBsqcx1glIQkk4DjQI
2aqCLbvDtiaqzdwTLP63IeYhQzFvSgwsIVM7M6IDbP/bumotRmvovCy4uH032kg2Xawwt454kJz0
rLPDURMwlzVMmVmVUihhCGzZDmUqgsDQL8xg9Br/DgYIoJbFC+7gf3rzR0zWbPzr6VTd0uGhtCdw
jTVqMIaG1p5USZk4xuz8acw6VGCcIyCSX2N6vvuAr8NEAE55CTy5oh/6yxCRsd1Y+i+j1bxe0pwE
K2LbCXcsqSbrP1NSkbmpl7yfyRzXCPz5RAu9KBIQfeN6Yo8nRitITMPiHGk6a2y9cyaykO9X6YIo
JfEU9bvPAIsl7NUhk/fHG/OWj6ioWOKOKBqyruLNs0qHw/2801p3fL0Brd0JcHqH8b8L7RMf9miq
9IB9lo/hYVy1+2tg9ucXDcsK7t4RvYMYLwsvQ9NDYgRM88XanBivZbJyTe0h7/mE2FeaUkDqu4JV
x3Wm7javvXf6dbgb0+n+d2YSVWQpOIJcxLZwywELSvkiEIjx1AWpTifEzJr8MnmhHfg+pQq8OemX
qUrKI8mqSXsu8QTlpu9J7n6cPv5fwxkHEC0trs7NIBiJY6an+A0NhFzyQXyFFnPHtvRcZ9x2Efea
NFdaIhFxvrAUQaWE9gyU9aLrGK6PM4xiDypo1WAwF26MtzGboJ9yYwX2/GSmnU1R70Eh9PLfff4i
y1sTBdqbOYB+yJ0JxXSww71J8cvtZlCcjTogMqesxYc57M+stBrx431sv7B8p9EjyTYGwLxXVgZg
IdFAwuxFI7NjjD9vS3EPpypGaFlpeCSUXdQzSCbZwip1VTs6j8qOordXRiYeDhMN9QA0TCcXCxde
Ba3mibhj+Z9TAMqB97lCDqujFXL/ibQu90pD6MHlnlivZwHaYRCVGL1/RODkhx04OU+jXJ9HrOGo
8H7rdAKqKspZ+7nJniiy6V5DJW3xLolTolmjHMkrATgRfTF3fWXoL9NbBh9Q68SCMw3C9u//QuPG
Xzh0CvJZlxiSgua6Tw+BOFpSZoENNw4e7hQN88PNpEEBpmY4ELalt92AHga0qAzmU2AlL4ieZNvH
gOEpWAuBuQi8nFXaWCrW+5B6mSoNgObJEocsln5k4TGI2urMbQ39wd6AgfDApdkZpEoCsr0arThk
ZXs9nVffXiwlZAHMeXqCH4ImQ1Wf+e2Z53E+NBja+AwjbaNFQ/TyTRResbzYDgH2EczaeFt/NnA0
7VwGq6WHtzi+R6xFxWhD4RMpfgm0/nMQgTvpyrPxKqRwh91ZHqzu0yeKWlcByji7MAkUfZj/JNox
nIzgnqQc6viTF7V32C6Vgq7zN5CN3bXMz63TXCHLKsU1IKePid2O8y0Ch//6zJSjTWwt1MHFsJzw
8vP1/p9pZRx8Cl50KyQxTHAwL/udOdw/sWQr880J07ctlR0DUphWJYIYVjtV2FrACnE1nB6ZQddA
hDDwrTSxYZPwFY5zoAxCEiZ6U2APqRVBKlr2hUfoI8M5zqQ34q25j9tHiMVRXuc4sIHq0dOEXuvd
IqUXqjCCuUHRJF8ndXeMs5mhhhYK+NrozxYN5cUfrv5UzEaARc9x3eX9ATGsh7tj4JNaLPvxXv1t
EoltGZiKNPpFQTbm7JfB2uNmsFNrcYa+CpkGbhybwkcalxUMgvkRn98MSvtP4IjmP5zW5zNkgg+K
74EzQvpdlOeLrwR1LAfxCO+P2WzJOO/3PXHd2HpnFNHChKn/S6YuI+neJIj+mChxXtqATKjpeDqE
bjv1tx99h0zq3C6EiWo8t8XpMW6u5qjf1o8z1vFSGhcx3sT1RtxAjHjziBV6yfbJMV6JCu9lg5eW
LDkdiJisIkZShCyG5wTWlRxq9Ay+hAajPKvC8ebN5ugEWkMOIhTDkyg1N39LQrz2yVEWpYFeD7pg
UsXSue9nWNLkMe0lcubFAuf5sk4P0L46rZc+DofO26ucH/hjmgaa8CIZNgmkRyrES6a3U+sI+rwF
0PtC+HjKh5DzHoKRJKPyFqxRyKklCgKDQmCc28AMkCmrzf8DvSmz9Iy1zhQ1/m+8gPUntqG19WIl
ctw3Rqv9ylpvDEwyJB+rechdcTWLlif835F560KIIo1K3xbyyfv0FouWB9TQ2utjdjT4jjqKr6wF
UcGGG9S2wvpKSZNi1wvRc47cDAAvKhDrAlabHTTrexwJht+aa6RZECHfMgqa0EKZjkK26LE0wA0+
retOJsKJV/pRpKFS4A/HGfXxy77CeNpodAsumZpXrnuItnebeiUMZlYvEIKJVl+4kZI1hJyF2REu
zCvwYqUtUE3E1icmNJw6R6WeZ9V8pEiWyAjB002LGHxs2omiIXbb/JFxf+xjv/FNlYGnMDmoDuD1
7L+ql6pPYQ7zbzHUwVWkKb4KBS5UkEITDgPL8Phwxv+76Y0W9m6TbEM2KdFBK7ZCmzAlpsQ4glGZ
00gZJURBTBPsCHSVyG3vqJI7s4Xi/J5w/qlOtT+krW6qMFmerDdz7l9Agmek4DYEzVDUoJTUOab1
PKbdGXnuOLegUTXftd/0OkVz8IoVhQKxTJ8hKlUb96xSiHNwRbZZj1RjfpviYaQ4ENdK2fYQHv3M
SlvGuPe5bWFBreTVIXNf+JxtoYRv5sLUXJre/NnnV6ZLngip6XrJezvBEq0woUWvs2VqJBThpjpc
UTaY4iEtm2Mx8QBZfFtPbs9KxE+4sRMNDI1PqQhrECQK2lAwe6hN79F2Y1UaaDs74uE0b0p1iUbc
jAbsAL0/RkQaX8xUNFsM9AVh1M1YcbzlvAiHiUINQhA/DrTZ5EKm8MD69rRi5m8z3UccmOxgrgGA
wf6OCZJHMWPCMg2PZqT4KOEM5rDyV1obs3FgymxIBNXcj7QIv96bQLH4/kFv8ZQ/o65wS/UvPCsB
/fLsJnMDMfFco32pMlq1SD4VC3zMVmdzcKLUlW/LSewJBSdDYsEOYCIYZCh6hPBxqO36qdvyQnsY
aErRi/nBZsavs4w7cS3GEDBmoTqjbRH9pjx7uxfsAtiVQkOR33Jl39/wbwTiZNk5eQxoC6uvfqxH
5q3wtCriVq6CAUvh9zr/AxWsjrEJpAI3qoSQi3l759pHUSmtGV8s+3i8aPemfBL9QQsdEtEwCDag
yLzKKviVXzcUrDK5KpxUo6HEb6PuZfNq4V3D0fJTf1Bp9vU0ZJC7Z3R3ftaBsuHyY7ZtUXnCF9E0
OXmc1Cxd1rVJdkIkDpBQ7sV6LykjMs//b1mk7m0YVOY8+3yVs6F5cZ/IhgZ1/G/RpaXjGtRFtZ06
L8Fyqsh2JuPrk8joAjbmFNQzUQ+ZjPmMvrL0ST2gnEvqD8XrkhQv6PIGTHbuJf6EQjckVBF2qazb
QH+o6VpuUqk/UiEmHV5zCJZQMDQwXUJeg2mjoJ8b4Y59kzzypMbDnTZElKtVwRb360UrbQ3A5JmH
1DKUPpybn8FHlQh8Ds8DC3j4EVtnmaMfz+iYuizoIHtghTEQUwydJ7X/GmKHqhXhC+NpxHkgQNTj
8VRvglJM1q8PaqwRFU1ucCkEQTCqw2azVihAfyuLXAk7TrM6UNU9EuqlkhBol64ZjPuAu/M7np39
3LgK07WAJlb7PVnU0yC5iQXFigoEtxx5fqMXhUPZS67KGqOCuVKrpspFn6rWQRsHf/otVUSs2KPY
iIRNG4PxdFoYidHYGlBeDNadOMpDWyGzR3GAlAO/8uN5FKtBd7CmgZCxcFMPhQpY341qvN3qCOHA
HCL6aIl3nAmK1FX+53nro4O6DvzqQB8ElOMGUTS0xGWXCYAlJ0/p2CdAHvMkaEL7s/YXP/GdTdmy
OMmJf3X2SY+Ms7EkTbykqXcxuqeXNcIPSIofVYuXxNmxN2fBBEFbMaVB/QU+MDZIiIIBnCeUbORB
wTBpy2jF4H/MuCA2ks8gTZa9O6p1oc1aRQbTdohh91ZXEYq879f1CmgjRDfTguYiXY87dawQyMFe
P4N1WDP+0yAnLqjJy0dAkAmY7HI6kaIoNowtImPrNrnwZHEwQp3d7yFK+jKeJtLeP+erG/8zyZhS
i/Q5mNIgh4xoLKNk3qWFltJCIEb+0KOjs/CiQbBIs/yISX9ERn8z+7iyFL0L31MQS8Dmu6I0RUQy
Ia79sVZMsUSkbpegmS4m+1tL3CQo0+9kKjERfV+VIyAxQRfrtrsiYDCFxuoa9Gj+FTFIYGJlcXem
ni61PVKDUL8n4of7J1XHlBLiLiwj9H7cIWiar2g4gZJnu0xkXPk1J2sAA7B9g70TzsEDoeiyNBwE
Gf+YTk/xPPTRevOlBoBDcNveTJvKgQR+n7TIxDzKaRveuGoZr9EkgygdfRa0P+jKLKIhWHY9xtFc
BQ0LEBpBXSOZr4yyydb5xiPFAeaePMbZPl+/M6P6/Nm4g5Z3sYTKLJlXFvsYCskrRbrw6xyQpDKe
V9bQmFtyFzKvKWVrUHy+kpNRbkl0BQEQiX9R99c575vsn5nNWqRc4/hMWyArpXW4UYiltZ2fWzIG
swpaTnUqx3Aw2jCm0YlGzkJNsX4O0ggxH2Yb3QJdeVUtJmlqoIDJYCwjefP/Icct2Z8H0j9rJYsr
es0TvoSpy8wQrRvNDbDZwbtXa2XKBU7at4a1tQEGHvYUnW9DyDrFTWFGnHCbQ64kCf8XQk/DFB0D
tECn8JzktJDsMvpv+LWz0xayN1GdLBzlHDgaKtJMzceTfWeTGrJfLgqDeLHwSXkPsJteRJlYn3Jm
bofIa6cKYtxgKkmVrPcGT3MDo1lBfVsgv3pVX+WzTY8wp5dsrnNHr4K3HdGBg/0Cl4M4cJYCgdyd
xLoFTeCGerxoEQWad5UmGkQClMEeMzgIG9MajCXirLT9b0MIZJvdectubXEIHa160TU9c57OD5yu
17z0/fLFOjNWx7sjxl0jtQssqenShs6GqmPkH1nSOcyoSrUs+rQk/GdcXwh1vZDoJ0P32XvSw1Xq
9xoKjDyDAbsy2MSKOaHX1ob9nQc82kHRozSGNF1lRTKXz4OBarsAJMoufyVacmWnXktm9ITGCsnk
C1RNyvL+U9WJk5kwMxsZYIa0lBMz8Sdf1F3yRMFcpHFJ/M0BIDjryRbC4D+kTsNbCN3Dk8HyYpQ1
KYZ5U53SpZ7At4GvK8CLwVa/FDfCLFdqSo/kKvJgI2vD9vMnoqoobyckdTcxj8EerSR8XA6mOr3F
KyOzCGGJce/NCx3emELQVK8JV82UQpQOHk+PXcc2vcq74asJMr7wWcZLEmspD3TkjDBp8RWiaCQk
bcM9Nq74/uWq5DrumFJ37dCqTVYbkIk6nSINM52+DPQQ0o/kXRI5G8b6sS+n9ClHAQoMuNgXqJw1
jo1fxLzjCCmcwvSdx8ZpqBAPf6shkiYRcxh/K0+H6LOrGWXWqfZU6bN7Emb1ouIP0ezLNsGrSuMm
AR5tgJLCgLq/c777WOa5GUjWTkv9TTvIQngIvgC2Uf2TkPXNWz4ukEdMNXLCommmve5LqGRsvTwK
pGAWVuQYJ1s9toWXTRVFhOLSpeHlrrvGZ7M1sYe1z/O1ZPC0YIJljB6TRETHYbq5z+jqPRyNx4OG
KNttQLoXAdly8+Yea4hGbQfweBKKkWJLamhKgweQj9XlwRoJslO/nhOX0w00Ajo/y0zKgIKjxzn+
6NlEVwanntDOZopmWaqhesfI5XtfcSuhSIUazVnh6QCtRV8DL2vE7KheGxY9bYgdqWoAlXMznRC+
nMjP+2UQWhSpLd+/bF+tBmFAX3VMs9mLR8a4Fplw/KoTWrpQPmyhlUvj/QVw6B6MMEUhA/dZcisA
B11rEUOTLTsNayDJYxNsoYN4dLm2B/jE2BAT93FNEoDqmksGkrlJB0C3/6v29P/yP9oUydZSHsHe
41t591ut7PrHwiLMSwxEb4Xpdhb1eeJxEyijkrdxBobBI4K0HO+Wjl79oPn/Q3i9LIsDj6GA5dr4
0I9lUHo4wZv+55z8NKxzMTGmQGoU0WCJnuoTcBQiyeS/Ecmg2IHlv8hWgbrpGigW+KF1PihKW8vp
PgeeEGKyjjNcYZod62yKmOJHZYX+fYO5KHxn+x9PUfys7+fJ6yEHOwIll0To9woyr0dMBLlh5vPi
vzvZfl0tHylDxOHO6PJsTDxSfb9fxt2T2Z6Qj6gVFGYd4h5R2mb33lrJ6DLyEphz0PPWQhY+KZBy
bZKSDPfPNYYQliTgH5SxGrlsxPPmSpXv034T54qXv8auJhsCjklIL2gmIYlljq9m0FsDj7qp8DX7
uZrAMut6AM5R8iLEq+45y/v8LOSqO/663RbIYLdADHuyroVqmtxfNJOPsa6/yGvZuEn9AOs0nhUM
LKmcCcon99cyoA4ai81427JP09EW0yIecnB2B61pOxEJ58Ek6LJkXl5RBdWZTluzktJHYdEskHp3
9016XDxFMkToF0uuNoFfEiw5205IA7gRYPmXMVomR9mdZJwWYztiUbRGFAkVwdGCh8yxQiSMKXbA
0s4rwFPftDQ/ouJr7aJXosg+6FBaej+U9eQqLrQA+9H2G8MLv8qwsQAIqlrz2C5s2k6CcIQxIqeV
aM+KdFqHPdp0KScZIpdgOCUjsH0s16EkqOZAk/LAqj7Nm/ySy6S+lJG/JYdzGcxY8sK7bYgMZrKS
eD99XSmkJUsi4GIuLRemera3dRKHo3spIW3Mv5IN09c/tQaYQCnDqZB+Cgsc5AskwK0twVyjfDtM
qO7uzkAPdNxHq+8N488rOOPY1iYPLNYcZptW6aJAZJ1dKS+5p5WnvrNfD2QmKum31ZLTh5ZPnbCr
4PGLZY4ekLKG+kPCPmFye/+WHeBPg4RTgGMOo/fCIVd/Rcd/9m4dWlN/+rIwkkO8vtfj/vAWz2bO
sRie2i/orVmoApDif9plhgjU6nNvl+ma52mt7OnJQwtYA15z9JgJ0UFUHCvNdUiBjHWyEmjhZLcq
UksI2nAspGRyGOdjNWBcRmiMgPjsdxLXQSzToJu7ERiCOC12MpEWvFmti18SiVwuchWH7NXhBT9V
ADG+ZUL9vLeBDQLj5KWUYEAMEAzCLw7VGCVgt9CeuM+xTDbOJadotXJO6KFeU8m8j1XFeglMdvXI
wA/OPSdUNk2WlTdiTFyC7w8+acf/ThnCSSmjt92LODd8MzgVGifpQQJ7ZBv+/Le6/23IsWKl99R5
PbQPkb9jim3IZ7XTQa7DOs4vHfzSeZbdZOdtGX6MudOnnJqOjsgI/9EeQdO5twjemrXYWe2YmVsh
v8tb4rT6KmO+NoitTMlSqTLT77TJzWN9pDpVY/xV2DIzp9jrmqqQC2cYzByztqSJ18dkG7UJRes0
mS/SKeYeCkKBfiBzfClx9Rw4P1rwPPcb3dOml57DMTKmZFaE/RNU3DQoAnL9At/lAjsCupmqzmTn
yk2TP4Oo3ncOBELbbXFpPfEkT2UpBOuZfono52m8HoCV1+dtAk4hPV5WrtfWhnoDW3drQJT3zcKz
HK1ztrJ8RCEY7W8q8OPYkKj6C5bdtOow1BcuxfK5zcNDl7B64jAvGuqYct/SynAsP5mBb4Jn/IVw
YVFQ5YiOnYBqvFkwEyUyCDd4xrCZaQ6wsSlR3frMsvZpGqkfXsCTJJ9D+EOATcmacydRbuzP/Bu/
cSBo3J+26rZQpv3p4Rdkmi5ECuM6gEsrfSuBhRgWgVw7yuyxykiH5h4hAdm7Z5LLyxyByTnQmeeX
1xFhUPOyY4zXgNEhiNvfcalY41xobi3Cdwj/FNMBVTbT5uZm+WjrkHb2gkBTzKl8PMs2w9RAZnG6
WuKqmQVsNVtUSNvut1hXq7xZV/AbLU7RbpXEltmi09P/Oe59Eo5YJIUIFemxbGxMaegrxcSZIrxl
cflZTZy036m7vlF0uIf4XQ25d4CxpXC1fUweUv4hh3iRrzV2FbyYk3e5TxOLQVRjPhAU2LNAGsR+
3uWiv7YIuHD/eHKmvkXsD/AX/VmSLQeGqG6z7x5yYcrHIt9zybc+M5xkZsFBau+OM1IBSIyA0bSb
o4OGw00rsZ7TQKOo/aVNwsEMQPOCqV9Oki09MQr/I6gPgmDJ2R7+OblBoBqPU4bu5XniidMOAlA8
09il0wiOLoddtgTkkOGJaKp/E0pXlmigJb14ugCSGvN02pjnYneobpFXfb3ftnZ9J9sh0Mn5DL7/
ZOEABpaDe4ROXVmUpxj95W8L6z5VPtDwEg1S0356zDWeN3cjDC9h22qInpgTGZsGCtoNrbURnmPs
OaLoFzPULWLqGSfxiM8RH4uFhfEYC6I5V830OnR3S4UCY7B3fbisIdm6PGTnFM9UxINyh2oeXH7r
swMuRhoC2XQDgv/uX73C8fF1qEWYlA+e5++t7aT+UbvwSFQQNM8yyJWJ30DdZ+Nefc44VfyaoTQx
oXn9MiHFX42G8qfM3+zAwp63TI+wqlbmUhm8w97K+psc5veKsG0qf0JLJoHMPJTMc/BdJ+EIKOko
Wcb0lXSEyJw0QHJQAnZUwnXiHM9teU9YDHAyQLIXl/lZGfMAYR2Yj1Ug4l7P1QO1Dt38/YSlbhng
Ws7gvNWky1WtHdSohHQcWSJqaM2gDQdADRAboanpwTGzM485IedkwRp3sxm4UUSRqSURKGbzNLm9
RbmK+72EyG8EUQvdxGNAHWA2CYgolXKTG4Ym+1BvuQLiAHup2Me4HncknOS95pTlG8rdlAKdqi3W
PyV5FEA8HxM6jZ8HMsBRU1serBCEz/Ql5PDbk210cNt+ZbZDcOvcrrEwlU4wOjM3HQyyC70UAkjy
1bx0REAdat/HLpjttylyXiZVuy3hpicH68J3CHuW1OahbYNKd6ArpUfeaj9Z7PxXGtz6MVPinjxa
ILqZ2PH/DDP8dHaU+O8+Yz1fs3D9bwTw6EbGSFYMdd/kn190683BFA9iS7oEwVdykOOdcUZtbZ+e
1qGKFq4AKwIsR/h+5ZU390YRPCmjbzy91341AAY/aOjrj4e7gmL0jO8KMJnn2UYDCJ1CSeBsj++I
YHYa1fO+YnAYfkXh2sjvocsH27FjuhxNAPyYWg/DxqsG3FtGC+zMmfXrQ/GfjgL0zr5Bo+wRS+xj
LT78bLxfWZW5JkE1cxqwWvRznpgPc3BIMZlMIzGAHDlOfgPwRj7cakQomx9HyQ1yC5xEruL+1vwf
KPrxiXKm3rmhWm1C41Ll7CiDM/U3Pxfnj1qOEAEZB6jXvD7xqTUqYv4vTsX84oU8oIECfcD7I/Tq
VXuOC+r+RB/5EoTIPWPGaNLY+TzM2T4dWcTJEdXGE+McjmKQT67o+rZgW848RLaCqTRWSVpunHhv
hg3hs9lWaMj4EwPtQUmyWQ3AE96eUQ2FYCkeU9wBsPNJdGgcBXizXgdn0CA7IfJPew51DyrswuKL
L7MnH8IiuDpterSZIYu6S0Pp+nQXQqv+mhuOXpsttEHw9qrM3+ZZCDbRhbZ72tsKuNDyEHoQ6DoP
qMBg33Xdf2Rr7U5bIRK96yspl0YCkPhXVi2jkbFmuwZcATPro80U2IdZygaTiesAv/BcWLZhYBEV
M0dmgFMygb3v+Vjbt3/1nFRm1l6Luh7o1zbdQhRBKfKGq/AWtLEO7ngUa3CcTQZVcYH2B0pGCCdP
nVhKkhaY/JI78n1K6ADgrIkn7xx6IILfAUTenp2a2H8IBTgRIa6zr0+SlctgvsbtHOfR0Z/Wwuiy
cKdiVSldXibeGgCgbGk20XP5Dp0x7A+wznTu6gLYxIftuJeQXVMymeTbJyGkjCZ7Wxta2VkPtFIS
AUjUZxcgXaHMvC1id9oOe8TCJP8mSIzA14BfsTp+JSwBtJdCfWdy1RfHcB8dz0K9jmGOEx062woU
w+kKQcatekRfKCZt17Xd1ezuuFDegoETYf8XxAkAloy5SRwinAbeYNaxxvavmIujFs7/NKhOa0FE
X9StAUFg+Uykz10h24QPl4LagTA5msaFjTKa87Ee7e9UVRQD1g28BH2kLos4NxA5f3onC57l5JIB
rpTX26y3egVJ9dVb4b41cgDqMso9cK+59OglGZVbOIUdHxbZCOVmKs58tvOuUsIvua72v+jlphK9
3DARKxp+BMBDcQKgVVhtXgO22CgxKX96V+3+WMTC8CiSg5NS93UKSl7XVtL+MlPm+zG9mDmvmmQJ
/wLoD0HUFMaQtGHfe4z/E8JTN5v+MG/wAfu+FCsfl6g/H8M6TtkWWU+W7Uq4uD58qqTGudy0670i
gVmFWujFucOzrlOs3p/ByLQC3vKpy7Z+W85wDOMca9lOG0TpxJ4fm3X7RlGIGdKEPDLkdiT9wsYZ
7OsIj5odWCdX1TNwCoGBOK5ThEils1M1iDdksnfhdTd5mqbKl0FEWWKGF6xzD4n4PpONJ8rvncpA
mskBqIwa8h3B2+/Ry1djs31NnoD8RxuwfDOzov3Hh5JPHZXe2EQf66R+mRgJYtXCszELA8TsnKG4
xxuvTOtOnElGRwc6LnXLiLD7ucZhMk3uVjj9W7xZSyrMnokgnQPmuUb9g4B5p69yjnia+prH3fDB
qqzvcTA5gCpFK0Gma9AE+xYAYYhHveAlRa9zbapYFmgY3Dg9/6YZj4g3ToM8Eq5Rlb6ROf3aPD0V
jYXgdiaDqpuP3BlwPffpv5mM7S76aRc9yEK7MgHAgNmF4g9jN9g58CHbUlB+rybiR/LnUKZ611fh
X/Uc5rwoT9PCn7kaFhfRZFZxx7WTwOosSozofxHhCxU07j5Bv76OPzEltKqlUVGAOiKOe+XJK3lb
4SaqD2qG/e5kPjnkZgv3KjOIQowrokvYsZM2NA+4sPaHAHik8JpFs+Q7EMbw5UwCcPE51oiR6Eh3
HHDVww9zA6+GPscGELSQcgRBPXzTemb6bq/vHL+cC7mFy8w4ibxbGbx/nBkoDvyf825fSg8VDP9B
1sr1nU1cEPKwZouTJZiMDwsBUZWxEo+jSzKTvQCZNGQtF+ouYxSM55tZEdbPzGngAoZ/oNJcN6ed
wGCz7VVY4fcFMcG9NTMQjRrLqv5f3T37nsbRrgrRPJ1u0aCz80BCTPxHsqgFiRDij7vsmRr7U0rQ
+cG2vtQaUiT1qO226CWRND/8WCGZsCYJSAXDaX+eMw22USnm7iRuTvZ+EHzRJdyUvNHbHLrqpf0Y
s5cay36I5/swAROnAcLkk78TEIXvG9Sv3tk494UmM+L3BdZ/KaNF666ky0JE9s2Nt0Ak5get6T1K
RipfdoEK3A6kDRFomBMZoENG8lGONzxLjvYeBLsTCCh3VMJxp5lTcpTmx1wulGE95G1qGxV8PARk
JOhAbhtBGjlXBVAqB5tm5NZv0lOFbWEUW86gheTxYuH0vwkJy/KbGQQa9ZKbh3UNSIII2t8pFbm/
GyIndQy6Lzjk9+dQSP7vLU1NWK0bYHNv/Zmw3XieES17/K/FgHV6dNkjtANRbxgeuQWsJDAc7THg
QsLp23+P96GxKTGxxIZ47MqCB/juXMfZhrMZktWrRnCO2I3G42OKiv8h2AFqEqBHraqcUHyxrE2d
F4zaLYohYm+DVK0QheMcb6BQ47aBIwmh2gi+1op6JAsU2RwBLkN9s5OReSjAlHHaLDNiKeO7a+oR
Bz21YH5dYm4abE7xvYM4lajgOKyykpb3IQ9mBDsaWWu8NCTz1JVh4ItYRFw3NLlbZ8tYyfT+qpiT
NRRBuXTlfL1cWuo5g6BJ1qnxrXEw+o63hVDr4ryrC01aoSyCWhoGIFM7eXkvudEQDSNqa2i38CEr
hb536E17sBdgIqprOApVcQ93a2Zc/9x8L2uqxxb7KiHZk6kxUOvxIrmPR+bY++Wu+6rbRl4eIuRH
+3YLGyg+F4ki68yQqlh/WeVkwHBtiXBwaQhxASUubn6AUWAeeF4Oj8Tt0dAcn08ut/YmfO3p33Vc
+I6JW1F7k+KRLOtTGRS4oPpi+q/lOivA6zzIknY+jpjeA1AcZQvmJeAV+zE7tFA7uLC1mctGcANU
u7ai5DcNUf+UMld4IlqbkY72N8JnLR1XZyojk4eKVU7Hc8KrEj9HEinzpPpbzw4wvyOpubKkyNTj
DMLTRQPoT3k/U3Dn4B6HbikQXMPyHH2U+DgNvXEYgCc4Sl00MYZ1Ggu5RZesRIAxQ33D6BcZbuaQ
ow38RddwiBs768QgeS+XekTX6CNCudR9VAcSaiyVCqhU3v7MNWNCUzLDw/ryqaprRRdZeO6Pmjtd
f+nev0bJTvxD2TR/huWxR3IYza4QNsWmQetGLTD6xAClb3yGaAP2in5+Att3n7GvWBtdlCuMGFHB
3bS02g09zqHtXUSK+D1CSYEAZi//DEW+EWJywbaPGvTaCacnfXsI/KsTUh3yEnisFjztYRzISPPa
Cl4+HYFM8TL2sdNLkWLiemj+E/5dL6BRg4nySI84T0nhUbU4i/VqjSxxRnkQyZspKWT+SU3B8Ls+
CNRxieNsT3HikTi68sEOFQ45hoRH9hw0gETa3kCurcKfg0i2lFSCLqUY+RyDuGrW1jdGQv3GTLrb
PuNJAFeld3eQOPKIzYmDiYHoitKKli7iA0YnJk9Pd0Q0Avgp9LqNbAXSPEGJP9johXOFXoMTsHlB
DR60EU0s+vs5B3N7bGzX2Fm9j75drBqtbRGSQVhxTA5jsGvshMTvcHkhCtcFz30np2MC82PzFZGU
8GaQkLyeckKWO2tUpBsUc8jL0HGrSQqmf/Mz+oqUYaWJMEEL432BVW4mDPUJZnHoFauIX80Fg690
DBBXiRmkLp4oNnAzyYzNiiJsdlHSMhEv+MvHkiPACYRcdLU6MVVZS8Ze90LfidhVHbvLna9QFBy+
fv1pPNS1TBg4FAiPoANMO6xJNddsZzodiEZyoyaVKKs109OL+6/QjkDSTN3PWw3TOUNbNaKda81R
JR2xE9kSmWwToapX48X8gWWooLaWDGqBzwF2pLc3mHA9xFpAGXem0RD7NAmT0boqOdyVkEkF7Mir
4//Sst9h09N+Z+hmSWNEx9luJzwZ60aWbt1Lgxp1o5Ou4l7Pv7rmdUz2Izy+yqTpSYsaHSKh2ceU
qTsNcNRMxvNQ5Jwb9KMqpNPKPXhjjdbE3ErWWpoG0dNMxvVU5Q6IjZGY+y9Gd66zs+48HtpGUSND
72wXfbafGsDnzECUn2hyl4aa8HDcPBbEmCvHsd/QuKcxR2pCv90GR2iyrQZIXK/MX0VZ5fSFehBe
0hShShfLLlzSv0u2n8R05o6GxeR0HL1Rv+KZDMh+tDrfvZHokFC21K3oxy1qnSgWwd9xFcn/MjzP
ZT8Xy293Dm03vGLXcJT1x6Rrsi0hbMwsFKnYOfrEB5e8TQ2ItvCrSrsBZe2C4GQjwpDpiINvh3V6
nEO8rVWfunlyO5BxBuB0Damw216cBAfgS+/2EJP4OBnji7Mw+4/HWP8ny8tGHRz/O07Ij6vEWvGI
ZP+FRr7zLRf7lPu+7/k1QY2CUzG65s9P/Wmus7TyU4nZS2mNt4i33m6NOw5OAjkERXbCAelgSffP
jkoNfFVCApdvwRBz2qGvbW0BbT0B1sxjIpYF136h/WcaZVVRtXrln4Z2VEg6bt7aUiSs1xiN36Uw
IVTjg8B9q5PaEAFNP/ogAqDCnXujfi+dArsYtfTsvS+6g/+7QY12FAklu/qMoRCE+XiJ1E/YLaV5
RMd78smoldlAl8+oiwSoOmWg4sRAu4lFb9hRTbYYOmswYn3Rwh57znauejIxXeeTcZq4DK+Hx7aj
fBrar9+Q72sqGhwUqBlDGypi1CLNaxUWDehM67oRtHR7z+ia4YzEAl7AjWjFPLCO/nTQnfVgls7D
/vrTcUmePL2Fqdd5bylFeQddn01WGDGYeT1j8jJ8d7/feAJlpju5Q1u94WJow5dqplGYefnYZ+HM
QkX6SAXx2vfsSS70CdAVcW/Acx3lw9ZiT49vED1vVBKRHVNXHKv6jm3O3ZEOkdx4deWrSZ/QyY/R
kQs2Uz89WbUKvHDk7FMY3Bm7OAh9ji+VbI8i38VHjqESM2C8TS/lsSh8qSHIfJ1IQQjtdZi8Z/hs
yJAUSf2PtgWlFaqLwRqK/6gOHUvF/lXmjGVAeKf2XJ2LuhU1TVKSD6Do19pvkfYipve208o5g0fN
xPll1KRDeb2AdSK/QVi+JXKNsQGrevrqN1jBto8t1c7DKq8GVswn8vm8eChaSnaEcRMGLQPDcWau
k3rUgeGRyPViXpatCtgEVDDlVJ9yJsCW0aulJFJLV9bL6eRh3rSIejSRkC+deG3wVJGWPaBn7olC
JQ4AdjZqfh1eWom3IcUF5leaGt1HABtgyyQCmmDhFVDFcnVEBPpFL87lgJJXjLbKRSz3zJpR5KIO
LC+v2Uj4r0h5kB/4Vy2mctv+CStQ9ylUNW0YePWTuk11v8EiPACY4zowFWT2M5WvP4B0Ovx8keLg
WBrS6CSM1c7XbjMYDaTrXsBRXcnCiGkSeZdZ7ld57mjsUx55TMzxNP1D1VPspd0BiG1F+lxanynI
W2C29daVuIlN88AkE4Q3MmJl/MQ3a64jP7/cz1dBe04sQJriCjD/NtCPn2J2mFoazYlvsUdoyg1m
qMTrq0I9igyEvSmzhfvFQpJQSYmrYrecMmbj6OGrJhoZ5zsC1JeVsJcu9SIlFN+k9vhkdxsZy2XW
4vT6EMBO3UzTKsxRqXfTHyAuslnNYKhkstcyn9qwQEq5LHE1D4AdcrwMQayzet4ahRVt5ZUKzsA4
EqjxCv59T0BUHR1VajIeklGz9gL7ShFdHEQH89PgaXUYxfB9Y2sYTcGJmA1RChXC77WUj5yEVeI4
my8c9XoeHyClDYfsl5Lw0h8DAuEzosG1NreHV9EkUSsatg3PuOLtn5FHYKhFBsNW5QqiBwDc8DLp
558wokLnHrNObkVTJxn/swSZAZPAJXRmacLackpAUlAkY9ZyiVldToT2rx/NZvO2Auw1kSPUtdRO
0MplzmckMntABSYxa3j0dig90PCIkfx1dC9eyTwZVAbrlQgZIFWLCcZGTcRlRXnKKe+PWyTqgTVT
lQjWsglgxyG/TxYKLKjhASdl3VHN5wQ1LNC+jKj+zeuXXRox6q92LARBXK68Q5dgaOrQ6q4nbbgY
NRfHWHqO97dVrZ8m/9yRrLmFB9dTOX1xOpdqIITVSBzYNT+pJUyNOJYgbsH0rYGbU8qLvuXwGxX/
XUYoFxL8aTiaQjqQ2MVgX3bGZ/ooWe8JjaARu0GzAIjV0nMGtdMTzDB1pBKSvNeJBI+doeMDnPZZ
mM1W9lIkxWkeDT9XwbyYZazfTET10uiL7GgrH63+EexK0rd5Nqvwr0O49DkkxHlJM30iFMiqk6WF
LBnihSFy8wAtzVh6eAjkia6/VBvzydbOe+XU1hToozdxoQF+gV/Lk3Y7zSRwr2lKlukhUiYtDmE1
Sdf7UUBuV7quZFRAnqF3fw65Aw149mB6wzS+5JS1J8HSARBjpu107IlSj/ee0Agnx1tc0cUvUjBS
98NhOuPiaISXjXDFGhgvW4sPAT9y77uSLbQ9EqyOBEn0vaa1fazWNSQC/gxMhC771y7pL9TOwuK/
HxcrqzZfWEGRuFi8mk6OL5DoPTkly54hkhFrwyKqSdFG2ff7xfY35boufGB8JJfrbjnouWvCdFNJ
J2yo5t3VjuI2OLj2i9W1yIRAuH7RcGwhhk57xTnDwGt7SPGac5Wfne1du8cTmXM0KIBHzu4smXpq
OAr0HpoBBdGjQV8pA2bsvdmaG7MTbXWGlNyee3sZQtdAu2eCRqISZdvs0bHNeqt1a8OhlCDhuJzi
WH//oDgTb60GJxax1vmEtQJxqlWHnN6rq8/THkFySUrmWVU4phd8ilvx0hgjbaYAAjnf5EFfx/YY
huCY8/ffQumlBUZWtQXA0rq2lllvnzNkGwehJjWIx4rSXy1RBL7kCHh/7NdQk2dQFS17ZHW+CVIb
wfghp6r3xzMrQH590mr6gwwlEqr/kxp0076e6/42H96D6IjrgyjFFXz6EwLIWTyU+JOeo7BfXw9D
gTWufuHx+ubcI9+fe+1tEwuNHNhWXXjzKanl+y6G38rgIkt3xOWXFKGgy0I6Y8QdLGgD0Bg+7WR6
C1CasWMW3BBcpD2m/ZvHX2FlT/grRNKTxXSKW/bdZ7h2/tLO3KPaeNz3G4MTa6OqTpbcqwQQkgDi
F98I4xicEmMI2UBTojGo1WYqmA7ZNwGbY1WVT2A5cMzE4ljylxylqQzohTESnqcGMqU0D3MPNYrJ
s1qkuFuynAtRPIWMLEaU+Zw/4uXoaK6zP8VHaBvBX+TJi9WbdyKZOudttP21Q5YLo8jjBnmFWwUs
9w0v9GU3+Uy9UOy3kkwKwwr4Fho4hkJxffCKWizM78/GpF6IW5iW38/lLql71ECdmFmK252boU1J
p4KURBSwb3gT/rtxESoBma/VXG29OMXTzk7HSQR5Jx7Vm5a/7rDODXIJm7K4baGe5C/+E8UWzJR/
ERYnpoTnlL1Ue91a+kOJZjNsqSXQQFZ3MBu5X5BCrunizrKAkK5sH7UI9uDZ0A4T9IQk5ezMAkFI
E4GdLoeWVIrn+lToiKu/QyThcJ6sGOcrGq6eMXuXqAvFUb5owX9u468iXv49SCPTSo3794rfpNS9
ffWu2Qv2nzRkutM9fPq+MfBNRIY4wUjOKqgsaaKpvk2cOGOdc1I3oCd4au6ebnpRutN+yS2fF7sx
foY8W0llbSOK7uIDpf7LWLXhd0DL4+KDWsqt0Pli/bGhvNk2R6uTVuavidJI9Ng340W7X3WFnVmm
seAWpIkYYeRVHrvC+9rUCga2HMDsKklZsEOIkogRM+x8AFEkbY0bC02cPolnM3asMJI9NJzWrpeP
gadrMwIoyar+VWQkDt4znfb4X7KzexuOAw23oEZYsQ1sQ+4UMaPrKvgKg6VrdmYTxUHy1OfvfQDM
iaHhU0UKIH0xbFPfqhJwCG2rUigOlImG/qAr9a088nBf2CcNLk1ZdDmMbOCyIwailCOtf7d5Yr/v
5c1t/iGaY8nMCwx5wScLa1EfPQiFLJ/JdOYH9j6XQV0triI2YagJ6JMgJ0ijSDt0j+tGqfu+C8u4
gddTcViZcD30nhgDMeP9SIGhoFwryod1WLV5dcSsIoUY1KVDNf7fLgMki3jPYGNj3ad7x44lKBJd
bj2g7RK4veEcDkLUsvHT3nADvH1Ock0dKEGETRoSA9CS9gjqJ/HDlHVri2op3aIQ8EADMZTR8hdP
QVJ13bfAIbjnp8c1jQHUUWEAGVA0Q2TRITBid0Bq/KxqISIZeEAbW0BsGqIg6shg1/W59XrtwQzI
FT/jZOBoytFFMRKnOVqtwgoGEVSWvO4b+bbbvKxi4zFxpYGhBNxdsry+z0dTCqap4dYgvYX8cS8f
zSaTmmFe0PNwGrYyS2kukRPGWePc4g+sKbR1K+Re27Sp/UxqZBsWeIE+3haWiNr7uaOVJe2tvayQ
3+ZVcOqsmK5uJNsEOJiMuLtxEoLTMIs87IWyDq0S3sMCHs8E9wvVJRsJiV87otYw6jLcvWfSkY+N
UqWEbwYmPb5pH60UrjW2+J/4jbvmPb43BUVrqclMD2tU0Mj63xc00RXE2eatIh3OVz/qQvOT9xXm
cQn1o93PONczaZfm6BO3zHBqD8aIQ20Y8uCkf+iASuHsTC3CB5+i3sU98KTRQVSb2qmfcJ8b5lVV
HZ2Y+j0PUmTpN6DwO3oE4i7a/ZWJ6IQsDAqZIE0SVCPeEPfj0uE/4009eRVvBmNMkxADOEKzBnQd
socKS6FYIaIiXIriJRPfFdNvggKL7ZDtyxkdKMfUK8turxHoMPEXWSm68CFWsXzYW1mC4V2YNVjg
kBOlHrNSSvCmK3y4SlGTW1bLg1nxLQlNdDiLTc70jwv8E8VnuajhB2ztQcjS9j/jBDhH/ZlsX+gL
KbMVe9aNNxaqjdaGThuDEQChRsiJmfj26qeZIgR+POb/25sT/nnYtl7FqZ+PFCbSwokplxAQoteu
aP6LR1GCv587q/DEkNcdz6w6B81tA2Vi9DUE3K/mW+hLvx1CQlt7p/xTItudiGfd0kZqstGHQBep
YMB3g1b5zpm9TF7hLgALnOz+hNx/uHWt4G4T82RN1Alt0mDIjbVKGqdHmVhtLAalmydLrnmohVzD
/BIMw0G/5frs7fuXZBgyIDG6Q6LfRsKKcuKR58fUbR3r+iATqpguLFk/bSXd29hlkY3FdsNDOxQm
+ZDoBOgHbfTFTxIEXzr+Pg13LxTmiYejgtBlyTMMHs+LWJxJZ+bq9yYpmCRXPsmSBHcUZ/Ua7D7z
nGVYpjB9qZStnAPEJs4qYKXRrm5uXrA+1JQrcEUSwgCfBSAzPR5Qa6MlRyrHm7iqswHGW6kEvKUl
bTvx90wC65Qhge1qNkpaiINg9ss8G+6q5JNsvoHBIrnAGXhxKKYs49nWQ9zYKLYChTbJ4xkBkI1Z
gaesss1+mEw1Cr2S83skn8H5KG0aOD2lGwF4dS3rD5n+dBMkFvYQdyuax5ln1bl1xDfu36GinxJ6
02xzONvq8JZQHvRrmwNgOnK/wWF2uEch9cCj3B8hAYKVUCnOOC3vzIrNRGj/ed5ICV6pR5O8o55g
HK2Lx5pWqKaJC7HjlXBb8s52rmPCyq2zPEXKE9siAW9yJcU2NX5iApgkMzFAX2XXOQ5fVROC7CAX
5tbDwImz+1XdW8sQc/1Av3Gokz4arE7a8VZ+/Jv1wQXwD+qIDkc+nIUJn+pZXbkGMuAxaAnFOgmH
Yg9JerTGpqKOiJ6IlGM3H7L9IBwFsLTWnngqbw29X9lT9e41nlitMiogVuU5kH/d/mF7mr/lsaOP
rkdMgK5JHl6UjfvrG9XoYU6LENbD2eI3mSKyaZvIkzasAwDV0CBdXJzfo48piBfP3nT4VRqp2KPL
nYLoaU2qZXkMTtzlRzH7PTW/r8PNFpTs0stv2UewwZdu/6DEzroctuWoW1filutDMFpzoQoo/2V0
PHs5wHDkH4MzH+u651UvCcOl2rtyPQbAN0p9ukBBQJ6EfmLILtRRud/2xZYG8bzdbV2zy+a8cAgt
H7a6DAUlIUSmMHxSHHaC3OX8pLmCquBmtVsOG9JWBdmxcMcUbm7ATmDlz4Ab25W1xDOZ7yJu6lFG
jVKuJ9x8IrPOKMvjRd7IvyCJo5wZFarLqyCEIGOovY/uRLqmZlUJv7Y30emnYLFt4Ll2dJGGtej4
Gps5hutTv7wOqqPSNViGfmNoqxau1gORadcFujSHWuX63KXtQTaatA4oLFgfCNUuJ3SL+Ev2zqrz
l0qLp0fxgvaIxw2W4XIM87xqvSKlyQEpyxH+ogP1vj6B+dwOliw8z1YXeTY9+pMRoINakTEFnwM7
uNHuKmHYm13ElQrFhKjvuHdIsUpG6n86oAWUcYCNoQM/k1gsGhfnTPss98PXBWeFcpAAXHUk6msp
jNHkfgyYQV5KbT5ZD7vxpeIu7/XFicsGjzwvvw93WOZG8kXW6lGI4XBadzQrUwS6SNJaoSmBmTOg
rl8Ltmznq6pLZQ9fIpfhHfriZzQkmpOTjeEPzWD8djYliEL64JCaregSLsO9QFwfOiLktJlPyBn0
DGNCaIwEtTY24Rzub1WY0trsng13enSndGVbsAYdrgbBRKaZ3hKv5p39Y1igUp7g2hlzpfvkYSLe
gMhCOrpQMDbPsfBNHtQB1QDLmpY1t+s9X8LwBW6uwBHfsXEWJX0h7Fh6B0Xbza9t9Jv0iQ2uISRJ
P2leH/Z3Ko2MzPGRCK1Rr24YXDJHtWrIkaFpb/zlch4geTHW5X0lfLNoRI5cJOefFmKWNaL0pWGa
cpoQhcg9ChK2P1lE3xtdDmikc02o58dYFleo3Ws34pWCqFYk5iR/BExaYDiESpjQSz2uudTq2iZm
w5zo/s1cYq4rf3HrqWscLkHtfNg1wByns0ugsOYJrxd7BGwjQ0cNW75rTPrOiGcXoPvzysdgM47w
KpCiwPhGxkhTBEm89oGQlfbv6qZ5xbpTVYsEXi39dg3ftECBBNgo/VmRhuqaELAQWIPLn3kDpQfl
t/a3snBfGE6DX2avVRz4ltyunIw32fKtNfhFR29JqhqLI2TywBkM9A1j9gmFqHbEpj/9nNcq7jb9
pbjL+bhmE5iUWZAf+tbKNbd5LTbKI6TcbA7tBkp9zfkjFT7i9weK4V0LnAnrRDB8V7VZ+96l9Dj3
UTaP8CqllP+99PlafgiaYCSdWwMM9jL0nySTP3y4Dk5Cx3l8lBHEs8CjXaylHKe/8o+7eRfmx4eq
3TvTAcnsTZ4h0uvBlxr9TCa5OUrFibNgdVEYQiJJcphXcS8xCbi/NNs8hM+fQy7TcrnTdGeeHdzW
IX/5ryVXDrMt2ii+dEL75QdOmM2AJkMtA7/m7Pb8bC6Kuw51+NwStqwkzRTx5rLlEn1rVjwWrx4s
mEi6VIWSpyTm9xYmmdgXCN55FEU0qMqmfjWQY1UUNTi7VA1ku6ghZD+m4RQM/PeEV9AjhBpJZuAl
MxpelI5k0wFJG+Qdet5M59aE+WqsglAaY1yF+nESx7h9xzxZ1GacInUqUMyarFdcXRAPveTHmkMJ
T5dG45a8ILzdVv7TS37LIPnMgqgZa90dr9Bsq5NcVF2TQZBlB1Cjx0RaIfXsdDP5Ou5XpICzW2sE
Y14CAybvcptoTiRZqa5zH1aTcI09WXk1bbgVXVykZcyxKm9Lqji5gBN6DAVDe0ae3ml7GgOj6mKi
zTmggI7DYJRIh5mibdeIV0GUjf+XKWiV/6ixBEwxi6WtDJNRr4G5RsHXL9yqkroGiMrKZwHVKbAL
RMu4KYbf+yqML9M3hf6+V68Rylb7XRBuDg87wzuOf5JCxAjNDsOCQ1Ihy4tJOvCwO1FPFcbX6GVr
+zxlIS9G3NAwFEsjMeeYbaDZZ7wqCcaSgQwUJHgw+Up0KBSrur8WeWnmIzkXOoqqF4FxsIDL1Vl2
a/RJN9+c/M5sWXVqeBr1ELccvESlXdWOK//0Q1e9uBXvDzB4701pQDpaD1yModysNfFLc8lINiJ2
E4WDl8Hia7xo+6Rv/2eyltFxSUUt0AzICzzKjX3U1Bh38HfCycUOXA49LBc7qvjHAgp1U0xHToWq
hsFV/z9QTutWwrwopfT2QjMHzmpUp/tsy7C6AN+QzeT7tPfr/Gj9RCtsL0QVsaJLk4G/NewF8HO5
lgWnye4XdSZovUUIM1rzI4Ax/K31fupITmuAGpQPw7K2riUKxDNoy2Y6SXGGhd//sQnRu0cq777x
SPa3HexRBE0f3gGbtaaVoGJDrlgm9vU95sN32aaLnHd3gaFqAXmlZ4A7eJ0yJg3c32Gi4dChverJ
7I+4MONMMULJ8AAns5dKpUIVljvjfGt8+9VBBJxh2zGShE8QKTHeypKzWv/AgSUu+/wFKN6/y3dC
vBB8RVKqH5KeFc6+dUZxw5NH7ZOMjS8ALf/Nqa3G5WizKJp2UNV0qA/knpa2qnHa7z43TF/UYgzq
dAg+HmyPSyKxxO+ww1uWQbpxmp9ryqw5RTmZ9Gb9oTl5guYUjjanKuyp5sW2GB3ygPUPubVYOOLP
U+TwYlQ6NeiLbyQxnM7JlDc41bFbj1c+4hb7xpjgcisV72RgtXqce5QzpKzJ2T+3MjeKuKI08amf
TTgMLsfEwEe6dwVo4Ith0hjRwmaIUMoGBM5sqqj+4r9ub+9f0oD4b3nUzeIvZjWWI2ocyAiCgunl
rjmwOZzy9MYOquXiiP3lIm67hNlz3tg4Aan7OdhXW2amgpRz/oiGqP0QbkgIY8uHPEnucCq8F3tN
/veUfQSu3VUXWSQs3lBEYZPEAL7veQ0H4fnr7uCO5f7w+X4maKJA/tKDJsYOCVJUnwuS/mMW5Iwc
u+S/lYa/HPWVP3xfncTMF1I6pwUgCr7ysEtYklkD+1wnBskor38dnHP3B+0afqaDxxArgq8W0c4B
/egv3oFxITRgl3rqYphzN8EEAa65peOeKWwOUAxuFbtKxpP6dG02pD/Du/ZP7AadmdWgHVTalg+x
vaQX75dI/2mH/YRf92AABFA0ll5ds5j0HfbUj2Vql0ktVHX3FsJBWxbe3WA1IGPsna373qBdOdja
G7Lod7GHWpNbPXb0z/6HrFPE/jHKOvKqJ1Wg/0JWuBJ0Fk0AIHlYpCwyd1o6EDzHgumAC7pejRS0
XEbHOb1MVgx9arXQ/2GVsk2QOIC23k8iWvlfIW0YoD79+UQPqn3Gd8w3s7u7d+QaOQDeP/QchNBH
P/EuR7FA621TeJyZvN0yKNcRMBpIfr1BXvMnlX9AdTYQNUxS8ysSzZyLjRC/SzUuFcLK8A0ZbwI2
LlYXR9p2WiZuvS4GnzQj1om9GM3kI9xRtUBjroN5DO29LrkSWR2urGxL7buA4fYgeZdr/hLbC5ZS
S0W3ZbEoPYmlF4O8uDnS/dWBrLdg+gd+aoRSy/Ek8Wtp69kT+/JstEHKgrMbi3XAoV/X593aLtnU
7igTpv5eAZCpVY5y19/iNjInszwwWjNjbACoFWREF3MyESsSgLj6MecfRkywRmOKXsYMDMgsaDVb
+OiENenp2OyCDpB1Ar406NuLxYxtzAs/a9shjl7j0Vvy/WrcLdjxO3QlbRggFLRWum48O4hmjTaC
VNuwXEhOCPMCene/JFub/soMLnzMrWMnkbsgaq5NgDNoSFnREjSZLHitBPjTtJAsXZ+19U57cHjs
hLQYNSEhD68PG5W9Th08qIrVsm6muwnakkvWo3VzdvMQK9o18VslSecAj3q0HO4iW5a5rpHs91BK
DGZ1Eb4iXJz4L+GlBQ3V7r+2ftAs3KljBaOJB7p3MQ1C0zNkhVwXX/oRBRDRFIHX1D0E2Pw4xHEg
fYB3ucRTMuy4XeNcuYg/DXn2oLJe8/ie8n5CGRRnlAJvD44T1APKKk5g4lyBrhH15QNptIUb1mUQ
Fs/U0Mp3LTYq69tZxNXDI5Ba0kY88yN+Ogc5+jNCiGScbe8I80mW0hTjAbUWf2a+0LWsXCSONPeo
48RMtHdjoFof9qCMKQBeONhhdqhmUU57RG6fTT6zBme7rwIz5jKGyHfK9yqiU8QjSP7dPoBWxElE
226jeECrrmj9jfZzVxl7rc1x25jls4C6xkLRXhk20eTYymKTjzeKwE8kDT/13S01g+hfTP/ebq6a
nzjUJnqCcWXH08VByyEhVHjiK9c1Sl5VRpFJmVK4OVl+mC2zNn9RzL//mmY1xwFhrnHBuTJbCPVu
UESMg/FAw+VUZeETaNJzkveTnKcOcIK2ifcMR4qfOLYF5vEm//0aR6RIgwZ2j6B4SOWaD6L+t93f
EKTe1yLMeQ4iL5gmMv8CjQZhn3yMTKGX+hiSaIHBFp+7kJ0myyqmmleaSvzwkmRAJDHSnLfFe4rP
kii4LWF1zr+jLHc6IUjuG9AmcQ3DdnIjLLDJD23zGwFk2JWb6ZHz9g6iWxQEmuT3gmFhNQQCoeGX
H4IrxhMOrpU6B3mtZIrUiwYbYnhYJ8upV8DSvX/qIJdW2KfpaVCcsaU0fevQIxVtv3yBJPRaCpuW
f0C9SS1vK3ihCQKkkAiWIu/x/5KWFtxZDUgRMmClpvppvvfGj1oAAqIw4DhirXL3QQkCL9WpzWwV
cb1svGOS/3XsRWEFgZNCFbTG5sSXsTkdbfiVOkr4+lJox23lpPYQV/GebTEhf181LxzPoknzudvp
E5KTsD6KsXQYyuO7xsFDbluG37SKY19WYAWU6al6sxFZZTIJwSWGdr4q2w3vhUGWhshYpB1Ow/GG
HH6/oWoVN97Lnxn53PdMdpwPrctVI8x2R9etzrsqSz616dL6/blAgjdavOIRFiAsVW4d6bKR2pc2
jrWx7ktYMin5YOQmQj86Yf3H3yifl06V4LuC7bdbRS+D1BuS+KFW8CZWzZ6+S1aELyJL+WgPN3kl
fyF2uVZIlWHgYFX80P5XhSMmEawhYtS+gNuxQU/9x6Ph1l+T4hxNR+hN82d0Gxj74MxnbiiBs9ro
yXaJbn948la5Af7JkH4Sa2wB2JL8Q7awp1akCY7ZQHs1qBvs8lCUuRuUh9kSz6V7fMW72BcQRl70
F6EwIQ08o7C/d90E7M6iTVactwWfVOydhrtyc4p1lUwLUuz8zTqJCr1g/qUm5B73eqsjuXTfdDWs
c5TtyuVd4/vZEADeUnv2FhPIHO2JuCmDo4G6IElKbHgAnY6xKHCxtEo4EUyabaQlKnMM6yVOskaP
1YkzUcUkXLHzbMCXpu8ymk+jYoCHfN/qt+yVeMLSqtqD7cfIPGnvaUxr8dGB7hxX4C83UrryeQtF
yXg1o0lxxk3PWaRrOg8zhE9bhpDqZxXugTs7W0OkLsFhm9DB2uK61n+qg3kLh8QxHATkDlAEVSWF
m3CbvDYgZEMZaybjmlIW0coUIdytcL7B5l8GCsyob+4OLBIOe7BT6v7RQKUyX0lEWaupBToNaC/I
Il8LDirXGfUJq5gGAiBhGEXlxy35r2WtHM2DwNeLD6luaQGlOybYus3g3jdqCpBdYdWG6voBJSQ5
z66UGFFUhTSEdUYKyqKVQAi7HOIxBl6HNTnaw+VHruVWKKJeKrIKwAT9qVgG/C25c13sDOW4q7sS
N0j/uCgU3Sxt5vbL5mujo5GfdWQCbUlVTU7mjxYLfJSgkAXvQ7cT8LtQ4rPaUp75HJN8W+rvmP9x
M/de3QdpY24S8P/uKb/HW3x9XI/bqGmMDR8FQE0A18OHIyjUZ2/iJkMs2+w95kDdbOYsJ82SV80c
L1MEsxQLn472sLBTAFy/7vwGM5mPwhOnGdubwx0iWVBVqLE+Th/AEYcZ5FZ/jySO6AUyXCFEe+Wf
kIb9Zw5y+WrvqyStQT6vh63HThfTy74ktWhH2X6+NrldjEnYAoh0S0V9w1y2FvVWoBX1rCUx12M9
WtfiFDaHcvKWLe+/4WG4MfVQaQbAGBkRyrAj4IQ0guh8DZyHKtSD/3I46wcytUGxVMt2/il/WyRy
yJP35Mp8N5YJTTXO+YMvLgui1R/8pRWrHrRhScnoufYu7GNd0Mh8RVx+AviHEmo7gRSNprgtWFMA
wZBGbCUQmAjtj6dx8P5TcFoi5gKHeypf0CFQyZQtKgMevDcnmnMBUIi+haaljqIARXoIAs28wV8V
uWP7aVs6L4QVds/zNqkL/nSRSzrPXhlGdaZ6Q0q/y4nuhJWUN3WKqYKTRgtP5Hd5//zhVVQzAx7r
bMU9703z5T7SeKW1wqL54+h6/9qgr3nj8qaAiJ8nG2sNCGirIeIKcx26gUOYqjX7WHWVvGCAXpCy
TDlKr2S6qkq2X/7YtjeB8V7meO/35WdWGr0hvRchmAl00Ku9E9tSS4cSbh14ZD9OP6adB0eqlwKZ
mtSqAVqBv0i1ki7J+GK6fSfJGsInYJL+A8ivtNjtYAWC15vyAz0gnGHef/D8FCIrCMz+kumaaKQI
uoLLD97186Ktxn3xkDGmjC3ZaBehdox+JCF7p3Kr2f47sGh1XB6Rx56sG28b6lL+mEqjs/5udHBn
jlgpA8tFFItNaIztqceApaOwHGsKoR5JyIzY18SLEHgry21Wy0R1AgduRmfDb/siA8rh2Uen4sPs
J6JusGc4dbrgopDqPPfNpm6FT673+QmcVSu2e20KyY0T7MQUnHK7ve6rj3EpimHZqBlvhnfTE5qI
Vwq+cOB5jOZNOJ3tXllgHMdWV+RUr+M51x0UrQhJOoewbvt6wNoB+IoUvqJN3usOa0koORuX8rzq
hIrad9Yibp72/uCugFMx29TI/vSoZ/qnpMXXny9gQc9aD+pdn6Vomzs0aqiLFt8pR9lRKzUURzdg
2C5dFvs29Po1RslpSN91NjHUmG9MoZ90IgITE9jkNAGBHKsjwPQIUWJo3nMsPBzV74MRGq3ZlSIZ
ld2xJwU4tLONJ4b++OeW040MzBdpWtMpXzQFHa11zYjXTfOrbSo1f8sDRa8jHEv9AMmfHI4rRY/g
gcT0z6GBoDAyLp8732es3ArPs/vzf9QD4xdHE17fjEglexkjH19SSKi1p9XVy8wNJu+OvO1GLHCx
M43EYAZypP9rRfYeFAbL7MfAppr1VGulEzWR5TjfUh247Ib61YB1H2DZev0KI1a4k1BManEDJJNU
lwHRs/f7gtVkL6XFBbHXhgFqRmjtbYDKPdl/Hz9b6gLh52lcNK25IlCgfI14/2QeSelAD9/Ej08/
TGk8N2pceSeEhEJVvulRyCAOpBSfl8QqKgiAsU920TqInMIwAhVckLrGQ6fUhr3tEGldy0YqCTCZ
enxO/+4tKfQV50vS5LpZRa8oOHUUmYu1rbAmJ3TPMDDE2gTpiRBc2B+/KLSpPC+aO9w8ZK8ryCmh
aUc3wK9rr4w2TlrsC/yOAMDt7eIPwyiPmYAGAgH8no46Cq5vYmdjGfNZsl4etP4aXmp7oXVBPATi
PXzsXsuQuD7N+9Cp8Ukc9SFqUGrmQt0MA3TpRnpS1Lqk8tETConOf1uegUy/5SWAG12Ksne+daFr
kXdId0J1gQaADJMTpliecVKFk2ZxdNCG0AGYv9yZC+yonpoKAKtBZOz+rK1t9KuzzYrsqTxsge/R
6foLdM9EXLWAORl8fog1NHfmCLzhzRI7EPqgfexiV4PluctedUshy8GD+NSmh+BKepeWQMNI9sGW
mMn2EFQ9Fwt4UBJs9SGeqYkDyl+JZc1/8Fb6pPb9jI/H+5iCu+7n9gv4zukvfmVLtkppehJV721k
YLGctgf1bUkLa3x366kJfzTPb+UziKF5f0s3LXKveswYHIyBql6MfkwGz9/VN5atVJybi2caeFGf
8XE7NG1JELIlbJ6DaHoIrEvVRwk/ob0TpV92nnq4HJ+mPtTHPvcsPh4317MWjaBkXIAtI9tGoXIZ
PtK4tHPatYT2kmNthnEtAIcjg0Kc0VGfu1LY3mHkQNfEUwg11Jd8wmBTZFZrXikigekbQYR2M5p/
TqM1oKJTEw7TvF+viOydvHlFQTVXhGmuWHa0QT7NMUmbM8O7A0Vxcxk5NTsdVGLiPoUbMvvXniLT
UvIh+03NBefNDG/WzbHQ8xXLpcBuevxJxDIEZjp9fuGNApdlIb+lJ/F4184UgSS0H1QKIY5mj6xx
/PUTGat7q6MXR4NYEE4S5t4aSVRFG9HVUNejDSSX2lcqBVUy4fJe3YPHLXLPjLmU6JryIA4oqSSP
Vl1KDgmmhKSI0FocalhmjkR5OrcPFkWfdBD0i4pNCbEe90bbQfn7AbyEP4rBviwkhJFbFxxsKZc/
wfnBCrCkR5LSPE8Bg5GnErnEkHF2VENUKvgbMj/uHrvkFq5Gc0KR67y79GGUhyoy0yCZddsH3Xtw
s/VCWh7njFb7+SIU+kCJa/gnVZ5iEpUBAuN3AOsLbVbVUueF2NdyOkiOd7pD4QTJJzKpZj/6zy+A
ki4mYreB+ynCPrORQeglPh79qLHRe2XFv5DGrGbvau4NUETlG23iJGw+xlW06fNXooPxCsJCgehw
jPxrPtDBX2/lS3Gt9+KX8FdZsV7Y67gWdavsSmamISBfZEUum2mYlNNK3X2Er9kxL3UDjOacZ5lZ
8ReYXqAjCBzrNZ3dWIBovPga764b0jBtNAkTv+tJyLDoQkXdWslvfHtXTKK4zIOSVih/cY323Zgy
Mf6RKyGlFiiVfF+RBWkWLPpudU2L2G5l2xAN/Iq3AuoywtMw6PIp2myVHmuI9xCZeQ2EgfvIuPLO
6oB6YyBD8DhGFevUzPR3uMwIVXdsp3g1hoJiiFs/julrQLpDIGcV53tXlytli9jyx8viDBdhQ9L1
jpU3LH1AZ3iabQSkoVE6BtAKHVdGJUrgb+wiye1jfZwfbq6UdjrWohNbsI/vuVAN3HKeI4CyYq/b
NUlbwYP89SvivK7ZeIhTN7Qzboa7jCkyI166tbmbiDKmV2jPx7mpDQ6lK8VslCtI+CBmQquCjqMX
nRxSvtoscZK+oStYz8kOhEtE1KobrIdr/zUz6DgIr3zV1C/2uUZBMBevGAW3QIywe93ERvY8T7om
0UDr7nKAkgvAXTokLSp7Z3Ne6R7EmSxe8SYaLnXQhHeN5euf1BnsDpm//zwCP7VbZ2nTlYOfdEF9
OIoNk+xEQnTooWqdUwl/JcFGWPcGY0EeEgdg6QqiMI6n1fo+1r0cROddzIrpx14IyqkOa7n7CLJM
3YyyAQaGfp9MdNHz1b2ARNmfoAlizLpw8S6CxrnPfoyOcvjw/XO8zQB97aQCrGXoRvkgblGkGR4V
5z8Bn8jcLO4fH1EfCEOsG0E7leXJdSgeTi7guE690xyYcPeVNb3YHpIgylgU6MuTSKESqEmVVjfp
h/IZGkDYgJiYplT9QQBVhCuz4p7oPsM0n/X1ymboN3AIr+Biq/9C0sGuz/3mq2IeHHS+HS7A4UVm
eBi2Bs56QxeGMz32gjPfRRxTpJFM81fYv+mdyCtTfIQNrysbtzSWF/KIDWVcQOSahilSoDPD3kMM
a0bvnsx7E9jDK5yU5vqyEBV/GyEWQ/mgZ3403B53YGvFZmtaxzsFPD9fHA8z5kxKJ39jCIUqQYaL
NnlkaZZobKAogLfy8iJGoEuUduE5qcHGxyazhJ43DOFIBRA1OY7p28nCa2IIA2Qi07+mfaqL4mX8
ke6GIwksaQiDGmo4CKpR6uG6qv+AiUfZPhcmTb6NuiwpnNXmrhbWCs0yS9oNPbYAqm9iSp7BlMMk
qUpH6arxWArcMoIHsLUTn4jW6LL2N4ayW2KeVy0/4NMGldGtbKxzFQ2V/FRPtI9p4wj7pF7+vCSC
n/d/AknmD+QB7JW/Cwe63ZsXIUMDmSOidRpSLIXZ6gtb7GP7mzUwAwzR8ryB1ZqUJUqRavSmPXiX
M3U5qTQ4/665SsLPR5QGohNYOBNuBqj7ufHh92wDHRM46YsmXCR5ZcR/5KymYW5sc93JGGFK5R4u
QRlO12pPeMqC4M2LDOdWEgWqZjnUd1mapoNxN+1S36Jlg4rTiqMo01NfhFUcSKAhMaB9QM+XBa+e
CPLNVFaN5imRpb3UI2OEglb+LI0Q50fLf1zqM/+2dd0Bz9+mtVkdE/jlOCqhq03q9/xDZh3Q/+9Q
25oepeyb9bv3N04UHvubuxMBTZ99k8lef1y6uitVGVHyaBEjVb6xcyRNaA6p1nMJEVw9fz1u4sGw
KKauHOAw+zKWao9HgiqA/skoyYw9BEPgcnvIzYONT/rrEg5R4SARFE7JJGH6D7hVIeLJH/fJvHqc
LMT6v5g6nYgaAfap3p4PKiFQfJoCFhTW78qy3uLu0ok3fGka6M6/E3aFEtd0ul+KHO0tPAxZ8S80
Q1QGfOeV2HBmEE3fpoMQosaJSSciivcQ0rRMIOVOTTD1Shvu1nogF/OdsrVQvBAPKdkOkzzGK19U
iGjFOiZK8CL5TQDNy8bFRCJNSlLsLWa1I+0L/W5/SQYKadC0+PwB35l4LUipPFa90kK15MI8E94T
GesVeTL6pM0D+zv2t9aaVP5ILBd4jKzG4tHbuJ+1WDDYYodSCkmI8dymCvpJLN8PWx+t/LAKIOC8
njWdpACXxFObOq1UdkWkVJsHQ0r17w5XdrQTGl6vITf8rFJH4xR1Z/D4Zk6e2If1iascmfIJBQKC
7tpYytKPXPiZE03axo7VUFRuCXjYAnrUbZSID3uQU83RXd5O80t6rNPdufVjziM/9PZYnPyJ5QK+
EbvP8AEZ5uoIw2wB2r/2FjWY6gjMfgMyp38/McZAAgvKBo3HEhlZjxH2tlCxjLaDaBJTQ/L+WjlI
pPczTukeQ7dJGqy+FvSJoXQ6Y72+6rOvZB6jPV48E9KSB/LgX0gl0hmcsJezhLDTGYa71OHIfK/m
EAmPLhrOhlrGWBTcGABqgLMbH6mhaIqYaXU4aMX6CDUraXxfPl3sz3tL9cCK/zBlp+IchdHT4LyK
cvBBu4Ulbv+aIDDcFpTxJsdNsbwgeXmJle/zBpykKl/kPAbkFxATF5itrgdFTDVJGNGZnholb2LL
aTGMbRLcn4SFvljMcMEIs4n4C8DDErSPD41mQTZxb8D3q1BCtNTf+XAKGrvvlwUjBrAi1G8yNg+o
zn9kWPvuDwyin5eljOuZXfE1mDcWo9TRRl0MBBy0qTb8cjJVZm1Mtwc6hA4EU3XrxMtPEJ7EFh9X
VG6hXsqaKaOm5OMMoe1lVvG65s/0erPFDuYfSGt2+xGogUzrmET6s8N9yNUJombh7va1ogAoygnW
y36aJMaNg2rN35viJx470tssegoRTyAotafc/9bIicohHP9BVJX02ike1E3hfBASLq288TKmZjyE
dUSayxlYUqYTC+HJ+zoKl0biZqoSLKG2htB/xq4GgoFUgnfdf7GMGZZvIAPVQ8puJ2862rrXXaLN
ej1sH2tPeerg5lEZ6pZSkcs5fzuY43rH4GclTRZrHbNTenc6vnXu0DH5WywuyWHr3myYFj5hoTGr
0uT/w6UDnAkuCxkXIoGjykggXBnNk/X3M/bea0Hld8noXr57CCno6dfWT2mYN+wCPXPtRgAyQK15
oayO/q9HcCKolnlsSQL/WRIhpJ6ZdocnTJazubMiTgx20pBg0MlVsp5+r0PCb/NOdT0zDfMr9yvQ
RvsWeQCoXKE9DLAhHhXVonGlymxlFZw2wMkvS4OMjbDREuj9hOTQAlpmBp+UpuJJ0b7FiEGAn4l1
nHZg3yDmf07nWshMnpN6oCx+I4Qjb7R4i/mu23mJbl1KxCn9XHjzXNTLGJhS/o8xS1UuAvzjijiu
2URVKrG7txF77SiNeIZEyHk9r+SwX1iah0NOUry8VpLZ3CbkmRroMzhsBtS+d/VozNdt5BD1vEhx
D30sYBTTES26mZ/3SOSxrh4w2pw7byM+WU6RjV8+LRotvAzCBNo4xVkhRAacCC18Ukueq/Xas9ui
SlbOyr/tXnt7XoMwyZPQAJeyuAQARYfY4hRDA1khYvYxV+wj0LdPElt8PAJcNk/XTR3dJkVK2ncf
IYtIZvr82qDAYtHGXvHN4l8XwZulJVbn4z6dk2o+ZJtyh4W1s5/ZADOB0IDeSlxhUipF0CAiSp0i
1z3+1BcSzHA1vuFeErqjs++EKptS3O+eR45AsqvMB3edTMOglEYF6UEM6iyKHfj5ZbNTVVrnCPTR
cIobpE5MD+aDVkhmMCrMrLRuzluXTW0WB983HLt9jsbKGMAoPGBaQjFmLAuQTZGHMp+R5ux7E5E6
PgetrfjoVk2gR5+HO4vDlKZopumyrKoqas4gHzZBQ28Gq1+/j3WN0SBqcYf/CgFi28nNXgD0BNMF
bHR5O/W+6FQLfikCIv7dvvmxkmJAhda2Zkxd6xwodfUoHxN9aX97o2hwhAOaPdyk66z0uZJUkSh8
Pm+sKmGf57BoFv6uD5FXUxNp58LafPDKcsCuYr0ExvYTqQWWKZwm9RV55cABhb34uuOFLHKUenjG
gjYu/3XnwkcVl2F6+AIgqNHIrK9M0ixbGndnQtXHwg3o64+3ajyJ3ubq5hndMLH9SgEqU0o0FKzH
tdMGgi4WPRFaRulVf6iA/W9+3zV0ts59AsBc/REl9USOBOq6r/A2gpuR4c0jloCrAUzl3T+QmHQi
IujQ/SMmXTducOaLTnkCts2WapllAYAbAdn9SMmHvjeUgjLpmbElVuRStDKuVO1cKZxR55QQn8aD
QyeBz85CDGzcs91TKNlty6MfODl8oRT4EN2rDwGuglTh+69GOswQo0p74+ok/8giOoMld/+Y3Mxc
NsbEEJX4A4FktfUYyOSZp7JWx7MXDPsOCSsYeaXW2UIP+wR6owJq4uhoC8ZZfkpbllXF4aHZzP73
x63IgQA/oI3zMwzXXFRZKOqnOrQr3wIb2B4e/udeeYqLjdPvcnL6bZDrGlJX3OJqc/nyljhp/aYa
/0Gq0/yTsoVaW+tX3c6nabs7cB+L9kClnLYjazULjdfz5YGo2pRU+ntwhS7TvlI6DUdHI3HBesUi
88kKa58sP3uyjNb8QuqiKfMEBppylFpQh/40hHz4AeCF1nGnnBm7Mt1uycOf6/CdNWRXpycTi8Xr
Ye/WAt9sP9Ujn5/cK7fy04D8wHZVLDIL3TzMXDd/6ZCG/SOrDF6VZsdulIyBW4ZqUe4lE5gJBCeW
xazmMYd74+Yd3YXlSQDZ4bXME3zbmm6LPnIBmgTkooKgHjyTc0t2fbPFhsT4jlDTslNHNOVeMyvg
Op62/KcegUQMVhAJ5Muq0m6QKQk6DDBgFiyRM5Gt2SkF5pbJ9hV9d2CFURJMOCrzlZ7GQfNQmlHD
ISCd2/hS0RbuJ3NeOfy6ZDNx7RFAX2iw8baCUExGZy38ArtG2zE4jtOUXR/3ehVbe9GlACfOEqjH
Cc872Y/0RRj+sWuRrr6d5E9j6AT121KPajumeS5FKa16svaEAIXklSlIo30ilbtJKtKUfPrUDmaQ
k20PmehNpMmWMkERPOrZePQuK9TzUwFtUW1kahnHwjQM+RwU/ZlbmUzsSKEWVQlOmrZ/cbnem65J
YIL8SPzecFy//Fkv5Lbrw9UWbmyIKPZzp5lCHVWx9kLftXHykfOIl57RGkMCvTJH59KHUjC65wtm
OnasEtiFAerrz92OeUuFlNPRK+XVhUugHNijg00D/2U8GzTOKe98MdjiYSx6t8nnD8sHxHlF3TpR
yRzW9RuJpf4Z8jA6INk4B3mn9WYOC1wo+YDiVCnJM8zpf79rgelgoV8YF0j4ylLgjtkAHawEd6VH
ICCvzNuss42LhtYJhHmuYAcJa10ZDOn9ylbkUlTO84t9efzOF80HaCILfYK0GkkglU4/lo2hFq6y
Znxl1SGMB5DKSN/idD2cj4jFn3hCBVigrhoLmEyfzAetUERnltF23AjQDlucSPgQ1CpFNym3QZ00
pA07mPYnHwuCzkCYK3jFHd3jqYlv/KaSObZi1345t7NPZ7BNykSXSDooebwHzwNJDwdMJHcHqRhB
mKoQ6785LNkbi9QnnevLyvHd+iPpEJ6TnD/I+tw4QGXZompX7qw4hqK2jN+dBE+P5ADqXwLDWH9c
fjQ7UdgPZyzN9u6b4GV7Pvs+z3rMeATJHDB2KhtgXrgVVUQy46mSFUBWK6DXkxB2pyGwR16+THvN
71HQQ1Rf+PoBRipdLtWSGj94aaUwZZUnEI1EavewnMXNB+/Epqi3eOv2eJHNtVkOHnlEyAAo+dkU
b9RE1/LMcW+BFvq/FDkhdKd7byhip/Wn92h0I1nqhcNkNCJvpGD5gasRXPkBzC0KozHwonGSwmBc
IGBIise0YtOWkZpHUmbGmOP+pmkG88qdMReqbvcrhm8qBTtGIkeGBoc8iE8D4grn8JP26Fo0e0ME
fQDgZOr8AtKI37g9Ni07PYRJa7KuCAnDQFEda4TZ6XL79IN+Fue99jGgiYoG1ZA0faSY5B0JdQJV
Xhuk/JdN3c0Blp85Vj+MWDJhKwUAzUbdf3STBYSfe/msNwi2dEWU+t1tbBevbz/Pg9f89uTG7YCD
wCdpU+lS1HPAi072uxYnphsSwrjECxH5NQBVVlX07Cn/JSUXSVvdRTJ1skv6iyoAmI0MqHwLVsvr
BWWIgJfq+2evYTE39q7fjsnylcRx3hJ8tUr5LQ28EqbM4+ih21NbQLD7b/uMC26ZfB4P+4O82jbU
umngYKcWULwNqY7fZHVc0bZFDh9DQN9/2qHh5K8YA7f4v0lCYIAwihN5AAyx2cBBzUHezidbAlpT
qqalH2xPeB+104rq79FvVS68MgWMZvMLDvSlkRdySqzGleap1OlROk//BSqL2hRmlSsCNJmxWsUu
h23QWvOt2pcChhXJc8IgVcJtQB6oCAojFSnTisD5INM8HTpvRrGvYA3xOaJKgJ1aK/Tbj/L7gpcO
lqEYjx0TfM6cVtREQT6vn0VUC7exEIr+fEuptNPjSSKs0jAzTgVmFlrsQXicQLn8j5IDiLU69LX6
TMGWzfi+9idDSQQdERcLVY2LQ2mxOxkjm/yHXyOJ4dehuaReG9rEBO0OVqiUTGWZcaCzTtsXgr9A
l2EutdFerkLdF9T4i7GaEWeNpfzNTl1BHr60YqrHxBl6U75n0Ix8dwK65YdIv3ne4Te9wwNZFvb2
Yb3nLJCd+UJjq7KIrjlFNI0V1vCY45eRzITm4oyK3fSRlEfGzZ22nC0GakgASdbcQSHK6AT6t+YY
a2ppX9KMU8SOCIoXfoK1fqedvD65gqWXwbKyRZ88edQi2KALPfdqs61JelTMFMcZ3jOfdrUbdrUK
I5/GHiOK1UMpm5H7fKuMnp67ILXpxyfkUrv719C7XhAK5P5Sa/MZeEOObZf7TM6YmQcURDKC4Bmt
ATh6Vps6kdl7zX5BR8fe+yq+hTsc51kFZDfwj4KOipKZZBOEzylW+EOAdanqbe/AkIkyx3Oo4jLZ
0nsI4XNJ71v7Iv/3GMOq3WhlaA3Et41uwVF9r7mez5NHTp5Lq97Ad6V3jq48wpCuMvXVg5qT8vnx
tnEWfosbajGkK9UwerPP+ED1KBzObBmq5E34B89i+hfrBtFHo4t8D0UE6jeCCKehFbK9SMKNHnC9
PkST4QN7Ch1ELadeLnLx5ginsAW7qNM2Hzio8ed5/0z46uzqLgqz+s1lz9j91mLG8gAG97oklEKK
P59wRyHBtVsqjU+rktDB/VE9/pE88UZJ6IYZD57yB+tzY89O9J7vUn+yqRa6pe5g0OEP6JOAWh2X
9VkecWOr3bFGmX+zhI8IbKlHxS/iDGsTpWmGGvtatmbGzPM9K4uY7yJO7mW6buD/Z/s0TJHeIbrY
rycjLIcaWVHSIceOfX2vR7fotnJBMoljOELNkCwGFuaoJpikrLPaLdkMLwqsB6bPpxFxAr7eJQJh
mNHzBSdMiGiHIgR11IBO4zDenocNyU5p+8bF6D6bVRZfTcofHoDv3o71q2pmornjcx8DZ+mr0pR4
5I0WUYyISNzh3oL1TJvm7SUpUyQKTjiaskjB7nLmiPCTQSgpj1GoFpKyBJT0DnSWc0+pYnn8C7ij
SkxMX+vVgwvjNqWUWtGZRgzYGFFZnqvckHIDf9FJIYfEbfH6fsodbJ/i4kRRbp06OAGGCpD+Z3Rv
0JK0Gz0zvel0LQxsLrlu3GyX/xObDtJrRzm6mT9prrrj9PlpjyZk0uumRWi4JhMdRSSqHDhkBLvq
lExJ6zKa7qHSIsVf+Ukco1wGUsmXI/GZTTYU7NTY0bdjNtEXkGThZO9bAeVYucs88wP6rFQm6k4j
o3hVh9QO0ur9pXsnRfSXB7z4yNo1oqgV84PPZXuJ8x3qNMzgGk14/UBC1lBIcMcH1z/eFpgfmfRt
GvI2uIshRd4MoWz9alFUtMEgPngwm85fS8yujevb9FONEXpE1WzHddGuPqjgSVbFfLquzQZO+AAi
OxkIpGkHDOOdgcFDrMSOV2rMDoFlIRQiFR0D5ieNZjVPl2QABg+YNAxovFkClzd34TCfRSk+7LTR
uad2bqipLlZWOSFYpgYQNY8aGgbqhfsbD3BqhfaC2ZHNnRP8wByK0/1tEE1zbYi36zgij3wQt34O
gpO42ZfgNJhsrZG0jjxnvCcCb/djOQ1w9/oUO2+pMpmDmHpuTkBsQrUKWl/2MwVmbaAk4j27eNDn
2L1SNgqZy6sYOie4CjQFZabsqeCQQW6FkoNxj358jg9dys1LCC9H8jN9Bhoag0YqCGOfkwgYYEsr
z9UTR5dN4+e3rM0wY/GDeumorlB6+fCZ77z8OCzhuS861idQfbCssAepBOdl8sMnJAPYu4/4/xrh
oikbObSa+5DXBpVEaLaO3/QUE3BU/BcQULDy+zocaHTlWrQYwncZnsfHFDX8S/P1Vg3Xd48zIh9Z
g/fvCLOkTbFFbXxl7wh5tTnSLGMYHkUBgM6LpnfnKajEoP+zGVcAG2KlbzPga72D5FXjZwQOegox
Iiw4zwQPnzO+6JoABtljd4QHT3D0uJ8ZLJOL0o4MvaH1vQfs1DsO1DCWP4B4roMa75YAw07vX666
VmvoRC97j3RTtKzF3cixBctmhlW+MtNmOoER4OxNU4Vcadkyradrr3QSiqNl5TUDG65vIc5lQuFD
YJm5oZyTlQy1/rWnC9gP/pRs5T2xYvDvVRawbIT228tg+3WSaSk+XSZtrQAjwFUgeBflILNOMxg1
vEP/voqCybszydGf/kKrXw4kFG2dLfIoaj9Xi1XWrQJix1DxNQmc7I22vP7DjLwBL9femVo3713O
oouqAraYFoxZ1aXP3g0/v/1GdaITBzlBGzruBZMoE30TB7Uy2hfFr4tMzQbutQV7dG+rS0RfcHTh
53+NqAwVPZakm2TMiWD8GuwO6WR/FI2WguSw92ldFgHZGPsCqc8NBH0/C5tpFWfI8HVSYXzvwLhc
Ptpexqwqnx6L1AFd5vxQ5rsJISBjskbdiCufXJlaFSzKJ9cmPJ6e1VCQguNgY5QqbvwKHjeOtIAM
KgI2FH0st4BkMfJlAsykwvJFgysLfja3dUN0+33U/hUFuQ0hNuowUnToZDFr7gmzmLzPKVbA1bZ6
PQSTjbc4qw4PLz7txO1JRIyD+jfbuWFKJ1C7GBpK1Ud9bX82NT8iWxOS/CU4QJg9xTZXp/IO4QkD
GW0XAwiYY5xX6ulCng1BSYq+gBZA0NZQRb6GrPOnndRYHY0+zQ/R1Ejvq0XvbVnL+GrYmujGZPpi
cwZRNbpcWwLR5uv8CtqLS952Tzbda047ACSVccyY9HGz9Y0IK/0AAf84aU2wjtloM+tyh137+kJA
Ov05CtEUqqMhLPhE6d9zjypbozKbDWw5HWLXq50uDSHmRrOOhe/JX55T0AZWOmCKGj0j6Pc0VmHJ
WLEsiMy2EEa7kRFZKLq2VHqprXNB064cddN+gQD/AgjUcSDHhTHCw9kCVFZeY+ebI+AbBPTrCKzN
z39AYQxvWsHivyS669YqKwpjMVlJhsDGDdr919039ahfNUMw54ALWeH1WTk0OqMb/c0NI1uV4jYs
9rD95Lxp8kTOJGvDx+XRMyljvjRlWNHk4ZHG62is/IySNlYiB5Wa36OOgtvdjYfzNRDcxeNKu5I4
ntaJLuDyjGoJabUjeWK1leJaO5Gv3MipPdJIAsIK1nugRCAsOWyEPt80nR/ldxhIoMFJyybUqu5u
MBJbzjGOWtVuSCM/Qh6C2DNa4Mwjps5ATszTY8H5jnIWIO19xd7zm88OckKStDf8SKpFT/L4/Kdm
C9nnqY0MJPsBqKjmXJNl6Ng/+CzOMPQRtRTVZl+f4B1ZYMJ3VeP4cG4JmWiMYSb4ITzfYZY0sSbz
z2oGT7WOVr26PagodTlypG4nHzXUkT6p9kR+hBqbq4Ci7oJuUpFnt4yUOl5fyx2qVwgTrDQqjgnS
MI+HPlEv0fcPoR6juAFtJkmmqBy2fB0TelLhNwLVzHM7asZqBpgX0D6Aat2tD7RM+ol5ghzbcgf3
aEFuicWLtUdf5NSVcIWRFAzTS+3PUasTrlRdBAm962AiM+f6FWB+GBIP0+EIBr66wAW5HfYhzVQA
KTEPo+IXwjfr8pxR57uZEB/gqMpOAhrGGmI5osLPP2+PvI5tgW5GsNxBatCU/+kBUMWDsEiYRnSu
g0GRpZAa5ExMleff0ZjOvscg64LMFMD0opN5Jls6BfXPgNNnNiQbAY+EHxydIP0b1BFd9zGi1XhD
caHPRBYWjfNMsg2yYqYQ3xqydoRrAHVIPoaFi5+29R6r6my5Y4tXDVZk0OGgoGWcplrS/I8Jn5Cu
Z5WhQvk78vPSLS3G5hpjfF+pXH9uynVIRKBCS8oe2IdSHn0pChb3LQu8bQXKy7vnGLvSiBWA+n0+
n7rpt1/h6/M2TBSLPRc73yZW9oXd7VExxXhPgT65nfJ1wFWVpUB7VAWealGgg1lOsWbtI3obDD/3
nHkB8taEzgd4LPIXc+6MTmk+8+dS+gyNSPkFmy7T4IVfAYSWbfwKOnZTqeZ9U1tmsQTI03Twrtg8
yb4M38bEeyJanrefupai1n8I7bbK0S6scsRvasCrc7tZhwgFwjOnVpv6OwvZMzNmUprsgfIP/IX/
ObmwHTtzzYv+W36dWr54ExkFAEz//2RFt/u2X9OuD5tGcT5RHRlPILN5eEXgzluXWZGWGHzhViEM
NmxtYvxNXXJ5leqc9kxZOsC0CK4pCXloW3TlDrJ95q8ouAJAzC/43BUJt9ugNZSNPabYuOAtaZcB
Z5zLutTpnE/lPV6c6tH5Ms8P8F2I7AYyvtv7ol47BdT+vgSiCoPuCmd5DLA3FrfBXufZ0KlwTKRo
qM1LrSszFfMx8XS9xjBleqYqb/VkTKvtNPx65Bj9/vcJpXIXcCLZh7D1p9n+tihR6NQaaFpqjEFx
ztHamIAarsdWJiYTanjEnyLa2cQlvOu/+etyoH8GR+hiqFAPfDYtbgsr2lqGCEod+hPgH1rk1Inz
cuPP2FbZlCj08TUxmGUK851J/ROrTu+vUAqolG6iiHOoF94H81P8o64fBfiQujOnWZpxYPfFEeTJ
WyQlaQIuf5KswySv/Xe2Q+UdTlFAHTBAtC962icy00eqMqXj+TgSkVGs5tpaG6aSph/NIQIBFOJm
4d7bPHOR+gDcE6U3ZA0Xm1DONhRyVKS6p74RuhKw73onvT0wBFTW/oOCMM/pML2ZWfyA7qWRHrrI
5lhHYSdDND+TdOBuHnggA8lm1DqGjQ6H3FneoaBTBxR1ec4/fyfMK54bwybkllHcwmTWgLJPkTMr
gkG6e4GpOZ+JsNvpWo/o6p42NYEwuOHQ/saKU2l0QHJ5oxwvEvNy7PvD7vpDd0jMngj2Z/ppEUTh
1Hix8JhX5eddy6KGu+g1b5wJ7saFu4OBfvW1U4LzLXB6GD36IDSJsxJ8lsfQo52Ksu1UKIonTty4
AxswzriccEyuvpMPoNbgdKDhr2vZhz8oM4ZrWdIp1NAP4NIEMgHPhvmZfiHmGLl+OPzM1x5XEZmT
hQyrMdAuDrqA4mE9et/lazatSXSKIhBS87UNwZ75tGog+eKgb4EWHSci/fFnLa9+NKfJbIwklU6c
Nq6PiDthsBi5vume8iFrJlaAnFNcMmSP1Rd2ILaZ9QihxrA6BlI+4nsDASVd+80nGjqSRgH7mt56
4+iUdiGaaKk6G04uiNTKVb2vyDBlLU583iwy5PwTXOm3L7hdeVhxJ1z5e2n490GC51HZ7JI489H0
aoQQ01iXU2UACYT81eSCQHgra5Haq87vpfOddKW/0I949duX66hEUuRlBRRMot3PsHaNuVBlabK5
9k7VbEka/yCNvQetE5/YszjPKa3xJp3A3JDjHN/sX8NWp2d+GQjX5VAHFgMZ73uF3JVDePmnZHqK
EBHGD8SjajQdlL8cqqM4SFDW0ZyhBPWdNlJWMcdV2mq2FTnBWKqAJmE1PcTUDYmkUcZ1n096WCcL
H1lA7IqIZtnPaJemF40TCr2hal999QTZ/R1NIAWcuV21ISF9VzNQqwa2RGs0luuAyX3Xf2tIu97S
KzyKW7ciD67T5mCT5nYPKxzLEtu0Bne+ptUE+XgTTgKU1BubL+6UbY9uKWhOa1tPLTOEsd1AETtz
op0dv9kXzGgY5jsfxNXPGxTr3mZvlpkTKMnVreaQDGcuyO6B3cEpObHTskeBCtoAbd80rSxqLSct
8gwuzXFEz9s9exbI8wydn2SBtH0f7qgDiF2LaZQNecWn+h9e2skyf6zR+ErHZwXbfuTIKFTBzbY/
tHDThXW/ZKTDH2JrCFPeShA1/RZADbU562ksRwaoDawfqd7qzhpfLUvQE4vf72RO9miyiV4efGeR
kwQAfwUx3VKowle7d/mLRITuOpE7z1E+2uqp2HxOaoxnIk4kASIDIHIu7uNIsHinbQkErs1FClQn
8XqJqaLG/yOlUXy4fv2Cyrl5sduhzNyszAJjPjU55OC96fVH3ZNC/I9HNHgW1yEdj/NtslLrqazT
VByYEChfze0=
`protect end_protected




`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
AFl2kw3wjuupeEJWAVRMjvI4n2F9ZwKYCyTdtTbrj99jYEYTJx3fm7Ch7UNHIYnYCZk+hug4a3M6
XIrSFOf3lw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
kJIX1i40eaci6RDbcVVzg1fYaa68r2QTZ19EbYvWyiO0MSVCOi3GfcyJJxOR52/mcv4FD0GrKyok
p1d2616K9ikEjuEHDsOkFkQxSSfEgbSNAEkwJoywFb1NEza/LgnXq4wCMserYGd0Ho12V4osIEdI
exWoz7u39lGc9ZiaBS4=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
2kMqoMFPLn7FsBBTsV6uCri7uN+peyfxKN5B0t+cAsrbL+lDiZoUrv6niJBSapyempvdNVVmTzxI
0OOKA0SUZL7oQT5S7r5QAMg9q0wHtWdtsxsKxFyZXOcUUs3IkLwLNJ9fExPXmVlCDUNWWyZ/Qtik
1q9ZynUcX4DCv1pUeRs=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
uW1nShxn5xYxSfsiNvMbC6cL7GFjn45B3GrJxFfTPdqHxW6l/7kPGVqMN4yc97bwWb5swAmg1/ia
P9L6G5Lmjygww+NIedzfhB4znXCEs1F+LwtP/Eo4UZuH4rQ55XUhLKrRNEqAJ5lTqYxfdIa1JIeg
6YgrU98QHKeOeZUeearBuTROZ6q9d2QFGZhc5MxjU8pwV5JQ++j3EkUIuMZJi3DVdwnYj2d1DzSG
tEt9nWmDzn5rqjvrP0c2GlNBg1tCMJxGfC7y54n+J8H6ETagMe97uL4QvKLTEhjArVfHkKedz6Hw
BLtL2VPOf8fCVrM+AsqxA6SscLteiE3Y/tcuqg==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
IV462y1jHGYFO6K2VU9zTKlfXJZ4kSNvewSr8uczSbz2qRhu1urkppbYmZyNPMNjUUiJfr+4xl1K
sPX+MN8CN040mI1y/WRE8sMEH4yPflkbYjeDH/AX8AZf0f51eUS3cIc3p5KYvECdG8h6xmZ6jH0F
7BqDcSAL8OaSnIetqzLPr2v1rtYXH+RRlVWmvCK2nFZ02kt8pCYkp8L5RKceyNIKFWCdOT5JdjZY
4tvHtPn6P1gVHsYV30mBGWhvJczj5zrLjwFlzuRt1FBD773q8FliSEnvM5VLjXeYVAshW6krIgcC
JRjJFfG2fLeH0eKFVJ7kqIzwNNYB0nt3Mho0og==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
gxKMu2AB/FASbqvyKO7D61/XUsdMsjazR7APgUWhLu8z6ePEw4il1OmWHsQOCjylECfctRxhrNKA
ZkqobGwUpbLybNlM8OLmxSq7gFftkFYAAbUlTfr+gHIvTw0OHQ1EytNPCAXJ3C16VMRZRtIOMhuu
qWzd7JSTNzsFNMOGqUkbAJ25aM5fSFIBT9RqdtK6aDtxz+XRgnizFyeXsqGdP7bY03KX5HgTMa9w
sW64LQcPjQEuBBRxSfYreUKE1jQbO9XuIjtoOmZGDsEtv2KkhTAdFbwHWRiiIzAO+Bx945pksp3X
TfC9rKLaXHs75mi0HkNR/3vshocjTDFwp+bJaA==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 122928)
`protect data_block
2tX3OrAL3An0C6eyNof6Kkn745C7iT2vQDuMKaih8hIfwSZs5l1VUtJQSpIoLvUVt3Lbe+SFdTva
bN45G51Q4qUhyyhpz5iXzFVHCiQ/FpTZ3j+tf2ItF3GOHVdpQqgA4RyZ2ABYQVtvCnYJOkCAkW1r
q/jZQAlTb1DeatJGOdOF7GxOnjCm4EAjW0ShPq+q127AqkuQ4GdqLcxOTak1KwcxLaKNLfoXDoaK
rmHEWUrIAc7r4f6a18lmwpWrLCFadWK8jFvhDZa47E0ILSF9cestu9lTf1N6eDFrn5tMIHVBdIZu
qjWoC2EN9VDkLR4SYcgC2+loLRlNZN60uj5YP0TYF2cRb1RUwz2GcBegMXLI2Nuj81ZTyo+w+ytx
eF4Yiol9GI0cgplP5kPP/43dXlsM0tU32YVTrEj3kdvau+uPQoLEh99+ugPqRf7WWNQloP+IvKk+
LkKUN6weyyUvyA1UEKnr/U3+8tnPWLQHb3R6V/OoU+240VW3y8r5b5QQZsuVgQdR49JwZ9vPC92M
QQB54Dgwfqux8YN0gQWBSAInxgkZZn83UxuEScRwEn78iqtbWplMBIbme2WVRyl/gBePX2WChcq5
WYh3alw2wPSrfDHETV6hZqGtQn/MhGg6SFyYBn5F7Y3/Tzh1Yu035mKG2TKemCGqKfKBG/d+iOeF
UAmTYN0r5EZtnZbgKJ8fEEDGC3hS9ScJqQvmJlEmOv1u+E2DEV/dGC4WF50FroGmLYxJyhqXAsLm
x+zwqL0+KqLQBqbVpaRX1CCP/Gl9wL0wyC8IB2BlSEBWx/KPfOrWTcIab14XgyoCgZ5zKgzYzBTE
+A6kf8Y4btNhSMzCjgaoT30ki9DPCgjfhQRZyIdXr8O6WTWzr0jcbIr12CjdLRniE/UE49XJ9wCm
cvPHZjfBZB27e+MxpTh2cXH1j6YuMarvkvvzxQfKSicRYoM5CuZlGxyFuDA5yiEiaTu2PxT4pNus
Hr4zY1EvCm5PKhJhrC6gCRBDxk9aAzeviN9pc+Wo4gLQKu0y0PA1Jk1ctM3ZZPOoAVzIVN9DDxoU
YFqvSfFteHw8jv06d58LuRRbaZjmslHh78pl1hVfvEuIWqSdxEht0hzSG+UjOH7oTpeG2U2+9JN+
UrTpWfURm2DSfQolF9KviCAaIZk8AgP8bZ1HN8podzXxsPyH3nCVfbfgOQ7xPbiYJIb71NsUNr9o
wMlMCEv5axZFWXYpe8k0J3/1xm+H7GtBDKuCQHUB+9fiNySJVFFCWa1t7Nt3jrbVXDWg8Kv9KngR
hihOjcbGyYUFPTc2+6ag2oTTOn3mRw9usnllxmQO3xUWO/tLamxFv/J3lMwxyQ6Kr1Qrw2UwZCwJ
0lAt6OYli50rJWT9dYoJPrOfNFze+LtiwTCQsw4Wvmj+vv3s/aBGy1AM0pG5Y7LBWnW6ivba4O9O
Z2pVbcX7OhIkA7rlkZvK4NXar8brE0DvBbl+6k+rCoph1NWoDXAytJ5RFPzL3+uqqRSZkiFqSDjl
smrzqG96sxlVQHS9FtYKup8n6DzCFI0ppXEZfer/PN/QY1xFFa3g3Z8cWiWJIESyycqKOecrPiZh
IU83xlcHYTr34CodGF36/ga5I2H77UHI/6F7uLoJmdVzhX2Ko559ncA1pNoGWhyPEP/ldBs5brzN
xfwTUDKKMRMFVs+eTZf3o1tbz26+uHvUQxsR1OwY8Suyq2fMUrTq5ezCWZ6rdCaJoqAfyjJNx0V3
BsSbc+WV9+p+sgxtBSNNRd2OwYKZVP+j/tq4pH8NOmZPwkxL4ZX6N5j4NCz8pwOiKmYqUFloe5uW
+IIn9bP52rtHJW07ZKoiHpx0fvqqryfF6Nq2sdhEpkM+67v78hUjh+391i6UR/7tQSzlYPsiAMeq
PV43LEo9JNoleXkagjos1iMJWXg1uIjAjYfGyyQ8OnbzxP6wTzS++ectsEE0D8Ak104FU6suboVQ
DjADMuoBpL0knq6L099T3ezhPOTMFJj9FFpCxcQlbYYcd3XBQWPgE+zPdV4V4kwrG2EHCofZIsL1
KwARZjgfIO7INBo2N6a419sFm6EUKrWEB6W+IGol9kL4QqX8Upeitj0hE1cGJwyhvPLuoQKubKHg
ovDhxjSYOIz01sIy3bg4mj0aLBAGNcSWUrQN3C2j/ZV7HI0i1TaZh13csifDCsmJ8aUWhXoVUWzl
W4owtoIJvML+HI1L3LprMYen9nzETnHNvdFOfpFLA5m6NZvHw5u8n0zhEcDbhJyJ75HYpU/aA846
uoWk8GvLuh9iQxZxLnUub521lJQeqMeuQD051Qh0Q4MsryrmT8M1sFwCUIrYU48jd7zMga3/Ewrp
WpRDA9pzZ4eQIODhOTm9dsnR2YjZgNyH7Fx0ToWMxB76NKxaAElyls5Y0XkeV0abPO5TPe6hWh0K
z3hI0uEtRU9P6+cKHLQIwfDh6Ozp7Tnyt1uSI0BOQWc9kyI3a9LckhSaLy6B/9Ov7GR/B4Pzaqgw
ppEBhSmAxznZaGGSGPkPuLmI6m6GXARfsKoYYW8P5NBZuCkOr8SBqc/Js7AqBeUW3+hr3MUddPT1
J6Evv6FS5Cd9kjhwOz4cgNjOSLvPQYN1JCn7sinNma1QC39+JcboQFyPFmRXQjuaQtLWuKmEP8f/
UGGuR95Ckhw3o1RDN8bi+MsmVQfbocDHgA9wLuN6Flg3OGvkwdSa8FzI2c2eDoj7imlxxk/lIzpC
dpkv0sm9LosjAjeE7/hf+Gwwp2Fs5RaDsZ5DA9TLDzvDhhkgVAdlKvvA1meoYhO5QhdT6pd74HF9
3Z3cDvJpf/sz5tzEUa3ae6PsSCkQ1mHyFKtGiYL8PTxPEW7seSYcB7qjNzkTP+dvjZiEXPQK4tYw
WS8hWWWf7YBldlQPapXzjo0XaN5kmHyd7xRy4zuHE/eMgA8vVzIvLrDAE6zvP5KGn80PuKHVRZji
XG6q+c8oI5KTsiJ5D3JLamaioo2uUdxN7ILxZSmXMLyb37QdUb4ni99YnADQpV82yM8v4RX1cYLP
eEfONU5VptuAIn4NVjKZhLW/zAm8RtdDmV/VN5cOT13JKWUQjfvk0rCg4Et3t1uv0ZJkSllJ2Mwh
UGsSVGeSJoH1BunK1xf9VpBFvO7wKXjOT7YN+V/LoQt0+rilzRSY+Dmd54ent6lSyEWRPUWI3Wfx
jk1e+kDb6XfyZa9erzi/QSvDwdQl0Fvon0rWv88Z/XCdrPXORH0fw67dad6MAsmlQQLtV2uabaXq
bSicO3HqxG953zbdtrMbJYeVR5niiyngBZdSLIYPwVrFmKdc82K8RZJ3XnTs8RFcS+PbdHRPOq9w
m2vS9YQvlpqngnTpjt+pzVJAvsFiV+srSj05714mDYnYz4dM5y97rfB/K4wAKXCuU7Zo+7yRBvHV
7Np8xsVxLCTF+GMa8JSFCtMjdV0k0i9rteLqtuSWsCj6oIDY6imJZQJ1wf0NnfFt86LJvRzWCtH9
HPKjaot0FJXVHlB31Mt5u81OhX3J+EU51soaf9vugSjYvIy5OFUoebEx1QXscOJGcWlShN/0CByw
O7WgEO9GheoRU2RRy3FXFPqgk24yu4HTNeyxV3+tUHZV76WYNjQl7t04zDzFrh9PZCh3p8Z8JkRn
O0Bsb/Ekb77rOVshU+k4C3jGb5ruF2zF9i1hIp+pp4I9lUBDGVTp8aoKQVcXBghI0PQEM+doD0Fq
1+bnwOu8UEsK7PcR79HcVcBUq8IWnhJ+1jbe6QoWGN2FfogIxq47faBWCL3P2Rv9214KMHh3Ak6A
YT5KVWD1OMUgm78aFC3FGkNpJU41m9Yk32y2zIgMkIvV+v8S0wTa6KhQPmwNy37aaOrv3Ve5+fFs
lwXJT2r4KamOyaYiYJLYBpLJXWk7FhKdb9im6CNESGSQKy6iJlcvoWm6U6si1REsgJ7giywmN5Bb
eJD/p9IJVBL9yZeM2kVuFMbq7A85AXBz2LpgsOMBLXlr0gD8PRa0rYb+ZaLCd2WqHM2GsI1fUEdV
JR3biU2+fm5AmRKcCLdhe6+lQjMggQU5vaSAU0zW993Hgkvx0GNd3I07oRGjyKw0mI98k4CSR3Zc
XZtMemSIZoI7jeUTBQgdIZKntQ9V0WbFqqg75pKlSd9P2f2+3j4j6fDUtdBwY0LRyl1IQ8v658kF
E9TTy9GviTqefxg9OsqUkEQ48ZpzWxx0abWlNWYIc0PZv4u63Y48gSZFC0BCFMPdLvMWuHgGlNac
O49F7X2kQJIRAkgXeS7Mf9mME5yw0qrhtd9u6OtaEUjyTfj9pKB4UUurkOOenNk9401tOQCdUiz9
rOLZC3/FlsqO8VUwRbohT7xuJkywhHDzdXaAmMUteWyM6Shx7/s7ECq9x7hNRymd/nmzEz01GGzv
f6ao11pkWJ9gnV48azORiGdo+oDTs9kkZ2SD2+N/ACFxqvsWDh/TNpgUmwwN5EhT56nxXaKDbS88
B4FRoCJXpNDL5c4AeM/9Q6pd+hCp4UsRJGrjKG3QxDDmEGqbGR0R0axy+CIX2azav0yfbVnZLWzC
VsczcXaNWoStimCygMBIazm4AiiVb/UYqH09vyW4fkhcyFVMIZdtwtxT/BbRlt8452kHdiC2lRYf
ChqdOZpKD7BQc3IvLT2XfnnLZE6wcKLXz53s0JM6Sg32dNf5eN0GemyKVFR0Im3d9pFgGu8xmu/P
st00IbsKQ22jcr5H/9AmBHmzU8y8oQnGAkgRKDTN3v9P+20t4djG+tWEdVbgARTbLbeQZR0lYvNt
FGuMujljdVLIFFcY/RviKb+NzMKrS7Auo0KpcUF09Z/7Hozder826gMWfAMfW25Rm2mIXsC8pMXf
SjJbGs2kWyKU6mwGy8bvrfSUElVhixKU4CYJmMn36Xz25APVZKPtp9+72xccuoPKgZZDUsp8rL8T
7LG41HVJ70bel4yT6EaGbmMpOhxazlpxh3yshQ9fnyvkhCiHYcNt+T5XiT8jeE1KdJNQr/O9Lla6
/1PYNRDcQaH1xFbI6ShIEwA9DVOTfQX4KEPd052RkWrP7+qMoMkgplbRvSVxxaWjBLxccRlG3nL9
7TeFnLi5+/2jLaUSJO86MOuMI81uLh1Cfdo4ao0vKvjXMYfLZitJa1vs7fTnFRp8lrBncAnHcZvL
MSHXglXKRFMXAKT6LZUeSzhiRODE/fvBYcDeBwGJlGdMjGQxX3JrKp9udGSWq6ZRm51fVhmusXUP
MlnjyBAFQAGGkkWzGlzecHTt8xPVH20LCK8AD6BPGoZjj3i4Lx/64b6/XnE8r3W8+sxOQNbI/nJZ
De2MTm02comRG+3P/igPVRoxP3QBA3npup5ac9Xp6kFrIPaPDMS+RSPb/N3bdzAjZdKYYKiVaRjX
LoZwXLTh+gRlyEpPaB0ncMsXX1H1/6dK9dqOta2ZfapFygKrj/+zORHtbuNz9XIOelc24kqkouQF
pF+BtoDIYvMjQ2o1zCSm6AdvAb6nnzcVOLxSuwG75f+YYNZ4imdNai9ZbQP4bvtwcBhN47NvQQue
ldlZ+MkTHKNJAnrRVD9Oy2MskKagrOGpM8ouNLUgf3hyJGBWN1C8ERyUrloVcPwnBWzNU9QO8O6j
vv06opQz6N1CWYEydYw39kMUwDx47Q70iQCxvBk3RC4LEMd9mRMU+gICwn4hYkl+iMzdDHB4Dxnm
5NH6uRdHCyCKOD3+cJ590k8WFIIpgAbZkZykuka2tqjPnGubHK+/fVn3BGtVdbZrT3XXX59TDTbN
Ln9ocNqg6Eh/kSQqOyvstf9iIaMc45MDCxcPVOKDgv+NNCvKc3+yQ79AjVbutWbf1TQDDPqnXC69
cYjwZ/0eHD4gtD6/r/n9hqzu2suaDZjm93pLMnEmkBj2EpjMOiCPMej+v6epBIPqIeMyO8jOmZyZ
soCmiBoWoQfCjXcHQ1WM6JuotLKM8eKVgC22DPoF7ALwH7cWP96VGkCBXlZ9K95TtrNCaJRf6VQQ
k9RmLoSJuEaFQQ4H+zpNI7wb0wSZ+9WNompwIoE8uYmdR2jvyHG24B3UkGoE8m4rnR1qMIeqeY5f
zWOOVfOZGYHQo+9oqFUGVcEUqP0+om+Z9Z9EFikv8XCV3haDDN8KqeAnKsj1dnVMpuYzh+lBwPxs
j8g2x4OUIcNX7eOfvR8AqQzqK0F+79t/GwdcWZXc5s6UrY9p1JjLdjIGDVq+LBEXp+VcNaKFjB3D
MC3MpKuTao8OnsRB7xQ7bBAnpaT1xCvluc/ctWemZfG/4EihC5ESm0sVSb7/2oYkj8SbQQ4BMg/S
uuYe6rUUgbPPPqC3fNWlxXoX8DS9V9NeSYCkQREfovHK/sOri7bkbLbygkCnxMrQAYVJocnHFLD6
kKOtIMX6tzpXxrASJ1Dok0R7UgIgunF8kWD+GCFWWSOVSLKvuKQZOBqg8Ja6H/5ShGe3QLGgSEWt
BsvP/nhHV9n6mQcA968BfiwtPvkNJ3Np8ix0PwWMNvsq8PVPIToSlGCOxpU40zQshHah3I/EiBbZ
/q+ZRiUFXOzqdplnPBUDWe6Dp2tqbZ+6x2HyI+gQAZlfhpbSturUu4eLD2p6CuzXXvQ+CP3DsALD
aL/wpodi4jcNFVgX/1tYd/dAU0SQBn2/svoaj+rLLuf4Neul8V9tgubJUpr2ufdmivLhDzaXbgGA
eOAzViBd61hu1bnQvt75FHsQ/g4cWxLSxVdhCM3+dFTP9PuNtJFHLkYbKPz18E5ziQh99O85fEgZ
B2CTcMREghpHKI4JwR1KlRTeQrpKsbva3egvcmYVoddz/J4bI+bBKN8jBEh0Ef/czNbJWubxo3gs
BJ0TRM7Fp0Iu4wDlw2MU0gNCmvZQdo4IIvtpVQkwGG3ax4Nb6tISlQB3GJ1/PWAEZ11SnZBRssSh
kg3BSGmuhDehYU4Y9CuGtw9aRMF57+PZDc+hGIfg9xEKnsdlKJa0AZDyEimsceND8ihSWRl/lAfr
ADWOgM3O9OuO/PepPFdf7UKBB8NZbJ/e3dm+5AdtEEFrcVGLKFoM3wJ2Exyq2kIfx6r5AqUuIEby
QTOV6DSrODI6nchpsi2faEsifAUQNXzNJ5qB2xt+5dEu8+x4Rid7GLFDO1vtbRKkcm4Zxl/1DmG1
mFbYUpUrJ+8et2XdDh2t+N0XkkODtNPkcdc7P1Pkik5n6WGqQhHgZg1YF+AanjqvcB+x7VEX65UP
NxzaO71i4ZV2Jcofqv+DeZDROHG0D8C1jXzDh/v+sf3Lj+iPF+gdy7tt5/2BhCWcWM6hmKeQF2cp
UwF2QwjdFVWyNTiKXE+90w6mwbCvg0zHzfynsuqNdaepdGWZHNANDHZngTcJWQRYGuhP5vnNmnKs
vv2Snm0Zn41TBAp4zvy1FmUwRz2xmEftUAbEcvMkp4CaNg+MjtmnaOvj3ujprn1aF8E2weYD/XZn
FGTJw+/TYg+Y0HH41HkhRhXaMZrtPvK11x/+6fqM4jK7M2KSv2EtFM/bxXplFhCEmFfTSPFh5R1E
wYJSnoleV0HAngbd/EQzi8wt6J/tWzYGqxd8Z3KtbU6Cs1U40VDfbmBveJ18DjEAsOMxFH6ew2Ys
cczyA4tiom2QprGADLhRxVmufr5ShEvdkgS2kL4TbjG8UZrjvtMplnvs0b5lf3mupftmllwnpn4a
swlXnIt+99Fpf7dfLpq74fuQ5SGlnT+nWQvdedJ28ZrE6YiLts0Z1HhrmPXfUXEw9cvSCNPpeIOd
l2lnFbjT+msAkotb4ag0tHr5G1Z+AofxnNuHmgbh1l0RUBotHFJEKOszjNNuF3Z7Ny4r5/PBhYVg
Qu4wAPNckIFct3faCtcGxHevP/lW2ZGjQ2NINm9Bc7cJOFpMqYU02a0p7+hWzDPb2R71lzZ4UYm7
NsymgpMwLAfASrm3gY6CgJOXTu0C25AeQ1BdbWGPxyub+GVV2x68hGfLdC2sL2I1A96rzDeCQm3H
6uWsDpvAOgR/oRxg2KXHySvqFkc13lm/+jrMVfZVZH7UpcSjXIN4IXG2q8Gbp+bXnT+B+gvmTVIB
L5BAsCHtwWNmbR53joLIugtskIuVQIyeUXlx410ZVPIb0Aw8cDbX8bYcfdEsPxl1r8KPJPJPk1s1
8PK5zW3hLs1QpImmieuYVw5+x3RfqzXqEWSXKdDqpxPa+3endXS5nyc7fILny/ScI7y9DqM4/EG3
GtYZiy/CmQdf3mhIxiQQsFwkykCRVooSMJKtausxwer34/8RjKbYtu87ngZL9/M4mvNF/HjCTH34
5aa2BPeUHKdTYRKj8w7eXogyjJ5lWxuREwPwDOlWZpeHwkcZha8/XYBwP0j/lSeJ8ID/FpgBIGvL
/W7h3qraxeCtUhx394JgsqBRx6Vu0RyUMupHRL1BJHVP7eCf2/2HFptkg2mDomRCob3iIuwXCY6D
/4BvD/0sL38o8ySFnM0svN3MN46J0qj6O/uAIgGXdcWaECRS6bcqDJ49L0mqhI4Wfv0ZRey17+yG
O9bh1uzKnERoAHyHaSHLoI40fzm9u8xpXcPbDyHxnruJDF1INqpGIbuM7k3sk/PUG+M3AEboITES
/5Le+xfFNFaUfZIKbzibTwxHIpuWN/h0SdqTu1z+mEKkqL38owimaNfuQe0LLkCghed4VhGsVUVL
+Cfdfvflh0WBHtsq8HlPQPOOfVrRc3kJ97qE/U+dEbma3EF+Sd4mrH0th/IHbDtV1rrIiMDWDrPw
Vs6fSyS8JzKjHMVdfUJVvJdJk4z/AjHjL2gcPGRO9Vjf9NSlKSXjD+mhKrX+N1wc6xsY4PPt8KpX
mVeL93Jr5rJortDkwkdyQ7KIk6ab4LJk1b4wTeWa+KONzjjFus70JRFTfLurzra6Ft0SYQBJOeSE
gRqrxZPyJupiRQH0jWR6eKL6WHD/5to8ylBnOhP87ifsz7k/seJ1yToPAu95imRiXLdnnsQ1IacY
arCfaWhhRgHLGUdb64/Gg/tFSejSf7+SY/w/i3zHdO74FnoOlxpD4XlhttBqPQ8/J9NKnoOYdR2z
W87Tq5EqMOYq6TXH7D8pjFFgowhIhJph3fGwxkPHnBzaZ0uvXmTNtdQdpmGBxOK7kfcBadelFQ+c
z9vtemJ0YqcQI42N+tAAPVu6Hpjoaf3IT0+2A+bU4u05Pw5MbniyzZ1fmyd0wzmT9ORNMljO7JUj
8UEGqQjbtbeznnSVtCuESBs3cSyQQ6DMB1j3CEAuJgutJBDNOhxCnKuZrtkrs8uQqiN8wRGhdCdh
PXMgEGF1hL86edy9pOFCh/d3FGB8o/vVzbFBBx3XBr+DZi8DsR7ywKHAVWi2chAx7ZwOSlA6L+Bv
xsVkYxROGMDxiW/e0eE6gz/o8bs/aUtIOBMXZ4pE0I0K1vq2m3LS7VEzOStCukzDKVc9j6mcXbkS
p95sNJ4P15NqNPhcJukWrqn82TAhwC4EszGrLkak9HrD7gQ/ISOVmcU8HFjAAhvFBvzKxJWJRtjo
pL13ia5VszncmoqLK2rSE8tjoRYHb/PoSIdGHbvRnP2z6lYwbk9DKpVi7UXv4mKEttAq7C8D0yw3
7sOLDxUodMN5rKnhWHFKZ4TwAcrflM9e0jubTtIFXl0d/TfbZJRi+J07SJ0JPhQVMePjvq0TzhG5
qaHprIFSBYIpJUma3puep2DqKJ9AQaajIK7K81P2AglKRae4VqLEIcgkw2Cuseuq9G+ybD56NvLI
1T4Jn/Ib83BGQD9Ma7x7WzqrXoscoqs3QKxrGJgI+KJ+9ZrtoTLcXpL8tSLQZaYG39CNM1Quy2J6
GIdj4VDGm7Znv8dYFmLcrhY+meQ/dw2JlXnYY4HKswAvs29tFkQ/VtTMxHzQGVW8Yk2MdS4hKV1M
gAIJT74o+kp7IgVmT2nmiO65oZO+dbqoGm5wlSSd2JJUYw3wEuvTE2wuhSseYqFwgah8Bki7PFql
2/fOtmyea+mPejTuP2rcb/6j8GRo4NbJ/aZkIzS3rZS87nAwd8GGI2Qecog8TH3Pkor/JoqLGRPn
/T5p8MJZYE+GmeUVjzSu7SFWqEddowLHVda1jnKQGC0b9MKnQ/U5C+/u3cThLRyNjDe5gYnzeMbV
vSR/zAtjAVzrJXEM1kFwwSw9FbOqIcEhcSY8k3TkN7JczezQQlx0HGlEXIoTYN3xPTqI5KX8ePLN
zEm6UR2zjY+ZX5pQBDMxngEkU5k7m4cCqK7dEOK4Q+A8QJ8Qy1XE5Czg2PYwuhbAW1AK2ZHBTtiC
9V05mPikJsDStjUCZvyP9WHVtQJ7hdX0krZO0cGdlky7n69tcYK5iDYj2ut95DZdAJvXIwFJMY4a
7C6F27Hq+H7cVLJqS4hkfhj5p86f+VqyDwIpTpzLnt3jJWicH55l5GInsbxVinXM+OGKQpLXtqsT
AfrGQXWKc7t+ut9dRky5OYVWFEmE9BSBNmoSKMfxv2iQrmEuC4LNikzwd5JG6BIRZaU+sr6UixXM
tmH9+z97FVOoOtq6WvMbYVMJn6F2cQi2XFYYPCa1SOYO4wWBdOr3r5grVrtyQ2kvoIcneNptQIBJ
stE6qxuozQYmng4cLKxp4QvNOKfRxcKiNmG5c9kexCUyPQ1AfCiDujLVdn5lUrNlpiStq7BgBGfL
DUyrDDIxWNgMxLMkWQkJL3/feV4izA1x1NRa++zWjhuys6QWREVVRkLXHl1nc2weJprmo7aJGewq
dIa4enXKS2BnoAqlJPJSLy5HEPl+nDRm4adpXnRclNw8xsCPDsVWjyZ+/u1zpmSvjaUTv8MVMBMz
2f51IHk59mhDO37OYw7GbJRNlWPVrsmtyFlmCXBKmECzkiLtE4j9+sDO5MpO7nq2gxBWpFa6ATwq
Q9Bk3cJuWw1RPe1GGr/wOhk3FezPJk20uwpVdJiKtXylIU8qXgec75Von6zgH0lXshNOt9swu38g
QIUmeauCtrKv1QwvGGZQGpfHP5LdiPruV/Fv7Ce7G/dJOh1n1IEbFvUcijS5efaNSj2mF+P1Bi8M
xogUQQ9VW/0RY8KJezHuho0YIBYs3PylZKVMWTToDYTAzM80VQ00U0r6I5izDJcG3wSzRbXjQOkq
ZBSKCwF/BxCf7z0xR8V1il+9Xp/MAvGXLKEiDbXJToYG2wQTOeclVeCDuzo1NfSpbhbHcorvTC17
OH+t++95H+qPwG2+CXv7un0/DOAgQcjuD3008RY8lKNkClyggOw8TvBIs+LEZvv7eUpGgZ/FSjL2
Eek0KDUNAQiPX7Q3ZvvnjvESXeWg8VczWLgH6voUmOoN4YhhEfJiT7E8d9irUoQUyyKqKUhLVSFo
Olx88QYk6lnuZvUdS19C3h7eRVOaKEUtPhMKfp5AH6XSp/g8WIXc9Em0tLaOqarCHBYVcn9B9NIJ
WTjpVWev+UB+Db6w3fV70SBs6PcTJPUPjIMMcTkraLnzaf/nYgTBfVmKk+gr7x26/4iDwRSqm6gE
czXUxzVBvRf53HngmnYgUutyVNsE1qi22mM7DQxS2o2QyZe2KU7iHPwLM6wHHCgR53zBmUS1CNuo
dGYpRHq7+Hrs7KrKBlCe/Bm6ztGZxFCd0qbxKQ3rzCn1jAMtRgX8EnIqR4dDRuiegeDzHLElkiwR
CIXqyEXxYEZruO61Dz8sJHIWaO3XNLe3Qs4unmNMNpra/ROFKsp5JJKVRXvKpWplBKdBW1wByNhA
opvBEa0pvReuwfJBt80WgYd5Sea5fV/tR2a038rWF3yiXsMO1F6JglcpKI7sI9EzsswrupdZGOOe
KXY3uSdPbmKTOFS8rM8wFvgWQnChlVc1HMOc4dVewf6PBHqIsJHxhoULI70xZJvYWwieBtmb4rQf
CO4HjqOVY1fDj8Gvfv//VhtF9h+f7Ldo82Z0cQCsBdpZox9Mf5o3dFyphInLDRx8pDsmbPtfh8NW
x+7c8V7xJL2AL1+FodDJLPG7qLQgV2WLH+Vh4UAnZyLT0wlx27s1xihMZ96a2OzbVaC0a0i/4IqD
DqlD0Bbpt8ALJXHxLqJpfeakFXr01rGbeEsu4U27GngmLiI7MCnFSdTkA5WZeRrCTY37+tbcKfSU
xWKKfFG5+09VCnxqEfJtRvwY+iZKeSDT2Rm0B2SXS14B/cGl3NCGZCCFMCyGn24sNGgreXs4c8rq
0o3Fhcbp91Pn0LzGyfgPOV+gS78e/u5zSeVPnX1z03HBZc/5HyzevAjR2PcTldM0t9Szu56Kcqcs
Zesn3W/WUglXKFanTJob2FMm0xreGvopg1JO0/QUe039QtTw1Sok4ghYooxm7Qg2w17kB2BqF3N+
7dKYOLDBPMuAH2hqbE0eMvN70yUQTnq3YfHnX2F5ZZhLMn0wpqJbzyBtJ0k71GZsNBWZPhLKTcGx
1dxR2m+gMjxolv7G9a01ZkkM7XXt4uTy4h+Rgogmgdn9ejWVmsSrUIbMDhH1gyUYUIpYSX3Wn/5F
vP7cQsMJFrh/D6R0Ck1dmUbNYUIUzu2G3BhB9bJVgeLL07GDVI/SpMOwltd8HFHJ4lnt6vk8+jJ0
SV1YWQijeT7Tzq/DlrSeDw9uVVKArlty3a93McWR5f3gEeBw6Jp/3VOID7dvMeyaT0c5CevkvPrC
Y+EeeuyNUTlxq/2XEC+i/1oDjXOw9B+0TG+LKMJjpPI2ArRg6wuiyG3jJbwhK/f3uF6ZeH7a+fZR
sBq/ip9JipwEox4NbMX8jMD0Vkv3cxjcwODT4/8azfuHuplmi6blcTBeHK/xlcvOYLW98XXMcRty
6KQNyy+8bALSIRF9sZnPg0uoztTunYtBB4L8FXnwP9ET5kqEZYTeYv5+tYBlgui0Tg4kcP/KYdFQ
X/45MM+zTZfh2Yc7ip17NN6XplGEBORoO+o3ebLgDifX4QMff3Vev4p5RZ0S4kNWV64JvvN0Osix
mDl/ftqsCJMJppvduFhbv6u2Nil66fFScpqGgPJ+ov1C2zBF38jA8SeSEFjzaHx3eVPXv+sheCaF
gj4yits1M7aK+VVJ5kJPI1r3JUb10eA71MQdiwT3zcr96XaFz60ea+L1WJr5Jb8shDzHZRO24CFt
0nk4hStYgEA9GkmbEAJsvzVeYZFWbhMg0rlo3EvXDqs8++FXK5l2TwxROpOMjL83m7XXtGt6U2PM
l3NLmPg9avxzFwsZz9S2u1qJF3wkdHj9Z4gzDpnRnyRnqtP2Ar4mrBx8Gf0n6LyeGdxUtiofW3Sl
UU9xY0PnspeMoa+kLjsQqBdPt1YepIFTc88M5aVPEiThBbmwwYU5LFCQFxiPK3GB9qzIEtvNoAAq
XQGini1IdRhC7W7MmkjIz+XQ/K65goNNkUbAyPWlgopDShOI8W7quuwqycqiqepXZPfMK+o5WLbY
+7lbH1+MMWnkovuMt5jXEIrphfkAFsAYEjX7qTwMA3qjcH4vhUxZJUsK4Y0OJ4o4QfgBTj74DL20
NgiS44Rl/9nYofB64BCSZwzAEE2Kgajtf2F3qwCOfLAE/9AknvQ+AjswiTVSOza3I/+EY440CDaV
gYH+C8ihZxGEyFS6vFLcpmL3Z/U6l7wQyUTQVJmH6H5MNtOAjBeiUvKOsBoMZPTN60/dF2Apedp6
xLCRNf/5H6AEG7ioWJU4SXAZGznPRYQ7TBa8+d+8euUB65C9GdzCzTkr2X46wK3ezR7Dp6kPfgxv
ycchB7dXxRdn3Yu8dmuHjwsOd3TORpOgJMAA8lrsIeAQQPSI+cr40dFK1OI3hLb+AcVxp0xkoN7/
1GRVUBx2LT18IYm8wrSvtwOhXXF1IMfWhme+dTJi6o+OIaEHcFyNK5BaXoQJ8MdCD4DLHiWYyJRV
DFfGcxbESoF9F0+ewjVeopXry64jqPyidMzZ9VZLXxSQrHcscKt14Y0+LZPLh0r1MUywOJpxC6WE
lVHlAAcCPwHy9q80lbZ1owi3nfzKdTD8XmgO6m9moeFQ5wvQJGQLI+/JZwbng/5oyBIhkPQpeUXu
PDFmxAGu6Cbc69a3R061o3M14qEQTIc3bWq1pLOhAJWHgbnxjkpyXy+1bsrXALOCD6IDd4cXU+fp
CKo5WHy9CmRKStGgm6Js39Y5db1hwwYixKduusIgPT9u+Qb9L992UWOK1OOwYvE9k+8oNmUxlX7r
ckmoqB8SfpcFe8iasULY8MEXb3Ez+qPJrgkyLETCH8kbEMxNX7yL7yq5/6qSJaNvUi9kGLmnns+p
/eXVCTmG2toPZBKW3W25KFikKsNlmV3RBDUbFzjqBScFpTpPmMai3zTGnvYzeypxB0hPmmr2i2Ol
8yyzgOwBjshqAs48rB6G/p/PIPDa8CzFnBLz+pmBheP86IM4IXXE9w33drdkd82Fcgz5M8wyPKlb
KU3CL/sNpDpyjusVRNaUPG6Mu2/AhzNotytVa+FJYXgYKKFEJ4vMGO1KF5LywtKiPNFyA+uaAiI5
lNe4B5CTXjGK8yLFhFYTD5vfzmfr7yrb6jH3dEXaKTWM/hisCLqm7p0BGtMG3+lo7CsJ87VYaONV
xiRd8/bwod4B3abgXW6GXACwWteQM4cNlU5bATIQwiczPCgBPFjXgdy2Q/x81CcLliYAGFn90KvC
dmEv3qaxT2LER0WcL7bBv0/H0wlOQvAiyGuTC8m0ZdYf1alEVWlf1hQ8zZOsrqNOCCXgJEwL2Myr
zEljoElPni2yOvlhfHiIDx+FTIY3z5mI+EOqSvF1x+6pJwM8deCDuwHR7abcyc3elITS6C1xHy+6
ZuxHH6x0gtAZgH0mh0QHQ0EVn9dmFyOkT/OpDtd8VeKK7b6H1g3rcR8OGHuhmsbbKYxKCw2Ngsi6
G8ZsYvybVBhbHzXtPdTKx/DkgB75hA+kell8vAS0TsEws5gbtiG9IJuJVMkquniQ/P7BQLt6Bi/m
D5YyL4ACHq2ldi+haDU5dmLe+C3dljcYATjyWavgNoT1rXBklcAcF0CJ0QUXJeDXPk7+WaNEXWmI
IJ7tmx1aG/K9qEUU6FsKCSTxnMpAprbnGuFUh9FijVmmrvQ6nx5KFphSgjKz8osVWM+YD8Ch7Esj
FG9bPgJDf/kldl+LcxnoLaq36f+C8tGesjOmM04LKnR2lnLrxvfbW8MJiaQlcvOu64YEglQRN3Bt
F5XSKzUngWPCAl3ISWD4C/tJjHMkGTEbXOH3qOVDZqJa/uhi/hPzRqLjfpy2AtaP0Yj7wVxRl9Fb
JGUdpjpVwhNbDxjnh8MMKTQASQKS8MaJcj/lD+/sHYCht8hOuGNeH4CLVhTWbx6BxJHcOzXsT0DJ
bX8i2GaqYYkWPSsyfKjUdMyBXBZvUCqCNCKksDVgxe1CqMY9kj703Nl+I3aV8GXo+DBUCiv/tArG
XwkgWILcNByy3ZsQdGa2avQc4prXTh4Fbh455CBIP/sl38vibxHCmYJTQAkTutIm7LcmcSkN11ug
WA0GEfhboFe30TTEseL8z/KsIXPU/X7sbvWTpb0Xoocpi0hobA2s9FrSZ6JJN7i4Cxs2auToc04C
kn5zjeRDBreHhU8FA+M5DlhGa/htsysnv5SlM1mA+fweBYYyZLf3OYMgD02yI4Ru43qPsDFThtgN
8fpx9DcEXa0g6yL0AdOhNh4r13sWwphWl01dBXxChG20oNTvknA/hCZNX8vHfspWq5OAGv6a5GIS
B7qXfCN2hhPGFOgB5kMjEwZHHmJNq6eavPwwGCoQkQhqBcxApvxv9vQATnFFb9pbVawsR2dvyQYB
EC0yjpDW/+eaAAJsWY5zI3y3lLjVOP396CWdZzLjFuNzPgyQkWqtoEhjJdSYcfmz8fVdp5QWdZb3
YX0H7074U034h90Zd8500HKBH5hbdzr5vYxiWL+eXH9TUexduuBGeV3LEKY7ZDi+g7gIkulz1jQv
I0KZEY7YWpkxyPDSn+Cl6k+p2b928zVlQGi+Sp7QY12mIJNPQXHW/46xD4RH7nFi+EmjkwdnPqhR
dr6PS5HguGVNGNbsQUCTE29b2meW+aZ220du7ErR191T/NuqDdARVt4WPzdj8sMEI1PXoVAwwhYi
S0x2g03j0XGWqtJfHhnLJEPiQ24R1GfPTdDH2NRoakJwDQpVrzkBiWJeb0YuEIMOracCIICQ2eEN
f7Ax55rjs71/Gd2BjEXg/MmU6GbOguGIJjV6VsNNVjEj6N/GSV1x9+GywDSpn4EvbAKLmg22DvY6
fCts1gTtNIJGTldGI5ClgEv/8ulbQtatd6FoEO+eBDFqqhbcc+AoH+6XeZNp/lbC21kVlhfP0/BD
9ZzHgrSo7+JcuickaXF2ZGbwT/P2tS26xcFQ9qDSkLmWk6kJ2lt4SoihCaF4/CFhHPjlDqc5r0j4
wX/TRA2hmWc6ScRUTpZsSldh5vwU2GoAhUCVUlYdqm/rco7yFMhg4F1jIB+Ux9Xap6HdFh1gqUcv
OnrBf7oYJ4FOFMQNRyl21RTdmjWymVAa9hgU9DyA4EdKzCSog6CMr8ypw4MET0ILRnVXhfHyZ45r
8PUxzEaaonoPCyqLBcqWBTXWxgoByrJaBqPOnKAiMcUbpCDsAMSY5JZ1MZN6WBe3al3Lg/CxGhEj
9dLhB0GW8QU2186n7okU+aWgzZ4khpoEuftTXaM/mGxXclSEvYaWvdNAyaN0sUGPT+8AlTFi1yGL
IfN15nfih6cbI4yBpW5Lj5BFlqtmEUsRPx428O+xmNlkZzhD9s3M2KuGW01iWHol7XLRagdNlkAf
GRkgLK9tYetOWo9q6SWehJUc88MyL4PGlX76Q0lVhc+5dHwZBKfoN+o1S/pRCt2VDed2pccshxLv
xhPY+ETz5Z5ykwcNz2JPOyHjy+k4gIBi8GR72sM3JaiDsXan9MkasN4hi+e8Jgx45IJDh/mildiv
twCP4WmJ0Uwn7aiX6DVq6vzsEz+PVyJjWcnLMX3P51yqpCXm7Go2EYrERuqMKuc080vj/UOCTc2t
iUkp9mWDqbi0of82oRtMRidYdUSwy+BSBO/hFTvIQtlW5VQcDyvfRkUwI0pHN0oPR0l12hYgHLkK
ATmlZSgZko+2quO7HQd0CFR04vXZXPF4QpkUu/ew4iNcCOEYsqimVB75b0ehKTdqZRUGHkofUVko
k42RwaTMamY4Ww4R0hZzJ2mrs8gNOQktcLRt4bG9opOx2UGlwE4w/88+v6obNWbcpbbCAp6x12MX
BsH90n67Lw/AJvv4+U5McU8D9bM/G+4a7+Le2XphcbaiXSD6h9oRDG6FNL24Vo0d1a7ZJ67qE1B/
FYbFfW5yU5zFKpJeYgITId9uSMZTHKER5uc9EeyWcrcOJvomrx3qM2/96/1f47YuY3IPrV15YebU
8L+BVk9D632OrOgnJ3O8UN0aHmEY5J+xjK2jRTqPPwNc/L3glPESfwQ62wZzWHCIO1J+JEY13XKy
NxAL8c1m2c8rplo6XxIrdaGeoAtGjr3PC2uMNxwlMaWc64A5xmzErN83r0CFRwe50jw2IuZTM5cj
rMoZ3uh1SKJlDOOcG/ybru1EhazZ4eioQtyv3Mcoi/9ajnWt2zUtxQVv96oUeApGv7P9uLVoRf3Z
UpJh0OwEZ4ugmMbbaGtlGpxrdtrkEsAIPoDz+g6M5mfkaO5LOv2JvZK/km+PQUKxWqTI7p+w5Z6G
BYAsXiE3I/P3wRnwl8ROmWsrLgUOrnoobVnIMAd8w4o3gEelKaIqE+LkAvE4CoRd2rpYPH5pKHu3
VocGultLxysENa2LkUbhDHiWKVHhp+GJvY4CTkspU6HJ3EBtisEt/FLQnk0ufzhl+mu5Kd9L9OR8
ZT2tTsfAL6WWMo4tUDXQ6rVPMtlysUYohp6ptDzbRBnd0aef66fTmdkpJJQDdJMFlfpnk0liAgdD
aRC0K+m3M/0X050mttaDrWtpuKTG3OzyuVH3fDlvkFVROmjjhiCO/nCAHOJ7G3xsXBUuSM1SVKDZ
4ewOWHJH6mammGagRkWZ0UF4zjMM96MYDO+MUtg9Pk1ZJocYMGRmBa9YdXSa2/NO3fu7UUxideOm
zFT7TEQ0KrdkTEsbDuyNJ40UA0FFpFyac/fA2OhQ3G7Ej4S1zjI6yajxP7hDhEv17r9NeBqBuQQg
siyUTTZ80uKOkIOslswYckue9G0FRckP0rcrBYSez560IzdkWc5iQg6MSk7cfZbOZ7AX7fnTPxNj
SRxOzad7Cz4a1fJYYrJCSShVSGVS1qwIsgWfZ7EEt8sDgXUTF/5HBKVBOcPxRPK6dF55jdZm7e5B
IQ9pZszbTMVsi9RSecJv1Xu8uRAbQO+6T4u/a3Y5uiqviFxcQQfy3yZqOUDGrFni3i2n2hQCMZ87
oYBYP6p7HdL9xQIzd685BR6YxjMZwgrp4lpVGvSjsjZD9l3nqMMqLs87zAH0c3741WJ89SvPFTya
iIxH9awkAPSKf/gaax2yzuDQJd63qJHh3nem+yQnrhSnL30i5wVmfhe4eDKY+aXqxEZkov75Pn6E
kSKHJp+B4N3YsD3vfVCPNYTHRWRSX6j8hylT/fTePtxfZnOBIGrqv3Z32YvUW1dcHX/aT5Sr597D
K01NByYc17HmbhGx6Z+QE9PuT+2XebUvjDDN+pnl9HT8ZN4kiPhaBejuBKItCegYlqXpwv1C+Mvn
f3ph7H4Uj/oIgvK9KQ4FdGsbXhYkTWEF4y+eEJ38twEaBaoPUMWtrizE7pZ0x5Yvbx/5wtB2b+r3
dPhzIUuYDTJMPp2g/uaYaJYXXvNZuWpy+33P7uTX/cgVk6wxdzrdEQ7AQhf9m5AHx3NUHFWYuVPB
ydhdJFHzasOAzwDfuGZBm1nQGT5tdGb91L1lenM7VP6fh+OOl8OhdITYA2vbmsnb2QgSyTF8tNM/
naube3ZiN9Sc+4RVQvd47CD7NOkdjEow+5Rau0tZ5X9Dn5oAKjvUaoW9+jMzY9voNFQ44FubvEa8
+xM9JhGQr1N7TtQmkPnUZYRk8YV4IADCb1vaydtYHLi9//EGzIn6JFzIY6uZ9b81j7B5FpHvQcLk
lbGVywwEqzP9SZSdb5SI3A5t6dr65tD2FQnB0gIzw4wbfwCLcT+Q1AB8b5JQKww95/h8mkH4/bhi
OPok36APl0QhxSVUzjfD4WTRiIIoSyATPUHPdqB1x02vz6ix8DUktHCKM6mHPVvdF8cuQYPY6Hzg
nxyW1KInyAWsRjcA06iPN7EzBOHVLAht2Ww5hdcP9+Mns7K2CY453B/2B5B9qnn8OtzwW+/DOakN
J+xa+I4Hpd+25sUC76RNAUeWThDdct9yinSkVbTU7q+c4najcSnCFpOix/s/pxXtsslaMM7VBrLU
2fIJ+rqANOhCPLtTuMCEn0qkW5O5uOz2t6vrYggdXeOIUPaqiSiy531pdbS7Lws1mqySnREojLAN
t1TUwGTqMx8St9UKEmvNBpkTub4+yfMLchtKXk4bOOZGk+cjzCT/EoLpxgyb9XlP9VoHUHvfaWJS
hIkNeYIdWYKz+SQO7qQD5Ju8xYMgoN9jsC9nahvSBLTaKVPFCqAWk5UlbUwC+e9KuErrHD+I2SN/
c0uWN8qd0XIlhfKd6q+O9W9z1EWGhy0X98IdkLsWUMnz8z9VAIJgHtRX4WOpUgpNsFdvbBlTnSc6
gk7XxvhzUjduQtrVlmEB/MSMC+fsDA0Bw8K5OAN7TmfPCW5muBOsRnH0tiYx2iEDyHkZ92VeGq/8
0ikJFS0ItrLK1FfVeMBzTW0G5bdPVek9BwPdfZb1UCwf7xC7mIUIUMY4f9Anax6ba8K5wxEDgGpD
nGmRg9ucv+M28eD69keKNNBw+IjBbnOuw/vS6W46xbZANEj5S0hBORv5hbPWqQX/gPgVDohK3oj8
D+XW4WD9BMxdMU3zrw+8kQrjRMTdZ7CzJPtMqbFm/OcIQvW+yczo8s4XXkHHEwooHNsqWZHbv+Fo
v8eXpizK4OMdmcq3Vq83/vk4SDpypHvVuqT+E/xoVHCxQjU9OoPrghSEis+iYPWkN2tkpekFlYht
e6ox2RVq86YXLsf895E6Hewpyz3bED+hukAJm8TtVx56t/IGfesd3jwy1cudwnb3P79G+tU4KHER
ZLMpayNf1cymO4rRTXp83AE97CV6C+aROgu05V6cB67xTyxP6ARNB9HoyKJWAl3ORc8bRKZ4DNzg
CYNiKWuxXPkjcqz2/hP3wpcqcjScPeCens5aHQdoWnR3/eUbmvlUm24atbvNv7s3N1c+8G6GNwoO
sPP/NTpVqROmksymjoquTjh20r5z1dCAiPnLHOnMFqth1SyhnymUnsTJpHDiQQVkOewqA6LTvnJv
hUfaVWqodidfaa23L09KJwsc2M4B3L/YZYve7sXy9LnU6/zkUG1PTyCHmJLbvw3BltT8rLfcyRBS
G2k1Y8y+eGF10sZecaECY4fgrdkMFeKseeV5IhKVRVXZe4BAyRvWNyEMWpM9rH1hNFjKovcIwd6Z
fQk+KdccxvWCn3m9TupmfkQS4oYq2qvjcgVvdH0rV1HKpCOF0WSDeu7UiyvkwRyaNjK1QzIUygNp
csmOGnsfMK6sEMQgqBDUXY+R+DL4X2g8dI3BjAs3ttR7OUPQnYIZ333W9vDL+kCrvB+3JksXgkQx
Fi9lHAe4RbwrjBYNrIIltFgzpxtWd53iQKVzb361fyPpF+/kchIihE9ZotiLjaNqMLS2645eSk7v
vh7cN+orqlta/1PtBVPkRMheTk45A5s+2EVfgwpppPc2eOG5pxN4Bzf/1mrKwoPlpB1p2WOoqB3V
Cfwx3eYiIPNTzWm/cCjiAUbccfJ4/c/wWFE7n5CWaFS/ZVq44N7+TwltBp1XAjsVJZ+GcXvkIDCm
jY2vPMKHCfm4RYxm9VxlC4fMvxTrfs6HbG0e09emuCsiz7a/EgIw4OJP3UPwtmzpnjuy7j731a74
bHT2ibhkywJzbpqa+KXA3Tr5esvty1c6hni36wzdM4IVrNvnee/hKV9eSN3LFJchAMAVnfNfpXbR
W8UvG0vdDcpxyUFkT+GohED0JmMVhK8BWcjI/8lXac+39GN3kZcsXgklKm1ty9YOU9Yj0Xgv6fQI
AtM98hLZ8+G7xmyhFmWQhZah4e5/n44ee1z1db5Vducx+SpCyTaWGdV1f1NysmnTB22j4A/PACFh
mBWzS/FAjqbyYuOulYTBEdNl9MMPcmNjWY98qPtsLTEOYN7nmd/jNcJ6nYSP666rl2+2pBQ6VhYw
sfgEbFHOq6Z0xF1gBkvFnC6kX4HCZtS5hQ03yY/5JWW4vUlTNAU2455eNGae8mxWymjcXVrcOFh1
+YqeuC3eNUs2hN6mewyKJ3XlhmEK54p9Ck+VMN60yIMFnwcv9rl4SmFOa9n3US5W4GloBjV8X1S8
pvzsKj2U7dkc31cn7CUy5rlb8dvI9PoP2H7GIDPoUBTDk0TlszDVtPzXspPbgv4Ur+VBrr8PIAyu
e2OSv+MUcS96EXiDL6PWnXu57ratDP5HEzVdQD+0584OyLfVU5W4DQZE2MRgl/rJ5oPJzb4pO987
cSqtgzmjFU1GzKhc66IqlECdiceClUyKa8R21KOw9t/XmnTmtZVyIKP7GZNqureUpvQwL0bLujDI
Yq3ZS4mXTV+4XXCtjSofi8ValphKFAQLwfFOzUK8eBe7PB5tipf4vaJ/zG04XH4Qkj6tsdjT/wa1
L92pH5G+moL8ESaTAnTRZkyIbN9RVlVejdY4Tdi+zDpkZZJiLkhtr/kqvu8vsF/iYyY+7nvT9Od5
za0QWjEIa3010wV1+M5l0eFkqM5tnihQqhvsPLVXUijfCjyQWAc0m8aUDgokRwD9WuYL+PhREivE
ngAzhs9mDSsHYRFaq+WtjGeHftAWM3ffFIaJS5Kk3SVPdJF9tTJ64cqcVlO7MSqv+snySiYMaXW0
oUwQ7H/YZEHengsA86+vWWR1aC3BddWpe7jJ5d0lqcZ5A/Ifpz8bK6T1uf2C6GrNF5DxiSspOJXX
PTPKa8kySDi/TZbQcaYnlgDG2HPddUvOYEbn0HJMFcFT7DIdqJaJTCspvAz2Hg7uQnarbbSpBG6z
an8siktZxUfFiT5H0WzY1QPbhS5VRM+Incup945YcMbsR9g2eBW6YEFJYCAcaKl484SK15OQ8V4u
ohPfFWH0J424MQFa+CrkexTAdR44RdbiGmw8wd0/259OOC+3jFMLb3JFk0E65A5H6RO6mYnEoW0w
e1guCWmn1ENnikWS0Rov87tWhjoCHy0cQ/ePmdobifk7MQEdtHezhKX695IVezfNM+HO2t+YxhuD
TtqAmZkAKDj5hmGevBdaSDscLZ/XGaxGiWVoY5SWyLbrQFbCeiz1PwwjfAneDsN950SySrkDorO4
OF7YgWUov9R/EU8XpB1oH0XpauYArVX+K5L+ZmQwOLK3xzIWOGCz+jY7FiPf/BDiunY4X2+ighAs
4rMTD7+xeR0RgNy/0ciISnUU+PUHPZgpIPUEF0ESQ9b7UqGwr1+fhjIubLNbNh60/mVA4B4OVwfn
aMs+rx2w/MI7pHvKj2pzDK38B9FkQ4M4lAOevzJ1f67KMcrpZ8ESL9E9md6QG0oVG08DwJLLXF88
6qN7uY/6M80AFSHbc9tTegNqWtolAN5u/RF961rBAlIZfPX2au2ZjUacd3gEU0rv/nfMDiT9d8lQ
PWH+w9bJpBNZWJUlAO2YCkPGlSy9GhEgDXsgBMjOBDwpQaP3hD1JSi/k9B4X17SIfacp1Fio/wK8
/LvXJBDxD+ugupD37QTgmadoodsj3cx00LZaW7Y4BgeEV5jlXzYnMMuDnV0PtpU14eHybBHkq8q1
wtoK7sHdNmMEnZjlcSSnVPTWFN1U0s7dak5jVf5kqq+uzkvlI/UbCozqziDp43XH6FKftFpzNy8Y
ItJw+u7bnS2td9Fn6PPO9B/mckzQFzLbl6AK9NhFvt8lwi84cJBeM9+dcw+kOU1rRcbm/WWZyG7N
ttjgOQWPzHQK9LjmOYcKhClKj1RiRh1nHUiFXbum2NxJKFlKZXVn+unC+IdZBrq3UkP9nb9rox7k
P3tBlflvi4pljp6K78D0kr/jh9FKf5wa8y8irzPyp/EcbhFkVq2Cz6wYSGJD8vGLWzpJoz4m7ADJ
6Wj65m/YrcwBdbLR0e5hFu6+MOnvn318uHGFaPJ1OVLtUPHCbgcYlC2+RcfxU+Bon07cPeCqMH4B
dl+J5W3oX9fZEGYybLZ7NcVfncqwhgsJ4WSBZSiA8T9DKKbCNLsc84mRWaJrcFeUiUYnGbUZBKbJ
aQ1CG9w3CVb5Z6tICs8pen4mNW545wRzRlNxGPTTeFE+x9Mvv2Vd2KuLau+UPCm2QdS8ZHLKsleC
ukSgtSruXoMUhC73HwbV8p4SkFkEiujSMZrY5HechHftWtKE2yGg09+qBLjIFBFdnkvdSY45xLtH
ANOUmy4wRuLBcIKPy0e08zY3SEe/uBg2FWwWSDPG8HNvn/nZhwZ0pdn7G2h6AS5ZNSfnJnhXZLq3
mK9XvLGsdrR+DoQ9lq7oITPq/Ds+JJgZmHtf7MKWuRLut9ibIZ410j+meScVBANHqDHwRuFKsfGj
JrJEseK7TIS/XnoUzYxKsb3l8mTXVlZxNi7IAd/gLL5VNHn4kcysJ2UxLq9wYASI0UAJt36B83Ev
cfk3RhTdaX8WZGQkej2AlMAKmOHjrtRTwH//1fYDMSVaY7Wa6dD7LHoChXzF/GAgVDehrACbCgsN
++U2mKmbGL8vue8etoO/O3eTcJrrSkG6DVJfCisz55b39wf77f8Jve7lflXLnWSN5wVt+sLoTf4M
GIptsAZFVCMJ8oCTkFrmRqq/gkisYylkQRGU8stbpXIzZbIlAT8Ny7v2u9bxHvK/456MYJt9Pjxc
vkWZLUzb3B6KKOhetyhiJ9MeTFlgKPVJ9VvsFd6MR4xIb42r6O6RNnBu9iynyq74ZJh23Nlsvns0
/W/86Jevgqny/nRBfOWbeNPEAIiFXf0LtW0/URpbk289/UEufcjlDZdH+Z0l25gzaaV+jzcWASAX
jPITSVm+Tg5r1i0NzXnWZ6P37O3UHrjpKOosxhgUWcDJMmJknfIsbFBbxl1h8MpuzyPx52qALAsl
pWskR5m/O8YlV76yzImczb6yOsdWbZZrk/oY7tEQgOIa133pnaq0QZtZqOQPZbO/dsesbC+Ck4zb
pnOL54DzuVvO06HAVcqrMhvuDm91iMjvsLmqzkofgSdoqNNCJm8iFTy3InIbobQhfHD61dBmFsu0
Z6V5cnE6OyAnfmp8agDvzr8MpiANL7/tuedhiq+cYTKHAdwqeHMg2Sq5VaTwg/EX0BQFoZqKZCgu
X/ZScitszO0buKHBhT/xa26Pnl8QUS5YPEX9w+oqrjXN20DJMiGfC5Dp5GnM7zgnoc5R1w/p3Sct
iqUyEQZtUUar6zWv1fN+m9iF/WpuDfg4BzCiztXN86E75hpfPOyepA/xJqRFNw1R7DOJjREM2xx6
exRlo6pZnL7+J4xGW43WTa6XCAeuKRCU2VNIEb/c20zxp5kxGuiU5WmcUmGiQGB/bWNtDm0F599j
8i7fVWRdZfyoxEcABzFhaOQU1sDxZUbJqchGVJoZmyiJB5kEnz4NUxOhDW+SfjfWB7XDgrz+pzVR
Ci5tM5hlarZW8zTyOYJcxaOueGhYarlqLbeb3YG2NJFZTGlGzCNhmkky6HmxM6G7CauD7gWijlbT
1aBGm9cavLZqhZDoKE5uZzDw0wZXIQQlvy6K2vVUifHR9K0t7rQVKJJhP8A1MYCN9x+Dgjh+NbtO
R/iXlpdsJ2q/vl3rPkopnTT22086erOKDeoA33KPb9qgxzLQPgoMFvAn4YphbY2Inv6BdRu/CB5m
r3WAW66IsbioxcMgeIPv/AL7gnEsvgnCigGTu0I7vaRU3+p2aFzorbZuUpgrZ1diusnW/n5rMLCP
kQe3R8IobnaaUwdk7DSx3iHFmXHmsNsCk9NU9Ym2FCOrrtkhHP1UWPaEE+rXPJCiK0HudnqnaoLk
np4E9mUA2g7trJJc0W6urJg6YWW6/czIKmajtjZZD7f3MHftGHRHtEcnVa1VtrVBOn4XU/mkM4A4
OmjDpaPB991nz86dNiE732IlJrdXEUIvwPlsIyS84dcuosj1e/kDgC/hWKvC1i24YckRqTJqVvLR
1gGq8ezWHeTYjcryUKnrL3kURbeKCj9qhgupUwKnZW/GlL3x48+ed09jQiT95bOLSAdjY+OGdm6v
AE8GpCwN9OPw89Vl8f3fUfqHU17cwA90URp4AxTmqeBdP1FAV1nCPmr/KbREm4qqrWO5GhaFrR72
rVGHMAWkEdkxC2cmiAYL1pzWcZ/JdqTUjj8IY/WcZhAQ9AZP2dNWOSNIDKigkvvzHtFml+h7oP7j
pt0W4JIQ23OpasjhQydGfho/BzByyu7F6/TW8YElPn98SP7ZAxBZnIDTb+LCs08GNlKosqhJKivv
+qEWKbLoIjIXa1lMUeKhNIMW2H7Zu48w2YHttCxDX7shf20vTk2FDBcWFg9Y81rrvt8E/jLz1spf
cTITY6EhjnXRseH/fG3MdmWH+A6/CxkWbatmDbu58BcnfOe12ILhyR+hC0oAIf4N41TDOhx0uunT
vymUPsQcks39NVsqbGvLtQ6XONOZ6SRBGDc8zr2k8I1h1tyldbj34VAb5+TEX00o9Pc0XlOwgTlN
8uExvm6eDmd+uP/QxBHWjhRC3aIHLby+5Xa3ms5n2enKjAxFdVu3qpWWEh3sLLcW0Hu1JBs/0KtB
+iZ7OL01gaE7aObBbszu55ZzDw7BtBl2iJxJhXLGfecTitVNN9VQ4OKXkdS5zDl+VBfXJV3afjxE
6hPHAGWu95A8VfmQ89XSk9eIkznoaqOCuPz4DssC2Pdd+HwrId92CpF6E/GhWbhENNmsyrkOFolw
n4kii1ptCcM7GMLi4u6RqWDacZTDqLE7hpG74nCnUQ92Q5ecmGPtZQOUs2T1s8T3NE2V4JzyZ23a
t7N8xRHzc/DBmqT/goXTyS0bTKJtzcGbjpsL2BNavRpgzibSFC8Lo3kScUxRc7LEwxlfd2bgNy/P
orRTzvZWItdFBj7DAduX0aIJX5FNEUe8C63xyPLC0w9KkekPfZa8RXIH/I5ZEu5IocooP+ctO0Zf
UwL9mzn0+3SRo13rv9BZJgAjgC6b4q64OA+quiMIlHkqSKQdGgFULc5l9uPCZzSxObLCvuGXbJg/
O9CXG+RBGl/zWlYmbDHPqhs352E0wG5CyMZvwQ3vtxGMkt1nvLm37U7GvKgYtx09v2WG8zyzuBIO
Sq3VcaXlZl1KBlM+2RbLTV1mn9SgyW7AYX+qMPW3IiF4z/1wf7/E3MbKy9KrIY22jnF1Rfevkegn
pNNkFQ1ZXnW+H0l7CZztEN6h/gAdvSHwxLnttvHcVVsORY4J1D+lwTORqyyB4c/TL9XYaQEWfn02
UYv4EmMc99uHhzfrG/P2Kh7HUgCkWaRGFM+0rmC4PdBauL1S7mxdViNMkd6pWVGEiLrKyfDzMV/+
LpIOhJ0OwALH2GxFKRG4mvdwcILKoHX8Ehb5oCiBPVet/A9/eVbu7g9NLasdT0sBksRgfZfhCh46
9SP8nFFzNYrWjUQdbj2hHHiP+xx78e9md5+E/WHQPQraOU9gNIjC2oV/boQSZdPe7zCSaQHKT77h
Yz3T9RolhFdlzGCMvREswZzdAyhNiGEE02lLymOttN1pxRHg25DwIQ4qqFzBL7r9M+7/vAPiHMmN
6o1s9tHowQVynKuxJ33FkjgQDTgGexTIl+LtyN/QxLXbeyNYpLc5K2RlB6HrkEJkd2YS8pyCO4GX
xH1FI0C+bhjhtyRRyHrJQWvBSkAclnxTsLt+Y/3j7O+4W7LdKK6dvAOCjdY8CZJh0BBmK+psTnxu
yyWJYaFtEG1aQIG9GJI++RNu0I4dVCYnrcD06Ntzfg/zE/jzXkrWBnc6s9hCD1f1DTKqGjK/BhUD
cSPq3U9u3m3CXhFYYYdckYNLol6+0pj43Yvf8PbUQ0fQBlb3f7nI5SWIWQF9zYn6plXdiL2NEmah
n8DZrMy0DwgGRBmVchR/+4ygpVOjOr8PUcZSV+x8Ec1NxQ23HrchbMpIQFWsgmTC8mJKb3NCN/9c
9XnSa3qGbLIf1HLi3TTONrlMFWAskLCtmAu0NtEqexbzV+D6SIQEIdg7n127MstM5MHnuexn8/xc
cGF/FEDlUj7Ux4QEh+tVIdFRiPsDov7iEddS/ypfa6pALjvYEwyobSc/M3shA4X7dOGVcuQVSfbU
X2iN5yLT7oPfUps3Dvxfm4nHM98csYIA28gHwz6YeyIFz8or9VF64qVTVYPmFgnbvAb5DavYMROn
wgzYLesPymKgekB9YC24Req0Jg/owGX7F5DTBJgAcOr5MycsBJgKX8syk5xKEBM02Xj1oAs9R0dF
OAcJ0dRu2ZC6EmrcUG9pvs2LfUZDPUFD4bifQ8xGaBI2Xlks9G3F4QThtikvSp0A+GLkVkPJlP0K
vZPfaVN52MrANqKk0VPuh2BeFHl+pcVa+tnA8PD0MOL2N4zwvmsiY/j7+Di6opbHqA7wlrzm5kpq
kZ/Pq9FDgT4XrajpVdjlQ4Pn8jPyBLu98krwpE53BF8/qGVQL7/qauSPKQKp1M1jdHs7NMYBPxnO
wCy/xg61ap9jvXzIwaCkxJZDUi6OY7BozU+zcwwKgeCU7VHZCjvX0Fiv5The7gXF7F4hAgbT73ya
s7Lzto5k+PBH9iFR9tYdcRglQUrdzIik4Xf7uenCv4szizMgEeK6YY3DYC4WnaVxHws3W1nd2JkR
4NL0/DelydGzIbgu9FjdJe0B+xCVoTo+KOcnAtXfGfEB/WAK2dm0pfkYMfOM0uutSE8v71tTE/0n
FBqdQximY/BFGBpa7QDWs3cIfp2gwko63tNvZhzvfn4BMyebvDBrCgxQIdyh4lkZAfYLnc52Sfjw
7G1Jzjzw//gutmzOWCHPbLBqAcbne+0hsdBTraIIiRoKYDfky5Mktzt7/ssvip0ojMGZZoGD70mo
h24GTc7nM9q9KqiBeIc0K9HRUyJjp3TGCF3gsapC+6oHnMEQ6T2l9yjLOhPtmV/fW0cvGYnRPO5b
g13etdyy+YsApzuLJdYkOkXBVb9UANiqaalvNVGRximyhxcd34mGpFdf6ZPFgc6aGydHab9WtGuC
j56KYjfVpL23+RGXrheplwKPPv8Sd0h5JjGZeow/fPTLX4DkWTBLcJ8ygu7KI9PbQnJ+OPfiYzBb
09urk9GXim4lVX2LwGWpv9I2NHnktmcnGHdbI+wMbHKAAqEyf7EYG8T4hEg5e0CCA41d9KD5p611
C813eGOH3ghX9SBk4D3je3vpNs2CqemgNhD2Np2gVsxc5V3C/kWk5myDOtm30WOTSwgJUHKRSN7N
9iL3qA4Uk2iLNOh6l1Xk8huAkyiXgAC1hr9B8BlubiPk1d8iq3JLsqq9T6YXmIga7UC6YkEpEECb
dpNIhTEWCWwFwyFx5Pn9sNf6UDnSjy3BWwJeoJKuVaycY+0zkcjTmZPnNGAoJBk7/MFEy4qUBQoK
faNTyVGwRubtfZtDPx4fO3yxhmfm3K4Fj6Rqcpmck2/fj3DXnj4Nn1DF6fHFP9Fj8vljQHwc0V47
e8C67irUSoOKFCgGtMGJbShdrroa+P1DEc5Of2Z/1WhXsz3kTNrpz5lR6L+B1Ew+ylO9/XMwXau3
/DKwmps6GOsIXzs1a0FRdms1XI60BTY3WW5o6WKO1KC5NuJ/fgwBGmfrShvR2hwH5gdU3dt6IgV0
2TeHCf3OggWF1pqVOLePa9fdVok/z7epb5uMTsSdzrquqPidmwdELNZzqk2OcvyBkyOvHa4BOfRn
DU7Sa5NSUam2UpfQlGy4r85Hd1/PlHy42JDnchsGycFPa7rOExbiGm2/G24qbKs4DfrlldGjEutR
NTuBmDLUKUdR9hRRPmySPPdBNgj8maFYSNVXeNSfF13t+YLYxaLdfaapWdfh8876SydlZV9TsAz8
7EKieySa9Qa2NNsMLe4kuuovKzwGYoWzRw9PLyBU3bRC3gkyBZe91Fn5OJMaIVQJAgjSTD5Am6CN
RNBI4JkP2pqi1TvZaR8jC5A3Un1xFAxIZ8yXlUiIeZzSn6AHj+xqw54P61WdUyLxkRalqJ2wTbOX
maEdxfXN8B5YcjfwMnmgmVOFC0K/Qgdsn8Gc6gayp9HWZWiEwqKv51WF/zLu2kdc78b/Hq2nwlIg
z6Dja4JBOAtBC7MS8nRQ/XPOXmJOgjGeSBtVMKT44f1QHT2bZqCtDI/zsEfW8jRxce/7pPyXcBdo
9HCFJXckXWPRvM2wISDCsxyZ/Ra0HSCk+n7dL3r973F4Qh1vC925GSCJ+cExRAgzF+NzNYc/dMxi
tQn/MhbNfCqAlih3qPLj59XiAOJfzWMLYB3MI68yxykXwMFuKaMp9E5rvXxrA5LEaXgxp7l51+/g
ypeYEpMy2oAq2ijO92LxWdnpj63n1Xz3X3ckTwQv/Fgj9diyZYYSpCtwyhLMrCVCYIJeCPlPN4E6
djwt1mc6ACYh7BrFxwhCtTYfVCtgc99yNxiNxdIllEQsfCM4mE833LF7IDl1XebogzI24SzmiiGf
C2P2RWF2itrGzY9enfN92WpyUdrQxW2xfXPCXS2lBLEBOt2x33S2i1R6wJWM1HUJu/m96sm0fXgp
PaTs0czqJzoayVtJ8rKE03v3+ANjqcu/f17bTB+tutBqkUYEA1hQBdGqVw70XzbMOISAja1mBI+a
QKOLojPuP363VuMbH7BE5cszGKHN6Ebh7hFVw6MeFK7qgxBYyAn3Mi031CmRI6oStOsmUlVj0aOf
SCMPK17EqQG3RuXmvJM5cssB9q5IfoYzVzpzcBOembvbcFy7J+HZoEbxUOvFFutPv1nfTig1GfPq
7VmEB0n32uD7Xc6ZwKkN/gEvOrLIr+KPDgXysX6BcvTyDdBVVOdcbsrfF4q75g65KSfVuhSey0bg
Bdenww1r9Jx960zjjGkjfruy+lkzF41mzHl5tLfr01PzEjepeq0w5/gxKARbd9n8kqZZbP+fk721
UkNElSwMqppQIWJ16BxAap4ycI8o7QyaFlfNoBduBj+3DOlzCwcl+nKvD9G4PO+t8nDblAEqSQOP
dFXS5mUmeBN15ku4s7n5R/6mUh18NpYYWgQZs/EQVDFXeb8cv0fIL5Qom6xDj/Pbeyp1oyQjD0Bb
ogfWLL5xE9Wpiq7cXmCdbkEXdWk/Yq73kafaypxVaivqLZidvth/OBl72Ni22qTuEptEKI+Fbgp1
Qa5eZrdlYna7UDJFbDlM1sU+qz9hawzmXDCgkQ8qKuq2nYbsmzIfZfaiyvM3KlPlqiYVl5q/FNbZ
08uD/fXvb0vvo0O+8uQZxqMXZHGu7D4mDj/GmROOQYIglQfW3sYoXmZ/4IUhrOfjJBWwb68ZuLfY
j/Fh51IyRtmhYqXWFGzJsShEE6e5ddVrnGpaHgkvFlT2rB6Qw9ddkz1Zrur5ASdV8AKs1vjpoPdq
oR1vXmYy53BM7oyjvhbnqcw6+hjcqtjHhZ78H5uA15P9LpDAKQ1ZDJd1iGfIpS5g1VsfejlX2tv1
QQ80y0i/Z4CGbBhPPNE2w3preDfO5FelZawNUBpAA8F6KFSHVdqPFPBWMy9KirGNm3L1RxSdyqYa
Sgx8V1W+45mDWiAQSvRC3ooln/MWLQOFx8X7+Mm6jH4LLFldJuOihAlJZIKHNbMdmbIyMd89UqNB
v3KjAwMAKhs1OeeKvx0OAMtFCVYpT39T3Is26iXIEMW0xzgn7EqcfRA9WtKu8KyWSYqZhiZH78Gd
YnzxqDs3QklnaUFk5zpc702xdTegp4QOhu0/gvxi1q27xSW/qWhwLgt2g6Lur1iPVrp2oLFg91ci
uUgVl6UOOgn3aBc+XD4sDPNFZUq5aqamqeppxTDoTMzxeEMQZSK86roSbbhgUttQbM+OynGFCUVR
9df6vjXEYhXEEfCCsJV78VFW3phDDcIvoPWc6ltNsBQu4SN5tXjYBcPM4Il1DhpL03qFYPMX4rIf
LbcNvDbGMuiFvdfkfggUSEuzbO6uQVlGEkaRKTQeklbxgjbWxekMUUf3FNKhkMtDNosyuEjAl/xf
96IbMKXfXTYRl/U8cLmpaY2Ab7YXJbT9WQVVc23otQc0iJurDIZcsIcjuNj4mqtIT6z3AZqbyUly
aCC+NHbXBou0vrkW553ytLYSh0bTVNiyvA8jTe5lF8bYqWu1y+Hx+LiG3wspz9ShTiZRdEqZAkLS
rglbYse1wPgLP5OvTAP9pIepYDUE2cPdtiVkTGPVgqvmpO3v37UZ1H1CMmckghgpO5hO8YWdczHm
rb8jE2TvZZt6dfBBA0Yo1SLTCXKOoy6+c7o+5nDh/WC8ebJv0il0Kjoh7yxH/M/6tAeglXFVwa4n
UTFD4ksLv6b1GdYNd7tHat00OiMOH5OusvyD/1X8f2rfkwZDOdb07tipNdBoq95H3w8HKVW4rN1C
3/ineM0gfBoliiAlDufP2WJfvlLMzl1owqxTd6c9+8GW0cUF/56xBJHOe/D3jqxd++5ErHL+Hir7
7jK5badJCB5tzojpYjXSp06JvU0we5E158PxrwtO5W3vRVnTFQtTs5wNn/ZUjgCTJ1ffj/hpMzi1
emDLRdLLBh09OWXBwe/Qdtb0jYE+uBLMe6uG9puJyU/K99uSEjX6naKDFm05bCfxsGiUCL0Mw0WK
UQTS1TBFynxuTkiuJ45jw8BmKKgesmxJ5l0qyrBCeq3xJnaHCaJIDsr013k0/CMrsAmvl91mGT/6
VW6V93nON526bywOiwH87h7EIuf2Qy2vZYRfiILAEM+OnoCI5VhUkzord1KaCqkvNtjHxgQM09pj
aZB4XB82H7DbsgE4rx9R4z+28DDLNUNho+xBZ6CEmIcuUT26setG9iokOj2AAMAmPxiZUW440nXu
X05/+ta4gso7l8OKz1rbV/7q1jBym0wq8hv4bQkoVUk48573ue9qN6/ncrrzZlIlx20+cwnRg0yj
HsoOQcgmx+l/fAEsUjVB10t33ogifIfH5COg9q3EJbo/D8HIOgsJNWWMYzin25Pzln/2Q4P/OUcA
eeulR5Urr+vJfO97scwcDwWFRyqsjqcbZT3St4vFo9uRqpJ6nEzvBpF/2DqAnx+Ebyxt0pAX8G24
W4NkzNyFrZ6+EOttjhSt55Z8EQwXDLNdpZm81CI32jqNk+X9gwjsxSl1g0LIzs3+8pOHMcaownHO
MD0olub36nZFCOC7vYeYCoH2XK+QiYK0HOAo0F1ssxSARx2G6Hikdft9zaovGWqFfF8JMQAgV3oZ
7vwe+B4ThPYup2hCe410cqZSwsf1TSIKz6Z/qeckwvyVw8q2xyixF60+YESGCef+pli03PNMfr2q
DlJmVchgkw7PMNahTkBj3ziPHymuaElp6jHkapFgrMXUx7xWhzENJnHrsqDcGtUQZS1K4ghF1Od4
LZDxgJpe0sCWgDPN3+3ZN2tjBj7D8WU6Om0PkUBUXrQGslEqYSQgWWs0bHO3n7ArmB6L/u8tEp7j
OQb6lH9uyEdxq40KcbTUo5vP5c1GerzZr7IImUARwiD9hVm+sUgjfGcVDVAQ/iIsAaPc/+bq1j50
/my9NQezMYEbjDiwVZe9+de0I9a4vHxg3olw4FsO7P7F2a6dRwDgbUz7gJXogVvoAe13QoJdeaVZ
8PPsfAhaKya2PyxBkBE7a92KcAsa5vSts/1OJL7txF+6NYeZNrDSww5Zy86fIt8EvZ7vMbV6rix5
4e8BtqR0Xa6P1PiYkFfx3vjpkzPm+hD/aes9LSyvItLwbPR63ZKxbvW85O3HRDDCX3ZbpqvUFxTE
4aeAGkPPzDgYg2O7ugt+X8jIgmdfkKOgyqORkdl5y57DU4h2HvCJa1KYmT2Ak2/MhENDrENwuJcz
v5k4hLCkK9S65iEsUjXO/zo4mBjWHstQtZCzFowWALg52u/iMMQg4IlO6Fp2u7pElv9qNPYQ0RGy
69knBDB6w0VaR9iZyf5p1ocdppFS+cilojlyt50RVorsnB3z3LTEsbPfsvAda1sX/toR5/SoImK4
rHKKi50xVf8VgoGPiVh7cyGCi6EecI6vltBHecSxp4tm9JIb0vEicuY9pL1mVeY5rvdWfAjr9zVO
E/SUP9NehYddOL/3466tuIk/ebzQg0i54Ilk62OleALWX3FT6hzSkGgoRt1PAFng0Ah+9PhqELMt
8uXTMBJbUtPsfGx4fb7Z0DES/S8kgA03rv2DVR02IatWqi24gih6QxFdcmYNklR1keEiUj73ep8U
wSxVbu8wEgRzsNeOMfFGyQibXjNPJPhHZw4jzguR6xo/Gj1y8s4A3cYbJ0HvQ6XmcKr4Sf6f1Lrp
Ch5qSPHjGdLv1zYnbuI8oC1a9Tea3+SUstfx/UlYPD3YxcO9YdNMm79iZmYh8ikTksBVU7oZRmQ2
qlpSZYpdfNBcjqUjQ4qRtnwNjlkqRLCdIuzOI3I2om67W5ir43ZhjlGhcb38ncc5lLeKUPCv3gvu
okln33rUxGSTBFH3VjzkU1lFNCEg2cFTHnbtIrGy1+daPEVdZZK4qjYJv0355pDVCbcozLe/P0yW
e4jbgN9qUTTqjI8Fo1iREwc2HpDu3LEzJmqflPh3I+MqUo2DCIbVlz68J0XN0UT6mRZo1nbxHBN6
bbfOSkNlrR2t+kZJZcE+TKJ0+P66x4x6KWakPMdQHm1L+BDNoFG21v+PpD7rae65N3fpeBrlQEfZ
a/1zlT1DN2hxZjDBRywPJ6Xg2jO8o1TEMwTr2bJrekoYIZrr1HR7sOqtdBJhNaJMvcI9DwUrqWyh
x15EvlKd5m4qqw57x1Pr44FOFEZ7+tiBHy9WApq9iUegQDHi4AqjZgZZDpy3JR1d/dmi8lDlYWDX
a1a0v4b8z8mYpSMyitNx8khHf7XlF1FR4tKPqzYlXO2aeLdxrF2e8hBgKruTHVU5+qXVIcBU0XO5
NUxq43o/YJ9IHngf33GqZrckf2Arjbr6n3XDrR7GFWTMpX7v3X1YVKOcnCMK6twoHiwWAHI84wNm
1wrNAUBfLaPiV8tuolWvoBVVM50ditQZA9gNXer7+h0XIsouxS1mVLRX2SjVFa3iaHnx9iAlN85J
vJNvEBI2rpjVM3Q6ZhM93t89iniVz/4/B5DMbyo3tZNEHFgSyNLACW0cokYm40nDZu7l/4EV4xpI
13Cjiud+WOu1U50/AEwyJrdn04yWydVu3587zdnu+uU5NaZ3aJlK4NayElmjeVX1AYcCHS/10Vhi
abAPPsUEv56kFlBQBGxcF5KaBem9enmKN0m2SYJlVgg2ta6nQmPo67WUqpTPYkYhNDA/VCDZLVVK
xm8KT9k1TuNiV6FR+xh7SUwGQdHna0lGPiTX9kjR93dSxlNN3/O4KNw2Z46TsXs3alhv+5c7Kmmo
KhJCPDiPzF+c3eMqzDC+GjHcvfoGwC4Ln9A1jNuqFRO2NVDeWKQOoVvfm9pM0jgPbxyIYH0cGU5z
SvKkxjKV2ISLxtUJzsrdXWERTEeNkk7Lc4xeTRxq5A9Hqm5stk3eQmoYhYcSR5Ni8f/8RNslxnn4
g6FS/HbTrIZl7Wbgu1gPB7omEJ0W79qOl5H+JSBHTgUbIGWAu5bde0B8iDpb2QvK1tE4zo4rNZRP
LNXwW1rucshiesWR5vDbU9/6ZlgJf+osc1hsyCQ1ra/EYmuvWg6hWXDKpps7ACM+fYb62quu4gSZ
yjZ0nibaN6i9Ei3kINkjT4ZEaAZ1OL0yJScM3x3E8u5AVY/mU71h/fnQS+5r1T/WB1few8jfbg62
DOhakurdYNRf3DVs8egCQKQGFckA4PPmFnhyUmIsKNNDNHaFmjRy7dYDCCKDgZl3J1PQNjP+Xs5i
rr5jb9YFjNb34OSFT07YACZccGKnD/3i5jpwHwAysrxDvC6J8yuqRPa9nlfj5J2WJw1tGSrhsClo
SENeM1m+F0YQBqfAgnZEDFi2Ps/sIhSaDxp9PxGEzj47st7/qCle6zZSgASlGHmJMlmbp+j8p2Zx
0O9MzuWITdieA172m2mq2NjNaH0mZ5opvA6uneXkYIuxDIbHcIVmNf6uxXGeA3BYpAK7hbcFAKHi
jYQBGfyOZ6/PKAfw9rRKPvkgWfdx+Fic+YP3C68o72f2LyBxB/vjZTrMS4CjMJerpnqRHofFm7zJ
3oWadEOaQNLHrpQ/jaJPcnfUhlweWwh2TNXmPjDOPhadSs4fYgzi5c0Lodpr/SE9XIzE8dgedV7k
uQyOKoBPE8+/q8atUgWMd+LQCsZslKbxoq6eLewaUB4cFw6CdIjTTvLiHlDi56+e2wuZcOo48Z6e
pgjcNC3elHJ4RGNL17ob5REJPZq1eNMp9xlLIJFuVaAU3ogIDi3ukItSOlqJrAgSNuRBy/7wpQs6
ZfG+nCARBM1QXDsjOngz8S/IvEr2j9BbMTQkcTj+8mQJX6Q7ZDfXddvrfUItcQ2yowlk+jGagIe9
kgI8fJlT/Dq3y2ltSnnTJsmo52sRbtL/b8OTenLP0A6ZDNnJagYdfzSXG//QLgwHnDMvCNS0xpuH
bhAY/6PUYAbIwYeGHYAltxqXjxL4h52L6Ga5mTeta7h6P9Eyb4Ab86NIeq1DvhIXxgd72qVPafwB
x/DAmPXH5Uy61G+bFmCIoiGDmsS666l36FjB+kgKdg2v3m9N7V2OdunzNk80lUuaG4mF7osGQpnd
xKoaTonFb05JL/LVQ3ktbUdDcuj+8ip/vvVdg2q+UdOiC4raTi2FKReyhio7TvvnMR+AaGqh+K6u
DAA3Tc9ghXnmM5SCIY+hkzdj7t1Ezn8uEFtHDECiSz9ETYWg5CJt/OS6WBNpkZYzXyyYa1DBJF3O
lUXoNWX70fOSQ4F9DC+OgJlMX7wktC39VnSWthaYhXvKN+dWfg+lICcpfWwieFdaypZvgyCSystw
emcwo5f0MFzDZ6DuX1YY1b3YarwBH9ppgaSdINgvcmsQcMLM6v3IfLa0UzU0WGLCi+gNK6DYAMs7
9jGSphPsa1gr/oylOpN1ZTQVbl0zC/gCSMzZPQbMldh2wQavPmUr3QOFNtUloQ/KXV5XVE4YxQhy
FSQd25bjYKi+FA0uyAUuIZEuvpM4xZGfFw1dYBRoofhGCCQXJIOSGkJRGR5/kgQpJ5i0F1eh9sBn
RDlSuNMi/bQvk0dN+2cq3umi39mKb+EwdBpvu37pe5N/YwU5BapF/7lymhq4QwlnlNcLr8DvfjjP
QfdnGGBkZn1OusY0JpGRIkUlhuj+6NqwLzhTSKiYWtzRIlu0XvVTLzVDGiCnkx+1A3Omz7/0kNZF
FtDce3GWCrfQn1noKRwKKVgD8Ia1yPS17vAJt6CJxlfRxnyLUD9qYBmD1pkg1VJ1msiATkCb3stE
U1kcK5FYOqlah4RxU6j90ehPGzAncfJG2i5iJwImE+FP9tzdvszqoB7HFonyDPCMv29CmjRt6pLd
1ANRhTiS56IdIDbaaJrGcAy048EdMDZ1wTHN1IrlseitZGK1bQg8XSLPBN5x91hESDuDlEIaWzt0
I0YHkfJb+HeW6G7f2aZwM5gh9+Ua6IZ2g0z1V3srN5SjEkOMczv+AK785swnqhSjGww2LpSRNHJP
U5P+MJua9YrXMLlki6sFjK4powzvxRpTIhxsobu34tvTaU3d+U2DpSzLoSVu6HG2OWslHvTSzd4M
JgXs7yfX/s3m1tOgZJhZp+qZyoElYlsEWxSIZpypcr5ij3MZy3Yqxuumlc3CPm2Jv6ADhU0Fm0BQ
P2JDSV0uU1JNjgbUcpniglq+B9aOJKvdQLzA47w2CxKkmMghfLI+cV2w0Aj6uZWor9CfKjM9atsg
h1U4UntMMMN4nFPw0hYAfGIPXMbZA3C6gqtvTFs94fr+Spi+5r4WE0M7T6msiGpaUQCgGd5IsFhU
M697gxo2cqttBkxrHVZme7O/3eJvzzUpAPFytiP67124b72Eqt8M9fQf1/NSIvgfIehskbv5JWsM
pTYYeXQjKYopGTTTNMLBIxGg0CdmI/DKhbiN5UXs2huuOFizlQZRgIyV3l+Y9pHvdpjpDFmjm5ba
gAWjn7ptYf5jlUoZPWLn2g5uOVGVNomOtrnECyveqsx7e0M8seSRoz5rSdKJeJsZu5333rQy79B3
WcqirUUPvRs4z9gVDsOP1HAF+rU6IaROVEAXkO6R24PUXGx1KxOxzp9cdFqjfUnxlSFo5G2d5WFM
qAmNl2aFIRBTZcQCgGmCZj3hHwx+sfNc4ua9BvyMdkRxxqvuOx6OYxCaUFlNaOIb7p6zgYXhVSdI
DCTkm4APPJ1eiXhzZHnk2NlGGAYSl5sbrNR6DPMVY4uOmgdPVaTHpKEd/Faqui7cN1l0cwC2Styq
yS3b8kmaeNv/DVEC7okiqrCO+SNVpwGEKXkpnEUTGuNK+5FJ3FivYLE5j3d+HTvjmnRFVHarKp7D
w5RqO9nAKOsKkGnnidUbb1nYfuOv9IpKnGR+Msope8QVaeSCahPFAG+mNZ5mxLWeq0FtgiOJxr6k
dJXKcoNAxwAhsMmoetmyhv1ui3PomkrHkLS6JVtMVczE7KbZEFFhmHvBWwSU7TItnAHi07J561ig
LDZhReFzaNwRhBlVeQjOYu0MRgx+w1QMeyWCyRPAxNciKKCiJ3JAAeFXxB7XqitH1kE8Fyjxjwd+
tWnN82W3CuByb2iGoKf0xcLviORUfZGByj0F7Fw3M7m9DeWIOATDOoB5irFIfTL15nNgjArvH7nY
VbLzR5to/uZAQPFOq3wU8T0OO5w/gvCJmsHT83w5NZq78MSRM1phkxhZ/DSRPGj88Ax99TQWlC2t
r/cQuYBTGRX/mQj07GrjWWAo/kE/E/yxpdXzDroMhEqD4VKXXdnSL1S2zKdK+Ucjiq+07bDqvTEo
JacnfB6bRnZQxAazd0/Do5UdPzJj4ZvGOwq3U2CtbvWjgdJq3bpBy1vVKPyD8ik4gzrbtYmUuWmw
DFN/tNlbQp08qa/9e0sVRqFtC6AdM1w2RIGspHPRDO4nsiWQ8AH02rNWsw7109FohsWg3cwOkenx
+YVktNCUKjnV/81l5RLFhITT3Hf1HNrjZBnwQQsiUiUlXzorNrTg4u+1ctyMW5o/v5HB+IKoXfE6
3wdd48lrIY6x6byDHeapcWUteJBmyms//LHnwacsc0IrfkRC1KPHwc1fikbn60pMoxrYITrpHylB
DZu5NvuPoCBYEFVGQ/oux+Y3QAzlVORot/Wg6BJt/E+v1dV+vo8KaMMhx3/Q7nY7zYHtHwTObKBX
FysQmv71clN7d6bFPY9AgTrLaCRnRyM9duKS/ofOLqm4RJdXqX4R/yr0MBc7IGteCFup9UNjqBDi
4FtJ2OsOS3uJyQASkfex3JfTQVACLHMuIOJWPjxjl1eQrKGC8NeQHvPgm97awqSVuZCoQoyTHRb3
1tprQztUS0bY06jr/BCCHUEmgQosDH753pMc4glDc/VgaXZQgIKuwzIIjp1Oag1iJ+FVshg/ZuR7
c2ybItXAMU4DavikNCwzsM5Tk3QOqjWEjRgbRfltumXYwHFRAn9NtjxsajSOTPga2zRxUMXOdNOX
0SR9FaTz+AEpVzE7tWP5/GkcD9MjbreuynRMlQBInTNxaNneeQO+qj8ew68zCX891phBvinOfkdx
tbpzusoK5myVLWCbRLe+RV43jJsxrEaWWvWxfM2LOlUNyQHTksBiR1pNiV+aTnd4nyozT8AYX36E
oECdF1HlShjkTiJUPc7A4crg5K5UFSfDwwfYz/39oLn0ZMroWr4U5PudH2P9Kl1Ca17NVfO7JIuS
cSeUhq+vDLjDErBW8jspvw3K0ECl1pc1r9Uh5vSGxGxEXxIVbaT2dC0yCRsVdWsN37Fpk+WL3g1X
fmuFRIPTAmQ5rYOdIaB03ziuP6/lBqUYXsULSRBMKB+jotxkMea6xhzR1r6P191dvHZzBCgtEnyH
JBWfKDm6mcN2obr2rPCIm8wGrwSynu/2B3pBgVSBlDKwBELxKklVzcm7pFz6HOtHyFPhQe3JzR2W
D3sHBahfvUqhOLQabMdzFeX2nZf9BgrfFeIjLcKSAwpHEMak07A4LWhAP+tTqavIopZuwFlYvjyB
rXhQ6Pf8XN4pk5xxqsjtqO9XKyJ687Kmt5raJ6jZ9Ombt+XoTNKiRqYhSxA69zH3mPpnavpTd6Jd
CCLuMnioKq/7aD49WtaBnbLqXetmNVlIceaDFsVR2/c7hDZ6leq6IIlAP9q/PfYKkowvCNnf68cj
WsoX9F5Bqm/6gM1apnJKX53OaHHGHqp+pBBngT+EgWch3JVNnuUBLGCDv5SWdKTpPb1HPHbJCHXZ
FrL8VlE1K4iwgQaU/NuEz6f66We6Tgn3ZxEyzKIzYLWqD3tPcySXQrAeUg+3B3cupwUFJt+Y1zvl
vPNYawlXpuhmwMJWkJIDELiWGmOD2BQzb4hTo3fOYUx6mv57SHQL5Uq3rFS7iQPzGjzYeCuGsb0w
0fWFez0Y5QA6c4fWtHxmCvNvoI8bmMXJZUV27m09GmZxT7vKDfIXakyUYOCPf9T7eQDp0GXqIBoN
IQiCcFwFngWbatL8kosC5WaUJfgK1yOlECxzYEZxG6GC1oYG9hCEVfUaMvrRHMwUQLI477VkGbXG
2g/BvIA8kqsVAEd2vkCdHPq1UXnxVND4hoLlNN+5ouhWQXwTahdrrWFom640nmfkLesfFh0jCURv
wqi4t9i0V2eIGc/w48aqXCgebOFUzfjQDKu+OIhu+ePcUfRJgoat0J389TrBBt9Ax6yyDrS756OP
lpdolJS6Jggkuu8VcnJyQ4XfOywwwQNFWhL0V87rCEELtSLdV9FIeHnBkyK4MUK//jf+rGH/TRGp
Qpf9M5DBsdsEMK/2ZdRpCjbi65Rhy0JzJNE9cU+wcGQ+BGaCXSfKDgOdYdfPl4UwbX7XnwYvXt3R
DPYpIXAOgLwA7wbM3Kj/trrAWanlNubJLbp8v4Plt56bvWB8fcjVPcSdvf5mJXI9uM1eJ3OArHpk
CsbitRXCwLM/WXdSMfF3jojEl/BACx9E0uajwB/mBNDNloxuo3yHXsgcV+5E8Tse8XIJvDotX73t
uVV9iTLj/U79RCYKS2qUwZgyDsVkETiyUTzu/nHZz3fZov/AFDSbTHdtGLSWxnZyIdQPzOzH333N
PKHI90N+31XOILVVrxQex72fXclUSxzA14Kdz7J5dFZjZQVRoFk5aizcrnut94mxq8zi0icZJQPn
m9VKqTXmljWw4gjQjP3EO94ioViFBMpTxGHNqUm6se7o99VUv9EdwgPoQpUh3LREZ6Z5X0EJnR4f
ES+DZXxB/zIQR6+e3LKL5ee7lyP8zEfTXIgJCaSvL869cWBGnjQLMC/ydL8osbhgN00DLRrt6/xw
sS+4S+KtMk0KgWjTp7ipx36IK0jMP9n0cLWgcZYNtAnlz0OSjmMfItlNciqg0jM7JcyvctA850dl
1FnM7UwJV6QsFzmjuAFSSX6sNlCEF40bxqwWel6IivhVMl4GDA5F7O8aOjQZNxXC73gSIzMT9hzg
gmF9X3HPWdz82ItMRxZZ5gOIsmXOa/T73s9s0K0606WxjSmp0fj1XziTy3L8mhZDqjcBUdIMdeEL
5zgQrj4pQhXrU1AL80W0RCm7pCvyj6AxIkpGmT38JGpiY720xRUETo6AC+H997ErGwg/FsNxfaHZ
Q9/0UrEI3sN510waka/G7VV4Ga3Dn8XPqYk/5bLyJyqHpcDOJhFUsIMr4PgBKK7yS7tcwsnF0AJa
X9AZYYbgrNvIVYnYZ/7Z9OwKbDnSUhLeqjQ00KO3w9XPsP7PlUOw606j/JIXSZvlyJZFj8XZrlfY
Rf9ZgCQucAcvy9rzsAHPtphdpsK4aau+o4+ATSWJD+oYgWGwlCkdm26/JKzJWwt7GyOAYtbvPi+L
dzjYkOa5oEHhyl9cyLkOoeRn8Ds8u9TrEPhz6uGTnJO84Ljfg0iw24qaBS0PLhppSff4wixBfEQH
keZM6u87KTJERq4mFRglBmBWFMCeEctXJkWI2tS3Z+3WEi7yzUgvcSmHq5WFW1uwq6PQNgz5NpEx
W1HPLNMPmqPyylNpetSbbmLWPK68nqbIXtefTwpNLkW81CC7o5GopaDnxcWd3Ql0MHzo4LWtEn31
931gvFq0mogS00WbbSH4mWavGJoGLiqLw7MGHTPj0kspvTFxUzFMERer1lSx1fY7FsFkGFWhXVHn
BYP3aMJMZ4F0/fMVQO8uyrBVl/BCKIfcIRhFYFyzzrxW0oyhLecsIyvkuIfdaoK+NzjNo8nUYFic
KUoP2vMBbGV1aK0cugSeNit/hUgfJa0WtSTC2oy96QnT+iXfOrtThR3ahaRAlghijbA+t1fzorpr
4BNGgIQKk8bAfPyRtEOpNGWSgzh6FHvRzeG9esH78P7HyXaWiYkT9pviINfYqnZx+9KatOZjwyOZ
zvvLZ6Z0aFPdlghaTpQM0Ou9egcQYusHIkirwMqtmA2lGVCI60ONjhAH6HWGWWfpCRWIESOUBa1i
MUsoDHaulojjKZZIOv6GG6RutqPUbEEPUL4wJYZoPn3FRJZLtQkB/Njsak+tR+ssXGvlqnY6wfZE
/7QJWDSYTuLrh3whCJvJ6Xw8qSSYO3/T5IJT66USk/ycrlMCxoVu8mZEdGIp5n8L9YGA8aZuUqMl
CAv+g2h9gVq7XYTLUDfPYWCj8cTKj/dc49rK4qdl+TgIbNUuZE9CRfnK+Cq/xJPss543BCgZMsuk
Nm0IiOtsjRNqREKvFHW8y1FhqIsJUNLhCN42lGBwqXuJuuC5xOnzfjxivX2bbydLp0gEn9qA+igK
x3nq6r5NzmSOU/n1PSN4XAVAvsWqyAAhMLui6KxR94LSpi8aK9sy8HAPW/pudK5puCI4LarcGpW4
WeaN9hPQ5578A757/5hFMUoEq9cZ8WFF5Qwp3u9jKElwRK6kvXJ06f5HXoogAF/fPycEkDa7osFN
bMQ3FPpPq7IBM1gsInPMMID4C9ywrlkRceycSiO8/QM8zTwmdWbzTV8ZMF0Mqt2X8GwOF/psMFib
YGc4SB7ncK1LOV1s5arOjVYahAybv4mxetLBIK2l35CyJIGFUmESqTiCLFko6/BgO5NdNAH3hJ0P
Sm7Cz13UvI1pFpEoLSdNWPHf1FxbhhNi6uRwslSBuhaIhKzAoDXF4Zyz3velBTfe1naxgrOpKAB3
l+cCKhuZIQxJFgId5hX2QWxVP538ZtEOjmNePRSHNdGMcCON01DhGwqQbhL7WIeqSMGPZAOn0HDT
2MOMgwBseI30DCoZOV6X060aDADG3G49r5+7q6mpqXzBsJkd4Qt1xHPtZVs5FJx6PmIjpEjOX6ph
TXUyyK2maK1O0RWIEQu3TtQulubYg1lUmZLwrN4b0El85irMvriIHq9RSd36YCyEyyc+6QQvOQYn
oma/Vp1olx0XhxCMTjzHHozK1kmk3uPY3hYnR5VnYzMMZoY7KO7BL/EMutTGEXGrCPaU+4upDcyP
IVzhbpfnUEWeWwCSEVPly/B1NxlTieV4MPgrrRUXCAQLmBuYmbDZVCNRQgpLkzqiGCRU5rvpz+eX
QFlB1tC0LRKzwioQxyLkaYsqH5Rmsw261eo7cq/XKYHn0wfNyCLguHvzm8S/ThKFOgkKkUo25kvv
/nbAd+UzNyACFSL3n3DVw0raHdddTVSUrqsAXGsnC9FWIFHlzF+BgdeXp08nC2bmlBPqTar++VTC
Hsi4zfcp9j9OiHToqz1opxDkFBC+UKe8LuV4mWbUuColx9U/kpJiZ96ZZu8VlzhR36GMIzT6kCAW
zKMqeMs8O+XLwYqWTS9cCYmCi/eaFxi8C4aYQWcR15zj2/4Uqu5dAtpWoHY0+ZGoC21ibkyQNVgm
k6/FYpoIUf2EmczHqy0QcUgRBM5l16EY36bnq54cLeuZSBBAVCLHZsQPgAJKUteo1j3GdoHn3Wrt
qrUjlVlV0Ph8cB8VZ2dok6V/sxTNFejKlDxb1scWst19IfFnILrSaRmLrMB+fhjiEnCsgLIQYQR6
2uM4Hv2cEhOMfcQobKm4cddrm1kZL39kXJtWjg5RFve+8VLlCJ3aqQI0VWVo251UeSjuji8nKzvs
9ohDKdRfua1PQjlKOc2FdHLoyvL0SgvgzpY6fEtrR7LT6OtswF/ZSCF1SOizDjgeooyRbHoxdV+3
WX5G7gRjXgKbvbGC/v3ZT4AmXsF8KUR3FUgQtpU1DY0U8U/0HYzh+l/EdgV153eZ6GhuuIh3dpWp
gsIYK7EcNSKQALzbB4NRGWpeSsHA2FapRakRqg1DuCRSEf4boKyslj17fBHXO9kMTV5hAxDcZtJz
Pv4DMzlLvH1ZxPEBwV4G4mAkxTq+u8JpDRFO2eL3JYxXRnsCIiEXasp78brXVCofyxdzwkzWGQ/A
DXx9Q6zvj5wtF7lqqAUG8l2QkVAiHtRlHzHMY5tT8vKA2bnhzuvYc2OrCMcNEw1EqTq0SGprq5SO
Zw7k1WgcG6dLctwO/xdf205wIjBkh4gekabDD1GIUl9jP+f/MeEu2wM3CLQTVORF4hxj3sSgRxNY
AFeqJkNFGx8rlqc+3b8EXFJzGp8Orwoz8o+HLWEX6+lPiba2F/QS6GOKcXNsO6+3tfe01hfnllNI
o65ctWBhDIW03wj2ZEwdR6grYgw9u+K/d/ZsrmF9oVVOFarCO+UKuBX9MbJmWag0jRR7Vim9YB1j
2spfZbAHqGfmIj+H+QwUYGNL8B5/PnRzODn1ioOz/tGay/2PpLkDGCCt302Ar2M5gRhV8CNYxpAs
sIumCfsQyNyWa5aq7AB5htKKZzUeqDeWlA5k7+E0Aj9Qmz6m3BvqNfoNMVuhf63YBY6VNhKtp3C6
0+rza9Qdl0VitzokyeS1Yn8nlf+L8yUDbwkfOCEm89yq19RZnL5PKiNddhKeny/msB9Q/2u85hcL
ArD2scFIYwXyN3aBzjfPF6WB7Z2FAGO1T0dRn0eUFTQIwl/akzLYzB54S1SwHV4lQYT2n7d/0M0K
rXYD6xIvFOWRyKG6U4W6qsM6ZkMOqMNYeAyUFj14obG7h7y3FvuoYNyA6wxuKCtNhzzxMBg6Owi0
iM0Aow7IZ8a526y4EHbZ/ztIlNqKp5sBQfM396H5IgdgyoplU+0spbrhDhpbJGD/W4ikStpSisOV
4R98H7H0Ok+N2OpTgDZb6en+fonIEf0Q9uryLE8/PUI3wg4hiskipSELcNVzXeo5JvKx4Y4/LTVD
wtDaKvIWcfVELTaWTA++sWUUEm7VxQR/SgS73tLESQIbw7LvgWTtdTFB2KDDNbBOkiYrNP8iXqKI
YEx7/FjltWvb9nFzgZJh7yeoFYjpUfJXtHG9zkwPqTOqBlBjVnCzFwJnJs6/0Xk94fJyzrTWZOcG
REHlke2vzC5XGoooa0k8UZ5Q6q4+2yJIburdGG0VrabGXeC+AQ16yomHsraNNVEfTloavNJt2qO9
sQsOhQ8Peyy71936Rz4FqcOOcITVz6pZ3PitjwuEWrFp21ls/W8XShaRN99hoT8kp72pDsJPok+I
k6ZzOir9Qu/tfTiIqxl51QDedfP0pDk0SrvmvfOe/7BIAB6ZSABx5S1SkRhwdbXmWumAUQgx8q2L
4CNQiwlYyb1YsG6MRAtKQoVA+Ak0Bj8l4JZ+JSjQ/hfQs43RJ7XVH5KBZ5qgTKt37Qj2j1BxZwa3
EvIdraYPccA2vvJgfDkFe/Ydp0c40i1NZ9zujIJu+z4sWqRKXvlcUWQNrxGJnMUdy1YgPaoGZsY9
wnizxcryfYeudfgJxRKL8mvUUXp8nkjP5T3lgv5lazviGZg+4q+dUCnZVZr5JJKOa9XZFqbTgXUL
dS5HfCy5r1KwJNYJmWIHtngGJZdxfJFMWx3uVY3FIooZ5kAuup7U6cdXhlJG7KCegnHFLTpDQ2jM
Vm7OaqWGsWlyPYPIn4zdpQ+8TyoiBkUudE+T7Adr+yWfByXYOWzmcLBJtYvZEXPII1yAbJz90LJ1
2OlZK9yvO2TFE++x/EyY/eV3syfsfzaIEY6ztw4OFG1i3Uha0I6JS7IShzAIMZ82iadngCxNJKnr
fG6wfjUg7IEei/Zk9MXkfIdeJxp6r+XQ4y+YfscYDJDquWLyp4NYxG0CAwMWs8q87BQjtHhAnHvu
XZ0VBZf01xuJb1eaLx+8QtSAC5t2NpojlAGNbxa7lLQdyWNUzTrHJEpJgxr1u/QCb7L9LxWWO7ZE
X5C5cwIgQ3D4v+7crq5FNdgTFlYClraUF4OfK2LGi91RF25hjsdNnBGJJYXECdT/wJlqe8lmepr2
yHCphXGBFAXKEv4xrX8owgwqgaydyFMuK9rvTSw6GZ9zSMCqqFPr/U5uQx4qJlnPrptH6I1DRn4l
vaT8c/UEFALjec79aunYrQXV68A7kaE4tQhANrN3WfsQJwHjLMFcD4xu2nI8S0jqJNb9qPqO26Xi
ajHdCDSIZNWXaYBNb3vE1/YjmcDm4Hu9CWVMkzhtvk5yCA63VRX3Z0SQYIgyYkgez82x5h8AuhTK
VjkF47JeFL0XBMLOuMzCd8Cy5MLWFaZNVi1OLxZPx1wDLyBMYxrVQOdlFIrtNmx7wh/kRdtvSooS
Laf8ukBnyGX95uki7wBGjYPKDbI2sNuw0K2GXvdTEXT95ChMvDiS0NLlEI3Yc/P2u789/ugTPRGy
Hha96R3r5D2f34k/iuAm4BaK8ZF90qtfmdb1HzABjzuJbn7k2zi2DRlZq7AGqv9XQJ+0XejT3FnY
3qJJF98niB8GAR+c8VoaWT8x+ze7NJrwMyq+AS3tUA3AcYQ1FCOHORiQQMwDsJvE4DDDOcVsvFX6
LLI6xzunzqSrQjq2jbJYrqMPeAK/GYhUQ76f31ExNmSga/5RHw4hZLWjd6Zg5BX/qUdtQyA6/zPN
Gmws0f3j0qyimPdtYiH6yMozogOxrHI8+rgrzPfKGNXsrrN2jLBK8d6to58chek0F2NbaKcljL27
zpIzjAK4cQG8UdME/4MSrRKUvJwpaHu7ZP0z5iI0j2FSTM0LBxl6P5iclo1McUu2t3orOPhvsxqr
HM0D20T3ZT0ldnJIPrBfGm3GxO+ElNXQVBjvvIV2BuQBotS6dj36g3xb3fwR7J08Vv3Nu3LavPRv
qWRFtfZ1ZGD/BqZi2G8HroGNLNsDh3wApPiaFgzoKFp6ENWBE71XvLG2LAAcW/wYlU6MY0J1aiTa
pdBQjTz/IoTR78oa0ExYONtF9KBIg3MYnuc8gTAvQLqzpGN3pQRBhu4uW0WOGoOdm2AW3Xx1Rpeg
uzPMMA0aRCvNkqEAEsE9GooRH7Ude7IAr+kyZTsmBJcUKnoIIUcCauBH6KbYrB0zD73C0vc7xFbN
2wY4oDjRvwT7WZT8EhqG7jrWQtuOpH4U6gzuV1CK3X9cUAXxZ5ZHZZOeAoRopy4NFS0HBmAb9nV6
hYIybT6wmqZDY7sQodSmyofQZgPvOuLPColqtyLx7BKKaB0Y6+E8aXeOvPMq3Iq5InPhCPlwuBRY
Xhp9dVEKDd7XuByaQ0MjmpU/ZowKzIzVEwALeD8iUYMdTQeK3BLSM0AKoXDTIjH1wws+J7f0ToXi
Wvr1RRtawsSbbpt55sv8TS4ctFR+1hVTmAnKbz8gW8Y84woEmBpKKqJ7T/xP7eAYMdn7tuzLri+4
NhZjQKOGxvNn05jPZGbvL0+i4KiObatO9UMSFaf3O3+d8j0OlSOX83ixQaLKs0Iv9YfR10jvGac2
K62Gf1XECER8M8l2jU5KsaJtwqQYifwfA0c2aVqS9fjK6mAyKgdzofMogCwOwMKWyq85fTmHREx/
JNYF5qBgvBy/SU7SvCMi+GCaZC/Jcx8xWpmWl/89nZs+184HvypXvxBq4X+HGCb8V2sTKFRP31JF
OlbJ4MwJJUoRQcGVdIVkIBl2m8809s7HFNb4h9tGcOpq3BVDYbfeEwaDQQZlNsFJUiBe7YQGTm/P
z6scpd4vxwinyLOnSxb/tfMWqa4X0qmw36FzpcUN2rv5eO/uGec5rEZTxtz0loDOE5fIMksnDLB8
Sket7UBaftDMl7PwIRnblC8hbIOd7oC2zcVkQtGGURBjdR+LNaJFwo+2aEl2dz7Obz9i2dgEFi9l
+9OJZZUtFim7WhUYpRRsO2qiUA1PqX4vQ06Bjps7BL04a3j5mPY9Tpb89NL1dNt6mus61FNY+XEL
sq7BvcZ+6LSgFSEV0HtBuLcPrCnJ3MDH/Qx23pCngp9AC6PXYO/rCa5xukqQ1G2pUBV4rD23CTVh
rKtyi0kKiVEAqQVIIg3b9Ig4Zam/ubZjw4IdrZq1sxN7Q8iFDu+/66F3pids4SUtSe2psaTN6Gdf
juEQ0sscGiy2oaBM87L5eMaFG5V3x8CrtihqnFwy7oYXYM6ud92tyMVxzgGKQN85oMVuh7pbtU9o
r13q4RUuEIuFnnDQk2K5+DOh2Yn1wUxOyi+RCVy2Epvu4R5bX+xdhJhqk4Ws3Nd+rXnCpATbk9Wm
c7TlKguaY8Sw3q4yJR8X4461x5vI06Jt56lFJloLXoCdOcthomcC7ja4VtCg8+NEiQE3/zlxYPLM
9IADbV8ecsxVr4oHdkheqN0/wHq3s4PlvZ3OpF4ytXy03UDUt3fnwW+VGf3vf4C0uYZkEeowTvJc
0tk7UdtpUchgJ7n+rjnyHMzI6K1bK8kDszUO9P/mLSB4Vp0kWIzlRp42UGj4dxOa2McSeeGYQtim
HoBTQqwsRuvOc1ODMRqhb44kxXeDGQZe/ZfxRcdgeFT16jsMt/rMMDwqzbb0/VwdsdzwomMa3ZEq
iZlctqcwNDeD6lQyxe5YKujqMZ3L9rcT7pEcTGPDkSQ6wz76EgIfoNIUTdiEHQoLkoAX/bc7iHMB
T6G9JFT84eoiU/8cUG5lRUkQAkJUZ+i4ncJg+hCdg/HZGX6fzKSmDnievOI5wp6u2zx0bhD08sbi
zV2DCO4rem6E1u233tYT19Nu7OYFFLi389qThiLMm+Nwray9NMKmA6heh5FglQrwdOtCuFty/fmA
g5vnXAoQdN/NXaf4iDtTIyTyyC0HX334C7kCTIgELb/78kmou7244QWO/TOvmcQOgNp2GYgAZwXL
7Iogk71Ai9ip+4f3ibhyIjzXBMpYagE1U4PtqkdXTeEuG1Q0Vh0SRZdycCjdiEvtSe48evpleGUm
tMp1lLGvaqLR0nw6tivIdNLHgqJiSLf1Zp3Rr0oTJSyjwd7APeMwix2ZkJYJl/JY3gp9LvI+2tG0
0++P+wVGhNf+rctxFbgyrHv6RZMWiLKshp3lDskHUWGX3WjhdkmcAnlkUV3WSfzl9R57uVy0QmGq
2ufwzHVl2DcT8tZb0R2Wov+20/k9HRg6dpKYGwarb2XluQkv+l1XJtXOU3owHEem2VVsHfI0dXQT
iVFdpyHO8lCZoSjoJGoJKver2LvdxrwkErZFPzVkr2VqMmqnZWuj/MvFjiE1zQ5XlSs/v87NNgsw
6gESS0TT7cG2AAVpr0O4xS4l/uPFbywUG3xN6hO3HKI2qRsYuOJ6MDYkRQslaGEl53NJkWjLcZJw
fWMnkMsrdgHNG5XeNnHexfGrJr5yR6f3kuzSQg97vnpfJCKFCQflqTLv0v44l33f8Zkz/YU4Yth5
uML9S9LLgM/hd/LorNObeX1eHaYWKgo819LE0jtreuw78b3elFEwT3qXG18ez994Dn72kuIF3thU
JHqS7OLp87VcEyzRwJrXvueQxq8uZ1VF6baJ+INT581P8eUe3NdjQryTT8jKUTJal1Qanw06D7n5
SheW9swezefwEFxLBGwydnZac/G15u8ct74NPYpvbTBNWuj3G4+hnvVysec2JiSQgU0AryLjC2xw
kkb3pbEW4iQVvMdBXqW5A5MpKI7igYGPVfLNdCfbMNIQGGIEcf/F7yCcqY/8HZZO8CiJ3+RqO+i/
13Q+0n+sjKiNZi0Rpe4uVXg9Ei+I0agScf4ZyKpQ4VJx2+RRKjqDmodqEdjrV01IRsafO1RLMEpR
7vUZ28OS8iM0rF+Vn/1Pg6R/+NluUDkXcSxeHghxaDTPBzbGD3Y/eMhopcJx0ybEKyaWb+cVHZV8
XtXnubFs1NadZKOWgAHwIourS9O2hfWTKMS/osfrl40po6rQ1uI7y6LFMJJ8n8N/8FifKRzoqhjq
vb1tkh5UJ+hsVf6AS3bG/bzQLaG9nuZpFfSBmw/SFcEH0SjCcX5ZpkOC02z6KlbxYLK3TdztNIMu
4g7Y1ORK80qJqTuq0ID9jPHf9TXDQAAYmgVvUwY7Ql7pbkj5ZAvD2ZqFqEakaYqSdvNRLlXukII/
shmeKG6DUfGf0XnyCBeCZOKrdNn2JALjHQA6Tei86fiYxO80qqbLV7EAhqxxsYUxNV8Ztu6LzvUs
rFt4JL2C5OxshRfaXbAOtcm6qnGYFsLMOrvi5DhQfLmTX+kCq7aPS8GkUoRwps38IW10RKzMmtTy
z5+P9EAMA0Dlrx6rUD4Cu3HbpkYV86kLVjO0B2p4j4LPxVnCFFYY/H7K+TiFF5m4zqpnpHoWpkTU
R9FJBmAE6d+bvru1hGDekUGouqjy7Hp1oEDPHMlp9oeSUSZQavlHsMHVz7n260g/4s6VkgAvfZt3
rYkn6kyh+YMxZUoGhgC3dInN0zyoCVr+y9knBeBTiByfWppdNAZMAttMfswum9vm6lqYmbao8EBx
6upqNOERVM/4lypERbvC9DfrEHKvyo5SnnLU7qydRo9H7UZjbd7R17AR/L9U3zf1rr/GmuF2Y++v
isevOWPNwdGVhqpfxUbg5XaT5X9fbkVvmWvW19V4mX97r8n7CFGVsVRnvxPj8YvIywqqx1GoCeJz
wKrB/RJIuL6g5lLCzTmCE7k9GaKUVVC1Kh/ha2BNBsavSBYP7Lxvm0gz2wFmPKmlgRc1huFkNECr
f5+h76cdl59VxVhX2hQvb/581a4eUMzuuAYMURujYwImFumzFtBXiOrF6j/xgYplI99UbSsIOD19
YM8MGNpMOOpNElB3yqE0pHsGOSqf0bTS7oEOD2dpG+zIo1OLHQ7KF0c95qnErBFznhdCdyaiZh2c
dEXpkT0+IBFOR7sZoR8vM+ubw9uFxhDTmrMtJc+0k2Hcehjq+Tj4GtzVA2zAyQiXe9TqA2z9SSYF
GMDj0sjTB55gpS+uCGFD5q1lGLahaY72Z0MeWA1bBZCW/JXMicC/3oWPUSE/XU8r/4lwJf9r5dK2
K9cpk2yXAPMCqHKbjypZJr0fb3Zq97ppS0GEqARHAYx/MKH9OvbMh3jRAeJ+Te5u6u6rsSZ4SDI7
sQ/uCfPPmtwBZP0/ihtAjKzWLJx3GObCUUGsbvV+buM68zQHpGhWuDwqSsO+QqpZelXT4RWqT7X0
Us6Ggn+KYVsSyYQTRwcP8OoN2h6ofFGGB0zc/XdXnhw4tnxlSwwfWVWsE4aDeZZ0uphpuoU6LFWW
qmOHxkkCpmxmxze5V327zKgT3cP78FsJ4Q2GFlMoJ65yjbOEcryESA4QYCfyhcAmw1oUx/Jy9tyb
jZLYm7AK7mp9tMjzSai4yF/kt8/YMIwum0BWgtZhSdOeJeM56t78UHZWskSrHKhGue+nuVmDnaYX
My4/mY/OoWYbVPZceE+8YP6bUJw4nX9gXDmQUJfOXDatAIuA6lOkLooyB5wQQHA5qTQjU7uvGf+o
BLZBcn/i+W9kEJS9sUWUB0TTC1VGaf3iHl4j2THvEJFSR8opjttQn+OUCY/Vda7nB3F+2NXHYGWD
enpnOM18mFgd27rq1m52D4TpJ5clPgBN1qzDhKAJ+CYA4MjTxigEql3Uczv39BRlk+/RKtXI7AsG
4tjYMv0DfzOtNcsBkvTs1C0IlY9gRQ6wXMkCP/23OwOOzP6Ar4HTJHfS4Bckgq1o6J81fUX/wsYB
5kPUQQH9OzjCPrwqpId8TR4m01egiyYFFVUfo6nDJmjvl/mCNTyJBVeLCxIEn+LRilST/tKj8glk
VcrtErLNVYcyMZ2pyOez4xUDjTOPG1k1mRTBN47fQDsJKczInLy+ZbFlM3J2p+WVe6olX6OjT2su
ubiD+Wzdhu+hRZnyn/YnbNpFl0sjnr3x+KI4CtIWyfHkCocVMG99k+EPSX9XGhXGLTDSIfXG0nFi
bFP7/BHWhlVe0FUZbkj02Kgs+1sZq4dTBIcS9h8FIjY3Hn5y/ES/mMqez5fFcV6UOom6NT+jaIdZ
6kVjI/j6Er7uaS55CMxg1Cyy5jeZbnq40RCo0aMJw7BAxy2/iAOu/leNto0Qx/TZCETKj0QI/waa
sAitcy1G9QkqwHPOy6XMRfQH1urNgMZjewDVYZMNGSkm/4SH2TGUCZWWiIOCD0sYfBVRTT3DOTDU
pKpKe3fBit5G0Oj0oh0HbBVQYPpwyQMP2DgJ00LN+QUlF4SwqRY6kcB9AQMfTGWT2Vmp2MHhxtTI
3Mb3Tqz+bSI2SKaHQ7UAug0i/XFawbELtkpjF8t4Nx9pYuo3YMnzkZ0sTIuMMUKWi/bnj133dFf7
apkz7QD3UcbA7cXQT4nVrjOMBFRd6Wn74lyLDWUnx92vLPh1Scwcg4S6ykyGAatPyKb2+S/JY7SA
jxyXXW7z+IKDUdOiaLu49Kwb/mHARO/fJwbBhiBI7f5y57wEgV1zzLrTqD6gpotSvCd89XM+aVUo
c9ikN3ukiuRuiB9040hyRmkAWaO9lA1bRoL18Hp4AMDAmRsgBJvdBZUEQVaovmXPWa5U0EMEMT/j
Ariti4eTcQcu4KaaJEMoJm1OJ2/8FzeTzXZqx0VM54HrA3uV1G/6LMnsxHwB+yMl9N5/m+kFH9u/
9vXrlMv3K4phdCK0+RUNU7oTogO7Ms+p8vccXJLf0WkJsiQtPkm+kenGPK+AUF/n0hs4lfB6OGQD
nroVjYPZ0hL9Rgc2FzwWm2JK6YEesSZIyQMJXdt7wNgHBar+zqhI4+iqvTly0otw7cir+3mI7HxM
Fmtmq2wpJISl5jXMCP+1NSslvVcZYmsPyjrqxEZV/vzWQ27rrQjmxf1YEYYiZX8i0lAs4jgrUkYG
7aM6zlPFSW11gsOxfuMm10zKJtdiuh+aqdlRvA5tj7L1tNHLudCB1XA8gC9d7+p1jJYku1PnHiv0
YP8RL4Njl6MaOXU3JKwo9vUp5SRqISgbRdnOQBzhEw4HD/oIwrvMiJ1EJcv/lw2UKpQ5oIK/Qy+Z
CSXBYJYC8Y2nhWOZcuMBn4uKP1lHibn2m7OlQjSBnrbW7A8HsJyGI96J5yy9ISJoazmZxOQPlE9O
ifY/geQQxxq9gY2CvrKyxjK/Fmea2keGrtINP3SILvFjtXxQCzaKpEtq27/tyYhHz/sJUWrJRvSk
Lw3HKpif2ETLzr9Scl6Yd82UCsrzgag9rB0IbLPzGCm8PbRiRLCFm6SZhG8gq0ZkrxbvrkQgpk8G
XqHawuIuieldSK2kvkCiyGYNMYSOLMiDDtv6si4wgjSzDwGU3MlUaBkZ+v7ggjttd2juvnNgqf5B
95wfIbrTmugYmRuQlVZ8ea0fmGosQz1st2jj+5IcdSMBtVIHpNnCmPfFkiAEy649IWjz8FEneX9R
HXYZ6jHk4RqywxSHn0quci2hUhDSIK1G4T6ukApAtnZXauR9UtJwg5RFDtQKOV0tfZYmtsVeB6yP
oLIRRtDoh27oSr4mTUwmpZLtBILd8NbGB0FUt0eUIcWcF7Qv6SPvzDFCTLvAdxUnrtEabEBo7YZB
yKTzgWkgWwmmhrSLQCoeVdSEyVt5iQHvcm9LhxAf8F3Q1qUOjNDApiW3b+qhR1iqgA6IrUn3qGKQ
Ro1pG5Yv3Zv81tMvosJYY1ppQguyH0MusWdDMWWwHJAL9thuWL9E5ULOrg3PyYtYOXwD7gmsgC/X
t5qCZZggA2mFSkzeEWiNmgPRSHGnYFDvsgMZ2ecQXIzNel13cvgglxILoerPxGRx3kkgjI9uJgOV
jVzhHhkC0/VLY/1WL0pac+Yw4Z+Z3dFtbonNw3AD+5Ypo6eqCsutdeuuSWqls7a7ybsK/ZhNLgfV
EZSANCvU/muaK9dF57ocUAlwybPsl26i8j1KZ9KnY+Fg2Xr37L7YJhGm4NyRR/o4xyBM1QyW3H9I
NWVzROoywwxNwbNmg8Xurs2OtJpoZ5LKd4AwIVY/u/oI9a24zIprwwlLT9VK9yj9W42neULnaUdO
8AigauPHkvIEffEIQkHsVlwSsbmroi/25zMK1djxF35zGAJT7rgxBEOMAh9osqw49xlkr5KdHmhs
pDF9Ig4QcbWMvAuRJubRgaZhzHJJ1DS+WDqJa3QcIZflJowDhvLdqrnxxKkw1LwiB96hqBO0k4W+
FMA4QHx/eF6WqyqSfh2K1sAVQt+cy8c8iwjf5ztaIr90R6jq1vFLUsStBYgZckcopJU6toPPhNuP
MZ2g+CarObV6DmxrP8WmEvzVanFGZUWXTUFWDpzBDBPoMeI42U8yHn7p/N+dBcu1S3lw/lq0tNMF
/tIUTW+mjPlsG++Qke493LNMTHK6y8xMJIfDjNM8aZR+uOPUUAerIq0hmtkhqzl2iZlD87A3loq7
mooCzGvkllDSfq0DM5dcXnk+n0xsgz2DW2bCeTmm9ZUCs2IXiTGC/y6Pv4p4ExdGCPS1QlxGnARh
dXDnkhi0FSAJbRk5EBbw6Ut+nF7b9r13pfOQp4p9f50rApptvslUc10wzP2KoMbWlMbCnEv90GYW
TXNx7aM/tbT6rcaZ/3jF7gwZpg5kx7OJzyUYcmhVQeNl5hDGYjSsNlRd6wfoUfBXy0tik16BV5sx
MzlT3db/6dMEeG3IM3N5Pcz9TqaSZtchZlB4+2QBU+4x0SMKdHOHNXRv4xywPrHur2fk0W2nKn0l
KAetzaoyqj+BNPYgzlF1uxW7GDH2SyZq769++LQmXuUndsvXoVVpUDAqyfAJ9f2iciIvuVJwo5XV
zj1jS3ACr85CCW1fnzLqaCvbrTRT7CohdyVW6KKML1K2SoTNIKcWJIgBKnzTUbgYUvi3gQmm3dLd
qWT6nXcFFnF0uVfmGM7avj2dCjXpSdlp3OiFLrp/UaMT5S9lPAZ9TRhaJx6UWBdxUaTYBCzVcoiI
9FNj0g5pFpyYc6qd8hl5fMRBAOapJBV/VT7CUulmrAktt0rFqbw2Kd1HQNp/D0/b+8JM3y++cLl9
wXFeaBK/jBD4brZroQb761wdqsmwWmYp5cicTLi66eQiKCO45C7FFvaXZiU7h6reedoSwRvGjcw4
xwF34qkV7hZsHeXWRfA0QpF/iR/4HamWiCwTnnTM+kShvXJYzKG3aCmqLYKzBUKEP0J8RgBJUi4l
2IL5BTElL5m46VGb/Stm3P4rxx1W2ibOeA90mkFRmnR8rGfVuEQnkyM/vV6AdrEgR8d8O4CMGxGv
SzPT5up26//76jHjoejPB9k7UGxfc5VHLNElq4+mi9Bt70++grG5kAGHMoxtAYRI4COV31S9cgBu
qnJhBRMWULaNHkW12wYjSmQnWI2NLpniQ3E2w5JWROsqe2du84zfjNsAFCFdtspT9sZOdBlA3rNE
MHx+d3aEG1ahWFIt2Kxo/J2rPlsjbDZrULT7mXjCOZioWIL/6xHwXEHAE4Dy4a/F8aLNINc1oMIo
JnS4H6mN73wGwQTYBgPIgMT244mD6eIGEvdwzYGyZDg7XHE4CHL7a+oILskBR2G/mMWzlxEqmTGH
lF1AoD07kXgiMk0cz1sJ5Xyd3MiF4AtxZUFh0eMN6R6bU8TbHDNNbHNMLpoIP1/a4wU/BnWfRYYc
8LViOcIlxiiWh3u1yhS+6KKy1u1COUJHlyXP4n0PBBMY7KCaJfKL00HuVsBGVNG+cJG5eAr5a5Yc
sG/Tx2y3zaWT0mWBMZKtOCtROJxTOMPmY11C7gtTwiXLC2rPr/GrTaNaBOogzrHF+sSkAnBd0WSc
O2wG4vLVGDfjni+Xh6zfbGtHiFUkRfW8NkYqaP3z6cV9efRoMh64pM8xPdtoBGLe/OUvNVCE+r/y
Xo+u5Z5UlMlsu8BFOi9KOSy+nomEDP+y/wClu9oANW/NA9tZsCacDkXkIw0Vemw64zchNNQza/2w
Cv33CwM+KuROWj7+Xrq7yq0SYF/UzYRo26dfJjA2KGnMBFdiV1AlaTuajMmpykrqkgSmih3fEYAN
Mv/v/Lo5X+ziiMvnRP1chn5s5nwwvDE7cN1CtvkZOQdxREw07SOkdPKh0J2MJkjBdZ6mnUxqH7UU
bwwj2X7lQM27+60ZfTTnrEQ987uYaQD2kRPPi3mqutdukk86syCAWANrOAVa2p9pA9Qfh3YXL4he
r++XX//DUpqdbBbxae/biIezTPloFHbMnHXh/3/en0uDDk6R3zrSkMSmd790UMKCqf3579+/1yrD
QwhRrQV8sfixL7dVemgNf0lcP7Q9NG7TCJSab5ByYlO1Xy6eIVR9IHLcVz548jPirMGMbLi+diiE
vV09reMrXNp8+0usR8cjeyuSekCjiPzfo3LxR8doH+S3NPUNzyiNUR/L45oK2bAVCzRJ4l31hpiv
It3nNuzBGfw8IyxxzzC1+PNra2LcATHeSzj8T0RGYx2OLU7fuqr9rp5U0mzumGraFCNjPyyh5jRq
GRJhvtmdfN2ugUN+vBzYtg9TbSuchYVJFpt2jJSk+URk33G2s5AQ1IvbkGsLlieaChOcEDLnEq1E
6wltJQpyIkPLG1/jw44muZGBGULaewxSWzcevbBc1ZyOjgONwvR2djsZ9QIpkagg5oTZCCS5fmVl
/lScBj7uDNZO9fBNGTq5drG6JM4m+E+wPH4lSs2BW85Ut/r/nJZbTT6nGzJQUJZbIGBVHBlcZqfD
EL3yg/kjyCdwpQXCSZmlDIVLA02ufTzw/sV1RWWu5y0v6QgyXRz7CkWFGOqIzdtoHgeobyOmDm+h
4PcGj0lENyBT0BtHsv5jCJj6ZzO4mEAJx9yr9rLfogkHDqnhdHWipP2WVqSAeCwPKUkd2h+WkmLD
riF+XSNqS4EzWN0ixwCjcXPoQ2sZfojoiDe5wwa6u1fx4PfSDF2keKtM/VZ0PQ7Tvv4FSWuHUiqB
WEPfpKdfh8PAOEUdRa19Zit1cntjuUx56MA9WMe6DUdxYVz9SfbGXOvCezPgr92wmR/s72IryptQ
g7SSNE+dLQLRK4yXoJLceQFq6teBnFx6oJNA3ODzJbBJFBHchg4yKQL/ill6WoJFg9hKGn/0eHN/
weFCSAyFAXR5Bm23Zcdd/K2zRGBEO4RBycFfq8oPtNbzk8pzvvHVzLfrUls1tXMHMMQLBP9T0xVp
ULGSzWSX3JrLjZxf4+HeD00w8KSWLnfbPMgboB1EbxEvGdUtTpRN4bZzpu+UpLpa9yOoTjbGLVXD
YfWvS9Qr+xbn333aGWjs/KeTXYtWhrS6VdrRGQ58YBc5nTKR0Q1qSn47rF4JtUqpdAx+zhHRD4rZ
Mf+u92jlwfajNTsKQua0C1/49Z1mk3BE+LfkVYCH0DQgMLoQO8wRc3UGbEem6DZ+AcZ4hKMeqSZ3
EYxELH0CxnCwCIZ/Pga4c/b/C8tfolZ+jvTOSB/+Xl3uykmKbOe2Te1P9V2OE1qvksdhZayTc1TX
2ku1+HB/KhKrxDYaabi3TsnNdK6rb7U1EyJtdCTXDzlKEV1QyaitDNKHb/9080VARMJHq5MOMI6E
c8786MyplkHGYS7QLe0QrWLAWq0PLlzgJTZuJupQESPtNf9DN8J63Gazg1iz1ottbO8KogOElAIp
2WdXJaaUWjQAT7Ho9TU3dL+DanbEf+Eru5UQ7aqnOxqlEKrGKLXIFC8lPWMEqdoEIKZTC2hrO/nH
xRa1LKi4bfO8HXFP89dveeFNG/Duh0s4qJfiVXP4v7u7+neWr/H4qEDElEGlFnFwlBmqO64rqtAA
8ET+kmp4iPLZhh9JaVw0ysTyEIY7EfP589UwuePiEhLk0xycP3kvdGN/PIRYSJakp1IzeZOXuMS9
oBLhUbe/IECzqnQT7qTUk2kEr54yx0dcJZy0SW839jP8+mOCJHy3LykWaJ9YIbONNDYR2o2nARXg
06VQ1/abxgFvgeNdEi3YpmIyFbDzta3QbL/wWDdzstcD2ZbzDrSHehDpzqmdRz2eFifeyoJX1cr1
iu14FdZsWQXGbgV7gD4D8EZX3GUBcfxTFuuMyKFXvG9Vc6DhJF2qxl7rWMl/9jtrg8o0HsUwPuvx
8wE6LADtM/iFC/8O8slTDM+OmeRyPCBNqoDzRObAmOFNgp4pKtS6TCIEaLSbh1nkFeyRT+2hExrl
TKK1FdUpwQaBfGBIRLp41ZhD67z78rYF2h0S9Z0m3iTyD5brLuBXgOXvPQFVK5KLqtvLfuqsakdP
tS2wihSTqnGYBvgVaqcVQ+AVpknBHYDCZgU4vYONWUbjxrEo39TxX6fJT9LR7Nig9NXKOWY2I5zG
rtpWjFb9E6eTJG0LQZqmlqY9e+L5Kkz3EuRFzJMjxMVFquvpszY9rvQQyySUdq29K8FrLU/RwH/k
GoNTeBfKrZ5pMDLUjEyHDpJM5ZKU5tYOTNchpVlH8Rk+JDPHqWwtVjsios6uwEw6ri0XNrxNA27B
129mcCDfGpLPrTHHUzfTiJ7GQWXfPcoVqHvGV6T5eNUGgSI6w5UsZ5raJjjIeYnJxtz2gzgLRlm3
+Ea3ivlr6uCXyOlBVVeG0zEl8sXIhH2a8v/+7bExkoyxYw0eE9bjfVDzdTGVMJERucjQrVv+4gyR
UsSfU7gXkljnQhsGT7rL0Zy6Ktd+CzVgJaU2dEZu75tfi7XZ6o5rVx+kX/Cd5PBsymrlWe+nqN7X
jImEdttEoe43AiOYiSI2YuPpCfhH09u/tCpXXicHT9hAcKMhXecyypXguth79YDyJYB5Y++IODnU
oceMo7Hqg5n38oDBazU5hmJc1SYKsrzOYT8GN3EfrG7kpZRETg6r1l3mjakUnKJFM+lOaOdhu+oQ
MxPRSpwyL+y6NYSbNnP59wAmLHj9+6TGgPiLwpKoVfQEktcEA1NOCvMef5UW1r0ZqHtThj3n5mkX
YbiN5E7Lsld9McAKJvfSdVhWLqOxLZxqfJknrsYuLmw07snD8XSa1bemphSbM5EGQYs81OBKbZa+
96Kwri4mYPYFk7qSgqk/c6gRLRKXIb5mnttLmo1KT52uUcLF4k1/QmhY0tXaUnStW8H69xiZoxW3
mDiwDY5oJQgincYbQu2ylKmMsBDF+bisZ4jGOoMrbqvV2ckjKtti9+54yfYo7dGDbpw8XOVWjlZJ
ixAb8T+eTVayXfuqSoOJISc3i6gRwERM6eHAoJC+ap9h0g0pYe5ZXjAqowyzA1ZDFzEsiDUj9kRk
7H2eOQDTFAHwRiADqd5vZwBtpZjnPPTdoq4FIGK5AY08s9W7Sxsk3DnOAKMvPlKdjZe3QwsAHsvi
TISOsF+4KycRyiy4u7fikABRsyCkzCgMW/BslvkiKBucM4jvJ8LMI/8pnGaBuOs/XSFFolvzsKoS
OJKqTuelS12cC53UCvGhYw5FKg25rloWMwHBg3QfQv1dTZ4Hluru05Qx7SmVH0hmiDOrr99S7Dvq
AipRB+1oTV41YjDjSVF58zc9TEc62wtqSOvn6WptHyLVKrqW+KMXLITOTCpQnl9BS1NHeBE3Clev
g9wQrwEaECEpltGrSkfvOotXOVB9IvePHdhbTdkbqn3wuFsOOiHNeeJ2Omex66TOASmDkBDW1J9e
xLiG4Uga88ZHLAf2UVRQpZea8GTC3Z9SsPdtFGisDMGcPOyhY3AMS+gQuiwikxOP0M3PKW1dufoQ
QGy0GSRaDFtL6t9uLZM8Xwyq9WXpUnGonrmiJzkaOVAg+VCZEGv1mNEv4SpGv0KDvd19EhTqbZq6
8oOFEaRnrmPa/1KmdxQsHxTQQvqwI1bE9GrQ0oRsmy59A7jAanuI8xyzl9qJEc4t9I20z1lUWEgE
nsrYJis8tJ9ayaVB/hzlaYYqF4M9wCn+YpQCq4HR9hI350sgs/45T5ds7gMyFGvCIRd/+O+040LI
nhZBAjjkaf0uYepqAqHBftmpuaYs4YPymGrWyDEPgmaw1eaqUqw2Pei1lSET4TyKpMA/YY478u5V
iyICeLMOF4rwPuWKiHUh4Q0hPqlu7yguUXdalvlsbMqGEfdg0BkzXKCmiRDTNlSmONYcwMC15ZV+
viyafyZiHcMQvhZmRobsbzQFADuD6ZuFiOIXWS+f3CwQv9Wp/KT8pZ6J3MlOZ2IsGzIsFyC8yqFE
m7IckJ+M4DraBqSZ93hK3rlopUAQ6zlIXEvet6d9iGq4DUF58ycncU/RJo/y3BIaAg3sjyf2RYFX
U2uw/Gx2ltHkg+yLRZniUieuld424/oXqMhOewoMSUGen8hFUUA6AjPAy4f6Ca3Tdu4n5b0psZxx
6xfP0lvDc+hguMn05Jdf9DefborVUQfMoabjPdt0BybXVOI4yb2jXeWjCSB0McHNuRHHAbi3LRLw
MRi4v1TDb8A1YbZTO0rBGDG3OeTTT6vKJvDz2Hzx9YstmZHNc6GKZ7KvspicEUwkGEicAg2mpc9W
uBJTm1MtrGdQtYJZ/n1SSmA0/LWfzdg82xA3NAvps7AXEcGnry7mGrLS4aX0rLL7e4g2C54jJhpo
A82JRNSNU7C4vKYNetVX20b5+PivbbaRJXEZtajl7txoty11zYXParjMZpsA4EY8SIAnbaKHzJH/
ij5eo68M6ov2hOgYYNwb6wlt+Y2XX4X7zU4lA5Shw1JwAKXG3ptGf9flrXkyPtrO8v7lpAGxCk0Z
qLXJbpxJI0fOY1WX6wsf0rHh43FaPOr3LT9XGXQowEcQNLJKsDw4gm+Meh9doTYdnVeNf7V8QAqG
MrvSVSyB+gFanU5evOR80md3rq8TRGK/rkAgHyLuuD4TQhTX001TFTMOX3Mf4k9k+EKrMJts/QpS
OHITmgpCU7chJwmw1j55ByZkV5OSRiqpVAjAebAjH0oIxYvV+rCcVlY9hxi8rNKkS+7+K0EdUpYM
bjz81RDCe9nvc3s0/Dv4I/foiR0x497utVyzZAg9JSoKsXphw4p3WcKHiUKdmWFhzeMFCJA05s3/
QMTH/o5D//UXiTaRsclfiLWqoBc2MTLz4BnaTmbaQF4t8NiFc/CaHII+x0miv6VQH4bhJf7f6a/D
ZRlcbm3F3OW3k2NOxsHuQ99acp8YnPOIbTuH0ebTMRZ/3SKOUfEc0+CO5zBIAG3D7E0s3fpaws1f
Y/hq1ojN579LsbbxSbxl89nHlpSm6cYV6q87YM3lU7OpfhO70XwOa9V8Hvt9+KP5pG164F2jvTuF
dr7pD6y073/eiOhZAtBUqZ9JR+2TyG/Wl87pU7UPFDapSH1ZZWo5gbXUgmX63UI8DvlldVfb9Phx
HEZG9X/uoFEul1svPUwRDVgniohJ+f32ik6ITAcVU2b9KLLvi+DvdrXAJO5cjqCvSkQzXgvAtSor
y6jD6exF0Ed7W/Ao4RQzLSs5Z+xQg4xXFN/OZ9cmZyMuDXbG7KWm137CePHn5ORvA/40WdcMZBXP
B40+NqxYQjeJvQ2b9P/EUbWBPDkLo/dFGTDhJNoKZrj+tvUuh8xCg1rIwC9ioTyaF0dgGrt1hRYk
V/9iyeGMTyqE0ve8NaOQhfyoZK2KgTD/ehhryW2c571m5XD7yVSrnoNjOouX2FjS544+OM/QN1Rp
2w6U7NA8tRorfIoA7IlC9CKG9pMG9x48M6Pt3iA3SNr1GFvye///PKH7jcv2EY3O52uYD+QMuBX1
TFA3WwIQiL/dL2mwL2MXHQdAJMJsorIyY5jQoKFJavMFVZL7Z85FWbjd17zE5EKW6cdDsvKwFejC
zeO2o6D+9qHkFZKzH5BbWQVPZBjlmaAOGN5ADF93CFVd3PKo5pd/s3/ilHyHLD+dK2KCnUcx/4Ff
p9wYzHg8XK/L49LzjQBwpeJBl96NkjlkVLkfdZPdXogpr6td+oSGjOP+Lt2LR/blFDp6sOfchYsi
8A+mraooy4VDj6j9BD0CaDQjYUQnZgO6ykXsP5nGBJ7fPrNcEDGCq/xH3KmwUNe/mTnxa1/XLd4d
jhSF6zFrONyWAxV3tdJW38FnjwqP1kv1LjoIoefAtqoOMRfJfd3pz0sPqPDuHQa2DONs3y2xmlyX
2eAK03vAwFmBRxPrK8zWH3sZUtsuHdc3P3kC+kdcmE/4ey8acVgQHm2Sc4xAoINxIKistnPkQNpd
dyt/NQwvNJ2+MXkB8xUiwv7EvMe5jMbeoUfpCkqKijqvwH3/rn+m2S8cBcH+2ic+6bBfVWERsG9m
VsLP/oRMhRiIkwv4R85sQtm4aRm46NcrvFlZE+3KhNP3cubfsQls3IlSUvjcn2qpL73Jcu0IZTQO
PGB+oHEqnFpOMhpgd6H9b8bAD8/gaFSP6eg10hedV07rB/NukuS2m/59CP0GjHcj0FEuPrh79uTI
nIDP56hV4xtk7rFGNs+UCKM/Vm6GXJBMBQIAl5Rtp+1Wn05G6dvufaa5NfLy4EAA+trzf1+H1XyR
uxzg8UexmqBiEISF1UQWh8h5WJOSPSIZcnpOUZgs9ow/+EziweRpwLzCTB7RJq5whuZ9uK80Kioo
/gJfJOGqkQx7iN2rquZQEbTi5w77kqk2faO0yAh+ag61fZi25gb6tVzdo7X8NSF8OitYRqTdlE1A
WuMnkCpN+cfsQc80KLKIBOpsyswzE8wCpBXAvqX41dHo0CBYrPsjmLTpBtph6XU+rGRYdMA0evOF
UKUdoUU0GII3ELXGvuwqKJ21tRQOKKdpkQe+Ew16Rauru87KMv/Wm5gwS1iEUmxFV8LP6TGHuqIm
rCSVaD6Rr0w3jPoQZ6g3IX9FYfqhSruHko6f4IwGfC7AO4KImusonR36qofzmE4Ssig80w0IO98g
Y/J4S1pm3AIF1nyFl8XlBkJXOCwOZ2aUSGiDFWW9bl4GikdiYEiv69JSuzet1Tzag3HpxHRbfPo1
W+P1RH4QJ+GJGWTnbHqmbyrGjZC1s9/Ly6OkoWyD2fF+gqPlaTVyVR3x1y44Skbucag+ah+rB7pi
0Ta10QnLkfGjaXeZBvQopGdL3XV0KGDH3Q/OL5vYCRS+l6j8P2oGQgV4abql+r3/Fr37a1DXkfNc
R4UR0dqMdo5DtmzdW0Vic4C0F2R1Frt7C0o4ddWpHdJ+0TGpTTU8ATHbFsoJFQLUo+DZy/0CU1fZ
1pIuM/20Tqbdq9Me2iFdqTtgpPLFA19TRAyWigdc3ViDFvYz5mVYyFZrnmwzuAWtwJ7gUb8vF1dl
iR4C54EpRGLow+4KnSUlO6qZf/R1emRFSVwG8cbG99VuX6+nCCP3JwNCpIYPTsU367ulb8pY8uLH
7kpuoMDGjHHhuUu5o7QPdKf7acyRc/5Hp64bpXw/n8kYdaMeJ95J/GAVSbb5nCjnmyNtF/LXsBJJ
kaWQ/v/J1tBkHJrTqcAVdOtJv6Z5r3MpBssMrZnk7tisgA5KEX65ahXvC6Hs4CyJGJTLzseDo2pV
HuhDYxTbhjOG4qNL95ffuBP0peE9mYUGvSsIeOQFi/oaqKYS0tvFI3t2xLftIdKMNIzuKr57Dq7l
1k7ZRGhFN4KvwZfG8CUXigBBkA7bF19JJtGD9B1PoKojBYeaYxjW1ixVC73/jUNBXabZ6umuOEoj
jhxM17drTqa4Tsn19NrsVn6UYdZu+hyahHINDDDW7a+DBoAOJJyP3US7JpGdXSmQmBVzB2eQFFv+
I6kguKY6E16MAUPDJqZmpdf9FGaQXLv7HrZ/ih+utCUthxkKLs4XoxWrjcnIVikwSlRQneCvLot+
KgeEblK0MxkcXCtAJG3otVGINZtz77olFSChBo4p4auFPfyd2/zzLIlXNHQv9rHyfEhOpdQC3EVH
Ob+FwCpbt3IIvQ9nO6Rb79DVHq7JbRj8V4b/QDGJjdrF459X22r3eRpofYSXdQpd9szHae4JYM6I
B6/BO4Hxu1BpbAy4oeGxtENvM7X2+wn6BlR6OeTnaf6AFwlGuO42UT/ySid186kMM8ynd4ZA8iKe
CyaVUiTNoOCDcFUI2dA9Kb891VA7GbKb2fyz97nEBEQ91sgkUkkM0i4JELd9S5xNhZfFo0ZfNX75
VUGtOq2ERhvXoCpZeimNeUy6JprFXTbmURljpdaCz742CWRfBh7WxD1ZbQ3y4dbewARUBATe0U+d
K2YE/e+QMuOckG3xFeCRfeasucire3TxcoNSLXpr2m+4s9JmR1QRej/E4QFA2DtPRLdVtSMspfqO
B+PH8ZhstRnPSYx2Qz7aYrftJJtxblA9o/zpQ4SIl4dYduOfyvdc0hsryxmnNvlq1H9PWJownlnu
Kp1oTntYVLt/fpBSUdldP7Argb+WoU7m5jtcZwBXlPZHfRBTep5MXsI1gcUw9VOG7YhhamsXgkbH
MwyNgBoSnKQOq6fLnRWA0qde5CVAO0njZPD6WDyVZYpYhKwGazAc5t6adHU8/R0t91Dtl9LDgD8M
poxKjYAREvltfua1FcDTLM9sgWMEwxaalj7+sZ8MPpG6IEfqgPynxOeKNfR2x33ZuGTaNn0g/bun
nm5gcXXkzwbVK1pvJrboqSfi/X0lUSuseN8vhqZfw8VW2tgv5XLAK+gdSjVj1dn7czvn5iOz8bAd
AuniqesLfa3sHD8CRhE2kfpWr6NdHnJ7NfbsqTAwJvqKl8dZ1X6pmZroWu0gUs9Xgxi5PyYUQjUn
l5bcX7OE9Fzi6ov0WiFagh7DRCS4ypaheOF9i/uq98quFZZ0bWU/IcZuvN6UCGXKFA7TBUDY8pEW
WjumqyEHN+whLzEBzNimrTWmYuMO6pLktniZVMo8v2KNL21Aw32pcCbYxyrYl+FlbyqdgtVFVlkg
w4MMqsA3ttUNKnrp29jt1uYCu15nh7U5Xks7NgnDfmNBIz4ERU1yA1pYv5abHN/MbvySZYsoVS4C
yIlW4lQzm7OTIRMA06DEJ3IZJPrhjC1jheF5Hb0d33kuMmwgxcevfpY1wXdg2QgLishXpK0s7OE5
Jsbo/CmvtbJIdlG7Y1MLJB8f158Ykc5wd6HQs2LJSyb7fKSFqwDWPYXQs4Nrc0wmu+kgTH11qgRN
7i+uYlhIVTW2oGpT46RGQ2BbLt3Tbaa8sjsu3cqSDbofeN3SpgA9Uxbb1LFcnpVo0tcIqI6dNzk3
8W9jfAU1bxHjnYMcuEaOfoKwfEkL1anUcXvzzdUNd2xV7xeSHFkL4FBWR8XvRZi7IEx8YVMhMiek
3adUHbwQK3dJjy9Xb2X/p9Bxl1I9D4f0NXAvpFKsq89LtVLoEg7TKuLuD4bWvcPLVd6I3SJOEqcG
pWVZYVgnO3o06DuVUaGKdUPR0gsLrX8VgDJL3m5/VLeMM/mdZNx+dssZeHtcowbSHDaCRpY2OeJ+
Enfyh5Q6Ig1KUl7wNLrxs+Wf9ACo0+zPnJtH80dfgWCxING2XzatW+gOj4xS2t0oDstx1B772CHf
HDTSP+0NSeRbBDqJu2JGGWsS9xPiQgwjfsTn9wElIspV4S5bYhx4PvDaG+Y1U/JV8oDsa2ZkOu24
g2p3WrSt/Z4EY0+3piN8eYQhl1rr7UcHUYuey044LCE8J2fa1fCCFELQr6xhWrKttD6URFPUnLXK
AxVvJfwyf+JjhAbp94nIq6nkWUbOYp8lzmOBpcWz4pJZBFR76ZCgwHk5a067YWZE4LkpZIttvneP
ffwvr9HJiNDbRXBv5kTr5YFFLxRLiQKNmK1o+qORRICClVhgGNLkngp1D7fd42lGMrs3LWtxO2lp
jxAIeF+J+LPZg+IC0G3lBk2Rgk3V86tvm3gMfWZ3VYmMjavcGCyQrT9R9dsGSWgDYpWGz3wvZCtQ
K/G+H/CSjxgYEoSkHEd5nBPOuZYC7CSUARSh1y9Nechv7OOLLBF4tz0uau471bRu0bfmImHRLPM1
x915qAcoomaqAT/WmzViKag0qiqG4ODznJCcPMBADJNRw1LbObxBnwQDoij0teFjc0E+UJNwCHyZ
Cq7rP6MdKezrj8knRzip1eNtuVuiGSG67lalR9Gp/X63FZVv3TQbzAh1NLptRKPQX1IEMdaACEjO
xYGvalBSvoFGjKBq1QbsbuazSX6g4IvZJObzTLxxdHqvqewTs6tAeHJxGJpOTDxcOsYfCYaBy/R5
ljDcxqdwylQU0VpDHkpXL66BxlAPWImzHGDs44UOxPm5UaOmhwJXsiK05/jkljg1ZB9NnpEdSMdO
Q5LUUA5uMjG8W6WlHM5uyIZsfnc4JWZPlze0Da58aZM0vifGkoZkkxwR08TjXtfkL9RrfTXccoiK
8ThqeK+o2O/4pSNKRgvknTV+zneNSWpNTARqR/rNRTHpSoGN0Cj5ZeBHfHHLvrfa/MKVtYVq+vYN
ocy7UNXVB145LjRyjWxnlr6aq2DbU8gHTXbvoci7BqZd0ogm5vFHlfk9ZghFBMSolRgYTIB12sSK
fqB0hi7Uj4hnHF7im2bKFlhfbb6I9Iy8Idi6JVY2Qu+lGSpdyXoDNl2CUP7RVKlwAHi57NYNA1Iq
dsv6OvAlHVY3qF2U8MTThvUXaZfWGbza0gEPb5v9PgfO1JeMKCWpZh/bUSc8xv34ZuvafGhZSseD
o1U6FN5/BbdDibpSfDJxW673x/tpskNIH2zoTJdBq2ExC5DUNN2QeI3dxYz7rX+ew1Qx7kW+IJbB
sHaKQBI55giq3k6CJQzXngxAniagkBfTCHTCiODfSV77qzMzRcvQ4F5F6djEPX1Z2Nt/EgOM5r0y
NgkRDMIBf7M8tXP0z5+UCy5Qij1iR3cuiwsh6GYFkEQI+9RTGdeNBr7w5UwBgtz0qXgXE/+kaSca
uCctGkIYMRdd2kPcJ53ysMmxxsr65Por+FJwfagnHB3Q/ThvfrX5+yGvdGLFiUMHgnvUtkC6TtVs
Ptzqulyhuj9Xuxz5HtbcK4sIMJdvxGu7SXGzxDbDQp03dgbkpOO1pbqKCFeW7d1JVhpBCP8bS/TW
0s/Lepx2028Y0Y3/aFm39yVREsmWCbA2hrp5lBV2RpGCIXHknb7zi/rZlA+6Cntplc0kv/WSBDeO
OE3Hlesz5W/QbSH+hxxdAp2v6XWQxqOc4bzpwkMQghOHjY3topIdE2b9epqtGapDwQoweBe5Z1SB
zyjU6nr/x89jDjKmrDKJqNcxyKpFVB7Tfl/LsPPdQpRYKotXBkt/wjHLylZhDArE0KJS23sRdBD6
S+kmOYO9XXWWJrNxQMJKnUNiZT7r0xo64VIsKOy/gBkdEvl9kTae2Cn2RDtnlu6GTh57AB7DCH/Y
t0gUoaw0knNmeyL7Bvw/b0GszC7jtgcKBcZTKjAp7olplQWUoZN5koVx2kmz2l/rZwommyBd8ozF
nkJ1GCk31JH/sKdR8JiFMrLxQRPR7X1PEEBjaYoHnJIxCUOHJFCEbi22p8pTu8z94DbXBcoTsnl7
KMcMI3hxDvfgZf4jmYibXZAruBCsLF8jmcqyvGyXF8L7cp4jbV0O1WB5jDvcKDZlUeyRUQ8aytWs
bwTvC2BFMLsH1EjgKwpXygbZN+x9iWoqngCkWzdXCIENKGJhQzTXbRHGfErL7z5IC8MmmLM56qRc
+5McRrULHmJq2OCCfQMWjkoWxaQTrH0iuzXO58RgsHolT1CO/o6PL09Yj9MSRHiVFiXODscZ4ruC
dzX0KAgC4IYDvz8XABOyEJgXSrhqQiP2/+JSfWmWhyqnl27ypoqarrscmF4w1fO37zSAcqPPuS+w
dmAaZXw970QqLQ/Cy1eeiirwQrI1gKxAbU6Vd0E3kDNGnk5kbmz0YUQBhA+MH/Pkg+08HdXQ4xjX
MnP+ayazCJQbB7ODPZ6movPwpqLcB/rt5K1ZhBRph8Omu4WNDRquRTxBCGwBvpPuFuepocCPjkPI
muw2SN/caJMH6HcxxPQWh3HrJDJ+fFwjy70cfx69Gtc1XqemaQOFUrlGGSXU1LP7INTVXz2fqDaQ
8LTMIoiYY+jiJl4/zQMsiYZ00i7ovasNUD7oQC3j3iYpy70p21tFJPPZfhyH7uSSoMM7jC+/JZii
qA+muYxrllV+8XV+6ma7XOPuTCL/MbgSzDu9CJ8KnkISVU1EvLHSCBER68m3ZUOmr80dPD6PYMKy
XgTiX2LV+4805kAI6BYuxf3m6xi+ygMEUaH+IrSleZapZMKNdXOtiB8UVhoszGSqALnHvlZYq7Vn
qrBgSDllvRYSHicH/5b3hY1ureYiKR68+GwlwaIcC5VltzHxKQ+iTvL4LI4gDa0o4RzceszpVTGF
4v6NoQjuD0+Jgpzbl7SrJA6A3aaRyqbnx7o7OpJTMVwl5NuzvLutQLLLkZuWrykjPxnPhWrewGMx
eQQ9N24A89SGVZnlDukc3t52itsFmFs2PqCWzYz8NrIYsJbiHY+9op6sH9gm/yL/41gbHCKC7zTB
fSacLAQiqThmyRQgoFg+1dPTFY3GLkQoZbFFXqp3SIAya2GxFLpD9qJoIKVvPtZLxz8T5e7KIPqc
AhVeIM1HTie3NaKrvQtIlC5m+UZ4W/6VLEsVGEdIl8BANsiQvY8q5GuvaDuYQjdyjKGvTcnRt9+k
QHswl8Lu2+QI582BHq0iMweExUm63JNA6vKfdYfTCfRqtAZXLTx8bGEH1mYrVa0YgMkhxQsq0VaX
ANpkFxwNqp+csZr948Q4uULANX1YjNF2voqdUPNJ2wnoyGHOGIPi97d5vfv8kek6y/TC8M2DJyr+
1pF9dsO4tBs3r2D9ccKX0pEalpbrpe26O//kPa6sdu+/hDXP4mHbXfC01FizvdibMonPe7Xbsk1f
yqFxrmfxPBSzja8WyLFidvkRGBThIFBJ7h4ge8wUTVCrCNYHabEyCIO+fy2mL3rHbCceUuqBhmkQ
WazNKMxM7pfQR5xmrs/aksmo/5QKWdktMh1MqcWDn1Us3UF03o3zAca3Nw/N+Z91leyL2DO9fFy1
V7zVNnKXmemHJUTiuclZXKcwgDJiH3iNDgUCt6gurPqWVRqwX5wKfilF5JvQkN5w/SnA1uAQdYf7
q3+z9T4znMM9kPl715FTXF4ky//22xeOcIJBH6oZDDuE+9g5IElo6vo7UDhskRN43IndkEKHG/wO
+wrmVgX1g0hVWfkO3zg0xsU2XX6TcOQIB5CxUTnKgCTQ8KoZWEHgdtH/T9qHLlK7jubOGbaUtcGk
MDjEohUchFHpPyaoETM/G4MyyUpBXW9C4j9NrE6rYnViwEW+QS8c8KZTU5NGrxR9eLS8pD74KdQk
NY579YDAB312xHJz1dE6aLV60OIzNqkioXtDHg6s7L4mbTVfx+YfPlekA6/L4xX9j3Wkpo1q5r1f
A70B/wT8Dbapcun1i2B+FYM4TICXhNhgGsJxwQFEOSBtckcUKaCfZ8nUlRn1UOtHAm5EW/q3ZHO8
lLrgG19zcsC4p2O/yR88pfjdLcyfpu/xiqdzNhrEMipxp84baZv17eX+WDtpGiWuFT9DbYOP2gK/
8ZBhHuycnl3Icn6RPa3f80fj9n4+uNgB94YLfCK261oEW7ISaE370J+uCB271CjW5EeEyHItSPHJ
c6GlL7ZOo8hY8/P1/Dti/Ce2T0pN60uMiwyqURXfBHpL5yuArIa13zsaMRh1gDxnOT7kmiSKxGZu
YZiEIP27yQ5LVQ6mFEEz2rj9xK+ZwFevy/AEJIUC8iVdnR5h8pEiQDAEOLYIiFme2zrB040ZvIpZ
R/pd3HWQN5DtoiU7LPjDg+Na4OAR/YdOaLlma4q2EM22JqLqJpd+NEgAJMpM/DD5vG3vAq9BpRJb
FjqFpdtmrKdOb5bP2O+6eKld3r6W5D2Qp+EERTV+/7UFkBIfT+wN4BO7qMq8/eW0uE+JWuKlo492
rgH8UzGJjP3sRjZrfPwLMu+vDbMcavZJg9i4pE8C7gDrcYDyygY76sXFE+AmVFvKjku9FbUGSUhB
SEPX0RequwuPZQ+MyzXLTkNRse2gUoVpFuCfnSw3Zn6hEtgq6ODxx8lR24niiFUI04jM0AHdWK6r
7KEF2EuUgc3nAy/OxYttT3W5eOmk00BMx3k08TZaaPLVPOnCRSirS2Vg+WRbuebWSn0kVrFmFvKi
usA+E17XJ6Q9AhgWjcLgM7KHQ/N1akrBIZH6rmP/dunl5vhLSS5hdsIL1rl7PGwWaGtOx5V4KCrA
Pom+qUYvtkin7SuBmBDT9WHRdle/vy6eQ3MYNBnjVrph4OnTRtR5gBDi77B+ZU7lfWM3MSdnOc46
paeoSnzl/d0/IVuNl4/UXb3OfWG0+j7qPjbE2sZhixcEBEkz+/shlW8p6YaFB0nzUKi1+qDo0n/4
JMQGDrz1ulInxFg+OuvOwK0mD+XzvVZgjVfv6FHwGk1cCnnhaay+sijFjAZ6dVRuv4TDNc23TKoL
NR7xDUBVFxkJYLT+Qi8ZdIu2jtAaa5r7etjIzoIuV8kDp2UNfClPP3BGo6FAiq9m/baQco9quXIB
fpMTWXcg/9HP+tgjMqPLItw7bjgx0dfjrcPt3GVsmgxf26Snb4U9LIASBXv0/PeZiglWtO/w7ftb
z0kB/h0eQFT8B9SeLU8zyMB2ep1OsB/Nb43LBPNpb8PbKvU9tl0FGC5AcY+UUdtYh0bWhDoGvonE
s6R2vHpmYdBxVYXX/RbgjuX+HknioOSeu1KU5as1O6Lq6EfjdXIQ9JLmMTqFUC0cEOZRRDMkIEyo
fe3+CQjy01Ob8owlm8jGrgN4ZmooM10SjJJc4opACSb42H0FMqLgHGr5zRRyQzqbsOBjhfc0caoa
YGCfD6qwfHdTTD7xEWeD75PWetXEVPwGHM6QAjmSwC7JMBKmsOgL4FnoDuFzYdvyhg/I96R0Cu+4
np3iOX6rd75YJEjjZFfpj3JthJusq6GkSW7C34kyzXOH0hKE8ydgulWwKXXXK1Ogrm1XXyJ7pK0I
hFPVvagy9txo3vHSY8UtedeftAdg5cZNDgsfg/PmE0eZUKWAEn1FKhBPyIdDojcTMjIN8o9Uvs/+
hwT++MckPZa/sjVfuY3jbhQqoNfBrRZophyhDs7nueJljPVMwtw0G38OacbqqDaAFonfU5rccXCY
53BL7epZyKZgYdLmr/Zbr1cpuhdADGtIQQMR6Jn9nrITf/WClO5glOHHRx2dqU4hxtKhUn4qZ0HJ
N4BYGyakcdteGmBALMRNDTrONxMkyYbA/oRQJXYxJiHI9Lo2BEVJysPP3JiGmIMuSdMlDAqu/rjy
Z37F/H60cI6Rx+UTrsUYRy9x6vJkObQMBLdyexcgDHWhcKX0bLwLxsuM9p4/M9gPZBq2Twqdzhcn
TOZP7Baz+aTOBlZypKgGulGp7KHYLa9GfyPnRL45aT3C+q6KYpE5PNjwBoSQ4R8DRc4mSa8djMYL
TkHp4cxtsxXdjVJVDONpsNXyk+CyFaLyURtosesc19HmJqBbvTii2FZRT2ebI9qH6O87Orw9Pgu8
OE7OYlTcpUgPT80kVDq7HmFMxoORWL1Snf/e/wzQmT5U2R4HcZHI5K4JfgSRknFJ2ypGtRgxpX2y
RUlUTWyS3lcYLJWKRcIspVAkDZtjVItemYtYSibm5960eKzm6K4m0aVn1EVU3+vK/9VFDAkF7IRz
WrF8T5tOu+SXxSGbgf2+5FiwB7WhYKWXdo3Im0mQjUjfW6F1U9OL9a9oK+DjR7zCszh9hx+1Rd+a
WF6Q+iwvruADdipZcWOD+S6B/fIVEwhWaLHq+F5fu/ePpz6crG3/il+hjNs9MOC/DCPiA4bGfwW9
wqYjLn5oqjpFOGyHG3O68sISQnEWQEsWnF9WfVQ8FZxk/zNh0zeKha92NMts2JxKXwSF6zYgZy2u
EDnaSW9E6Ki4A6uAXGQX0xq6hCbkjryZOxsb0G+P7qF+AgGCtGkO7hFJSNDxP7R2UzVEupf9ti1h
2A/ogElyZthG7OfQCcYUtK+1uebEC9s8SYtJSPZtzjhCr67MtubgutVq7RbsIX2t7YUZ16LDiCvN
O7Wo+kdbALUycUsuDOjbUnbwOZfgRMDO2apJBVDqrM6pklZo9TPWuiYB0I7FMIdOKpgxX3uYw4MQ
Mt4oZ5XCudNJqUr8sWymHKRveHX1uImFV/0QZOAZOivOgajQ05lv1gAONqagGZE3xFxzdwcP0/Ni
lVbt+RY7eIiBUlJ6sZxmD/muFGHdzZLlQZkr/zvGVw9TBpOZLu8hVpD/VhVDjzctys4NOL/HfWB8
58QNs8UJIkvsEzDhB1bU6eMOmd0Seg6NFILE4c1jxxcQn7so7T2hAzFxL1oNQuFjYBQ6uPQ26ztI
QDuvW6J3wE9/kAVrucc8EMgaGPYhZxu634yRaatKZVnlV6RLr6Eli8Ylwd5mnTreaFk7d04P1EF5
rl/vh0ccUnwt9WF4PEoHGoJPwQ5tUsebM2KzQ6Rku5yTpHtjMg+KmwhJ7aJ/WmPmDm2fE31V/yu6
fZVzP2xoOY/RV6mlRN9avyGHTSMyvRXsiFakAfAn02sYi+C93HWgr3m83JIHZDuU4uD0LK+nEnuQ
LE5yd1RjVzP13+aM8D+d/C/xCkWq8m11XvEf/UFIy/CDKpZBAov2QVb0dUzkIc+Dj6QBRg/Hh+6H
kBAyTXtnpipFEVec3t7prGTNO58erTrQyQ4fgGps3wU0WDibfrN5pxdUIozCf+mIU7XFnOK33WsQ
TnT0YL4vj6YDXHXCYKvv1XijVhYo9zhJ2CdGfzd8u/9OhEJiYnhceMO38TyoDrtYSVp7yPex4u3c
hHH8C8obW+OF8CbjYj0mI8qmoi3tyLICfjCMHZYrMXHigyAMeJgzODL4Vx/aaBHnCexOHwSxJM4m
t229JY9JJ1RJyNsGB4TGPrTVfK69Zb0zyXXAAo96pz0aWLomUYqOh3acyO+dvTynl0sXusLTkUY8
RtW4OyIPWIzd6vnxjBQSHdqF123XIO0NjMMF5PMU26Ktm6wzl3E3EpAgev6GXMkcSWEfQc59j9sM
tCK+uAsIHjtlC3NYwN/nv8h8leGolQDZIBAcJKnfW9ej3JL1hTXQ72zOhC4OjvVfdBZx8MWDkD1O
7DmvucfKXsst5faBt5CVri5d5OtIr3Vy/xY3crhDNCSkJ2XGHHHAe/P4bAwHO2WPyajVMuK00/6x
7JWH4FAwvaWirTo4n9N7XLxwM71mvtde9SSxvfT+NB3qmf6gykoEygTf2h72hXPfgQ/NNmX/wEZT
aftkCToqCuMMAXaUXQMVLCIqKo2h+nwOorshfz4mIptulry00RocMaZJJBbK9RS6j3yajNf7VWYX
8bf0cN26F5t0/Z2JtZgA7GP0/VYbpmGPCJR0uNkJ53Dv340gbX/0zExJdj2RvldtUe7WKMvExDa1
qxfsr5VMFHihtpb54LgOO91ADPH6lP/lEFwJqTFvqlNqJ8bayOQiUFn6vKjQLcu7swpqA1LhQAlg
gl5CUgWm3BP1AljvkUyT+DSUQLmRIL6csn4S4lP3rMxQHmmgQ0mUIa3FL1anUbUBg4Rug9QALzVA
nVFwoWZPPb5/8x7ffRhH8vjrG6oEANDDpl+wM61tuM3NXpnc3OJ679z0vE11FkjXVNqevA5eLdMk
13un321NL+yXvwgouU5hU5neoCVB2udo3Hy2lYIR8lV/S7nIWapBQZmrnfUIKJYqgKDsaqT+y2bj
kMIfDC3//YdU6pBwxfKvS/P3W1xpvWW40Qt4Df3DhTM9UNdJaZFSZ/VjVbbUnZrdEwg6BB+Eyj9O
ciIfska2qct14/rS1hAnXCIwv1QiSUcmmf1eTV/eXTTfqJKfLH6h8olYsCfdJpXfuXtHVGAPKy+S
js9izPfLOV7tnEdldSAKXi64pcw9JaEbT/2iSf0QpO0UWtj9xLLYC1fspgiZvGtSJvTNNFm8H9x4
TktO2SG9eIRBBCPihZCYphc1nZOUK+2hWaMHuguv+2KzK0ZAbLdheF4Q8i9zG3QSgcrXY1zMbeMl
2b5oHXSHoJBDrjYyiVhC139IZN2G9CQNk5+azQT6R5dleKDVxYMGMBTBbV5D9hrp6kBAs9uvPjWS
ZB8wsXV6upACoUAZk41WfML3NAfHuXoaDXhmYDx9900cKkcwWcdPfC/XtCdSpV5n5eVSReme4ZAE
0Mt9UrAhym+pjK3lHoRxcy3VOh9lbqzb8NmwEf9lt9kVE7btmRmlZMVT5dNglQ21h6VLAiQmhzsW
fHBKa3Plo/05c9MswOlbdSawhdGSqj8QmPTNu1rw9fNDM8a2gbVSphN//Y6a3wWEhKBqJZ8JNNa/
yOwTxyjj260MoALEqZK+Hq8ck7h70HAdHyeqYoiAy/ESlLTbTT1NPQ9zGxtV19yp/4wwkA61JJEE
E8b1LTpJ2k40VTEcfmEDyWreL7PnB0yp2vmpn8+I9T8rgX3rAncNYI16jAtV0CCuANYYfy/TbqM1
xIu4Q4NCZPmjLwsDMmqn5aP8npE81Obtl2aOUt1SRAlkCPN+fLipoDhpJSD9o5kWTAwkfzZ6u3KT
e/grjNODcAx525J2G4wTc4IN3c8Ed3kWDfj0h8sHHue+2asJYOyKd/SnJtazFVektglQrFsXx5jr
uie2gCzN0xLR5zBpO5AjcrfhLjWLoi3vnPkGqLxNaUlhnP98iq/CC2SjaTfG0QUFH8kfkrbh5LYB
H+6NTm8ViSlB+f7uNA8EAXUc8Q2kigoW43v8cXEmLrrHeH1WxjHeIuixXroFgdN9BfixglAwGWz4
/wfkupM0Egcv6FsYYAnrfriN9Fv/LvM/q3DeZEvpLrmu2b6rECVNJg6a6KBB251Y3qDCnTcesutj
UMXzxEsVXoexLiZtym9SGCrEg5wJ3EeALXRBcMKrZKwgsRTFnTeNVAidNRg4TvWTjPG6GYvGLBwM
IH4r2klc+beVAfgUwOkMkB0b8WVfBKR/+ffmYNkRclcHa4EbIdrg1P2/8VEjBShun2TurDrg5Fgq
4bULgwkJUmN5FHqnwDSvP6J4Dygs2lax8eRJX5sjZwfyGJmMApfrkKi3cCS6yHuYq5hLF2Dnn7mb
8y2iEwfLlNQzyBJl5Pc01kliifmsDmkHkIQci0WNtRfPfImV7VuaAfQxjlDCmn/GRNZtKHSnXJFU
Q1NtfR5qKGBHGyKbZlQjPiloj2oLVeToK6LKL5hI1UUUG9GPHpO0tWlJ2mE+ot6SpVEA0vdskWFH
U2JzpuZ/arS4zlajiSKi2bWpbH67JlRLMtfDxuMekY1glqEJ5uhimB0I/MOKHKLEtrqJv8zERTc3
0PolHCgoS+JH4OS6z2djGbqdRdYk7kLd5AimGs5sifgpHbqVl9lvqsoK5Jp0Hg2ejjmvOwDAUdEO
/M45O/PsL5Pqw3qjoZ6S9TZQpmmmm/XuV3o7oPrH530AZbZsB9JVL6BDvWY+dqR6TM5AKgVGiHdt
WcXdc8YFcOFB9UgEArBeFv7aw9FESKLvw8N1N5KVfwKz5q8IoM8u4JBEfZ18T48lN/uPF4y7it6m
t7KpptpOPmACyiDvQd0tg9n16AIwO8EKOkb1TXLrKzcktd+b830uv4/u+zyL6lVkXQkixdebTqSF
ukCUzmc9YDUCkozSv8rpG/78JkdJJaxfk6XrlH5TZJrYiXrHdKni4JvkWe/wJBRcafonlneCSfZs
0YTFYM2E/GG9GC+7dtVWU77FAca9HX/rKT6kD36A7xXXAFkrzmKDEhqdfD7AIef+Z4BF2gILlHFe
23SNfjoUsq5ILHqO/o6n71DXnNSgHa8iHfcre6Kwzk8YTiTz1S+lNRzf882CmknX6TQ4DUsg6cbw
HMYilWVpjgfKV2/3iqwZiP0hMLM9YrrwHYo/RgodBdDk3pAg8PAvBg+We5Mgx34MBooYyL4gAYPJ
+V6jUJERVFZIO3C6TFpyrC9u+GvGWE0GrsGH6HPg9XZxvmY8b620VcrOBaiBCx1l2BG2xhQ5yrqN
E/bSBuoJkhNXSWXdzrZffvppfNIX/Fsnb0gHz42+zML8UeL0GrV9/G1E+2vXyhGkgq54jmF49AVU
QL6N55CBPTIe8uKnBYgIAyKq+RPRhSYe1uOZUIZ+OJv2rKxyfRMAwIRuAvzKNO6TrgGAD02YEb1V
QM2+0t/6Gu7b2aqx27ax9PMTaym1JQG6og19xHIz5sR9c0U3L14yuGeR+1BKDebHMITrHbgGOlDk
bDDetDgJh68CFuWEUnCKPqcoX/PiNjo56mf5xXHzsf9+tJ90JYn/FhrXuMzcSSRTyiU/bN6yJRFC
3XIw+rCSME8BcgrMaA7trKMD9z2JxRUWfpp5dPQOwqKLAklmkUqh6jif8kDFE7Rd0ZWVdQQ4JAup
grI1wzPDJeivU/Kbu+SYYxdbNMhQKARj2amaqqFmIdKg9wZ1od7qzioiYYTWfuwbZfTB34Cc3SDc
WpGTi5TEqTLsuHHuMEMoCwXwHKVDj/48n1bEhdHFm/nKwX2/zI6Z2AAV37kc29OO409W6jrTYgbw
WTl1w5OAwiFWXaqlTakxOas+5TDe37IRzjUpphc6nn5EIoT8N/WNg/hHivkoo3pOIjreJ7zZTDsG
o01PQ9Raj87oteadLtgSA2g0Lirju7BXII3fN/ScJxe+QLfmETBPtLd6qQP9bMOYjZLFldw1FhN/
fcKs9stmLP2Rdp+VjIDyFkqzaU25xYmmWVLgLG2hpCoaEXIxBu/Eu2ERjpu5gRIbbqIhjNU3f6sH
QOq9Ai5AtNd71rwhw3qKTLXHgIfof8J2j3Yd/FLA3hM+Na98+rwCwk3xC/UunXUryO3qQ/wqPXuC
NhOZGIyf9KIwcEqQ+c/+244FYFHVahCfF4RjlY89X5dOas1XwCKPwyBce32nKpd/pWEtZumEVXnU
o1XHfYVip6Db/qu5y/eQiHVv+ligZppUMbxCqT3F5vBj0o7eR5A5yIWwLu8ioRYhd4bHDJaGRTbH
xp8nA1WfuxAGYxXqb6pCKgxg3BeI/UUXnq5565B9v/fHEO+qlJrBU9wYhsnqcY1o33cU+RSNpK66
72gwk4e8TTX7Q1l1QYzfqFmLTdFDenN8fCWLdfAXJxHLd+4UDQ4VogL4z1T4ub6B9V6nMg6n7gQg
Im08rYik9G2E18k1J1KEORbb5H2QkEPXxOBmeY7sPMnlkHha3IyfIrndToiRZW05UpTTWPoNLdlc
s1xVAgXBcPaztRReuDcaWjY+hU3wsdF4fl7UV8duXkMhZ2C0vxitEX2mP05VQAl3U0170a3SPCTl
G7Wgr4d/lNsztJ9dDyQNyDqUTxkxDbYPvzCq3IPdVUCT8gICmAQ2CZYLQTBKxnNiJQwxG2Kkorcu
mNsspcsc8464RhU06GMAQhDW5yltnlctGTDX/Fft0JUJaZHJuPOHhlWnDzNiAMHPKhj4YA/7iGYM
Od6vvvtSre5hwW2kfMhYwgHq5SJylVnEjT5lAjBmfiaUwJ855ErAbBgFcCukrYOp71r+jDucb7Dq
rGX7gT+JPXZQfp4t986SkbrIsnq3qyztiX9OvEU4oLL/cFQ/nU0a/4qgm4te9G6ynJFe7CBUHz/k
0gvG5FQ9BCSH/WvbZNaouZqSSHaDV8QolNmvJZcyaiw1afLprefmdLqAmrfwPauJMKbqUSBpdf+u
noHJfpVsJspV5KgQB2xXJ9f2emIq/FXWHNg+2OA5hLU4/2dKrXy94qviQYoRTXjy9+5+M4ZmyP3z
a67uJKMFSJQbqh1hHT+gHNSh16zhGqYoa9iBTR77vsUsMmt9UvDV2IXTMM9hjc3k5xitPRE8JCMB
pT46k/pxzCFzonlsR9y+V/b+kTzWzryp4/GZ2QM2k8PKc2A/tnDJiAbmQPeex7+5jgT3syfD4U4D
OVdmoq/J0EZGC8Qm+0uJ9mrae9Rn/b4+Gnih55twSdcSeZYVzmM7oDtGZaBPrXBRjWTxu4cIH2Gl
O/b8Gx81MUV2Qt5DaDc+3DKnd0cOgHmO5ROsaOEiLXug8El/loP7iT5rMCEHQ4Syivf5tY1yJyuY
dGrLut5vSHhALvAZDvFlDtoA9EkfUwnahhu6eJC8McdSf0wW7+09Le7WcyHHGBkFLUNPwyxUTmhc
vYW+8b4OXmulqANWeOb4k56kcCr2gpu+f/zO09puuz9+rEb4NyEjFqUWirmTZFIkL6rBbc/hCxS7
Onuxt2TM+F9xhy9DnNYyLq0aF91hcqjWnDqngueoGs+S4g3J/vwwJQIJDua63JPTUN1sJ/lm79y6
TK5CnBNKbEnN2NX+P8rf9Yv/+SpIgQ/bjW/GIL4+uAQVY+IvIBfu3dKZzdYc7R1xpconWPOMX6TK
DiGgngnN5VuTTyXUqWSY1k5JULGPE2khL0i7+U2bNtYmQRLKBigfFQFM4z4iVDmEJ6EP4rvgkkOf
+UdBBWAHMTzyUaBDX+5tXl7SoFgOsPwGmkjposYdZxwyQLg4vwmCmYZCn7IQbmz+4s9BgH3zbZU3
JJ1PNDZJ4kw3CJbe0V2/+gBbm6CWe1oDSdE11eXccvSSRdksrF1SukAXURaxB5/OEXr+Gesx3rlw
5uBO5FkarCees4Q4BfLva3/bZPwfclNKOZz8Do4HtQwe7tp/SKR4p+pnXQiIHIQpmtjoJASNDsEq
ck/z1IFOmSX4+kKmJPnJcsq0xvz2eaSqn5gerUfV4UQk9pkcvs8aiBfc0Egsf/fsjCm+yqGvVUuT
Ep1h7j0/jxGHtXEXU4c/BfWLvZQzTNxpt1WqKQpBrd9k7/Bdzrfn9aIk06akBBejX1ihWtlQiZxt
AgtPj1Y+Co8gMjmxiwFL7fUEqXwb2esY995aTQCQcLOr2YTlO0uuYNlo0mkh9rTc1Y6Wxas8IQRF
ycKl54XNLcV97H9b4AdPM6k8HVIFR4YmYiACcgJXaP4XIEOsmM/E+6UcJgh8aOH75wVJeKoQQv+4
Rt/Beqz3ywchnWrGk6hDxQRp5Vxh6B5r3FD7YEXGtpSo2OS1mpk5TuiIiog3o878wYJCEKtrAIpZ
gz9POyatmcY7ql6NKXJBpWFb5I2V8C3jiTxAnxLkd8d/o2Ig3CyM2Y27QhrIAtlAEy8lfdqgDLTX
ug3NPeLcjlfLNr4v1xL5AH5qMFoSmNpjDc45lcZrKHZkbH3JBsmOv4mg8/e6HPIGqwtf2ETulLKn
qvRJpvr9kM1zSWzsQPxjyvWaSfBs4cUAtNbdPlqZpPr+G1jMGovDBZhWEJoHKNkGKit54RLjvRCZ
Nd+CbiEdo73JEywmFGi3HL1YjP/3mXqUq12mUKku6LYUHK3IWCLjqshS29GwpUbDltJpr/7L5BzP
bmusZLFUbSPZY/iQ7Xxtq2u3wVC+woPe3FG1fz9bBUmBtAAyiipqveqs6bSN96rQd7vHRItBezyo
PBcDeLjWZfwJcsYM8ozGk9wJIPzRIfoPJJ7ul+bnnteABYRB4ww+ndAKXmCVr2WcEMdtDFJ/wZwM
x3QQj7Exv0FApHquSTV1nEfGSV6aOsS1+dmq4+QpNLXiEv3Wgx1TvgMprAkboo2RnMWRkcyTAPN/
vMZQ1qhf9rj7Ibq0XgE0rfInEmx+nvQl8Y/y3753mvKWorara15tVC9yJWT0rCZkwvFZN1fmWcQN
GSiVzO+VBgGMtE1JS4l4YUgEBiMe5UXNm1LkDLiw0DEFeBzfQCOeo1UKmw2JvUmlXguW22WsWgc9
oaV6+SuWr1lhmMeEqN9l8p21vq452M7t3JYIKiH1dHqFQErcOe4j/rE9XBfDSUs5E+MwCUW1zIXA
RJMVge69bKMN2XYK0X8z2KZtRXjakNQnhiDzMByTLDk+U17Af5+gw8hbPR38mR4/b3pFalgxRuIr
PpPrNTBmCswFT7axSApQc6VCryz+A2b6yeYvNw29G39px0msV9hICaxpH4f90peyBi/u6tXEZOHg
Oo7sz/ByV1zDseT9vCDtLaafNBoD4IQGRj5rU9frfaisd+6YBjfkBej8T9ONYrGq3OGLuj9aGjIg
v+ZDkfS/xOWuijR2iiRiqrxhVNpv+vr4JW43cd+uNrc2EH2PcWt8niPHQC32nAFqxqaLmfGKbePk
LWg+q1puQrjhUqjvsu3yIWaPvAJnObGSkbooRigpzOveb+YcvBvu4EtRS6EZKSYbj4HRuB3159MN
pYxlW0wWDT11Xg5gKMYIyfHyvYdoIietaRRNzQlHcjhlOY01luKclyikWG64pQVtVKqAy7jUmSM8
/dmNo6h38allc2yWErxcyGD6vfrfp4QDFKQoNuOQZvtrvH7SuE3LznFWn9TetkRgYnhz/IsgYmLO
a44f71QvbqZhrZAyWBIe5B3KhZWezragj0IB6IPlf1ZXZ+6N6cwlySchU4wpjXZkcfHmBBEsri9C
dAZ7PXbuEuktAVdtLaQM85eA16sgaAKKUNammYb/gooEr3z/PRBXwUhqXnr4N0KzawBXvCVgUoUM
5DYaZwRVTEYK6WrsA7gjpJTxePeiJccbWgIi2rR2KVFANQ2dERiHXFG/w64BID6qeRKNX5obY37h
nvPqCZs1LXmgJHIVXNOWTCi4+JAIskZ5SI40Y3yV386tWYhLu2WBThD9azgaNGYxLD4a50q3cZ3q
mmRKMcGBVKCrISE5+SgxgXPy74GfwwG9V1JmfKSTZsO7tklJSzj8T0WBoBJ0szDDt5GFOfy4Yro7
7pSaifcHX74yirLy55KcYfVLj69i8G3F5vQtHpU9UhTu1/EmswzAW6K/eYuL8L+QAyuF7V4itMFV
+9AZTC0L56ruPmA0t7LSrFfR2PXPPZfzE81BhSOf7rFBXfcCBZ/BlZxR2kLNWeU28x4mN+Ex1hu2
/jUmyW3SkurExOyBFMsbxd8WqD1/4ouySKfcQgkrCbP6o0/jrOSv5PwjpwHrHSN1qjMbs7Zp8WcS
j69NHtUf3d85YenOaxhuCg8Sw6vo/NdXBjH2rGI+mtSKE1sueBmnAzSD9fOPw4fJ28R7d0xxm3a/
kQfnIho1u17tymjlNXt7ZLAFy99suCa+vM9dpT45kt8WNl89A2xOQW+Bi7+3dWg0MpFO91h0XtML
iaUrlXqb/DAD7oz6ca9cnMBkog/tPLhQdBB8qVcbROk6MISG49IA8pL/RHJlPJaCgepcjLmdLdZH
9RyO1FTIHHKElEz4//l50o1sScEs5TldOiRFhbU5sCw494D28QlsAtV1dM5x2hrzYzUy1/wlP/fS
8nXFRgE7fLzKQOrfjo914VBBlEkXKEXCNFTD/V89PeGb/YA43euKCP6pzacf8Nlb5T7cAJYGO5dH
rQUfvdwATykU8jqgl9N1RHfBnJ1t9o1Cl9GqxHBbm30eRTKiBbWSD9/9qguVX/nMvCTdJI1mGT0/
qWPWfJC0aoU1kOpuiPSyLXVNg6cqbRzqAjSJCiJVh5Z8v24E100kRUYZOL5N1OfK2ZDb8OL/GJO4
ylbmFlw2MAQDYNP0smRTOHSmNzS9TcLYsPavx5yvXF2jtaCxERw25rkpuiv8xTKWKm1HKwtbgIs0
N5mkQpGS8jJD5YzbhmKnRgOV5Zj1niBQKodlLOiDlHr2l5jKTQkdDA1ZWtsjdv+Pj/5Q/+6uxIDB
P9yk2nDNCu1+62Qiea00L6AFnetVSF/GggcpMmkh7+rTWRbODGMiD526TiJb3H/Zx04CMBLFMvoA
ssUwMZT/PD6+qNhFcCitbwHHMHFKR1hSXXvbySjp/eUgKlDlQqT1XLBMwKn7yGOuVWMRwa/zS7hy
z4iOrxBcEv0473+rpsQT8PMKTgdc8YrWwejAS4I15YXM7aCck3uzn4gZkND8nqSXV+XvMoXjzzkm
P4gVgeAinpq7BEFjGuTsNRWXSt+w5WTR4kZCrh2dkomcg5surh9GUTOl/5s+NqEbQNZ0MFMFYOej
/Et0x7ypPSxajF2rW8iHnj6ZtjKXNZHmtTMeTGZsrifbX6J9kyFkWhyxLcgmlfnD/qdqn5Cm69vi
yBoYlOv7osal1lC4GmJZhFzuWz8f6Xz7UuMtMDRuAWKEcBWNFB7OE6coX1kWNEeOC6/j/Aa+Hmpw
3IAAZGWyMd6xvZwUVqQF52lCG33DkPSHT65HcSi6Tax6Wse3PtyuMl6Q2HBK+0kuGrGWOI82q57f
xJKSwf7aLrG46awXlET8IBidZzBtpR6J1dO4uQDl3Aq2mxi5ZEwYgApuDiVCZ3M4VHJXeM7tjWcO
YhYw62jvyabXUVpwdxWPKSrTA/s/WHVXMuEBRbdGmEcD6Atjlv9uERwWsJMb7QyavW8Q91qjgBOn
vyhGgZg8VnQ0RcNez2qjwDRe4GwG1GajQH0/RaIoRNrMiVPRd9j+SdPCXDli3U+Opfwey9vOKA/z
OElMVA4aVpaW7HJ45XZ4KW95IAGqER4i6mfIHBZJsbrh/pp1AZWV4NXAZvvGq5ob1IU8iMsAs6E0
FLv+n/8t1ZcUsAHVIUWZ+nBROaxqaljaWptp+/tm40XjmsVFQI5A44B3VRQEZtZyrxBMFWhtv8tD
hWAVDS6qg7IZmyvE9B5QwZCFbNsGJdX/scXqMZGQz106+X3aagssqdGsHEx/yYIhIFpfoMuPXE7B
VdqDjsUqdnVfy/RozqQMxwskEL6RRBQFFmWF9RZZcbIm5Vr7VPZ05D09zLcxBZY7+8FEgowinXCn
8VCZy1aGtTxIITXJGFP3msBknrNyIhib2BJ5xeZqePfb3YZH4Ukwq3WAPd1UoRLeMOvR4bEPHepr
whhKtjQq14R2rWxD1Xs0SSp+NMCRAB4tU+TroDS1H5ccuJScTboNwkpZts89VUiq4AbiJQ3cgu0M
pTRl9pB0P/ien983gMozver+XGseiPzFzjReocPpPRIvUGOeKAg7PBMSOzHrenqjWuoXAwMXUm3o
HTcJ/9ihe2gMhTVTIweZRXb/+HknBSNas/eRchtzfoPu/exavLEr6Il5NbidIwohfuxo/wJyL1G/
xpuh5euhudeNG0TClHs0PTPsUsGdkAFiptsaoHJLE5QzaOYPfdvtmh42K1QAiBu223F7ViAhD7i0
twqxSPXpMJWw1eCQ+vrZZ3AidXzdCeIhnA0KgNJWijLKT9TBm2LleyesytCAQRGn49OtHKaORQVv
aDRPZhJL9VP8ExAGNmnl/LJtjbVKlezewglpXX/0cm0mzBQPF95c7fljPm+sS3HZqqpH6u3NYnf2
yeW/mWNPEcgKsuk435p9cHw4Mz5lkHOqK2bDJtIRk+q+uZumo6vO077iVR+RZlD8cqVuzvyx0wRT
wviDQp0iuSVW333+Hggl8RckDTa+vyK+lW5v+sObqycwLYyKxAuqJ9CL8MhRw4SEVrP9vkC8uXZx
FoC0ZSV1DTuW1iIWWMhvVij4DViY7MAJ5K7N98PX85tWGLqEEKy0vopB9jm0xr4uevlPWLGK+q/V
dYIZ5DqFft2sD6XXxSxHslhoVGAzYRF5wdy1mOx5SuU9XxgmP2uo4We3g5i3AfEJ7sMUMec1slQL
bmX1ubi81pQ97I9CWGR8pHkkNOYvIX+YrV/X9vrOGGWgtaSrbgz0qSVVnz6+L0PWtWr2Jp7yUy+s
bOG5Ms9A4FSpJB9zbl2crVArDf7hyFvnTvhllGu1aMH1gM89IIc8pZk1+D+HaQp1n1oN1/+z8ZkZ
khRbzOw9NN6KwYwgyOOto2fKAIh3TtoYfragH6RFxpJvKCSMIbZTC+phI206n5JiCIyp404LcyYa
DN6oYXmx4q3cWx8ns1XgW/rRmh8DfZ/E66GL6UiCwXHXxQZOFzjXccs0EiLMpkOfBhzhrkfzbd6X
oi3g6tFAt/EDFiO4CwoWsPpOrizwwL1G0O88Iv8DhQHWUhYUS0kOTEp+mV21AkpKFzf9Xu/+8Fmo
dUb60EEiRimKqqsFMeLQ+yI1Pshm0YRaBEnzu1QFJfqWci2zv2+WeOaUcTEPPEE4deD0rENWxktf
E3118xm47uUkm0tlvMFUQODnS1c1uSIVlbbbBhhS1oeGskQIs9wZFD5PnGhj73ibhTLWlDilgnNA
p6H2GeajOOnUMC2dZrCPgJqOvAycxU9TNe9hJMMXMo/OpIylYoIjR6nb3e9LiBe7RvZvoGaipQ2x
a/ZpC1E0tSkTCkEqM/N6oHwsDWJMJ404wIqlCXWRWQNksiWb0sk8x/DZSUDk3+73TviaWR12/Ucm
KkHSgLRzQwvvOOUDxdJ3NiMmGI2/2u2CLXQ3epk53HUM1tsBnSsq6/888gRcsGXYti6c4bVztpVN
Ag6M+YhQ6vpAXGbNxsEz4x2lSLd3PRuWevGVCqNAIE3MsH9I8qteqtIO25GHwIQa6txcArbdJJDc
fZ5dX2eBseW+sdd/2Nrwy5cgnDSUqv2QXs6fwhAGl97c6SjZRwOn8WL7BnWq7M7WyDLfemz+RRz5
q0s9Yop888qlUfbrEsY4QzQQV3BC2PeicxrCa6v7ssCyDYY+sAosz+c28MJPDk0tQBoea1BVkWtX
k5o4AMNaR5ryruwUPJaM2C5CP82HUzE+F9U5RJHAyp1bu9C0uF2Xcg5WRd1PMzpEdkzHSnMK5DjV
QQMSSqiwVoPdyNzhjfg0riqtV8wyiu3Hfhv8QGkxCl6oSQOgSZlYPKWgqIR1m0ZLsn4MOHRg7SNz
tS+Fz/f4fO8THYB3R/e2pLXWwcPTC5Gonhjk8xW4/HzHySEJa5fdSU1zodp5x54x8g5b/M1nGtHA
LfGB33TQzIClWyFcRVR9DDCg824fH+S8xpfXC91xLfIa097ak9HOJwW5uNhQwhV2Vqiz7W0YXCPv
Sv9Sb+t7vKtaHfJrYYUoE51iJ6zwZ63Z7xXSZyfq1ZicC/zXTbX7aFWVzmwcE8rAxbbJB8fk/e0u
8r2qFuaXXTy50tmdkaNl997WhDSZZgq0xq2drUSdv2iQygCmfwQM8smEGYQ2J2gIQA7mu5WyXqHQ
8eueSZN8d+ezuj6KOkQtDkUiW0jFw1Yz80LFsoabZnFve1WysKSPrYQwLcnvpBPn1YZBlUKeUft6
YIXsq3maOLFOp7dBYFkgbg0Q8Zv5TeXGWr/bhZNreH/IU2Y/be+yFygdEWv7h5jzKKTxVN/YHHRn
K0KaniXu8c3o4wCwwO7M2ZATyjnFPJr8BtjbpNqqFJvk1s37vm4W7PqF5ewITjQrrUtAFfWtL8sf
KwpoMuM+p90aM6KF/gLbyTP/i+Z9PHYoabuEyuzyvWqwgYZHHb+3vNX+ayktUlO+LAAJMni412xJ
n9zXYB3l/EvSxCCO0E7GBddnJPPM6Ix7iK2MKisWv5f4ImdujSaydtmrnbiOpwDyl3h/NoWLpXWm
lQhkpb5ii9gUN6YrXbmkqlAGWTvfEEmOzYP16Pg2WDvB0bWh6oN5grh6IDDKtzF6FMUoc/FTzJX/
NiMm/PX4oqXcbdI5AcbEGhskQ0fRzjxD3bKFJT0McwgfguH2FRWERI+JTzhlZlf7b0XA7mIYemvc
qUsJexVcyaKJiyT+x8DfjuJ/Mlj6EdqHpx0aQpQ5/xc4TAExa6A/PlSgQ+0uWtpl2WV2L0Cgwhhj
kPBEhAOVqKOcC2x3GJ+lyi9G0K07NdqQYZa2ZJgPcFEgnP1/+9ShTvUN4n93XustDs7/GinqPdiY
FhWWlM5HXXzqOZ3huwzGeSpQL2+lbvbdJPo7fCPDGkfEuNGWqI1Nvcih/QY6c3/WTMp+5boYrL62
aL9mrHgSYuKbvfyD/Me874qqs/47pnPm+SjYXv44jKNw1CoxF8FUE54kFs4EESA7wE2SG/4Iv+rG
UxEKfwiMQv0orG0G1PHF5KPlLCkjWvgTS3icQamfMEoBiZXfJd6D8e6LXNWW/6kTQnygK95b1oeZ
dVIis9Ac1rL6Fd2O7auBQ8BqkrYXWHT6RoKxD/SLui4vbc9Mbh5JT343w4VZaXSMnLC9jRhfE2To
B779vktG7cMemBuAPLnRBDQ/wisbu26kiHTcz5AyuRi7eLUKAuJJeviLZSf+fpqPBClbByHn4vEk
S/AAW2AVoQtmL87R2A4G49MGPKd5bvIaGynt+/QajkzkpbbHdBkmH2alAp5qZx3MiwB/7Nyb2lYU
wHCZAQT749/bAl0OQUJNZJyGOrvZUcUlLSfHiw7yxUr07ZIB1Zzi7iaN46XhRNzzNc2VzZiA1I0i
wLiU7zptqkqvteiloGbvd6COELOdAFPvDPDN5C7IB0sC7Hqe40qTZC4q/0yyBlPV45deRCQzGxqI
wew2DC4Oo3gCwEhEUe7GJcjcsj3l07IpKvq0tDyW7xd+ZeCy2P3/I2DDPWbPotrowbVkaTx4FxK8
5Ux9dD8OacM6VHBxkfR5vMm43beScva8AyRMm+UITQQq8f+Ozm4SGGoecTbeCVDYBW43bS7yXb3s
LkNTLYMbN7v5jlKXw4dE/cogF44hYishtOHfNn9rmld2E4h0+w1BdhZhxrmW5Hhu6AkoENR7WjJp
sjsP8hSWrZNJ0Bu6H+o9Hu1BgJKT7ksL/aCL97pP2O8k7BUqMWS4F33m+P3o53tulFIxd4fkbrVF
wpFSod9UZHoN6nooVbaJB0Q720bqAxQGo44fetXDpYfH7/mU2rx7ZtvEJFt7xphRhowwdkgDKCtm
hY6dRsHUgb2E7hab9k5HiTgAAO089FKnav5/WLub6YRTmLIJG4kYXOtsXykqrGO2S9f1NGZp77oA
8/B4nZyOv8hw+ozR0bHIZDT+hBhJye+JKBwj8w6Oj7nx3lsOfQtNfMxaKbvL249kBqd+ohAIMicT
nanV53EfTZ9EU4RZIxCQ8/1ukZOlN5Evs+Z4udqOOHBrARdP0h6WBrPOZvW2rgbuPClbRP/It+MS
oCAYFLQaWF9dzCzDtqFmzhR4dOrc4xQVYtEdfLOH4+fKXaLTpzsrMC6KRzhw4kry5ZbgGqsh/6BG
OJeuSZFSJ8NFj/vki24uf7Y/LIaEGAx32FFQPhyvhxYxl8lXUrqvYD8UgvaVA4upnrkUFJRyVT/W
S5OIEnACjQUWPWlsEngsRMzDi0kMNHRz2nwyo0kffSH2e+MFa6x753QAPOV/I1NbAnE8Gfr8R8xt
0g3y1T58pNloT6wn3uPDwnFEtnDCYvaENWrxEFuYXs/vcKVQFxHJTAjGN6BK7cNA5d8S/y7ThhYK
EAQiYdUvehDE+JKQQ/lecWrBspnzLHlltJWQQ17uiFYpzXceiOvu/wvZNbWY1Wm5tn2/7CsqSOof
l/WhYqIcrkMZh31FSDN1YKg0BTzNWSKWoxCAAHpeZ78+/uMVnRiG85tPSGJ5jDeblol/u2DTMSlW
Z+COcpAfPzng/zypR6FZGL6kW//RgKjsdkALZPIJ5wrOPC5VaNnPgSJT+ejopGoGIqdKwpYhqgs8
lAV4BGKeumRNaNJr23kbQFrGDWFJlJqHO7Qw92S7PSnRoSS0HGR7QIsNbWlbghbpaJ2/8o7MnnfN
bNcts4xMpjWx+By3wGdm7zIHBmzbTmlw0elBmQKkudszFk/VZraVMns0RBhcZRkPp+LVJyAgP6Zm
WFbew0e+ycOvwS608cF8X5PFNXSE1d76B4ERJs0VNrcTIuMXNofSPoM/dgbliDk82tlOsGqOyKyP
59G2lZT9rPhhEb0l/kHggwXhUExpGbiEuG780tJAb3unzxcUYDa1StCnCEKO/OInJbopMF9TTkXF
xAJ32pD6XM/+iAF3fUrFZ9QMoiGAq8DQ7MWWSoe1MagQlUdbLlN1Rnpc1ETsyp9ZGi1BIH96fy2+
FWDdnHbgDMLiGQpyaeaHbYD+NEh3xYrRElryXN1uaJVgpVGquPaWy/Ov08SmzedawCWmPujx/zYA
dLq9iNYU2fgGIA8+Yr+x4Z501kxHcAFpTJqioH5RfYHyxOi5OkFjEhKjfRNwRTgCqZs5HimE7/eD
cSMz5HvXjjC6eE07sY3cnsL+ysmbaoQniiuDzsCUm6Lw5wCo6FSxTEx1OiRnEFS2GdDiCaqsh7hx
TnUdC62JPq6ETWbs5y29l5nG91I5w0RmkTX8SG80yCOSHDzlStfxlf+pAusCvPdD+jrGjxVSSA8d
QF6ZgXYmugdJtJy/uLAfjLMFhht5Jwk+GG1snMYa0Qbj5nxF78QzebYawb/pKWwjBPArNwQPHFEx
+08LliF9iy9MhHeZJHN0EOAef+b/dKxZc9UzC7uf/pCndtvSIYhA1gUcp6AeoNgITKAFJQSkCmp7
WbtEPZS0Zj7Ln47Ysk1ZVT7uz06IzsH+fW3mvVbHoghi6dpVjIF6yYUGqAA2fXS61ge8+PTm/EzD
GpuTmuMl1eeGpxgTBkpbel/OANmSfE3N846k6u5jopKJ9D/ECPfcbU+zx5CkEji6SG5wLKs/iCTP
LaMy0zA9E6F6d2OGs0RhuKUPInQR6VjL8xWW/tB3kY2aB2o+rydRRneTyl+g33URezhIgbP4FtGg
z+7C9VI7NIZRUd2/ET5qVaHWSytZ7322Q64ImIQuqwDzTZtDeGR2o2Uyv9xOoXZZAT6120VaBJCh
gWQV1jCVtb2Qu8XnTliRfqf/QT92ZjOEH3Rzgu6My3ioy2CSBjTaGgijk2i8/PlDqrrR8LyIGTqO
G2ZvRqvO9ZsOZJLHD868Sr3o55lRmvsIqd27EYp74LUjDMYYLm3ZzV4HmdpK3cEEpk7L7ZTN/6Pa
/9iEHWK78P8vev/6wj52u+OiEHAVMlhSpx4+CDzB1KxQ/2oJeDARVNAW+MGFrrf+UAV9eaOfRHg0
HyPHq87XWyGU6f8xDPZtHu1q65/jcBvZ7Fma0bdNyHJJeeHJcrY+AARUGddDazVu+u/b8JRhUAkd
mh6c6MiKeomTwwsTcCkDIhv4eKY8nOsuzAA/ykYNjVYKbWOtDcq2VKMKFYnKiJFPkfX413yz1uxR
u9bjIwyVc+D/xp0qM1bsEAIRV2ii+ZOzfo2WhchqjU2vtQWntFTaXhnfVPN8tYd5Koy86+5xLoqE
uQXbLDw4QQMGF0IIT8gcw20kGttj95lJyeGaDNwm/3FFY8M5sQ12DVn/fmzDS2mw7/wnrRLMs7m9
LuET+DYRlJtXfxToeau45IJ8+XDKOXXiJEptit3pD5tx6f/DkUgq5Aczf56bFjxUa+g/E6Pfcr5Z
EgcRWIe5kD7ACUnO7taO5OvL9dBoF4sWNZ5xK1o5HdUC2dE5b865PVRGCrczzAtejafJBdH9AHeQ
MLGxsoXqfhutUSNsroBOiL2NOrxKbl51lDNhl+vSVBeaz3L3wmjr8auTlQRYumZi+JYqarB5HYFd
y4LBHv3ba54oP/4lUkW68KXr359PcPVWXA0JZ7VsJqB4S0/pX+IKe5R0xDOTpbbODocnREvsH8ii
RLFcpMfjFcuSrn7qLYghndPwU/JJ5mj/BF3BifR0Q+pVQ/oCFnYDmJCskwFOYcHv2tvXTN1Syo6T
lyfBB8dFy9D2pLA07qg1wNgfjV/OQ+6uvcjDWL5lF+mr/5gSm30BWnzNNxvSIl6Emo5ked3AF7jX
a3gfVVRz1OWL+a3PFZbGAcHqDuqpwDyt/S1fKRyZGPHPfTGuUTTTiZZXSVi/AeOZXxnYg8RlsgNT
x+rnCc3G7U/U/LjaBXa4FOqm6vRmxvMA78f6az6IBwK7E1yamarsCtA55NWqYBMmDgwARpu5A+Vn
3fX3MumPBOwObv7zMXTmOZrn70wHOZPYdAjLMyh278vKHjkkzSqGLnolUZzAF0pf/ZnvL3/fS7gW
03b4CMQccudpuN+CjFP1PacJn2uF5gHsreWeKtwQ2en512vIk4yqC5Zl4q2OcuCW82NkYQix/coa
w7qxs/oDYFo4fMI79A9Sgx8fyzKm2ZSTGHoU6wpxAlltXk2gNiwiQMMWz6vAZD3EmCYGWvLg14H/
s/GzORfzuLVzCGjtpWwVdOaYFW6xqrv3+PkaHcHfSmgdk1Fo/+dw8qIi1MM2adyFIjSo/Gw4vQmp
twS3DE18tp6294d2zVTAM9EkwTKCeNKveMeQm4dsOkF3cU1yPxunxhjR8IBkInXMTp2tcl6UwaJQ
EkT9mqEJHg6v+QpOYx2s4TBdMGtTmb0Pbp5CZNl0iFrwzG+HFd72TjxXUxrOqktiKgnfCD1F5wD7
rlXSpFdWwgtP2dsntKMh2So7LgtzBClS91EKqkWCStUzVVrh2kcB+Wu0vuEka3IsVfmJteBSKD1n
8R9e+wWwgQ/9u9v6X1qih7N8maeHPckx9/URoJ3BGTuE5AEE7+JWIp6VdDruLcRTalSeMQ7bqox/
6+URn3nuApCBksQUZuCmQkqV14qWBAlE/HTPHRns+rA2NapMA6psEW2yzenct4nGA2K6yHU64VPC
Sy03dftkdO+fhsn07m5fxwGCYAgovEql22xpg7XUd1UlsJ+virnnPkmRKG2JAUtqLlIw+HL0/7KL
Q8ygwUVvwalXygOmI1xF9Kj+w5wudANhJxDUb0s8kkN19gOW4uvLfdQ/kvt4qVOWxO5tYdZD9nlz
vPBSb0DE9lNcdRk2gBRz2Sx5ei0Em7PZCYIgQUrUbLT/g+ES3dh04V7pwN5l6GkO//5Bzla0j3wt
wNgvPEVQatS06Wxe/iqXknUEF1mS7clGnLz1rFf4TF13sps2EfmbmsNllTMkZ6NVlIP64KpbgrA+
yRXZzIvFaEsR1PsmOKdHnVFIFzE4Ax7glt34ZRQipV3iATgmSgDvsQJnB+tPL3MWNReuhMte7maM
bfJBhBqsk22GyqSoAnZYvZtYg9UWR+DaLsakFbIkil3D9P4E0dODtS5OeEfZVfj+qQTOOLWcgqXi
bc4/2QcjSpKaXHAqZJUdl1bQ1hOGbJG8wjiYvvUfCyv4ASSt9XdA9dZrhmdEz7v6YmTaxME+KUF1
Uk/OaJJSoYFDkm1dH/fLK1BfPChtGQwGX47V49gRGt6BBESktf7qX24hdH8XM+l77PHxPn6/aJKS
fMcNTnsTfNmSe+3V26LUGgK4xSLNqdWPxtTVsDpM5k7aXI6gTCiTbAYmn460t0cxTXeUBXOpt/qn
npvW58cX/MDYDyaOuEjYm6I/zfaZTV4hBjT222RzB3NYb9SCqY+lSW00w9xGn51S7JImDjFutE1S
53qC9btTEOuxtNGsu6/wKqpbMwxLVRQDj3w1X5tEnLiuiBDY4W/ejzxk4J/oL3kIA6759oLNIdVS
PzVoZpRXvMM1kSKUWTVTqTVJY/GLOimaAHDyhjxREi+IHbha8AGDONuPkKCgzbbTE3iOOcOAYrg7
LISKbqPswoyFAlUODLCFQXPkSo1zjuFfGoKdKcTuFsG2Ltz6YqA+dh+ia8UGFcuf8/dmZq08VIsx
go3Zaibvc0Ru4+WkS9aBq8t94K3OTTtefwoPeS2dxLGEySkSF+J/e2j/o0Q1CW+CXEhdKL1xlkAG
5meaQP+j0U4HypABQ+1W5g1am6odFGrn9lFx5K1mw0BrYMytBGCARyScacE4xx6f/S6RGD1uoqF+
V1KCp5hYLeISKpeuNu7ff5VkPLYlz/rQQYcQIHZUfCMGsJ/rqV1B9Tw/s1TbT8jji/RqzFFbAN4+
NOiWU4CSXKJ6wXFNz9FJOHsB3esRlt3jwOLwDXB6aV/+7juRUO7UEuZrlreDwUG0lsYK4L6ZFWGA
4VDSV8oLdUTpfhowsa3G7B4KFXAHMZ0JmbZOoY7hz2W8DMs9u5vYdwJNMW67IIygN6s+JEYtoTP5
GZIe33tIqO0k3HMQ7/sLkjIJToRKmcVsULoInB5wnSZBjGGvLgm2/iHogltuWGpMcTBoONYdvlcJ
brucSqWJjx8ycyeZQL9ZwG7hsxI9yCPvoqgVBtPbT0OXxvORUxbjRB5LHXsPm2E/ybSkmK35hHEI
sdnEzt9RlvqQF7YqKsMIHyP0d1QThy28tMrIlpeRkx2MiYy9k6Oz3UeWXajaD2RRoJqCkVVRbv9m
m8zEU/RFfUHkK6iDuHP0DLOyAZEIe2KUXwY8vyxp76B/izF0j4GaKkxrdc/x/GpblKaFytL6GIsY
+PyjqM7m2x93W43ZB2v8/+a9wZTIAi/ukgHy1Vdt/WwYxbCGLn6s0NtrPRkNc6N4br/WHGnz7FSG
UYutLcodt0WUxK7A5JGipIwjEFTh1TEBEhBWwvkGJFSmsVLoKGxFLa3d13dC48Ob3Gh6cCuSVWTS
BL8aEIlCBvLRDdhtHugi3G8ADaESarfjCtprUTRxT8vni2QkuDc5C2TJ7amClcjqCixEpX1JHlC7
VvAsk4G4zQ9fNcICuj6RfsQzfn5dOnN0+cC1W4aA2oBA++DeOu4foP3AuMp7QzUfwYivyv6E8NqJ
5WpPIKcmwgbOJUt08eWbIW+NNvBuc/JGHTt09RSGbZfFKAmsyQVmZq9sUvuF7Le66FhKe636s7/j
DEHxNMbl7J6FaSVl4Nrr7MmqyF0Zq+2N4uZr5o9K7wLDVZWOw67PaxUp2PcP1HD32jnhJaoR4pHE
Lk8coyShlkKG3kXGEqodFAy236ySkozW93FatntZsP5hlItpOk19bXx8ldfLJ17Utr0uavFc/7o/
BufxHBg/ggSbJHajVTKWvvFMIQ9V+FboyvF5M3jkDgM/vQGH2mg1v3epGtqRQ7j+UHSxtdBohkE6
58yFnIxqyTI6r06gQMhuOFUV8mZU7c0tMXuaTosI81RW7HetisMWvxGi7tx8sH69N772X+39QMpq
pbV6p+bx88LrUEawApJtaetkZYGp5rwPeWQ/KuY9yBaDCEkS+SV4V1+PDOSyepyJATx8iD4OZ74v
deLOVB8esUi0DSZIJPM8GdgpnoWvMTF0QVKZskALtq1o5UqpgH8KtQ5krwl7oR1xsZ3LNbU7fmC0
btxe254u8GzMZ1+gwvaBUhazS2y6NLyNJ1ysXNYTPkA/zk3xw0VeNZ6B7Lz92yxqJo6Az/lxZ8sE
Srt7q2aQD45s2p9LHZCxwB+q1qYafXbgnwc+4sLiKuG328MyTvLZCE1qfxQ60sB/00PDdgFivt51
nqmlZfNlWkIr3sdne8jLBvDV5Dxw8oQAVceSkqlIL6VlRTFrt8/Vnjhb1+CsX/xY7BaE4GShgLNE
0RBxznjO7Ji13M7SHYTbz24YiAbB47l4zS9xuygVMWdRyRTHXHLhv+69a4QJOGPJ6cyB4DUD9ddz
z7XAjn+7ZZE6kMmHBHEShDcPR5leehv6qzdvHX/mqWzu3GnpD3IVlIL8sFBvLQcHGgC2HQ1D2/j+
oudIFK2H0MxYxaFyUw+wh2m0z178+4Y4abbpvBt91twFuswcMPqd7oTdGD250YIMlvMhIcB66hd5
ybOF4rGAiKjqvpkqyeVqlPDR07xLH6ypVhdfFff5LxD2UaDfke1O9x1n6sMeGqb4V1rnMumBfU68
0qel4byipHtTwS/qS9zgMPn32pTbRnM4x6U6AI804b6f2FQKh/pNs//k7Aboo++fgcaCwzIJrZGk
0Z/aHyOa0DubDZwC7tdMMXO+7yzSeLGybxe9C/J0UuwqgS0aMNO9ZGfIK3zaKFjm60/A/JUOdkuO
yhUtx9md6U7htH5daFDtRpt0Sqvi4SkceLH4qQwTouBrz6WE2RFj3qalZhplVksRB7ixmalJzuVf
FtHMfSXRxtqqcGBGqehDkjZJ1FLbwbvEWjOdU9R3BPkPp+FtAVibHGUqA+UwGy25hjWuMKC8K4kl
RaAVd8mdC9Bhxk2rnIJQ3vny8Jgv78a8YFqGJlTGTwi/+kuEY3s+xrRLtCHN3NP/u3Jz34ArhEMC
PwhKY55ZFFuKmXVYH0DCQwdQe/fmecn/eDP+7haVAjxCIPIlRh28BVkeMFSqPEMGytTpX45woX51
qWGFgKKq7J2NB9RefeHgwyU9CjpP57UJNzXUPs7qfi/6DLvbcq7nGSDtIB3pqhvl9S+wWH/ByTNi
y8mwvcrBy6QHd1+jj5V0gkppk01MdFRE82TBC1wIGlQ4vK2V9hVjndGnRaPWxgcbj0VIFlCWUo9f
vOcESBdDSFdmyMIaoTUna+RVn/4pbrnjKVp8Dzbhe+pwTIWcsEtv2dUNZPqFynnoEC81lrxlp5u+
2pzEShQaciiTqexlK+SCxqceDVwXE871Kgxy8QtMsdUuQNGA6AQ5Q0/D1LSr+a9QKLB/Kfuh56uA
CZvL1kxgZ7X1CrnI4r87XCkbbaaj9jPeOUDMPNiasSJtwzQ+7ZcSB031KvbLgrWBvx14Sb3PBTSw
Vcw4ZNabAPOP0Nq08erA0ITXJVPLCsqM47WCTa+azHZwKvrdcho+NiUWjf40WS/b7p060JReRb1E
Uz8eISZ8ITRrYJGtVjYZYUyJiZqkRKg2Dbk0lmQPS9W6SMVwoz1XaAHRBvzeqZfZQydi477cayi9
AT9+6zRE8pIowqVpaECO49ZGBva1DZjtZzMBLTepSdOF4OQvpBxH1CyWQN7hSnU7mvbq7NX54zg0
t+Z59i1vBiCKKm0safaoz9nKKR2WHnkTiSjMScDJTa8BTb044PLLB7CvdUkdzgTSJmJDoDZbGtZv
IpzXjCaQkJyaiUtlqGVJsIe11KKnRaqCzMxEB5rO7fPiz5RzL2PFXZzMiJc6EdxHBz2En8Xb7cjz
ca5blBiAqcTFG4IxiREeOV/zDKH38hpHyKKOodpEKP4iGaObS2E7iT3GedyZqAzEIK2713SU5eoZ
qR2pNx5x6OgPTmr6YaC5C72x4qm1gr8s6p+7Oq5+t8fHuz+LhjVXRzwZnlEpNpb6SLToRcC1WcjZ
pxuAxIdnwu/EfJMvxhanSIulTamSxkYcAkFc70DZ/6xpURSXRILQdW42AvdTY8Gmxw3qPjMVWFhC
uhyHuAJ54+WZppC5osVdEaKa5bi8IJdI7kTog4p61NIWSPQpq5IgNCrzwTX2iIko4ziu6XZkzerh
dMP43pJsXUp/Rpo35J6lTO8qEs6Ps7T0pVObNvoVfkkgat6nf0AaW3NX1M6QwFU2w7mN/OlWN07y
mN9rsZf+N9vDdX/jH3iHgnm/3XlwOOfkkmP0LP2DwUBnDH4k+X21K+pJis19UP/02MxgDvBeASg1
bb5BB6VLKBklAQN4eSF5QrDDJULhSOACGitLAHDcEXlr08NbgjwymbdTAmlmJ+xSgkF/Ggi/4JpH
fkCpY3Wc1659gZkzlB3CKxGTYm0QZstRJV4klluVZDjO+drZiDABBl1PTiPNHJVAFUB1lGDf7Zun
rK4Y9bzjAp+HIkZWfDiFgiOM7yKPD9PylqOm92H3t8jmw9Fx5ig3OKUI4MuJpi9rMeVUbq+WZBl+
1p9bPJtBSNT3pXD6Sii7ip/O2vCZPmfVTakFIVhtqNkhd3Rc9QQzuQvgwDp29v2YmZKkusUSY6Ii
BeJrxbdilf05QEJlNv8THaMZN4g1Vv9dgIGN2x1mepVszicenqImUA/2qR/ts5PQHICFIpPAJbQN
gp1eeDH/sbyjHdTi5b3uQbFi4pKPhkNLronq+u/v4B++ZQkPehWvIMZLqR3UwwC8AH/61/p4oDHK
3c9TFCbJLtZ5+cVItdG/o9wMGnLNB6aC+W2HehtaBCc7ee6B2r3yxMsjr14cbvO/2NvKR4XFoI1e
4XZ4Rt6gDSU6jlaPI3nzf4K4aJEELXbITLwmoINC4+bnbvFSub/jYffo6GtYDtuC0dcgHp9DWYtq
JwBH7XJmULEPk9/3BEC3NDl3w/1dAK9V1KCdTXwIJpsIgOnevG6wopgaRntL2+0Etp6Du92erowJ
AuXoe+1hmeDZHwxFwfQrw5tMks5JFL2iRsnOyfU5/OjlJL3TnLUNmy994Y6KGkgispIOKciR1T2H
E9HLqwIz1M/1ReaYKRDYec/rk8p+nT/Sdmwj528yvMQcc6EGDeYTDUguni7Af+t0ADlaajC/nxNk
Bdwv7sQuQiaeZWrXqyrsidXj6pCk6fds7x4fSpLQG7+PfthYTWcgGCcc1GvbCzzr4sYY7BqY7gVb
k4rZ9MfpJ3lN1PYx4orRTdDZzmWAydeFtahzQLgyKD8bpYUVwR4pVSmMWaDwSPoZc1NAZoMZnM9R
AqGj3Zg4Q49dqL7rDjYW+8Sa3XTQr5ugJ7RB+M0ONuB2Hce1VbXc8pAPcTqsHkGVOq3cL0LxUPp3
63SM41hyzjwvOH1BvRhM66HLoDFrV6A93roZPgD+sHpD5esUCF7bXcpJlYlNgoOhLvbSHBH8mcIG
xfcUVdtrLi6AuKdSJ1O/ieECDUI2HXUM2MtfANvFBSleL63bOLEiIoME7NLX+59Vpl7SGisg2wW3
iT93L159CXrmnOMipKuZaxgjk62Hcy62JNUYtC8/OmHqRuXWhrYx98AHcvUVF/XpzyJlk5e0oXub
gxXJKisBm7ouEiUIVdMfcdVzs4IUNNWpFnWSS8EIFm9bWvFlmd4WZtZ6GMbUgOxOCpZbr2AhRNCw
oBOJ6WseYAJ1iPoGaf+Wtnvs5Dzv+sCu1YGV9haCYvhEld8l3vHbQsDf4ObZR2jHaQVkzrWIZlAH
9aopqMKDQ7Fq9pnsbspiB3/Q75pXrwcuwkMSnN6WjUva8Bql5EL9UajGQa+MRNfJfG800aJwYIS+
u9WH+Rkqszvw2VDlcDpnTo3xKrJWfXV8jHyCap9kjaVj+rXBTBGu5QW9Yg1+G5FUjbS7pk1jpJiA
Y8qLzzpxSTAWHshiwguEBpm98brGmadAM+5j/sUf02mjmAo1DzLeeD57m6X8YJ7LFoLnuy5hCJ2t
5ksyDGDUmVx4RyMKTfJgL6u9SvnziYMemS0ZIdDz0Hv36dyTHaBvFaDUL82WzTABYXnjNyDTyHXy
8dzTtj3ZkoG1KjTqfDxi/edd8uBSx2Az/x4x1wBC22shaz9g0Vwv1XLcwCH79klchFCSBcnVMinx
DRYRkH5AnTzkiiAo/a36sNGo00ZvAaL+cfQMjw3LBGsV7w7hFnzqDLuxAFBdnEyGZ4TF5+xp5LYD
etmzjhPEqRYByDoY/xQqnfGyb9/nrm2o2XlwSKnIJu2DlW+sVE4+/gMXKvPn1898iyYTkbjXBwxb
CRuNDnTLZPB1eqm5OLKtQwVjChHWGFOMFfnLiRNx0mnGLn7pBldpBiQ9Rv8ljps5z6FYxTAGKQ8Y
b3dnwM/S9A3kSKK6iuLUmEE0xQk0CEdpgOzz0gPP4MeGkC/xzbdtXUvbfHc79mbkzSMBrz1gsGyH
QOD4VtMIIKriHtuv4ujZ9e48cky4HesDNb2lGoEcjtSZ+IxAudJsyfYzlevWe1n94qSeb/Jz//Pi
5pXIcK1KvlqRE56AN/94YWX4w/yE5ZLisxxUimC9L7cvKJT3Dgep3ic7W7kSxJovnHPVBReDeBuA
YdLiXPdUH5/X9MbuwxH65d0/GcPXpH9yqN3Q+p7l3Qud84F5Ow2zjzG8E0dGvudBFIoNFxPpZzAD
HrCfZ1f5l3uLfSpubWZ6Zk42pVrZ1513G7Csp5MUJVWInMLeOYC6beTrxO+pv0AMVAfETgpoYyY4
dq3DkTsY6MG/gD9v6apuLLEg7ufmfAtZyoFqamuRBBpL/a0YVVhA17Wc46AXHZjqfVgmDeOzO9ME
0Kj5iqoUsjfPGnySYeUhF9hH2jDXgd1PiqzgeG4urbJzOH61a/RcOq/MwqIpvpsedTVbE82ETt52
s5srVbJ+h98JV0PwMxi1bLy5+O8M/uRr7Ru1I7IcJMHs7FR2o7YeHLnmmAyTR9OV4cEHN/+OPUMH
T0924Wj63LYzssOesU79UdtDt21SGhdQ0IS/FPgsOsOcoqgYBeLUov4XEmDHb5u3qLf5kjtI/te0
34ZOHeeGqG5cN9jA+8vltivKQ64+o5qSawpuEyOm4ulevyjMuYiaZkkMF1P4ysDAoFplyXuwA+Yt
XTkOrB1LSuClR7u334AYW05GmLSGYVi6u/znSStBAUoS2DwQdJnE4rRKFkUVxEwRBjnkkdZa2bvv
pZBiAAixWVFuGQzFJRosriB3yQZ+sZ+aBsDpDNvca1yOLDcOh825bvV2vzlYeuTiGv0gjB7TEVdF
+c1Joy/bVJiKsNxJsEwbUduGjFp71rIpD2Wdvc9UJQIZVNfmMcCy5Kwfabp3h1tGGvqMjuPqtz3r
AOjJD6uC5WPs7NpWz5ezsW55Efak5ISA1PvbvVH7S2Emf3j269ZlabPL/DPVej9aAD7wzi/59FyU
5TbvwdNNgvyFYxi4qh9nyrlAAEBjd1lEok7sI4Ad5fCM8Zb2NgksNj3RNcuqUItQwNuo5yykhRAZ
lhkMDNwKb4Sb9TfBSsyUiRGS2XjBUqw6Hjna0+UZOoqsQWzIJcGK/f6GT8uEvsX3EStSTqvaFrst
orju2NYl60iEov5INhy/eRmItQ9UWaxqSTAkPhLUZbRRwqL1Z3jJYbeU68q5QAWAcyLNi4oC+wql
McnxXxJ/4Pe9EnCP6vdTBUumViI36fyn18Htu35JkHECtdhfqRiwfL4lVSPyyUzoHT7a/elVHzL0
I7+gaaCosRLzzzOTqd8c3bFJmFAn5jJB9ahmfnfUhJiu7/jqug3dDk5Uug7xKMOTUU9MCzpYfDNo
16ifXRAMPfglm/tByPYIbYfD098pgLvtn0+p7UrJ9U1bw+RaxE7kftq3Wy77KYS6gp+US8FC8m72
qxmG5M7vOVSvHVlR1pYJ++TJTM+JogKSF9I+mzbLnhN+aV1pytJquEmKy/nkjbBMd5P57NyPS9Yr
BhL+1wOUOadnOItIFqX888yS4/f4S+SDhdaqsSdvATNO18JIxazC+ZtUsdhsE5kT/+37A6SVm+/A
7ID/TlfJWn934A9MeGcHBZcOvVcV3OaKfPDTEvbBPmWJy3ImDFd3hyJ2JBH7j8ys529dPoIObKWN
HQ8J6sttV1XNbNc4n/c+6byYVGq8624dzY7luVhPFyWMxSVMI7r3CL4Us098iYNZ9afH0ij7XVod
B57ztLlXm0rBbmTwg9JY9Fx9wZWLP78ebh5AzlrBiNdl4lG9ULBvvF4fp8CP73VBuYj/3kbN3FKw
RtRZ6IPeBesolN2D8cvBPyPEdz0cb08qVl6Hd3a2GQ0FMrkWbgNd2SKA04LS1MINWpr+XiT7aCy9
jSz71s8cq0Q/DKL2TezTPiiOlQDhpIOZpuCARA8UTB4FNc228WHkK7XNrivqH6Q6m1wF12PeDXL4
pD12UbQgtBlKeguOb3G47jA7zclqAZARLcMkAA/wbqZthmA0dprUbZF/0oh/685D9AqtLC1Gwe4J
hhzAj0ab/cd96I8YSBzgI/OyhmDMmKH7HEGjejx3jly1FYk08eLCPNzbmwKSo5L/z/catSL1+2Us
lenKecEebDs5GFw2tH6LQ02R5MIMm6TJ7ApQuTpGyO9mK1ZSCHTaXUzqSqsuASzHtOtLudKAFL1/
2pLPqjuHhtSaO+uTI+8fxAArpB0wM4E6DB5AJeRponfZYcUJbW4U1sCQeodcRZ2pKe7ZEAowaXRf
tB1MP0KM8LnWmjWBZIUPIqFv9dbF5M00XGAe2yFa4mUhSwqyuJcYfLIGb81BwAQG6BbqLCpUgC0A
WLluSWb2VYW/8MbMdkv0isFYFt2dM6z+LFclxI/CA45lrmSybgCeGYaL9gw6I2+HlLd84RcMv1bW
/0smEquFyrtGiI6BdTr/5dXYdCWq7DuYb1iUj6THe5qxnleoHOn0wF2iIpAWTPMy3RwbUpG6dNr7
hykNOe7N99cIe+ZRGKlNsxG7myUg4zeCgxRetisz4j2VHCbiEVNnD5Qx/8Z3Sl06i140qyeKb1w7
LDbpRpjq5pmzgBpYN2Aec5tgnD9FBc2nLIHZu73i1h61kGbWdzARemZjEKFob3hdPzRifLMMUlKR
7neHh8ChkSXTYNj0RJgPSWcznrMXIaSifKgZc8pXwa2HtbRZ+u7DGfeh34fWxVIcOo7BhKX2mdtM
v2ZJ/psSlcYGT8Ogpf+RfpUntr+YSb3rO+pZV/q4Yr17SgpSKvTKAQxa3W3LJGugJp5ToR8pmLSZ
8aRrFIb52VeklJjZlc4ktNDCHAGB4uyPnTKudZkk6xJFd1O3i0aroEupvhiCLRr1hV5NKjPehBGJ
/JQNqOZ5jVlsisVH/0WpQj8OeTWxues9zxQHzH52w8qpZEYqspAbRAi3OQBj/4RGPJuHh2hkEJAs
tYDfqxFbygkZKe3BUJRU/0IVQJ3Om24vhpCp0HdzGXWl7pMwiU5XVvoiQ6zc7ucV+SHSk2lag6eG
4Kp9D+Fiuh4RadfWLvzE+H81MTPRS26J5hP6+gNeOCIBF7DgSyGgppjFLty9Wcc3PUhyzKaKHClR
7g6ZF8aCsmAu9GyIbZ2QgLrai9rEHXxJoDKYU5N017548ggQ36ig27fTXPi4HqLH+eHxgLhdTXXm
f/XBX3xVVoFnpn76YHlgt3MeUYQHwaJ+2oCU3RVe7Vya1pS+/TBDq4pwbHRPqH2Sih7KgkdEwaCy
hySJDWlZn6NJAEyBBv9BavMu1KL77u5fGzQ3Neh1seBqLcfocsDPbbNfC74Bzjxk6HYMbJBWarQK
OWhVvEXZZJ2aYrayp+iJtY3agu/fJuKNphRMdifLw9oHpX6mUFgCyruAJ1G8E/zPUvwSsdjNYyAc
kgBzVwQ/UqAjIJHYVnChp60fPd/tUHP4TYoQfxoqi27uzLlHLPf9jRdfjc8vYBQoFH/gA8brbOKl
OVPF3eBDVM4yt3gkzKv67rNK592e/kS4l4J++fhxgznI3KuiHxlmNWTtntxf/+lDUXxnmLD9CElt
OkaGiNvTnK8FYp56ZengXm0VJcxehaNCjv7DhZevLJ5Aviu332aqX+McqVVtyeRXIqyA+deRf3Py
GCYqsaBcwBzCLVceIGH9K1y9hT4bsQ7v9jiqDg8Rx5w8PJETVFrbyv9n8jpVyWTrUIf4LCqFUz/6
pgjN/6KfS9T6sy4euBzNQ1bKzpDHhg9CepTLmGL8VfzYBi3CxtNGOX8TlkhtACJMbboXmocVGYsD
XCTq92WD/wPgw04MtgIMnZ8M96KImTR33zci/dzkl6OkbEDmIj96T3SysrQbouPKGiY3XTIm+M56
pJSGgIRvnYdrGZHLx15n+XMaAdP/eRiZjipXAh7cEhb+O/v0C1lK/vdrM1z5CB1wU62Hq+nn5Wu4
pxu5dS3UknZfxlm915xdNo7MQUfYbtTkGWqOZPTSfTWv2hPxp8DuVqCB52jUcDxTdBjeipH10BAz
UweHGCmBCewzsPQhvAY8eD+OrBxVozJ3VzRsM9/A0EDgDBueiN27xfuuT7gihavkMI6q4cLkE8OX
IY/ViHvLz+Hnt6XtAsgBcCU6QqvG6PnynApalE/P90aFY2h5q/dMH+pbxUqZ29pbm9hXlqs9J5sP
KkwcdHwjKeR7YelWjNzGb5JbKG8OXvvYQLKyxhUisXBocNkn2gs1Mdi9Gwd+Z0QoNK8prZS3gPIU
qiJExBb6f99EKp0H5kWjO50ax2FEe/hCUONyLQS76cOUWMuNWtm0j2iQFIk3OKgRqTgf2KVlZazz
yqJYkyaA9iVzI3Et6twSNAGlmqRpQHr1RxmI6yh3fDlEdKVUdtROaxaRzkSXqCv0DaBx7wcPEHMs
sjvc85B0JaNCythFvEWkPGYoMCqyYwySK42eFADOdvsCMHcYdaJC/UjbriKrx1yUjPpJ7yT1hNLo
Yoi5ss9H/jhEKnVMuFW1dC4z5+3rJdN7B8KO5/ocFpP0NbcC2MkSK0eLZ93arMAVhg4TsVQFF/ce
4tLPn4jouJ1o23MXYD8RcHLRtSz/I+AzrmtuQnkpQIltzWTq9cqjI9v82HwUOOCieWl5tNhNCuC2
vY1Fwkyri0GyQYVRbxwGjRi6bRHwM7hWZT1FEsCwX1EDC/bNLxlXTN6UapvpYonDwFuos/b0+bzA
qiGHYEKo6Rc63QtU+lVJhfcdNtn0YJhyc6SLVawhTE1sor83PANnSZZ/V8US1PXf4TAgWkhcBsr4
3hN2AT4znqV8OMkkilJDMmfYKuT+jiSxPanhYgVra5IF/tY1C44pzIu6EJ2uImP+MvaHiQxWcSOv
M/XiQL60VnQ8HIlvwHTgQn1G6ruUqSut0f+ySc7uI1XTvf5YV6aLIuDcWmU3em3do+HZLBJeXNdM
qLxkb0fqoV9JCbTw0Ncu1BlpZnbVL6VyU1MNkc5/5ccGt0RcourmjkcgCKRvu77DaMNVd2pYQ1rp
X7IUqZmYQUwNkRAu3CyuR9KJ7c3j1mPRDqUM6eZQjozlp1dGYIEq6dY9hDFtZWjrm2hxXp5Xsa2V
WhvB63X8wP62HVM2sXjoRWSHnC2v+owVj/hbB3Yzu7SHrNOHft7u/gaHHgHj7Y7MCus+zKMayFMF
wkMAdnMl+gL2i+SW0ROPsoZgsQnmSDSzdUCNneaGeZsqRilXU+dp+4fKaPZpNozPf3T56WNbdpE1
B3YHt1qUo9JDqwew7Zq7JneN6l5Akiry9koBNI1fpmL+ymm3WhjKq2ZlVLJrlNz+KLeuBe2nCR7u
7pa3btA3H9d89gG2gcngdhc70IVKCWxnJFIKCnTExU7OnoYmTTggvC2HF3MoX86owI0rNk2DiM6N
EzyIvKpui/6tP/vMKrzJyvY3adtNL7StO36h8VXP1F2Rq6KrAuheozRp36vIdBFFWHZ521o2mYzR
WqKZeJt+lSnKC0IfcZWlzKNV6cNNLE2AmM15H5WDALuix7HIerKCVxcimEQDYsrJXaFBU61anJha
EXFTuSOyizaPQ8sFOExWurPZjzxIWgo4XG03irBokQtGKRtpBgJRz7pzGlZnSOUZ+LaPQf2RcvU0
WyZ/grkOxEhto5/hot92N5NVgSxf9lfpg6IpquVOc7vPVovbBRQ45jThMdJdvrXJeb9eY+cCptNx
6lKoVLjEZamarOsI+1JO2m4kXmrwos5ivu9G5ya2bR3qYcevVdd/zkgvIs2dGHi6DUtGNbSwTshT
+EnCoZaO2wRBnjwqR/dg/qkaUeVhJs7sI8SdLrL7C7LZb2s1PhDbr9CjJeAenYa7KTFgX2+ErXGw
SN/MvprYdhAeXdSTgcxC7lMyoNfEIJJJjDPbEO8IauLf69sN4iOfUBxd2RUWKNNkNMYOIBG4PpjN
nZrvZ6k/8bALkaUE53Ay75uc9vaOgilwkzbBiyoK+dWawV/t0bbRgbb1TdlbmzegaoA2qWI4Kl9z
Dv/SpTZjdIP3DNSu4rq8w/C1JKrxACdxYRL537JHoVsPUPSBMyH/BOawdicCdUlg8IPdsfdOS+hl
IFpVVyBj0/q6hcGGjn0dfh+tqJZA10cKn9OK17XUNpBMP5OG2ql8EgkatW42HIPEKCSEpL0LeEsc
v0g2KbX8Dv6schdwRa1Q5ZixgNlhhGWQhghcr2R8Ygx9Juq5RoF1JUAE2AvCtvI1AgP6LZVcRVN/
5+V9huo5RGrzq3gj1Bg+Wln2Yn86f1+kSfBB/kVkH4YrBdDTICT/XgcCga5LoYwNTQvjKWaDbmH/
JbdkLWQy7VKI6N/TD4k18xOPSKpoyGguN72vJLYwxzSUYEluAflukF1/4jPDSFnZ+NSSyDXJStm5
bmkISc9f5Vq5mtj5cLPEuqnFCUosHHkWs4cDXLD95VvmZgWziM/kmmyk3+Ys14FUz3j6YDRz4JL2
jbtnZnjTd8irxHkm/SiZRTx80LNvirx9W2lneK5ompG75dtO0tSz/tH/sDCFZoD2QtMSxD7FU3o8
16I6gLhvMLG7q7+B2tNB12Vm51zrSHZ9YfNm+vrDqWezbRdwEoR9Sa0xz3DbP7OWNF4mbt9/nZWQ
ytz0e3lYiBXCSpZhMDEGse4Wj0hndr2XWm8QbXV6LyeNKpAJFwSr8bxAl77r+P1aiv8B9eoPCJmk
3Lqv6EaVtBfmxlHHoVHI3/jfpdLqUrj4XVSuvP5pexvj3jvu9Ec5UA8KN4v9PZHH3uTvXcyBFU8q
/jiWS/58S/MKcPG6nRqF5cC5+92vhFml441ISR5koaLgiNynS1ZPfEm71xXKqZlaS3XiFlNViV0t
2Om7uXGWMRAIedCUfMXVrv7IcJ0wBAJfQ2mjMa/aQNZ/VOC0w8o9rtrVRhTheqIO6NIqz8EXUAWY
7mcAxmzbKIgy3EpyUBg6qOegMGH1sbG4c2eDOfWwgduktvd6fHRwvcd9k+6WzUenxchuLSLD2Tjk
X+R8IT3cl3/JSaFEXgeWmZ1o28PYFS453C/LTiy1UFHXqenxC80feUqft8jG3gtWtmpVjCW1+xtr
Cr4dACMYmh8ZQa4z+QK1D2vWL7N5nZSehBWYRmHq8CptgQ7l801E8XmU5BXPuFGrr4lsHfhrY3SG
APkIGlC4ufVItJuVCQwFR4dlAH0HkopiCHinDnYgt47OGkid/BGsl4GxBZFmDuBrANWRnyGB3pAg
dO5pzgk/Bc2TFWq12kqlUJ0vFNJxRIdilS1DheuJn3RspTPspM+TxzRqabX+nkIW4of6ViJ7DkX7
UnWgg7dYfIUeeaLGUtK2wGTicoytjas/d0WzwUIAEmzjrapZiHt+Qcg1L7T4SkuEiy0YjG0ng+y/
YnQ25K8615BNMEj6I3TqQ9UfvMHB/Jp12Qr8TpvPiyMyMKYP0KE3sJ+3IqwbVT0BEZKNf57xg0wE
HOf1Lr+zj7lhhVVUg8CjfIzyIo3SpqTcUmUvEFT2hOpoS6kbz2cYUos+PVB/Wu8OqXuDJcnTRGdW
yWZXqXzCZfqqqC4LNO6HNqDCKk5TWTgrlvZ6zvFvJCOw0hCuQizZmml8QbfhrsAGjAoC55qa206m
sCORcA21cPolBybIaiMnQkZY/NxIKZevGTxOSsT8JxJbaQHeo0fDg0pKWdxjCgX4NniiHzt6UqKX
m6sLazAYhkTf2BozXb0OE6wbPRaaJC8FvoC0gx4qFo8YSZRugSd6GMbL3xhXFNMMuiNmAKqBrEwc
tuMFVxth9DyGVBQClAr663x6XXLAgFAyiC+qof8B2LQfWswM9LDY2WzCXi68vPCMuBwU9nhe10TV
MCue8luez35BZ1+XCb50qIBrjJJWjwytd4pLBFA9eko2WXR0ItM47g/1TaQXRCB5Ucdr0w21Le3X
+F1FmbsckXGU9EitTWGmpmSKzk1FfbnV0qSkES68DoN0QZahbIpJgrPfZJ9BxouB8qS5wc0pPnas
e/JZrbh8C43c2BizsgME/SdX6MLnPbeKtF8N9gHdNAqxF1hrjKc1MsPXSP0EziW98yROL89imRrA
+JuiNp9CW3zxVR8YzbMgggjFYaztqXoAnDiDgIXIuCLO09Ic+sQHy1JQ0UusXxIHOUkwVvdPSzCQ
Lmb8PxhtSHFChL1fosuKC3SO7+cjyV2C/DpRPwJIwszRALqLyuX57v/ilszYJkRVUdrxlh2MgqVF
aKmjK9Fld+IdzdrdU1I0sk94fiynLrj9WcZPuUiw7AQPT8u4WbBiX8rysf8LOo6waUEa7HPqay82
k5vJI9zR5M/ZJLGhKHq19PcqS1j2KCyrwjjtrHUwTr/DoItzU4fafYM1ZvFeJwK/8Qd7j+TjHT93
oyoHkY0GQHFnDdYosy4jRAoT9ubzzTpif9hZhAm8TFeaeYa50JvHbMwnyqh5A0xv/llChQBWAbgg
GldYQu4kto7gU9RHV4zpmOW/rpr6Q2GaMkIEIhkua6xhFqqVv5uYusZeD85mNhuBae4K1TDKwTi7
3Fd0zHVY20clG62e6ouOiTqvHhaN5UC0SXbDaAZOwiOeXmv7GB7VySXOcp+4wk20iQJo64ckqPaF
n6aZCMUImcTUHqEUKoBWdPg+6PfY65xTT3PcALkSju+8Enb0vkpWg55Y5G1wHd73DD9xE9/KhSyi
z48h7X6T865kewRNmq63rpYtGyVsPn6r4GvDZC/YpS4nJc8v3JLkwxwoabSEj0TwF8FNygM4Y9nt
GEqUMCkbjxYrVFRAjswJYi8y58+QtkFPbZFfeiBUkJk6lRB7VJ8bOTAy8MIs8pWN9S9KO3P+Gnno
kOYuo4pRVVtNCY1rfM7Jjr1rjzm0qaZtnrUYyhzsmxaP3fyLIYtmG4g+YjuZ1STVrclaYUO8csw1
kPk+SjX6g1g2UtE/nuUZRNZj8fyK84i8pi4hEX/6hoBfcap7fErn+XsikOKqff4b2QGbYhgQW+0m
B2UcC673RQdnJW87ZcfeeTozW+KNq4skCjg2OFmno6c6YnNzx3/RhCk0aNxTV2W5MjDv8UcVObPM
Tq08NVk2JhWCm8qOYjZNpGDlVmT22iwwB0qRfGy9inJOR/nlrehwocFfHOx9z2dmZ9ak/YwTyo3h
gGNpbClBKU3u4+mzClUkwemD47HxG1h4iEzOeTS4I6Sg9s4QFz9O7CJJ0oczWMapaIUJ66NtUWi+
ZcBLS76R6ARtBzxwlzTfu5MrCFhe1WC3YA8aBx+3NofRs8hArJ2Y2k8NqKvVeVHDG/+8XZjTTNF/
FEyz2eL5t3amvVr5XHFyrkNVZ7KDrFLVKg2KvvYhHkJbwu7NQeBolYIGcWTImDILa0eXrLlm/sQa
Rq5Glil3bVdh0GBVKqKE/5GNh9TlihUxnVtlaowzGXSZvh5X9vc/63XO29d3552GTS7YLYz9Hxp2
7vu83Ln1X8e3E0L9di6/HlVcV0XapgoLQwd1ddRraN2WVAeyOvSjrQVFTG/J3FnzBmq+yp/oUKrg
OdgMhWOkA+NM+fH68fQNpFjHePQ9Sfjm+tTas4Lax5DFepMTD7xID8/UY+ua0fQHdbbGNM+mked1
4goBXNaEgt0EavENKZqyu08mxDwPhiFI7WCyrxDnMo98bmtbuEKkhwi5xHGRmmWUHD43M5QhoMRM
jCIsEYORxrf95R78BGNW+n94C7OXQYR0YnbE0Kvmf1wKDtrabNGO5OjqfE9JV2LKEtjL8cdHCCcr
4rpqwo033X1CuTp1iSgUjTAPyqFGIOBGNMKrZn7pheevPuyR+AnvAeOnDmOBaUqN+dDX0Pw0YZEr
Rl8yMHA8eLy9Rxkj2naeF1PRFkfshs4oNEgPr0b/BhCYlQlFb4I6YErQqF7Jp3KSsNXPKvnoTPvh
mXoLxzYrpjBWfMIRbTGQtlmXbplgvpd8N13Rh/rzB6PZ1uH1USwBte8YF9Ypg/nFTjcNovoPVobc
+Smn6bzTisWbZJpZfHNqJFKvsYZQe55MVtNbGoFzlrsJ8P/aJW89sG+oVEeNPUo285cgZfrcQa44
abf67XTdi4/LY72XaQRkr7MsjYkIovDtnxoXPH4wBjTHwTCn1tt5M3n411XeE5EJUcsDApLmHTLt
EpX3f44pbpY51G2w+0c+Lesh/nRcF6lt60mliJ21M5ZftdlFbrxuIvhASxbxYclCQ6OUvQwfsrRD
EZMZMjzaUwk+xGvEgKL7Y0DSVCuyKPlr5zK4+WBr1YFR+GeiGLhR6pwAttkLuiIdjS9RTX5Qauxw
/m2RIyPBXPchAGY3ybLfcJmbDNxPSM6GaX98+Ku9etUJmkhD+f3M6A7YSGAHgPmLAMGcHQLhkQto
+DHXEZ6uv6tsKeK1Ge+0D8aVeI3OhczlQto6UUCIHAZREXLgjHENiqE3hzxeYWsPSYkXBi7Owwom
4JmuNs/+Lp5uqQG7qCiUn1ln6aW9wt6Q0S89FSeeonNwRguCb/Vo9wCqakvGfmVC3WjjhgwnKhYo
Cz6P5GUi8u96h6TLueIkRL1NChb7w8W0DT4Ho/JYdqFDI7mDuNVJfLdPbwkDy6NinoN8cuLVNd+Z
JLaEXtSNbUpAI4p9JBz2qA1k+masuSyehG1a+E33H7IdbLLz5mQVk6zQWT/eK022B8UcYWsLP3Mg
ABID9UfUtl34GMkOm8jfD9vQT6nnHU9cyUZnrdfqQ7QfUyGxnbMI2bmgKImDJSXeai1grIP4MFYK
5uwFz95GHwGqAAoPFKei8jvYHKfa77by9s6Y3hrwNncws6qRL2cdClANsxAzvDygk9D6cpP4JJGr
GBFSHldUxMYClZYtN3As+aSWGSx78SKTerjgMFIMUokRcx60UZKO6ReI/wOyyUs95WE42a/MMpl4
yuwXypiiA/KqIHvPWeVyoIGerIkS9bI/6hAcNyKaixIqai/fyX5VDdmSZw30g4Qi+ZOLM2xtPy9Y
uwmYuvsSid3An38MyPimeWyDHvKYQrxaBZbrOjAGVvya6q+SaVyOdxtc3Y/XEfsG3G5kbtwvVEAc
B5q/xiRDwsrRk5s+cpRpwreH9Ko6cFKjTdoCKhw9WaKcyZNd0TX3TFONJ9704nzIexezm0c76Zu3
V0Io8mt/keeJdnu2xcdrerOBHIiIjUjBhru8QVUccXi8rgZn8xflEBZCwkFnfP67WZ3KpDIzWH5L
gemgSEskqeV2VbR1TuqWQYBTvfjHJ3Kztv6lkxRxOyLR6VtgoxGqMIbF9u7upFddopkJwhoA03Y3
/eQz6X9go7ItXGWiYO8DQAk845c3l1bzU1KHUNLmWQJXrSSxApCpfxB8rzcot10dVdAPx+uEQEFK
1S7BPMZnnWX0WCULyWOKRsBRipBmuSIfD4M9hud+qgSxqBzrDfi8MItwOVwS/evGtkg12NWYVA5p
ZY2F6UJLQK5aVxRwLbFBdbV1r3R6tK6IqjjFgkaP3+Kwmyx1pd4h5juy96CNo83ti9aQhn7dY3o5
OB2nXM5Bqqg5QSav0iFOAHP0xZifs/beMDs+f5tCKOXfoUXl3iZ4MWfMEicV+E9ncuetCGpPvPYL
nMPHziaA5zRRNwW5pn23VDHBunIPmYgAqiVP1OWhcZQpNWuKKS8OJpXcbO7Pp+KRdUwIov0L3AU+
grt106FYu7LRiH2b7LH4R3Tj/F4VCpIz2W8VKNuGIVP1SSOESzMLeDFQAO8EMSdNcGLMMBeSDfgV
l16kttau1nqiG+sXdyf73uFok1gIuvjORq2atG7Ot1vctsAFNGShPQ53wFhrzHE5rhxjdxaxUZ/j
qpKdXkB1NoL0HbYKvSLVPA3z7CW35RvraEjHo3rWetcO3Nn7dxrjlxAIKmC54L+sHDB+8oXD4+Ad
HjgZSNzmGHx6OpP5Kak7O0kz1i2q2elT0f3qDHpvcwTBiAacs018FKxTGKTrgsI8BFLarcpRgj/i
06YShc6ptwB7Gi4P6rQVnrrBA9FiHb/oeNG/f6EnqgiX1eTICzPEeplufdApqTAN2udLX2aheMtV
yJMVqNR/o40wPk5jMQ2GR1qUVhMpClP68EOgIQ+UseVYJNb+bTVa7Kk2iVShbB9tHYOKcUDRNMN3
AJ9lAdKmMrKbtmZPV5QXXl7mWz1lLdfLCG/edd7ssK4MQUaeHiTqYyutDxYROb0yy8K3rhB5ZFRJ
YaUaj0Q++i2OYHZb6hWh+z8nd3s7qW/qlbRj/5AIGjFfLy9V5Zo4IiRn1fEbgCz1FaIkpDwG0p77
WuHiXvG6fQlgnlYYg9j9eoT+8euqRb5ew2N7h8pRrm7vXJy6PTndnkTYyc8u/LwYLWzWNi+vdk1K
46zLfPjvXEc0mb/wUBwbjSdcqu/Fb18R7fGiSRBhx/+hBsfVNFQdLml+3YyLdrPc8vm2McsP/vVY
53rI35DXO9WeOVjx75DA0RkE6BWmqOtCdn8YbryiyuiEEu4kcRsygt+3iYI1ialqkeREuraMy2WB
XALOuB7Ot7wLAfCWOdN5/F2TcC/+N40AWq3lyoMb84H25U1UmVfR/WuWBrYnBDNLIt616dRjtl53
bmJB77q7j3VZZde6Z27Z2o070eKZpbJpD7V8nXfdjGn0yxrf5Duh/xbJdrmVdJNeILXz2qRJJj9+
hIJ7THD+5yy0RF02jJGoaGB2FjkhLHWbBcyzucOGYGbW3DhPdEtQWVHQiK47VGZ5a1REI9/HzrXl
vapSYj1UHovtIL7zluV1Tgsby3LVBroVK0NT7upQqtK3TXhHU4vpVUxLgp7Fn7wgdf/c8PXF7+ee
SNYeq419al6O07Cyq8DRsmhohHVqymkvI5kvY+xBJwDBeTh0fzcF9djPOoa/3brIfVdhtvvKqk57
O519JzpqJTPTp8Gw2CruiBFiGVq5UNl8gFwHGBl9msSY+Br8fkNy2hadmqMaI86rRyVb4gZbIw+v
QA12JEspqj9r5ZQaeMquFudvKjT1I27Id4Y3fWG1m82XffeKfuZApZ/m3//TPzgchqqdYZyaMOoH
2bU3xTEsQ3ubgt4a9Vidmta31gwjFDFWe35Dsspp5f7mxkvfBl2oxN0Mr0HHKACDv4e2/G1gJkUZ
/NDZ2RwpAtHKmeCOuVpuBrFMrdME7ecW/nfvyypMGzfakYNd4Shb5/t86Flcth6R9MbzsNcT0mTQ
DyhdRErHaU4FPPhTHk+Rp/nZcoOaz3dPMTDGoQtnCj9ktdvUuWJsgILquB+f/0PMjCxBqCQNA3G/
PEUG4X1sEsoB/+H5KLKl1JAcfEtxucDeat6YOgxtZ1Ja/zGHiE6yhB6OhrG1Xcq/N3495tVeME+E
w+08fjslsFcYmFCHqr6R6mfBy+N6EoPFzOjR5LmlsNctRqoFCc+321sZxOSBo77A99wWk0a3t6JH
B+biRrFwnB8Sup/sKPWu61/I3RmJH7/SEe//+aMmg/bD2ltFs3dU9aGiT0JsqsnEmmJw6w6pzw7D
m/HKkwUJ9pzgTD6wrS6UZLyfOLS00H/XndFILUg3IpAIYFyylqT5uB9oeUneryTs/eJtJ/DYXoAh
RmYbfjmK79gcc3wnYwKM291sMsaVj7RsLC7L1HCt4SGuWlh+lqeBcJZdQGTHMvRJnjQuMMty/JGe
25s0+6/f6fvidC2XIXAVqdgaAAQWOpLQvGLXn1UT7sBbu3N2YtdAiQXWjhOqLl9YS3tfe+IdAnB+
sYh+BIhOMCGTF5enjmdPX7JdOTQVal2o9iYjdSOQzhtYHHoKqaYmD+3yHUgvVwAQttXqwjiGJJsy
wztqmJI2FzoOthx8aQ0ogy7KFRcfIGj0iR063Kz/zV/0pDaX+u5HhMq9b1sjgf5cng+69XahF+on
mAE+WgYdKkbrOH2m2oZYR46K+XMETlXs2AXJHbGkSrcAeLa+gymVfIZ1GG1y+ssJz8BzHwWw1gOx
RAqdHeWlEY9Nk33s/AqgZ79+ItSCpkEhZ0YZBNO+4cK9jn6DlyGoOvYqwwglrHN2FQnPE/wyOkEL
c5WEM2or0V6icmJzyGZNQkuqZo0OSvNsGfG/QChj3kSPd0Xb/wKPICzEBcmeWysMCUDDlAa+yP8L
+Prx660+cK/nqBviss9Z6xUlv38mme8BwnAX9fVM7Vp+fEUsHHD4HOmIUZOxApD68rAbOEmJRaeH
BDbpiTQxi26bE9IdVMmP0D7i8EaJrQUBAjCYBSLec1BuzSbAxvGwVcxRpmmTHs/mtqdTC9lv/hrD
P99Xk2nzMC39hk9n0iNMWhUESxmGqmQB6uvoOcBlFgEqdeuxvtHS9AhGCMFxWtaEpGoWEN6chfpD
zBspplcVJjTYRqWmsPXxkW3ryxHtJLQrO7wo/BhUEvtnCxTXJeHpYyFitsWbgI1DqxtH6Of31vJQ
6wWHQkhU6bef8Mylfqj8OUNA71Qsb3iNDGw+CW/5w59xkvD+gREOiyaICNWBTxo5H2tZq6X3CfFg
RLPFbMuqL7f9G1Q/3NNdPBKD7uA0NojWj45zOxCkRFGRs9Wotvir4Vn70lqE7gsderwZDDtlqeFu
MrP57WGQP/HhgkCqapthcwx9j4xfOBiCizFIftF6bQEHLAFtANk8pfSOteIfp//yu8PgvTqRT6/j
HNK1V8wuwMBKW+DUFr8y/I0bpFbs2fn95P+4mEc7Wtv3HoebLLUb1yvqiiiu+N0XQ+9pZ4bLIq8h
lti4jYHo1QjnKSlwyNcZ+5N8t7GeRmkyNs4YuhPZOH2xKoodTbhNRHfii2FEBhoaLTz8HDVK/6fp
+F/UXmXP2YGUW3WZS0c+Sz6phHEzj/KvDN3im9lOEmzMxVX0wN+x/GqL8m1pdkum7ZvWOlCulWxy
uwrRB1MVldwkM8OtGWimWEvT9YvYOo6mcrDr04aadTHz/VjvIS3BAIMUygkk0SGL8suXSsW1K/b8
DirHSByfitq36nLPXWRW3TfS8algqlUPDSGrNe9wG2uYEfi13p0xHEJZpXd9WitFXyBgxnzntXkH
0ml0ftFKU6FwpqRX8qMjgZ3ayFIi+ie26G1eY67fqbGzS/vSbQzFikqWlsqHLTnpEDmJ2CgQ2zpj
3Kh1PcGVrWxoH0ZBEJUIjfPjLgysSHhw0oDYkqAkmmrRvUSwto6AhoIu8amaLI8IZDBnOqHPKl+J
adliSDRyJ5pgeBfRplWo+XrktefOzxlWbwjBtK0Xfl/53EFZ7GAolpHklfsnLA2xn5Rs8GdCFMxp
PetxpGa9C4CKtkB1rDehQvLzwiY8hqzHsFEVdhUKRI92me6aewcew3dsI/zWssUncDGqNNnZi0g6
8uUOaYKemqSJ3m4uvyhhaZikMu3WEWaBHomG8MsgXdaHxWfqspF0lvuWF7qPDYeB8o3Qqf0pt5m4
V6eYKYPntzdBfM0RYzzgtAIhUYcdn5ptLhq8JycmUiC8/+YDLyjyF8KOKDYZHiiudUDa1lbznUr0
p4NiPgGZTgdWOBo45d1rFM2JVkUdUeYbhtp39mfUAqgJMBYrOZt7sN2d67xKOcT4M3dLkGIfbkfB
S2eN1vFJOynUGOVty/gvcjio/Izwqy1y4SHdegVDdmoPyh2fZUBgIOJYMkfRX02l84e0faBZEp2e
KjexmCDQ3w0KWkYHAPU4LYbII4hBADQ0ANt4Evaf0vLrEwP2a5IZHSudzVWIABkwqc5D+7H3kkm2
ZqcUg4Xalh4jCCB5k6RgZ8Q4pXoAZcQpBq6JeUbW1Weob1+R3UJ4aEdn713kF5XHT+Gu5xKl5edd
tY0+VF+rxO5steG08lqcl/kGlgcwdjqGol3Crj1T9N6VuslBXh80+kAWPUkeFi6qNA/qCne7/N8j
9Q2tXC2KXxzsnktp34i7jGyv1W5D+RS3LqyXFhdxOvkNs1UPRYlXPozErtwtm8rTUCA2UgH770nz
FSLsy1399N3P6qSVjp6NMDZp/QpjK/A89hbFh6dUjjNyE1kHvF00bpQ0RTUOryg8JRm3x7+XEBYf
pfOZOfR8RTNyOZN8pCEwxE4P/CWrT9VoRpgpjcTtZxlCuGGwuRKEm6qOeFNlJyCrks802rXvlCI8
XSUifmqhD+ekSlrDz8N4QuAv4SLFCFA9FbHImJCTk5wxZL3hhSfll5CJHG6Sr03zJUJKp/guR8Zz
ifs5YZ1/rGhhhrqWjQKOzZsxuBjvQD3TfAl83L7N65Ftm9Bqn5JRzj/ECejikbibrJAvnb8PXeU4
4yAVr8MYNDD9zblW3hnuZ0GD7Z8xRSSW/wFRNHDtlNsZP49fUWP+83gWtrhQbjAAJ5rBAV6AGxnQ
Gc3EongKeg4QNrDVvEBby/0TyGKhzzuA+aH6ie+wVxQCJArah0NBPkRmAYYNp+GabQmpA5FxCMZh
uPcyf4MzF2Y1S1xRelOGInt1WrRRGmIUpvmZv/tid8Ri29Ku/ogkfYQNkf1W0BEz9i5b+V+OnXXG
SjgToBe+nBT4b8NU5LM+a261l91Vlf5COKkz2/7USF4YDOep0GGfb87GpaB5e0LUIcrOSoLhUCQT
l2CL24l+mxOY7/n0P7/fJt/LFZ7kOZznRVNIpOhUgEexKtz4vfiNEjclvoZ6GwmNOKbEk1MYlJ5O
pW8AtORL6hrdx4xmGMSJvFZv4JXttqppTXq/vNX95AFMIY1ZTytyX3Q3Qjz+QnyL0bu1+9kERndb
0XK1jYwJaGXlOECDHexKA7x9d/sDGIs5w5Rp7Y7h1FVr+tVK7eDjHxSGCa1Xzxn1mcz/NZ+J3jqv
OND6hawekyo/ITFjztn8kRjbGvygxffEtP1VRodiuZZ7v3ORoo7nNfTD8ro0ucNvygD3SH9lc+Q/
wA+wl7iPTyiu7Emf0h0QQYjKMbX3/p070I4/FXWK7KHwMx8u6fabUPuKgpHL8XsEmKorZabPLbmS
K5d/g0o7rL17lJ4KgB+JTfcLojJx23UIIiSVZa3X701iXxkZFZlUtMiW1aLGjgHSwxwBRnHi1kLq
j9mTWjwhgEN3V/UuYHZpE1yKnHai0uZ/IZwJMknSkMwlUWHJvkFfzGJapadmib7cuFOOV9fWvoSZ
fmsrpGKXuzrDa0CzQBZgQHpMmXMbPS336/NrhetA8B/97Xwy6AHjlbke5vKGNq0VtTEyi39fR2Jl
x1Xd8aetOVJejJu0k7L+oZec/2KyuNPPtObHKHS+xfrl3XzW/usUxmtdPkd/wDGCMTgVVwFY73Te
AsT1JwnzdvE8x6Xq/YXdU0KkSowMhd2oSqjW3V7vGmCX7xQFoOl4igOaAl1MrTHfT930KkDl5e22
kEUIwVIG99W0eIi/3pOvNAWn85NyFj42wqY2StNlrLK3uDZ1b/iiHsRqebLOlADKindfzCG8+mUj
cq0f1yg7QZXLLdbGLZ9L2a+A+MhJVleLdTYTS7IL+zp9K+ZxB34hpzRLQdbhkuorW+id7YDpG+yv
r6jN7dI9m+Rvn9978vTszQqlg6i1G7mdJMIQYkO8KDt4PqwGIhB2sidOCK2OSpJFbkT16Sk17ODf
cCPLV0b7eIHY8z+uyS5wGHiK0ojX4ZmNJCwTMci8fIKTk3NP0zd/rRzaNpbrHZ108tvUe9UrLqof
NE0IDc8XABpmk0mhIjEXGldZFAdHu1y5XJjUakiR3XPxnKwtcpe1K8x4pS76XE+O9oGyDIDoUPOu
L9J1Ah8UsUb4sYxWpmxpGGKZdr1bap+A+cG5XCGLuxO+qYaVQblSvtDRmHNt3urIg+1wa45iZNu+
C4c+AqD5Cvob8eUfvWnkkQbxYbH6bsTQgD4ezuA25BRMPkMkHVCEb79qTX8imJdz+ZJOZniJcknH
XiPsHBdSXBZhKyd/nlN2o2RHMfuwUhRuF7CXUK+TMp8r3oeERso1J8nMtkDHze8a1nzhE22l/Svy
BPVO52M2hCYMYkZci8GyfYAYRl4uqbPRYgFDaxpDA8Ph/X1GOO5nvA77Y/0vJxKFE42oQjHpmnHk
M9UC1WpWg9ewVcrjnJOzxghdoSQx1sZvF2dVvoWLrClTqTX+qsGsXHJD59AaC2m5s4fTbihr2ujn
gwtWCRoIwsfCilWK8NVsX/cYZfqiAvp+eanZGhmtpIXPKLBhQzGcwiF3pivnfdrvH8SZDp8FkbwD
lG9SwcFV323t5mp1IEkA/CLJ0oSh/gnQgMPNyU8VnstGgy9ILSerFl+VM+USxljv5DESzK5Meh9E
4t8+1uec105L2oc9vVAduASujmelwnXRBZXXvL+vXtDNR/IcX8FK5tw3ycLxzMcyXpGwDoXx09Ld
B6URWbQi23E/5NEbKEi1IObPlsoRj3V0nZE494ahDriWmZEjsygvdUEXGbbm6ZIUNH0Po3/JsxTU
emIwYy/eFtD2nBliIgWJao+9zm/gQoLZJzwh82+YOLQ/V0F8dq/RNr+3EXWutuRwDc2xVlwgYXwV
1ch/FUy6B3531iPlgpmuWFQAyfUoaa/Jdb7P+mWak5CmGuRMPGtZmG1CxDmRXxHNZ4kP6cu9PvQR
5dU8hxvLbd6A4Dczyglt/nhyCbVYRPT+j9zqRivXKnkhAcm90oFqbfiaDKANYO1R0qFvLDsSmgB7
rWG6mYfBB8NDVy2OZTZC+E4qr3pqigekv3bNtuQ3yGTtQWdBAISHUqiOYwJEmuX/7qElaeSqTwNz
iEFNKS8Mgddzl3dDhv176ztuS8RnlUO4AqbyrUj7TzsI+IkCRhzJL1gC/600ST/slxdwQawb/4tA
EfUEXUTBd1VsASSozZLrizLLYSmK7ABN860CLfC6qstnGOl3C2eIMfJUfL8trOahxUOw5RwjSogK
7beWZtnA1jRWXmxjduYERsst2C6Lo7vrFkZcynlkw/l/0qqmbO963CNsBhEBB0zzgT2PVaoVmjIW
d9xCiLUsyhSEFc+WXW8c69LYx25IoZRkwFNkOG92GWc5PA2kJXpyEXc51FI/TfYyuikcgHJCJ7Jq
b1GV+LMZxIK/3Iz6Irtt9lps8YCpcu/4spn2oVdUOMhDDbKqUh1VBFcMTtK79B7KoxXK83QA9L1e
nVScO7rGHxtetBO9DmHy8e0Oc/Zp3yfxYeJEmvBVo8UhonxOSlV+vU/pYCstpj9AtDeOFV/wajrA
lrgw2JUcWt6Qn+oe0hc54Ck483aHWlnvnr+y90Eb6TNLLaRrGHX3zgaeiERBJ5PHDoB5M/d4YWw3
NE7BLjKhQJktF2c8QxC2z94pkarVE6RWf/5HzPngOJKwGhJPJi++doxSprPSnzf8Ij7cVtnCRw1m
IA2jndcA+gT0moDAA5MdS8xsgfcAxyBV64eikgVa9k1iSyCN6ugsgRbTI0IfCZEHo8xhEpBzgii5
S69n/LZ93ma7RSToji5vTL3EDopkWR0dIUr8kykSiiEKBQPg7arW7EhwuKA288uF7Dp44WW1oAzw
i00umj2M4mkbWkWUbKqmEjxVMk5A7NelW1Bt0bNq2QkujwCyGkqg5l1FYorbPHm/NBG5NdGnvgPR
4Eo+JZx9zyV9d5VNKBJN6X7WTDy4F4F5l2ms9NHD67p+kuglolMKUbyOqaeRKnL0OuWbQ0PvoH3E
S8RZmVMPPCYCAtQXLydaG8QQPXY6y7IUdXRhpMhUfk9BNLoY0OzR52IjH0fzQF9NUOkUIuDGEry1
Iaz6cBxvJHQySy3vt1QxbjDbaMpAHVYT0s9THQSX2hlRY/sGLnDmhJPa+zD16Tw8FTZnG7G8VtpR
9m5/bSzlP6bdRo1wetn0ZsXUF81NSPcITHsVU12JzwJgnmKNWxvUnKABkKBMnBzRfMYFNY4lFfUE
0ElIftdfVpVA+CzuOmjWPr0fdpbAnmn8sp1j3jZjDciFKsX2hloIwel7K5ZziLRDBtKaSmem4l2B
0RMRQWegTZMir0sDZs+YvSOTLhSwH1Wie3UaQ/jgj3I70HoWtsxLRGXj4yvzR/pcGQHh25UPbZHy
8KdZwsb+URduglslq/hFJCRb9TNVbEV416P2dzEZ1huQi15AfpA4KeNmQWE1YWB+vVqx+iYizZM4
3bbD0u1F68LXWX6ChE8WEIjZ9w37E+MFns5GMo77sAhUpaWQR72an3UXHTWA8jNzifaAB/SDnkf+
6wSL6u6e6yxazr4pfDtnxgSw3MVQHBriOhDfqcwqf7Hf/jMsR/736jHq+PxnKyCLL1Afq5S8kZ4l
qKjyb+V+zxrn7HYjrjFtuIKaBiyRObRmDM7Uby1ImQmpLxdb1IVjiDRcdQ86dpIuezTVSVFvi6hC
hW9aEO0xIH28Ig1S84ISOoN/RvM794UN8JGuPHKdAaZxA0D+uCZsuZdzyd3+hK1f5sZIMOOC0uk/
AHBipNDbvuVtm36pvotX4fif1oq7IhvjNPLSPyXW39VR5e7/XIOzrGZYjMSymqarXBvgJHxUn50+
uY7mFAR6UrCLqRLxSSZZIsLcIiQ5eI2T8Eqyg0yMmOYA7vQLQ3KEU/VktAW1MQ2LKboSbYVbsAxo
SGUHSzn2/JY2xaXnWasdP98K6J4XrM0Mp0W9NSlc0Hd7tvvVbS0RJ3zRVQpQAA+Z08AdrNB/gSzG
/pTJwMtTuQve0z6x/b+Yc2qJ9JbsmGK1+8o+HfeVwRxlHnP+OWDxslp8Ci/9Icn0Cx4tbN8vzlPI
u01afTWBoVOMf7LxyQvlFcw6UkEV3MZrxT5N1fKeLylDHsL5lfWRaOZv1U2Pws3TQUmgi7jRKsk0
bZiJjMBacgtxiY921727tuesr7GuIwYuSdkLyx9xOpBXZlT9PrNd874zEaKwx/3KqV+olp3KF5p6
3gesVmrg76r1DEN7a5v6EONlNZ/fSi8Ee09e3CkawZmSBxivRyHtxSLpdCluwminxwsRDjLgmkAA
aFzY9KiDpMMz6YMeZQiW7i5UoXRx/DaEMAOoTWT3QRn/g1i637u5+obQXnMhe67da1unvSobpD34
lDxw/eHJHzJSKmjD8SoXqpAcclKBrVHi4jv9otuFlVv91zF6R8cFzt9Q4ZJ7SWELfiRms3SQGisl
uIPM6p+CN7UpkMhnTp8BSArILbVqXrVOILkOIFADqWq6xGDXNuK4qGJMZ2Thkfp58z5Py+lyUpX1
/6xjaZFZ8phw/fvFIv5vuiSu2k4BQ+CxPrW+NM0A2OVgIm6gFBTeGkFQ2fA/nIWTTb6pqRsWuh7n
3MW30WnitGct2MScsK0eFUofc7x8A4z9XFztvijzuwu13eEuJKueSk1vB4V+tepHHVSouLov/jFA
ug513IRfZhI+JooVtYThopQam4/I2FqyUTJn94+iRSVqLp7XdWG7+DpALTKkNMMBcB849M0KCdKh
5GMtycVMu/PFCV77dEDBNjRd+AGU0CYNrHykotz33wtw5A7h8qQrH1pdhh5KFl8YtgRtPeiC8JQQ
qvMRbevKCh3f4NDIxTP1/oYWpxd3XYQiomCu0vdC/qSNyOWmCGxpDF1+PaTspkVO6pN+X01Lzdo8
6tkbP/x8sPidSpyn5SGQDlamJaEulAzptx7PejoLLRxDs37+FSiOm6F7SJ6DhVjGkQSKlnyqZ6r6
eadlXzGsmlYjUPTUKuNb+t7ZmWCEFOcisJDl8IsGabsFaiWjl38bJWWLqldVUfz1WwpV7JVGtLAw
Wo6oSJuIg+GTVbxa2Vyot/3duT41ksoVlkAiT9Is8Obz1UgGHFwUfhDWkf8bwPs2XHx5ywpo2RkK
SJhMOzqiof/B0QXCaStgfEoHxPdwWvBnWzRbnZ26JmW7EG40dGWk/3ZzLnokF8GNOBmojf9POFk0
YoeG4bO4RPUQVL0yrgOceXtJyXQFy5RvdTtFkWFbpOwXQUKwybj/mDW+AeGMP8xzjdDP3NHcJsUS
7X8gVIoHcrZLrnG9bZ2hJ9AxrdaJjmp8vH/n8f6z8uQP3V6i1It9qKSjckYg/jFoV1sEsOga4xJg
/X6Zoy6gtyCpUA+giR7kL3hmmX5r8XXRu6nkPJ7cJeQoOmvM7UxVVTCx60zDVM2N+1IxtuGD/MOo
kGzB6J1nJQeF7ObUlmO3lHVo2JW8PS7oEHMqgLJR6d6egdeHbdd4bQVrEqiC/MiXIJEBkRmYoRQE
vdwnzlwpXcQaD6/3PfsyueI+0ICFmDM362+efew7UmiwG8J0dViKvZgRd/FsRCStDanF9PMqPOX0
wj4O+EsGgATOZvM5fFwBUqH2G7plY3GjVMz+m2nEup9F95aviaKf/sTAoa0PotpKrVQagR0aTQML
egpgX8/6YzTGFS5m+Cn0lwQWjUKL3BxaraNQDWO9g8ErSOGjrPki9tvleTFj4N826juT2gmdNNJ7
Bb8Fb47CfZ6xFMcABctpywjeG4nk+TI5k9zim3+bhKHdB64A8lEB3LI/EoiQ2Uv9X3fLFSqG3e/f
yx4mwgLtNLGLdQhxTKft5tvltZY62A+4fF9fisMvqUxFoQDESM3aobFIyazdVB4XOu4YKUcFgjsx
HGrc0yZI7GbiJH/N61gIinKbVB0K9rLK00J5SRvwCH+z1xBWz3nIDC7Splf2Zz0MOZuVIpQAa1nn
YiLk1Xqy4ZVnYiM9z+h2zYCVilhLhKdIBRtGmdBYTTVYN3zblRrzB+0b5d9pIzBWxJzSflDDzoAF
AQd89vjjn22pRyC57qReYScOMowVMUWohgMhhNfd5QWn67/D0IqcDP/m5v2YElI52W8mJjrZIA+f
DzCDYDLuoGSleGWu03MWZ0JWXHlnQoNFCAmpicuJkesc7CrtVqite9MM0WUEDf2e1B6UAGlz1BzZ
64KKigb501HjXTdtCigV0ENii17ytvd4Dr4GKC64oq0Lg6vf4WvfqveDSYg7eyeA4gn4++ejQPrv
Bhr6zVWhppNxadNQVo/OxgVgZzhtgNT5lyDFarAPGrGgRaeNoOYHdLJS6zbPZ2RAuPduDCW1Knxv
6JnkjdPzNh/3dQnaGMUic0BfUPqEWqqTjrMerorDmA0Eo00CqcZtasJlZ/h9OgbK910H65Y884iR
0zeEvN4znO7hYgH3exfq+TGPZKBP5dhP2NY6d9TH7MMA7MoP6a0RcL+42jCccxSl/V9Gvo/9MW8H
ZzWwTGWd0UtxJ5udWcWoxS7RZjx1kk05+xF+eBHBt5NAAqt5XWu0HDWngGAooyzU2wRIk0e2UGSh
VvPEHgh68Hs9zlXBZTAewpVoz8Rsq4QX0+aFX4BqRzwP97ekmS0f9Zp6V/4A2bQcmjK6oO8ykJ8D
Bk1QnNH+tb9GaZ4b0A0FXlYHD92JriWC5hwQDuC4W+QB4rUCunJg4YQLxlQCPdQgCKKOdXsG4cnh
W/Ato7EOAki2QlBiozK4voK0eoNXMfu0ZSAfyPNO4Wkq8LlKnV7u+nuNdXMreHCTKffZ4RUmlpy+
kx4sX6u44mAcMCBMw6YxWE9aIFRP1FepvRC3K0e+S/v7vybx3s7O+Gz7XxfuntbyLI8XwVfr0yWl
EZ8/W9U7VirMmvKSqHqDHsh6tlSQoMnLSeUO/8mgrT76h1wDO4AauO0jFoPsxK+Ez5TpF4QQJYkT
UHlb1/ND26n6zpW5pD1a2dbTZGqLNeFb4pbAUfAOAy35EFwEU94uR4skpBlXBfksdOzI8oNXh3LB
Ii831Mj3F4Mwep8Eq6avtVP2kTtnpHkht5SHj5S/PxZGuDFebkRYZ5O48cVQI6zrce6KOM97otqq
PRHklGbiema2FSoXUFTVr6P/RmRzkkgZ1A2fQjOmD8USmERCe+Koo+D05PzCB7H13UKcYtm41G5c
R6OAM+ybHBU3mkz1OyyvbTW+oQkHp0o78clbbN6fIWzgHahslBxDAlOJzJyILQr9MHY+Ulx6zF36
tcCLgKtY51zO4wQCbcuDpXF8RlPlcNwk0tct5VBoSqX8a0fDwfZ3igIqf6jqYtwHoFOSC+SvrqEK
cya+RolC+XmB0iNgLShWvW3c6IZ73Ofxh2tcJBeOD4UFs2Acj/GBKQe9z0KBVvggaV1o86a4aMyZ
aupqXKXwoEYxw647c2LeOrWctfZY1zFMPUFb/G4c5oX1l2wi6xD6X1rrUAO20xRACZ0VID8OPsiG
EnvqdoN864R7LtLuxBJwl0tAPro4b2ej3N46Y3jp5HvyG+JU87itgUh+07r2CzVikLg4TmJtn/Ou
Vd8poSlCGrAaEz4jUnV5PWTuwnWLY6kBxUY454m3kVfyloRoYB6CmIeZoa/frCDye7cWPjqF01AB
wW0CL18s6IkPwLh04BR+hx/2ZkzEucUSnZxBwCOgwGX3DuKms6mIs+UmN4/zrTZq4qqCgXGh4O9M
wqBJx+rslvSui45Ik/+vhj0Kiyjyz9E06RHje4V2/MAMztE/PUTLOD7Ir6Ww8WQmsZJZRTFlJ2pV
pzcBh3k0O4OYCkeJMVhsVM4+BG8q6n10yFjZg2RrGZgX7KqGirlYWvLyzVYQB0ERV8LUJ3dXyan6
TcaaoDSDy9i2iGLo/76B2/a7Pn3KBXMXrpO9+2YtMZ8AOqNLB7xprVzHMSe5t0BA5ZqOqyCK/20D
80Ubl7LwTi9SPTnhRjWKyM9VbBjwNFhXA5K+zVkIk5C0MobmizRWllU35o1z0iB93LgGKWSWQLN0
NhKXiISDgU8LLtyOmA11cErO80Vm4OUhpErQBkkKSri3MPW9DPwTnG7EgoDaeJ3xTToecU/d4MGQ
5iqwo0UHRuf5KVTuZNyukpiG1ZjKYENSXG+OgyW0ik1cwSbYoRjqSgJjLWKCjQZhWrl0qveHvGQc
+YFVejQfQa817uH9WtIyEClKmo83Mu61vaExDsFxHXLuzFw+cqWmSQKU6147IE7VdR/vEpR3Kppk
YCeQmMZ0Tzfp3n2AyGHeHhpg0Xh76aI2UbEsHhflQN4bL4wPkgs61cytQG6rIwg8HBIX+sLxomS9
kqJlnZIv1MKCqklViTno07gX3LQ333I2EzseLMPaFh9/2ebspUDVcOlPvgQUKmyEZDvBzDJFnUTF
Jojwl+o1iI7vf15R4JNakcOOwDXTKkYNviqklKnwOkKObwxscxkPNCtP4WireXuCBdWLQ4ThYEV9
g1Db6DJngQt3JBXcJA6XQL2say061jZEX+k3HnrRlHh8orUDgksweZPrllUB34bNuFZzPQ/RELUC
Q9xLCvdLbyMQsuq74MQy/FnmWKbnFzFBjVEYK+6krfGO0MSYA33JmJ/7wp5QFHejC1rBrdKbb+WI
klsvnyzODwG9S75Aj+eoh21Phz/4V6p42vYg2Sfv8Obnn59Mb78WmXeyJWBPCMgbGALny2uurnox
jX3SckBktZspXd5Xwfnsybs/8+vuVw+AdLjULL03xZRkPZwLuOp0NMq9x5qHw1ppsAZriNxo6Tf+
7ofQEJItuaqXL8TqfW/o6qo5HfY79BIXZ3DaPoXTuS2oRGChciE2Wh4QP01A4/K25+nfVfmszEu9
Ox4ufD6MmXQJG1vfa4Z1s46bbXrA+6gVyn3p7fiZU68DRYrWOe2FtAmDIW9gWJkPa/p8Hl3LA3EL
XmRAis+ZFdsmZObq0IroeCWBSXMm+s1PrQUQ2wofEn0oYcGIOtYtflNeIpCs58oqsCA5rotYnFMM
aRj+H48TT6O7WZ7PrSLuXlkzQtwI0ad6ZIyp+gu1kgb5Nr0sb26ejCSukUZni55nR2KAsz+A+BB4
eTvX7kSxnk9pypr/FPliN7jclujKeE47LnuGn/PFqZobnUhkF1tTlI8KPWz+xk4VlV+fCcvQKPRx
wpTF6UCz1ayRz8m0D6g6RryOyE8p7k7kJg/w9M96lGDB5GvJaXtk66SOGzzo9lDeG41URLAGB53/
v0PUYwJIuQz/NEKR1dVNzZMw2yhQfuXA58thZ51rKxFUaVcnS6LIP1niBOwy9jYdfWDguP6QmtFI
6xMmWcSbx+Yh4PmMsyOZMuL9qoLLEr62tgtWacyfoOCZocN0jpZWmjgWUlb1ZpB+YsJbqzwwLGzr
4etcgjPEKiSm05lCTMeqw6VZpMSp6eJH+4cZl1u3CmF7fxKANPlH55QjlG+smgs3bDNlVADROO1E
DaAVagXJpQHegoarsq7V2u/jH6o4VvAx/juVBVfyPEOol1mF4nyyL315x13gsxzbai0E4+BX1j8M
shGW+bGyP5T6utHiQds6CFKg18+l8TwwVt1xShIY6iXLyRZyAaBvoyQlCGvbFkMlYLj1MadRqRB9
YcOlO0p5mIrmNX9ENJpl5ZHmL2ZPSwJIym1uQaJAq68vycxu2H+0mH90wFdr56W1G/txsNzeCncl
SygkwHlE7RPvmd2Q889CizFnTOUSRsYJviM/eRGtr8byNXfoq+DH20gndEGhl087h4cKOuOnsl1W
AvxAJPnNyb4PES5EdHY8Wto2QbETgq6V3Co7bksk0sPio8Vepcvz6WJ1Qwp3pkg5fP0+h0+SS2as
OvDE88n6S35SZGUinLhewGy/+3W7PkeQff+SWCmXjgF9YzayEItfZBzk3O+qObJax/hsProEmYbu
OxzqHWGGcJ+ZDLBaNSjdC7zV1lz7vmfaRJeQLQCR30V3hf0T4jOZwdLT0RQNMUG8oOH3ArggcYFK
UoPJb4ZPBNrSa1HjS3TtLCluSAKHWQt8scDC/8Dp39a/ibH5mJvIKLR6AJuARhOYS7F4R74qbLGl
3S1RhncBp+qykZBLGCyCaNK9O4JrfSwOFnUOwOG5TZ4BWZ9NaPMjQl5XvYyBDB61If7ikjaj7aWY
Wor5HYAy+xFSNOdW5J/JhuHEPpITQuIxX9r9rhoiIXnCE7daklo+b1H2XlYB02U+J7F4oVyDwpkC
XF1kBaHNfNidzBuXTi9GVYP+eaW9tN7iVsqS+KGh9jIOtlXLwxnp+B2KSsgMGwl+LiQWh1k/RnJF
347+Bi9FlZi+MBPg3G2JvwHi8qCouIuKa60herwwlwLOfDDDS/ovjfNWnY4Xs8cKtVtdiiWftJ1L
8UarpIrppJMjHfwvbsKXNyJLKwMRxIbzY/4nkG9MJPeh8gTdGUxeBPKAdL+1ypZvaWaec7jZDxga
Lm2g1goSe01K0uV+qaKJOhnt639X3VXS+aKc1WFqbloSikOX88Py5AlvRKHJi14M9C3gPDOXXvzQ
JQVIT20+8ogbO5y4u74t2EkgBFLO/WKlT5Jj37GKavPY9jrVHCjPZ5Ino7nnlTHcw/pTEcIKQ1jj
RGDq1621Zoq7eOWuYBq1EUQRXs2Md7/71PThO78tf9hrJXOPomgBheA9Ozp0HnDDprBmfwD+WYII
o4Fa3MhQ59f6nOeSSoUEGcX5EAmmr1eFojXci6p5inQAX4cTCkj0rvFbWYwHEyTPDg8LouMPn9QT
FVaa7AtFbld0chUbKsp+XvzAPHN+DIUrGTsFUHyC3o4R/WLrrrJ6JcUBRh2h6ZCx6kR82r1RvXp7
NyCH/PPSJfpkZ4lztHpG7BJPEEKimcKIjeB1IOrRTqiTeUrxjzeb/7X+n/skaKBsjoSGYgUnavRw
7XoROURi8m2bXqoehrvbDymoemQXlchxTIcopsou9BPQKtVWog+1dN2jtdE6M1NsjdshmVJYUg6n
QlkMlvKbO9aMBEqAcrFyIPSSxGGrhoaNG4uvIjCFoxiijP6sZKXm6AKFpd6dcDx9av5fkWICOmI4
aynWsonhP1dpHeK+66IW2LXabaMX5Z7VNLD0eQfSlegbA9cZCUoUcbE5sACSInBlGihKviFkLoCE
Ay/HLdh6v/4a6v2Vy4onioNWpBUldQO+MnauRb6Yk5lzTseCzuwa+k+l96zLYEELSqUPpIf90XvI
sab9P/7RKN64BCJWL2Amljwp0zGkqmc71mtwGloe3IUygPw87qppVLh0tDTFJbbP99UZGH8sFcEY
fYljajOLqpqywDJYjEkg3SZ8eJh1V0QaOjW1BJdYKIlxF17lWFEo1abpORln3aPLmH8n1km47erP
3wLDTt8jT+P7iIvpVGOsXAMCatm9GcUug3ddK3Z0CudYcdqzyI9uHrYvErLjjBao/FrmVvAfbz/S
eO/fqWg6x5RO6nOQrxJY7nCicFMEy8Hx3uHFY5gTju93beL04ZVJr50F2jJqA3kkTO/gRQgqESck
GBqt22WTLqzAJTabtp4EeGD3XqZJkvQtE6b5hFaH0UHWE4bmxbh3sCfLVsADihi9N7Pbi8t4SjCE
ldYC2jPAqr8wdAYUO8bdc736h/9ZP+72bbHR45MUyww2tsy3ptn3RMqwP8t6M2Fs53vaSydMA1x4
Q3Zlnpm+f+kmtKdPH5DQWGdBjPf+0mifiFcR2RQnpGSM2XxD/KZA++9ZoCCXwM2LutuhXu2F4Yuo
D5P1tCCDTtGPs2b+Tjxj1t5pw3ZNG8A2TW2/EMvNSFeYinoTdQzc3vBQuBo5Kk9o3kt6SO0zV61L
ha2XsngEtqFsPaq58ZWrcC0ICCOhAtqmdU3pTEXAcxO2MWpBK2Zx92pvkoKPmFishn/lN6Z9HyZI
9qzRUjBEXUOoCB5QxkeCYrUzG+m0KHAu9NnfKgTM+UZ7Y6t9EKrhJtiRhWcefwbOUuaE6YHjYPKT
MKF4HfYkZ0FOO6vrX/21CYs2yodeBiG6HCM8T+afe5QQfxw6Yuc+UjF1N5jZ/lrTFYdDjNGw2um5
MVWh2H21mYcspKaFtGy6mxgT7EAArnh9J+yklL3J1Bk+X7fxj96FCl5DWAdQTrcCZht1ycKKbS4/
4N9QmXvIJXHnnCglbBgEM/GtOPOTj+gQxnpeRUo3fVCXg3ped4qmta5tUoYr0we9LLhl6WLKxOub
Duw1+9awUQUa1d7VeLsIbxSl4EQYVpnRXpC/AwvkwCPKZLyvL9W/C4xDffE0JbZ9DZvkQc6vJMFX
fJQkX4cKBgBaY6zIR7Bdc+Reh2pSWHU2zfx1Eg9CyodAXhYdVLO/taC79vD2XmBXjHABUJ+RxoUz
83slWqkhxCJ+7w2yc75jwB0HJrM5mEBp6f4itzVhUXdRmNOtRbkIlMFlP/ECWo3Xg0sxqZ/wSzgj
IuLWr+IP3VwDJIj4OMeVOyIBGFuStYPXGq3nrOn/SbKjDf0YzEMJlXv0znqfoXcl4k7zFhRqPkS3
zygSbJnrTxl7gLLnEayRwRhg1DxIwg7K730GeFL2nAYhmi1tMiPVrG8/1XL1P/HCtsTy7jxll0Ly
mLJk7Lu5aV1bp3a7HXoC9Q7MDgnovSlHny3KGBT8VKfgv9RBEqAp07LsUJ45QXCDM61AP6GCo9jb
O/aW/lN0FVo6ThNde1GP+NU8l39Y7+bBSeG3EcpYyfnntlaP+T2aSAuR0uxKywjfZZM8wh6rOQV9
6ppt2hOQ1TZIRgKqBQ+F5LKBPrihFp/vWc1fdvP1aSt23yb3DlLVPZhAexTtD39FsRAWQDlQy5SB
oD8LSur1xeVESyK8GZVaUD3BY/u8k7PrY8lg/GzPH6ysuQBqULdlNRYXWhTYlQKOtILe/BZxE/8x
CfMH3yWyMwhsJuRLYzV4BArmJOSHN/3bmsvepDwH8aq0dGvzJpEps8RS/taBdATkBvgHoccLnOek
Yp/QzjMB8J8CNyBIpz8bO/pTBsKeTfvuE2U6o+bOtw1ha9OXf7ABOtuxpxCqsIzGdQ/MVEFjlzHW
urlz939fYutprhc/nr0fa8NyA3v+sDfGotRbeMlaUs9OexYIJO8hyh7HHRv+8qquNpF6XGFEl/cQ
yx4Vgmlz4T147CSVTUROXoxsZu2RGys+sdiJpFohYrWENLiJ8V+TLrGAwcifP4brADuolD0ydxsy
YTT3j/5wiKoTB3KGkH7e8com7GqYxIDE3O7nvX2QOdX3HujhOfM3pdu0y/aabNru6q7YP61Z7mon
mqg6x+eGtZyT3IIU1fvceI2Oy3w9pLlPNXZ9xPd9VxGHfIHAQjup7J7UStjw87gPXkY1WYdt5kLN
CyrfsJ9BTFBCJJMvIL0O+Ui0AafJALKi5qApT6ntLDVmOy6BkIl8sBjssQ+7VBX18XKqatlIqOHD
x7aMXb2BoDhG4iqYDRcKXroqcc5LT+AfEkKBU8jNS8yQyPMO7ahV9A4BsnjUR1qJXWcyYi8DhvMk
KG8IenMh1WdC8d2rbKd9ViJ2GZFt1vMqA0WDZhbBuB3JE3vgo2vZH4KM96AHM6ghYUzSgwwg1waw
bZ9SkEasaYDSESp3rs0JBIoqkUJU2cJFeob+0NEKLm0ky7/fDYCQKRhVwagA00mfByPoR1GiNl+s
kKIouOX+scF6+5HVcRl7W+9NxeXQKQ6cgFbQY18vMCqfIA2O6TPaBUus6YGHxuMtSErLacn1l8Po
XOdQq9uFpDIFfVipRbY82C7XSQpcUdMFvPtqDW+Bi8KGGvBVK2odz7mXIyR/CHRt5cHWB1fnAGSY
NwcMeNvRaDq8G3TZJ1XyHfA2Xl0Y3+ezB6MYd6riITZi/r5H8YKnlsPAPkYv34HBQ2FHKDeWv++h
HXXQfqe/1VYsQk60uhkKg7VjOglfpTChlwJWR9XXXbIqycg+kMxTuqY6CKCiv2ty2dnJiF/+8i26
Okg3IBZC1i8Rv9Tu6Cp0aW6KNUWQExmNHAqmeIBf3QaLXKPPSBKiSV8YFjH5PfCMWphRCzWivo6o
PQ0Dbo4guVDZRERoJQgU3tuf0OhGXNw3a+qOF1rx/DD3dqMWQBItL+gsRdOpGi1z3v7/xFKYc8UJ
KlN82oMH9wvIVXlePdcAmaCxCqz1ad3p2hfrLWN/0izAx9S1JCiQFWp1DNXebMy6fl/2o6d7WnYC
qGVIOmyj7FvKPrkvqcsvSm68Eic3Hht3Dlx51CyL8AuAJXjgoHmKxVp1EbgiT9y0O9mNG3Lonyvz
Ee3gYfc+2YVXtK1rvpJ+rMvTKkr/zR7/yRdYeoQQTvqZP/3NYx9tfC/4KCoxanLojfNk4meyaIGe
ZD3ljHfltfHsNbBHhzkORhi+ucYZThTEfzoQbPfqE8UHKH8B7q1hkEXORIRjXMS0gCUd57ikDN27
BBG1owm4683/BSYayiKTrXY6TxMsFQUNAfpCrxn+NbXO7j4tuD+BCC4W7IZY9ZhTfiGPP7vNlkye
/Y4PO3OzrbUOXD7yE3riI/yXY5cfyioIRs1zp9w9y+3QBMRAnBg7ZFKMJtAxIMdYOrXFQDC/PkYB
LSo8+5qqC0cvCNFdghgGNF+0Wo5Hb00mWs1cdKvmerWinehVo2CVKMutVzZwvdlPDjawdqlEM91k
d7cMgsyOA7qGDRv0ngjslukpHSq3dkR6VGLJ/asmmvAsllY66s6QqwC+ClBuhRmfr6ezA5UyBA64
M7itb5vrvKfc/cBX0nUFnwXhnOki89EuanXEUDW/SQw1yrtaO4krQqfOkyVqrgWuyCZUvrasuh4z
uHIzlgyha/UK2PnaqVUD/qB4qIbok2SsAU8NnjR2cvF8iLK9Wgm5ElxMiYjCLYnUOETN5EEEFFes
3o7tzt+G2iDYcgs7j2MGqoVVUJwjw5fCDSVjwqq/SxvpIsV55PBx1i1BzcEA2mwTil34w3q/W4Qm
2TymAxwE3a2qeVbzCUYIRUR6ns+ABFz8UncpwanGMz11SzYMZVKgSPSZ7LE1iYsIkdhtW26Pg6HZ
7fVIGSuVopbqGEK7B2x6fv9DyxZEHBOYtK6GIAcmwVdmF4/jI3KAIUxlplYiLaqfAFP4b8dLagiP
01T5FHA/fLE6iivmi0qCUxnoPMtkk3GDiFItqqYffNvwwnJMHL5kEL7naZF273eP80AeO2qyCCD6
MTmmbpFtEZwzaW2MHTxWIrA9tXuojYaGMhMaiJpMPyogRhiyJf74mxvN0HCS57a/8XzApTgC7eL5
vpiV+t9LVqdFM2VxPx7eV1MCUV2R8rcRso4/iS0wxLpV1/NcEMqjzMtGNgw77TNrZ0NpLevw0kRY
zHpM4TmFXthQatpAq0ddHqzWV2w8AJ6C4eWlq0huRJqSkpdgAeNbjjLWUtdHX9kDoOjZrS2JSIFr
w8ijcZYekuas3RX3zsvBLDQHL31C/fM+UCtmCYYoheI+vJLpGstzDoSy0pDBvLElpxq7Xj6zRRGj
7iBQ3nCA9d/5MqQizgVaTnqI+wZHFeG4AJirr/Mvv1gNUGAMYfClcDGp2WZdm/2BzliitOveU4Yh
ApugE0KLlOFcDkwmE/l39XHGDeP++9XJE/E2n/Hwuig1jvSel32WF4MSBUUUpw+KCJhPYa4Mq89Y
Knceh94JM0/o1p/6UrOqGlJ5nVPOEddeK2otZorUV6dJNc7heCHhkJSXXqHS1x1PHoNkEBDPxk9j
4P/CD0cQ7ReWXU7lYRhSZ+L119TwIe8/IDsLP8/xX66V8bg0C8SSjWMMmM//mM5qmhXH9ZWLubnr
MOUQz9W7kU6ZtK92fR8dIQdWuVnJY6eATr0fiviAoB1qo2g4QPVUXavlq/7k1SAJzr+z8O4RuZI6
m3UUnQeZ8enwvgTDlGIqv+8uot03Ans8A9FJo2C5WbqXZMahfzWsi1r8/XSMiVCFyrbY+NDMRZ2f
4VpmtjTqr5iIdKKFodOMTN3mJlH/6o/8kTMhJpt7kYIhbztL6TZInIwvV26qlkFye/n81xkmF1dn
vnxnhyKs19XMrQtodnLw9sY6TCHCgoWheIf6eg7bpAfr8aOAGH2/zOPUVPVcuSH6VdUHxQZrB2Jc
W7NyaWGR68qGuV5xiWn+PTDzH36cpu68iJmW1Vjb7ZMtiZj4ZNw+v8vv+z8rt13VLWMdBrQIlwjR
jQ6aTuxg+X0FX23kpMXPzyod+a0Hv9WoeCPucJvlaGBLS4/pCncx9DQOavT744C5sf2BXgL5Og72
Zq/zGADWOENE1AZJbBdxlUo5BeRznfMJqjR071VZlc8rEGsLH5UNouH/w+CAlEJbDDIZNvoBRstW
cDzB0zJjnTGO1i3UCI2kzBzIbi+DTogZbz6L9OyhItT/5Jl78m8sVSFmxIx+y6adeJs7Snp7KJu+
pmofLJhOW7jl8DWcpqV/HTPrMsEbxDbowzn5f2/XuhWERBU0htpQnnBnjd7imnrUdenSn4bbrZnB
6s/q1XSIhOh8twfa1O1tlWFBZz3EXIdJJOfM4/wtqMr8XpHVhCsPXZU9Ib8FTcGoxmjMvm4s7VOx
piFgn/N6p08BnmJ49VLpWpeX9vABmHQ3qcH0c21ty9yQ1Bj25PjJIfKRrPXseueQfH2jPxlCCbvm
Rmc907uAa7W7xRmdoj3CTkklk4ebjaGBpnt/iun2JR0sxNJAikUn5TLtTMedvtayta+TuNIkhGKv
CL6rXhp8zxyMflT5aWnFd2IWPwPyVWaMc8+4TDtdyUfuoalt53/Gg7H2lkQPIVGzpuaWBEheddFL
/osRP+LmPWdaTNsRXTKn0puv63ckhWSOkk+O8UglB9U/fOGvZc0xbtwowMr/5NbFzdXC8A5KpKkw
NOVUDmX4dnwFgAjwfOyfFyuZqtDTUW8GqoAcA8zPyL9mORm/aO/Lx7At0AsM3fd8UZ+DQKPEpGU5
SXx6k83pka7XyOJyefxKlDDxAUnBOs6eSsqAYkGr5AkNv6gts+uVnBfdr9xiUwPxBXlAkrsi5UFh
XiFV0veMSFFSpNBkQ8V3aPCIf8TFwhQurHLWM3P+MWhT4dN5IBoYcOU+0Uc2/2GKbinr8DKom7/F
5pR7fDlZQBx4HIC/5AdoXl23F5Vt2JnVC3rpIHDfgUfjOXQzZR8UT3vcIs+xEhqAY9eA9UoIzULf
e5DFzZ+oxlpaZMcl/wImlGOto7e9txiVjSkL/KXqqeINUaygOF3mnYvcgDLb+fmT2Kt1xv2cE3J2
BR3EjzKYDDPSbDVlU12o4YnT2A2+LZCVX2E85q7xZViE9pEBcO/ZtPhwEzlm+FvkK3rIHCGdWUq3
aymI+Uom6J/EWoqRy6f9hl4zmOPi+2KR0dM2yFP3D0z+1aZazLXCQX9Rutj4fLVGZj1cymSiL1uE
nVGw3y5YPCiqGgvtsRY8awSU0862d8bg/vz5iFNLczAPFQ7QtDtrz1AmrNaijnn2/5xyRToHD6Hf
ZW7RP4ic1WFtzabAI0t5GMxIxAroYUQA5EnppIPAh4Jn5sHr3f99mTISMh/sDCW2sKqFmqSXJtue
Y8q2GwHhY7Q+sHIETJxwNFrYAK8J5PSaDyLwhGWP3svStd5W8NPcSL6TnqjPwZl8y2HHeaXQQSty
/hOcOh/43SpMjJNGnyJhO9cl5ML9RRusD02iR7XyJEwjoXwawWG/gmgsyl5ZIMITvZFAjh8dtkAC
i19udqHSLFYcmBk7SAvoLtOLVOTpp9vK3rF0Ssig3d9nXN2+EA80ooEJPqtJ71FluS+hGAsznrlA
olwQmJlwnvlqFGyp9e+MKFAqVfG8nG6Kh082FfyHFkF2ULHjZZJKtIqP45+z2/RMQL5uEOo66s3p
uhVGBjL7seIH/vO8bVYf6/GP/QvOJeTtGiTavhYiy3WoC2nKIZW/id8a/tkhlUy48Np3IyhQtEoD
P/q43GUlfm2LdftMsRAuNdVR9mepBW5fFVt7cO47t2oQx/OVUiDoTO3PGpT3PzfmCkBm7z/g9Gvp
c90GtUJyDO0xpvbyDrfg/V2Cs9prmiyqwxDffz3YDM8kYELEr8Ye6CmcQx9xExJPwEdK3q2h8XtB
BRROOid3NfcjTauU35SVlDAlMool/+jAqQRUw8RnaKu7oa4I2+a+QZ0fqR0zO7t3slMcea9cRziL
aEde+0NzHhyffKQmqPH1aBH1fP6tRFN0l43yxUPB7YhUIwFUFIBtFJIpyXt5CJuRKimei3srNTG3
1GOmUDvAEYMy4R4NCz0LVHg3T5XhZPXIeFg5MJfoL0VeanuPHTSF46NqbcKPaFuU9Ii1sCm6FJnL
HriGWzIzZkNHpxBDXVPFizkQtvsfMVmHD1ob87S3lyD2IJ9jPihMzaDLIqwMFgwjugrmVVU22lAc
AGVtvpcrHOQPmypjRO+Jotbs03QRTp6uuOvBxdCTvLI7wpNR4qvtvWGS7bSpKjI1aV8nw+OrQVnW
BVxTvvf3CsdbHEofwNALoHn8oHbuPxrxULlpHmFbksRtcNZDqK7XfOYppM0td4+hvMT+BWCq+r5B
sLCZVelJ7GpbLL75REBKKX6/Grc67IX6cAjt2rax81vSCEH7C0bNywNenm6ZvaROSMjHTQRk4p9A
xyTjK8SWjWLBdL4i9/tOy80NS/qPgGVB1toUGz6ZpPLvNjKfhqZ3ExsfkSNVK6RAfC5Y3FFK6fWL
KzIK+6bcNN8TR6IcKmZBpNOXjlFjCi/31CSgTeQ3iIX6DPh6TSYvzhzduLqCymx39RJrScvRZQif
5bC8Ke/lu3KcxXqFuMUQR+Xvlzl02mHT7oflUFxjeGRcy8SAmQKo26wM0MscXWGBk+rfCcpxpR1j
Md1/Lg8llwBhckd5KRd3k1n4KPBIVSo+jWR1DcnJYgMeFF7xf9L6aUzXKg1oYhaezDcjtBKXsB5p
DpRWVavZl80AyuCHydTT67G6c7pbtBnDPbuOnt63rBGigXAgItxwa823/X9GnJLLuc20R1FCKz1n
5UZnwpMt75YVIvFmCRd9vMY0fwjSKiuoBoqYlOy4so3w/LQhXC46mpqTfmCqQDNfhnb5gdcHNjbM
XVBgPeOUxjFTQP9UcK5YF27cV9u3egUoBSCWL7JuhPLUdluxc9qxkils1YPgAgeTKNMD7OvRO9k7
zhp3K/aLgOujMFxDiaN4QpLHhqqzVFGBbwK+wlsK4zCfggJjP4xu0/cr3vDAlI6wM6Y+QdVGS8Zc
e0Qbkdyf0cGG6vy9m/pCLaiR9tM1O/GIyNqHXQFjPTGPDKdADmw4h2blJvyYpCBq2uqp+y/WM4kn
v1/YUh+ZFhEQaWTD5JzAIQYqD32QMO/x22odZk4JtAqpkbFPWOPYfM4MG+lsvlgphiwDqRca5uNo
Q1zYdD9a6rQ6IowiD3o1Kx15mNf7XBlw4NiCpTxbafuPe2TY1+s1tSD9Y/nDIOhlc0U3Fp8QazNo
p49nUhW4Dl/hwqBdibj5UwJmlFevKOvrwIFTFvMWCEIBrsLRKYG1mNGkQOv+C3OW2PdBkRCbnJPG
7hpv+bZWK66T+goUu5WU2jGWuDKTCio7qX5ANcyxdjOZtErYCTnBWZTl11JMWxsiQUwVAvbAay8l
73jdYJ6wiRGGJpoIocMaEJ/r2p8ux9k3Odh+Fwya4ak9FX9SFosFPF5wwL4xFwFvKek9R1cL1tWe
XHF6P+I7gG/RKTSsJt+Ep5iLdp45gf3pxd+RwXk33n8XmJgxnSbjTXQpk4zOCk/Omga/qvFE3hHo
bHBBPX7ZPfFPQwcw3bopeNqV0wQaimhvK6uv0vFA3IrRgQ6yVXGvMXLNEwExsKJB6zjTrRTmRvNX
fRhq71XMkJ5VaS11tsTDAEX6N8n3E+3ohsASVFuxOb6T8xDQ5mSrg4o/09NWjpEhy2v+gicBkreZ
FqlQF2klPaXbO/Re3PEHTgkiWFjssQHG3p+VdyI/VP0oI6jQGI/8J0eYGw7SFN/HeYnKiDGs28fJ
vBfyOySqxBwnDD9aiM5vdXlMYNv3WlI5+YnsRWOs4J9wsrPY7976q7rbYQjw8rsQ9KrG2nUCT7D/
ho6fP+AqisLE6hY5w/q6PKfpLuy942/3tRuhhqCwPsOkazGYaIp5wIoIQE8wTPs/a1gL6HveW4kL
29sZQkCBco1q6kLLEyKS1wzgoBxspJHXFKXbBAyPFyyNaJB30dsV+jTbOMxXKDYerXpYTDTu83+K
B4C7K/cCOAXc5w9mACIVUma5ftHgl00xeQO5aO2vNNV82xlVMpkUzkoBt9nz+OyXUi99ud/4CZ8W
Sq0xLvp+GSlLkl8MTTtdArptZ2ikrhSVtRH6tr3t3OQTvoIaprvEtJqirTjgNrd6LSrSqlhVlOGu
VI3Sm/zyVChsblSLBC/NiUkLzy1h4D5n435iIIFJGncuLgRb1gz1QTRUsY8XTDmJIvF1jlnis3qB
88PRPANEiwTMo4aI771lLNxiITqFig8YyfjV2yzII4AUOXB+PdPE3ki2bYmW2dx0Mjvg8yxcRENU
cx0aAi6+L2oxa6HKHjB77VI7Yxur71z/1KDVWdah4x8FFBSNr1swBxqUR4bdW+yg4Tu4UqindU+x
mVT0nysysQts3Gadv3m0kLlz92FsDmzpBkbZ2J70suG6uusEfNP1oAgiA6QIu2acVPS11G6qC+Ub
B7m1pBRAA1Zi/oQeYHxyt/eeQjG2OsjiyFxfflj213rNtTKwQ3XJa6nRqKBoE3UTNjG8Q3I3dAiS
QKfx5jho2tiHXkX/4ILPKbvlz5sS2D/GuTfm8PC1HTeuAxs/rOYtEEwGc+9d9vQiqKnw9weKAnWw
pobyalsFQH5gkUOeBmuHXi4oRZWJnPzeeAnyr8mCrX1hFFCg/D46OUyngnx6mVxrzAjB4PT751zu
gtxEHkgm29wJNKdcJyptTfHWByZ8SXFPwYxaCRZ8ijsuwvpDmx6GxRxMxpUJp2xE+71mhFP78S1n
GCIss3nEo/XLNlb23rBbLOEntrbqMUW/e68HmQxqaJunrk7ymck0aNnRVVXoFSf+YhCQ17yYrHBr
w+3tfTMZoRsQNYyW5z+6lqGb2bEbYavWlxJp0jQyy/ypTwCd1T8Ueiq6VffSCTKRTWJjxeWq9eez
T5fjetE3mpuVg5qeBQyeN7a7JtaT9W3+IW5YBtA2Tj4AkSKmbTp0q7KhtukRaNHMG0XZJQB2FI+r
YIOpDbSm9T8/q+3YwSJq77EyqpaspV39ZQcWEayBmVsyHPBmPy+4AnT/sF6DebTWKcIURaEcPAHn
kUSX3MqH41vdTxUbBQE6DxUw/WcQ/ziUpxUydhauu3AHWud35OOBTe4MmMYW7hgeFfAQppUWLLPx
4JSBzq3ajBrxmJwqvElzSCVjlxN7oMqzC2nNa9Un9+MwM8osjzu3LmMV5l7SKthf3hRnwZBYnouO
Y3h3to/y3mZpBQgBdc+ah7YdUfk4MjVgNkDWSeCex1O5mkbXNSsih9h+vjgW7SftSwx/azQH/H46
XRIbXPc2ljk8IN1U4UE+vp8/9lp2pPUOP3bdl/WD8sguxpSLGo9LFzH5/PbB/xWtMqBRZEwLIZiM
6kBC3rjZ5tdTwEtKorIALHMoKL9htawo3w4hthCXq0ibZxfLPChtpx9qAVvJFcv9rToj2nXp8PEs
K4Vny/oDoEcuu8N5DtOAoktbhbie/9su5RQooG4F2OuleyJgNeiURbsWC1KARqKIdOSIXBh+mASa
9oxDISol03I6Tj1b4tsui4U25jiP36nwfuTKMoHGSm7oj28bCy1okSNcZkXEMDE2xIyGKWhn6+iW
++8UMAKL9q84tgtf9snSDLZ/V9gp1bVBs0LpHed766D1yXxhm6oToO4zcUgZOa8KUagYWU85kFw8
FTgYJdM1PvVs5u1kQZW8htb4Sclcwqw6KzHLb/PuBPId+Uy79/eCZ7jdK/J7JgaqtVMYWWEgDaUA
2vkhtALs3SFaZlYW0jNTMjO1JrGyp5iwY76raHJH0OgIlFq9MhPSjWOOmLlYUkSwC3Iz8XPVFkkE
Y94O2T/fh/M8Y+wpVxDG6dOiD0snyt2mS5Bz2cmING3QsQW2VSWYcT7mgTvD7ac88U4wWSwZNpoT
VJWk8Azt39ugmBsBi5HFqwYVCUWnPDf6sUXsVoR8SyhJVSzqi434tMLMzs3q8KF1oMrINncbgJDp
Hd87/ESmk7z/BD7X+Lzh/2OScQj4SOWMaLHfjary8CEKi16CjfTcdTfgsBq+yI6ydv5lHsv9SZNy
zW0IxM+00Fg3IZ7nSACygpZhLJtO1N9JaXINcG6nTzECJCeN3WPssR1/QKmJ51ZGwHw7Ia3uxMhX
zcF6LHBlN3o0xkeoHiVyOTmKpRUb0JRFVXXxgZg0t/K+ifekfL89ADpR0YGWWMXYNWETDgLLJoTC
bzeUXrQlTtNDIsh6+E/lBaUQIXjXKlV5vnvKpxEIi+cOMJECHRG7jJwdI/qmAU98klJULx6x4vc4
Y3QHNxl5oDccWMQS/nb/nN3ll2DxKak6Os5/ypvgls/Vi+SaYizi5mYbasrNJNkVBoevEU8TAqRY
2E7FD7g1qEGQB0IQNWU7ME2nIWJ45tgu/DxcCbMmLauHV9DgMrCOv1oRiDqyVG38ifCI0em5+NAs
lB5DtDWZQltgVIHrgUwE++el0IwGNvyQ1W2EM8HsAoDGkBk3JBvMhqESdB6G1knHhs5gM0GGU6da
5A7fokJhFGEx5Ta6jitPTUs0O1wVfe/UP6kXYKCGA66v1roOzlsBYEI1Us2DaF4HkguRB7tMLL5K
0pj0A2A48G/UOpT61SUsXLRjKf7JvsxzNX52XwU59PTQ3Q/geaOLqwWfx7CD7iQzkqe+CxGhwETe
+oVnCPXMwHfrk5WFMVarVklAMsjFiyQwCXCdjujb3QBfCHzpNUJzU+ec22PQtAH3jSmqwA8d6P0t
cWiDOZBMxWeEaNkxpmgKXcIz+/Fd5zDeOqeBowhp7izCfDcHKQfAdXZrBIeg/880Q77S66ePAiog
85qURrEGqGp6C+sMdmmyi84EZt0/GOvmEX8whGJYAEy6ekPwyK+g9Rjba4/Oxih/ZQNmWJ9PpkZD
aoGjmqKSPOJEfFV/c4ewXENWdjOwknP7fqHdIfY7cnj01+JDErA/Sh7O0hoSgHwzo8hbGEtAJRZn
h+go8vHlkT09A/GBLEi9vQ1BlZmzt04kL4Ia6Dh9JPdUItKkIO/RwUMX7Ny2+50ak03wboWbAdQ6
FbkJlAOJ7vV4dWX2jHVhJ/1Dr8Vz2RbAFWAPdWcYzuozwS1jOjmmrGTu2kxYh4CPGRSySeodkP2Z
XV9gdKbZbbDijw+p2Cjt0uSIvgtdprWLXhJoFyB0jeUZ0jJBLKPNgqFOfkDXdWAqX+/+oxaXqPQG
V+WELj3XH70s+jN3qhn4fdwQh4My27JUxXluduNe66eHX50QmURj+pdt0AyRzdMhmEauX7MONscK
TLWmXhkxVrlnhUq72JwfA5mrpWwQk8fkvXg9croqQKC5Rtq9AKKkPo9kMyksRzb/Hbi7PASSFjzS
Mw3qBDKTJjOuYeMHCR8jkh8m+EOY6l6sZUhqmBpOAZLmgoKkdzBl7ITwPZ+1adarQdJsfo4DcC+K
MZpIoJXiZcK5W9fA8RseaQjks6396g8iBUYS/2AszlWdFobtjjezolB60TTREVAbr7NRTwrSZBkI
5lZJYCJdH3/HBnGmLSO5UA7JoQf2dbjPIK7fev3+loPi9XoR8gJl3OvmlYoMDlzLYNWj5XaL3l15
PZHz1EowB1MhcdOctUwSDyZM+IqrmNxgYu0Rxab3+vKUU9HLYiP6r0eqrL0wJYrneYzRcYfxTpJq
KjyQZjwnjUVUjXO13B8/2YyTUr3ykpL8JVXA3XdLErqROBEUBMG3tMWzcopt2JNDbgyq9pjco9Sx
QviyyYPooxHhW6zmOuxnGFQwgUHj6zXkeYjFO1F9bqQRZ77hsDIUDeDIzJpP8xzmTqclMEY0gZzb
WeBRBcjXTXDWPsvv3yHWGGZpSngEj7oHsPkymFn9uS4JEU3/pjGUCOq8RHY24extsm6kWU+5/RMQ
xak/gOM/BvKzJBdm0VmhV9eH9aZsrOC4u3J8BkLYQpObleyr7tiWiHKXJ/Sq0jZyTFYFeGX722kj
BClbQ6SUURKuMkJs1bIFwReLnmeGMOdQQEeR/S6+tSXlnlL2s5zbg575DMlwUZqyyLsT6/XFhbuz
bp4yxbZSYDTULU2+mp8h+hkTMy+wFD6HMXuWqsD3f8JQl3cDjUw7HMsmOKpJ4l9XpdK3vp2Bfqyl
097UdZ9h6B8bFVFLwswlMXRhnYl2keeEJ6NzPh6G8QCg+BQcWJD/Rrj0v+ACSKafkwuNOGXozMJG
kwqxWkyWU1QRcy9RegXn/ZjL+3Uv91YloNFNE9W5eZDUW+7321z+5NIqVnHqXg8Io0c4JFL8QvVO
nt1O4rZjCgq6lBrLDDBEV3Hyqv4kGPC9THEJ9VggKNblrvQnduKnr1Ky4L53teYxpu9eXOpwSMpk
BEbtHrZa6W2UdlX/mk69S4m3XmQNBcH7AAOGM3QYlaYJ5RQVbiVa+Ts/16pL6LTFjxAJkFBH5e8b
ZBY3Ez6vXFkoHxlVxn7KpJP/+A8+YzJVvYtsCx33YeNqGn556alfbZROD5Y3Xzk6gqRZBE8OPuGA
JM6QhIOQ360+SJ2fLzw4QQzUufHYCcQbm7MvpzpPGeQgPDP1aY+Y8TOXeylnHF3cegCcnp9gl4MQ
GGcWZrQx/9P7bL7UOy9tCrSzrKVzxeZulVaSKZsmb0XVJr3vCqGBQm+ddFJ2j9IoOQoe+zYLO8EE
6tENKztHVr6fiLyD5nFNb2TK6PKWbMXwGwLxtt1KuLTFyXbITpuB890GB7QIdOOBRCTRPWlDySIZ
lETDfRQg8ENYAoovuqm4QnzbpvBNyyE4ej6Sfc0yvhpFNEBl9DeKMQ/WtVv7tyRCqQpB2e5srPWJ
m0+QDlXW/Qwc1UsFw5GYYfszQKcD7j94+6OSqCHEsKoMRFXBp7JLiu3tylV24xdX3yQQBWxmnjSv
gLvvaE6YSO5o0sO8AxER/o1e0W2asYPsiwDoNXgIXzqzhHOHakU0vBBg+DKkUm4pXZ7mQrmZLUvS
AlPB4eelqiTv1Yg56itEWO7bjs7tD3aWBZ6YssUkHzn3ZcF5Afj00GiLll/RGLooWillEMTjuqOC
mwaszvZM+psk8v9rC5GbfbqHX6xDYLDsmIAJgz/DF4nIGQ29Dt1sfNPScY62FWPLqq1buqn2nglv
QB7lPsCh2T9O0veWmxTShZOMt2DqJq8hozIfoJnSRlYFvbHem22zQLTnhTmFuBWZm28AfPV8QOki
TTzmfI5hLwr1pIqyp6HzIaJYIIv1TJmsPR0ud+9WJUiQbFnPSfcYVF94ILr6u0QghGYtTwkrSfKs
8724ekU8+QbXStKgYl3PjAgKx9Hdf4Bfq0TImgOblN7T0F4GUna7jWLiaSK7zufP7e3TaM21tAcU
nbqNEE3gGv/KyRrytF1pdX3t7dFyVquuW5o7vILzFPxU6OoBLC+H+lMJ74buAfprlaCXneJsoC6Y
LcrSKNy1I40K2uqczvrkLUsEEwCqNsineLtX0DtZtW4Q4RprZD5tmIqgnfbqcZN0Ifz77eOA1Fmh
FHaqehipWo+xg7jO4E2Og7XT0sRrCQoFIHi2JKuuFs9B1QCWWtEcQiYegnh2pSLh1KiJccPgeqW6
fX4iUhc5eDQlij84WQWZVTjPdKrAe+PeLx5LlWLo4PvoJsaPXs0Wz4tOZI12KGkLD+5bfiIpWQbW
CFU+E0wN8xBR7cCrNIofrcbz3BKjvZfszBOs//Q3RtFN/Nhcud+5K18YRO3MLiewueVP25WVUkE6
ClbQT250h3/xhPJDeDBCXSd2sKN2hatG5QHU/HEri3TIL7T/JsnPcCb2TVdwjz1J5s0NjVCq6bxK
dSRQ0q8wxP9NwJt6TPsPYRqVql4cTGlM9kjTj52tS3ogZcajoUCwQTpdt2OHhalN5JwG4jLFyz/5
JKH4unIwzRJ5CCicos7LIYqiAssOY9Y/Al79UoKDDqri1gVFPeLi+7fYak9+9p5BHlYphad2GVMe
pjPqbzbDWBpBrEtgaNWazmwqg1LNbhN7tLroGeINtp3K8k07g1PtGWNrQ0l5VXzIiXksDGmX+Hhv
KEH9PfbB1EqtiBoa5Kv4wYzVzy65ZXj/6TWPYP65jVOUOthWfPzijxKgygw2O2cF57D7ud4IjljW
LEvAU1UJXNVwBvApxI/uW/h8uZN/5+LSiiNckPQnc40qnUw2wi3hdvNZxxVpFJGcNdg94fJWIgPR
mpKhllRhIx1Poqnp2Wvc7WaIk5FA++T+yC4jIBXYJsTjR1zBLwcMMzv0+VQhF95TVutws7xlAW8P
xao+EuLU5SZDI132s+gsKCiqM6u9c75/sKZL0vMOdk+O5VZNu2yVb9KBaGxSJ9FJgkhQJAQ1A3FR
7ZPlwv4fQqtR8yctLRySGY0R5zZzMVD6lZQiQ3E2VyoYii+6Q/jIk9Got//qM6KWFmizq1AYYTWU
3mZ0SHRGs8wTtPLN7lXXIsmOtQL0MgEkYSTstoyWB9ZgRWXM7PavM/zLhPfLWKCTu+CVk6pOcHrD
FQWZvBKeFVXXsZTrXVgYak8nD5UatxqQjpcM+9AHxNQp98bq8NcpNGQlKT8xQTuww/6e827Sqgqy
OQi20xBCJvgoBGrUypFgziEQH0rW6SC8HZKP25L20NL9o+Ap5Y1wN8eaWQKmwW8z+RTa2qRnWn9c
Z4MpHbu1aFbcmBE0w3rSFaMFakuvv4VQcfCDsOqwy/B48nT5nyYm8ODp9sxKo7gjp6/cI/1Dnkqg
T0K6uh04uqaWaH2PWkurf5bhuVyTB+D/3Mlt8DWODO6ngiHadbw5IkTzYXty4UBv6oqgKc4k+o9s
Z8g3h0qV4xe3PAvCY6oZ1fp3YSBAsiUlVruvR0eoYYH1NWB+GFVE7TgeMO6Zi1lybGYCwAYbg7ga
Y3uQaXJN/vwaE/N2sRCqlQY+poLw7KpLkKyMLa3OhILVhntGUWNRsEVrlra3nKkEOs8+FehkPNNz
RZgNa7s3ntzHRo2SZuxNTTADcYq7WfryFvP74ZWLNsFb/m94kIBeeW8AeO/Gb4bOW9viRxvsbGbI
Sh/LbU1bg73rPlo1/ubWfwah2NARGjgM6OOsvkIRrKSOlG1LC1+evr+dYc6PECqwwtzQtMXFfKHt
VGbB/SLBRdlo7aoyRr7htVYTRiDY1SHJ0CvQg1oo2zc8pTl3DGQeEKu2qq+tZn9xcduErYIHSeMe
NMxzkTSLSPwsB1BbLy/ktPOlg/zD4+TM0bbG0BP8s/aLXWSCUAqI3nZLO8buWNMyimckPZL3miDI
+ChIWI1cZQ3xihd3vD0pFMxsEDzZKxIRejlEcLJuQ91pEZV1yIgqvxwTAB63ivpriDhTqAUmnWPt
qQsANAyX9Yhk1U97EER2NF4bbxLdArzIx+7Jq57kOq3Xmv/FSeycudg0386fNkumJAyK8WgbCxPF
PrMe3EgZNTFAI8VJZVxkb+NYc/9ApeWTUEjELj204Jsj3l/TP+WT8szE4Wqxb0+GEPpYW2aMdNhd
FP9UMAv77Yl4U+WFDA9pTYFrKsIE4rMRxBv939ay4wCPQb/Qqd2qjpAQADNgt+7sT3ftjqx7aFaS
LuGMnVddFRtpVbXBT/pdRf2L6w4RhV0/tN95f3qoY2ieML0acXbR4JPg1kQCBGVJEnaTRDoT+3hg
4C31SYaF8FEOqr54VCADwugl8vgvoMvWUDsC8XrKPruWZ4+PmI8BLjLJszcq38QJctar+eoPKRLz
ca8153lUF2l2mHCZEv7hLG8C3bDYaeDSSjcujmWmz78QF3As4PJPbcIiegEtuhcms2gyJG9zK+Ag
iaUrW2VzJs9iUZsE6MUY4/Vi/NcPGc3ZC9OT0yObpR37tjMPMVH1Nw5x1FsRlMNTtAkUzt3HeQcQ
HPyhjBdpLu8dCiwgRnD0dc08B/1AQLGOWZj8YfyKY5IwwGrGFv4dWrcNhQswb2tpLSzl9VTz7ASu
7t+V3AuO3Knxa4nQTYmQPkGNXa3VW/FWAApKBQxuOqhunpUyVS1C/wksCMylEWBG748WWgX7+BSf
hQTNFOzV3koJMcmlio7agfuzMqPIATSn5SwYgwMEWRthCVts7hzd31wIohZ4frZnWW0YN7j4gLwt
4chjphmZu5e7PaA9qDhvKwg2U9Rp3RjxZH6hqU+TzcgS+KqlyZRNcv8Fe7r/p949KJF6Bphi6l8d
WfSPKjs4eVhbIWjgadnkQP8KQx9Q0iSF/AIORErOMYR8sAqZ0f0jsChrylJ/2cg9LCJgK6TmtdCC
8/3DrvIAXVB9WSYLXF4la066p6Ouu8xfc4lSuawC5aXqs0O2/aq0Nx3O3tkl7TB0pHLRG5wIhgSA
k6umt75UizJGtGPIrM+E2FrQcaJQW4yzb3FUWe47/wrRfiRXGJGAg0f1zkiAXDV4mELctYJcs1GS
u4d84K8fS1j2qSQHIzKjQX/jtOkfdO0steqSzPGjne8Rqh93PbdW+lwvQKemCFR6JWuzZ6sx0UDY
9FOAav2YkjluoJLqBuS6frfq0Ree5LHrNJdNImiYS6hC3+Rh9blB3/jrzoymre1BVCkZ2woi67DU
n4fqr0D0zBzX6gEBm9W4PhBAzJX2nOyH8fjiPAmePKUlcxZGqPKOA5CemHVPUPcM1Ac1E5k5Yt+X
mWeXYBfNvaFv+aeO1kLitGdDi6ARStlrX6M/spWyfxdGxZo7jBFzPusfj7iSf7HPTuHinK+Rvyd6
8MFC4fhfHE5f7pcsX085d0JYoAPefDKxoJaVJTlvdQfxD9mbX+H3VboK/8FoPOpIMe2uDr7QC2p/
lBrMVsKEXOwhdhCdMH8eVSey+r1yQ07uo/WkxHwbjWGulQ+kwN8OtIH08Y/ThSxoXqsDkF8/0HO4
U8H/XFeIDQK8+gTdQo7dzYQog/9f2Gxpz/NAcfmrXMTbyXfXEyzDoQN9D/HeIkv1+abKmtlD+mYJ
MGF0LSfJzK6XTUVvvPeClagOZjPdzZ9Bhky4v6iOjHyDfLW0t1MMb2+5K/hNklZHaIHYxyvK/dkq
BMXnlfgWgqQN02geYvsDFYUOTruLPU03HIoA0SHezKEkuz0bYIoIVUIL89fl/pz7FqAmQj6AQEef
MCXn3mr1sDuWZyJIJ42/4DDL7Hk5aqM9XaU2tT11LGi6kPl1tE/AxHbQbc+gUiPXmzmNoDU68wpn
9CtG5cnmjlJErY3op2F2fRfGc2WPWkOUxWi/9dqakCwO+Rz1Ld7uTYXyHaiRaCHyFodY2u5lbGGX
wKqUapUdvMwpaAyZL1Z/+aoy9cX0KZuRqiv8L8fknjw3Hh/2w5VG0omstUQD8nkhmzFf/AoJ7XWc
bQX/uKNuOdC1qxPCJInD0XizoH/u2eFzChVqZpDS3+p83ZCpfsoZZMh0++OoxzPPmURWYtpoP/q6
bt4GMLQdXGc1A+mr3VP0ctPfssB8MK0KOwmN7+A2o7LJH/dipht7aA6femwGjBnaE1oIj5xeEDfg
6vWuZyBg92Adrev6HPsD2OE1s3xl6kXlbZ3omtoYOHvrNBGBFE70iuiLcwKfktCXCSsMtbPPBfjF
MdZJZheVf7hYoiGUu+kDC3N7AyHubi0+d7ZuGvm4lCazIq9EauMFI9/ROXom9mJgzJBBIi0VUmP6
OtDOrD0NIUwoSjVPFmMUnZ06ZbDqy4TCZk+NJ0dqaEXnpRU72q98cG1hxDlLXTcoephr3uzLHLrm
X2g2UlN0+IKzbVK0MDiCHoLuCXIp3mhcJaiRj7smWqcmzbZ4W2eB5Gu2meZzflyhUsBQsMTYEL42
YMg4p6Mhc6bKoGSxKIdiwPfgb3tjPOPNx/a5gk683CN3854VSClVndH8fR6URREW7C4JS7ZwEqfh
Qu+DBtqZf8ZqV7m0YdcCmeXVQhQvau2ec10nqFO6VvysjmjWR0EglLbh9Xyr/Ia6nKmryBsVdnzL
6BOhXdon+eSm3N+7+A7FQQG8fZltWxTDBd84ko1iHqkuuWlT4gP2J680VyR66s1Iue8nQ4Xlt40R
s1IfgeVXegqvWl1kdJDhApNT5DRP6EXzBi6pSaA9iCWJw6ODerMzrSEWTSpbCl2ApAS63uDSE04V
PBD794LhZhqi9wFa08H1GTYPeq3Rrroe322EU+O6T/S4Br8Iro2iTbe09wDmSLOOxVfTU4VMVOT6
rXo7X/r5b5GbHI74wfiL//tHSpD0GFl+soCfBu98Lrc0NLryxym2BfVhdCdZI/uadGsUwfrtdn4t
L6PEVbWupRFh89uoLN4n43dcwokEFCZ4bARZcG4Wh4Iige9wiwelqC0MzWvJBP9xnfkqHABHYG62
oR+FBOftRshJhKJPyQX+KuxxDYkFxNqdTz53PYwbNOUGGSPoTeCC47vpr18kerYSUEfFcbMmT33k
RVBQ8bghopCed5FBON+HT3eACwnMfiG2VSHND1G/F4/8DR31f6Kf0Ppr9N6CfWwQ6MXzNfZvsI8g
1liP8aiAnjjR7vLXq7ie3I15uWgAsNrO0v4oQFkJbVc8Mc6/hdGVTnLEubgjNVDhfOwMrgud0u14
O1uDEFkEOSToW3fHyTMv3aS/SUEt/gOFUxpSxnCOjP5Ep1Cbvz5XHqI//XwEMLRWyI0/46gpa2HI
fPilFD4mRTSdrumqaIz7oP62QQ0mKUpsk45KQ35QSMK4RF4087G2PUcjre331FCo3BjLhMuQ3z2s
pKyLRcsnUqB4hXdaZ2q+GELfYUK0dw/8P16pG1wcFaW4D9mHkQPfYBuBzf6o8a0J6m8X5ts3e2kW
c2lEdnmUku633t/YrSPGuN5rB3U6f/ZQDII4fr6vbgqhhXNpaDW93/wm6wI1pKTtt3s+LbDzcDC/
T/ed5ZccJsAr/H4LeiWzILZUIS0Z47zSdV4vr1fVGnhZb+b/JzfWmmmUCioHsXhTBn2Gy2DeXJoZ
mcgKQdh9ZScQ/JF7VTfo1tlqwncJyzD6TvHfh6WxahJEAk+jTSp+TjSeFCJkHkdyQGLU7TUumLhT
S58jlDIrmO1m8Sn/rV4NRqqKcDmew4dTE53LtZHWWlNtbb3pkOamZMjsPqZdnEMY/2azKrktGyyE
WuCs7qxqmWsKAuwNswfJVnWFZOKlUB8XbfU0VnTbz5yuzSZDzKjFAFTNPhqPeB+cftwfMvV/qhk1
9hF1JdT3fn6EAgKp4ffbpX6NoCHQd/oudo9sAmahkGmIF9lbqYc7hXoLW/+l0Ra3Kt7ROxja/VAW
ZCmQS/hd5WaXXuFOqt3z+s7yJf3DWpff6MlvLSKFtjmB0bm4Ntz2CMSbSA7v+h8ZVnB51vhzSKNo
2G79ESrnkf9CZfPUHTdVgV62upZQuOCv6vI0BVTYIlX6WMZAPLL2DpMkjcPlPwuhwuxXB5U/kqmd
go2Fz3aK6wE2AczrUpOXFbAJY7mXWfEWDKgfwtL6AUgJ2j/rByUFkpBOAKp0P/nvoJ2qBgCi/acr
RkZewQjoO/E29lo8mZ+1bQy31qeTklXTnh9SkHFtwhMzeJ/hu4XsZece/L/eCA4A7cneGbo4kZCJ
Yoy1GyjXN4SKuuRp2nP5Vc3fQfsqVV01bqwJHp5udDo1SuYq4tH6+dLXQl1+Xh5Dy/5lGw4Ftju4
W77d+3VuAxZyWlKZIbJseZcirl+oFl+TlijKenAgWnIax8HxjCJN/mnbJ49T2jgULyAhzuU4oEe6
/OwpxvDwpiplwfdaOmqvZu3ilIVaq34tPAf2s/V/eK4hFJj4RLpcKcSshBueLYeEhlC9s/S5owjH
zOSqBW6WZ3lGgvHDSqvxyTfXbZv0OhVxCsKkHldNybit9NiDtTF7wvsvgIzpnPCCjc9JNqiqWmGQ
HPYctz8iheVknIzy3ybi3ho5hpna28BppqhG6sPVadPHvjjSJH67dDQTTNfnMC4s7jQHQyD47B5w
lgwcTnsXa1a3yigcfmiflsIB6NKcGaFqsYvwabbHqSZL/BV9uLesFIcuCS13TIGD3fTiVxc43YOu
r/pTccMzLor3m9DtYYZPv7HYAGtT0XRxmazTnG8BfMfIVfT/0QqJBGpp7KJP/9Je4zG6B0ehFlKc
OcsuX4BDOqakoOGl1s9RLKmaY4pbblfA3Pi/ENaJ55cV5T+A7f5Xij4j8wmSU4RxohTUl6TND3H0
RksbRE/Cc7nNyn3bRzcvWjJeEAl9eTOA+y5vbqeOg+r7NlorIwkUayHIPj2mthfhnVNqaLZg7bK8
pqzXfFrJMDeOtKauT0tbydnujfkctLzDYr/SR62hDC6OKgJsQ6mOOVwqm1HUJY4LsmQjYpaCrtrK
EpMv3NKTW5aMfFoxQeQ29BjEHzWNwFfgcIEhsz7hfizIsVWSXaOL29YIq+xSgFLB4jlian1VRJ6u
r8iNASLeBQYXR20B1kvRCEUfrjXjegxWwXkVpgLQXoJGXbS5H/Xa5Z0kfkYzEcWEncgQ0JHcTdFi
KRGpMfZvRBrYVuzku3zNVu2kqZ/w8dk7JJGbiGFUEk2YNyeGxtVEw6SGezO/Ga7I76OM0rpQA2ah
1heNBh5KWkdoNig3E8nRzkK2NSfp04EFbx1rgcSZn/NSj5Rf3qEV+t+oqopQG5U5m9rnSyUlSjc9
ysjWW+QRmIyU52v4xMhUUVB2lPYzpGFyJUwB7QDbhk9Ce6+NY/s5uKPm1HXIdt54oUvCK919wOSS
oPqsJuxiehcn9rDobiJRuCk7do80vmbntCwIM9VxWzgJ9KaYWQDomM8UeTCHYfXhvOM9J4UhceyW
RH8vfrS1C929DUwrOe0U7JM2T6x+um8GVZkQIcZisQgtbyIWZFd7b7SLp4YrIPSySsSok4T/ecfn
vnkD7O4oDdT2EDmJ1+mkbg7IoPrvPKjeE65wSkuBH3cDdb6+e9LPKFOSeL7JosNjOJFzXXvR6+GB
3ARujF4QfUCRdr5iye6xWXeCz6H07WTsdFKVN5BO2g4KutdPxURMLQ1VamaqBHR89sY0dwN8m2ia
s7NQNHdutK9nJSPUAWi/LrFsy2dXaZAOXsmqA/3c8ep2+nRG2yK4Eh8804vidPqEYCRGZwgJQWgK
kj9Mo+JcslWi8rH0I/qqqfR/HDOsULGQVJwkSMV2zuDPMK6oSWJ80TOwAC4fN1+wz1qo+vb1eBGc
TFZRyhayuxcX9jS3Lk1JRoPfZK714TAhsoZO0LDiwglo8S0778J6hGC8uCDoGN5j/Nx8WknY/YXx
glGlXcmgafuq99GpDKM9PvlNzuMYmXGGTQZFQAPqVx0tmbpiRXbXSo+MQIREl1MlRvI22ZUUfIxK
2sXUQTOpYqrt7qYUa7Ll0slNnG7VRdemIID6/rqLa7YDB9CjqE3pPqQcG0wK51uRC7LEzLUswl2D
qG9J1Fq+UHdBUT51bdhKqWrMgpgAh0pbf5GeFDEV5LP+HEGt2ducG4jPQiDZIofD+e7tvW/90Wbb
AgcS+pkBxK026rZOxHQHUnbqCyn0AnWzhlS7hH0Vls0YfkRJtu3CPCyZ7IWyuFzJZCymKgYz7jsx
0CSwLsSgzKSirAP6P5Ak5nPtfDZBUhYETZE9htPjPtKriUXP2y2vyHNa1AwUwUJchoPIoyYs2/+c
RmbWfew1fK6wfVettFIXDgZzPUoiYlr4sC2fVrta0rMSxJ2HnjCjKumyOKC/0Z0yFENVhZbRj9/3
AYlW2S1Hh/GFq5Y3F9eke7Y8ShsHVTvFUB5/vPquo5kPcCWQNkTJvpL2NNvVZa2J9UUT+d1MvwcF
YT1zdu4AxmRgu45lEsNlyxZkKTzCTzfRYivXHJOIeQ0+wgEvZLVzuGyjC0qq6rX1xG/Jznlpuecn
FgNh9KcMWyOVxI+EbQyM3aqldJjO/2h5mPyUw20PxHB5cvFBvPRDwvqN2IkunbVhz8VkZK1WSjaV
nfOEjJ8UKoh1qwBH6Bg7/wEhklJGxpZjSLGcpiomN0BlCaQ09wIfjXewmxVb8K7b1uCIVT0zBHcB
ZNPHWcRCHYY8/KL/hJBHLaxlgSTxbMTbR35trfAylLuShegsQDd5zm11Ga3G8kxkky4xkyAtz8Li
4FzeVR5tls8hcZLs//0lXgn6cJWYoQS5yySVCnqqHZMEtCGsJbZFPvLcpFVKA0CXKS1i2LNs8kOJ
rH28QCsSaNoBtSqavGykLnSEgLNMzF5kz2mM181C8NNO5/5dlDeNf8sX5egidB8F9+k/B05WherW
rWarcHYQ/Pfm1fe1gLoZ4LiFMS+ADpvJ84T1agtI9bLyp64lrpQRYKEup2H7iJ7OZW01f1CD1fiJ
Mb9CICRdM/w2xMOTkFkxrgh6tOueGfPoDFYoHudp7Dy1eElnRHbjcbWYhbC6DlZ2bz0pCgC2Cg2K
9+LY+8jqABN9HQ1QTlhxW+yt5bm9Nth+JvtHY8RBBqhxN3wMGntSEAZDw8FCcp/8jDmc206XYBEe
j4LNe6CDmovwR6bLv7sTh2q9UG1s5UxRtGZSJjWMqv7W/tNmDp2T/JUKTrBD+tAIEjZPaMJfopRJ
zrM9URyzg5tYEwlgFQfb7DZACmq0mRsXSVSPkccXTutvd5IXqodFJ/YIGL1e3/XrZjS2qiGVvM+L
+t66aHfkJzZ6ZqHCzzTrnmrdioYRTBEJiD+vfHSh272sswMfyvgm2mYs/FCdO18Hr3N3TlnftuEM
zvdw4i1yBMV1P0jwDooW0Vq9AK6Z3i9PPGokaZMPIvL5IbAE34mmrJnyVBwp55as9+YVacvw3yA8
aDkDpMSMTHL50ORMU00Sq8rKtacjUD9TEEW4W7DRQLLzQ5xzZPyXXzKANmUzmecBE/GIkkaPTkbe
oe0+n8Ij/SqUIa5T8x5K67TUIXTjVbiCoW5QfyMTieb1U45mXCxRJjUGh4x2bHhLCgT6IPeYTiqT
vhVmI47QYMNmMxr92YJmKBctfI3Rz28cSwvO9GBYbJOoq9QCNeBTzLhliiIE7Wbonz6DmdwWKRHK
fugDcECXKir6KTyMIg7JfT/LBB++SXUJutZ/q4al9o4Jma+7S+4cjoo92jl57F0QsMOc4f460/RQ
ThMu60cQssCJalyKdAFbWitmy5Dz5y1RhR72Nb/YCghyqZZStn9jsW4LqMkx1YRc/3erKNwGZw/R
ZZ8xKGbHFaSR1ebbBHJ0FjuVvuKWFYTeAO+N7sjH3ryjkTisK4EkajlZqbhp9nt1ft8Ch7GbQgSg
yQ4i9QGYfbr7amXDIbpGfEtOVKi87U4ryLuq9ujWUDg3tSErD5AGQ9gFiA3N0w6MNx+NpKE3bYs4
B/fALX87tI9D3d1kjEPpLUhkPw9fmW14nrhEp7eKLejZQrDDXhg/FNHfZJWm1PKQLotiJGGGuvmy
AJRT/sTKbbGpRJw4SJUAoRfdcNikjd3BVmnXu+Biq2TFqOlj8FbJRBd4E1+0VyZUVK57fVgPXI+N
fH7cAvngmNFschCKxFS3JjrapmomKsdxTn+mKsEF1sluYoBgnJOQKdFi8LD2puOhJtWNvgy3uQHb
AB2aSh56c/3dDrShMkvjYTL71LnNen71LX0UWETIrL62eQ9TlIZW1hOPibkRn/VAAOdm6VT/yKGB
i5X4Yd6HEWqLQUo4E1wZGuwMkDwHTR825EhoZHRPOxLwJKAXT7gfhUfzT6KGe2Wi+Jx/kDpsaH4i
kRjhGfSMGr3/g8MikCZkN7NEpMTdt25p7xrpa7e9b6GWVoTkIlI1QF6sQEVQ9BTH2LzUrJQqf1fQ
FtuTF5uYDcIp5Fak17httocBFem+Bz0JUWfy+x/mp5qmGVyux4dsSdW5TvcMPeml6M0IRola4kk8
rB2YLqqv/5wsM66ljCjA0mbOR1QOjvFU762a3dTRh3WVVjRmxJ9hl6uCZA/Egx6UwmULcICt492+
4wMPCcLR13TJxGb+GMqK+cC9VRv+kExo5Uw0kN/i+zZ19T8qrylQBkhu0XPt8nfHwzQFPstFaomt
B0HWEeyx4BbmKhPwwUjezQrVfh7l6jrqD6yRKy/uy/9MQU1xsmNS2WiDuZbVYqhzTwdgrOguhDPH
ylJCHNhCf0GUcwBE6/kXSQW95t4CfsAayTs+P/HvUXzGv03wo+cH4xsppKcNHiHh7MDEGYDWnNNp
V2Yw1690WeF+JDc5Kq7DrGuuUxZM3Mxj4YMwkc1phj+NsiUsLOGrdV4Pbwv+mvkgMIDnP9+1QIsk
2Sz2yViGhBn531H6gUn7ujxGq2amhStVKUd98ot64DHdHJqAvY8sbY7NwOXot013WJk+5+m2A4Wl
F2ycAr0BiVne9qv7o3aFZ8hcxGojR0vhgGbVK1iUeJbbg/Q16fzdhlAHHCj17JgYjM7v6ezoMmVh
x5+LWpU3YaCYCP2w0YMgYTDX1CI6F9vQWRHfYL6oo720ZEWUO5JLQqtSiO86shuO8RUqeyeTtLQ7
D7LfPUOh1G0Z6cejiJzvvJSsQvGnzJkjyx1pW1nrgjQE5ulkqUKvEHoIM7ghG2rxTYV+YJ4urZu+
ptmG/hxjX2uzIBMSI9mS7Y2GVkwdR772WL/pkiDVgC8IKxXNT4sJEsxANhON9QoJSwI81ycI1GOb
BKu9vnrhlgL61cZjhZR/nW0k321ImYdsBX9pJjL3Gwo99CUeiU8pqfJ9f5QmESlqirROw6okeL4A
+wsI0pPqrC2ZgeO5K3ot1sRIev9GfAo1dhUwHf2pYx7uNv/OdDDg3OjKbo1TPLCdbGv081Aydg3B
q2Ha3yDdYT3rwi9WjETv3qBB7Fhd76cX4e/ubjQEQOtt1Ulv/UwPAyqP6zk9TJ6EbM8FyTRSmL8J
lVhELFOFgliwDOKb4LE3SoTu0b9luMdYO4/lUTQYvpZocrmn03WKCjYMSptFegpCBSsL18VpHgM9
pN3eEGO/A5bCSnjlEe0ZHsxCF9ox78YtRdX38BehYwSUKaqd0SoYvIL/gHUlLB6PSZJp8EZSHL+O
AQOk4SNJV/WvebVtRDyS+7xst3O9iOu57RGrZKv7hH755o/UB7qPujSjvfEthR2z+Iu+9kO4JBXn
+7LdxZKH8A2c8G4RjPuvkGsE4u8S6LaQgGAScS18AipRgZLZPOQTiWHuG1BdhifvEjYmceKUr2I4
aLs3vWsEeaikcxVP10aSwnJwDsDNLmoIfJkhX8kVQXSamLZXo6JlIXxrYeCfzLg4bO6ckSZ/36ql
QzJuE3VP/gY+T41HDVSIUTQw2XKQcqXJ4b/DK8o1dGLKKhX0jcYa/gkuyGAs4JJg3nZxO9n2sddO
F2v0QdQrqbRf8aqdP75vlzjQKJjyL0dsZtk4voNXVs7CDUybIT0J7/1V5Qq6EwCn4CHksKHXBEW4
5edOl5a/2Cpi51oRnRUEOWNwyloFD68ecesUMx2RbaCg3nYJu7fFdf9TwkBNIavclTN8oSwmUd1V
w9kyJ0ddJt9AGGBREzPj04DHq3BvFL5/doeT8Z8/DTwonUz5QzvTxSZsIamiYBfYitBKVDdEqfiv
avrCmsgY/hkfqSKQa/kJCejDVgbdhsvylC6PAYqKe6QlKN3gm9QSDwrdCq0qhoiibH85SdxImOzC
PXqZKJW5E1FI3OnnqykE7JyuN5GvKPZgDKkXNmVmSzCIftITBhk+RekXdvZQfSePO1w9c5qmsIOU
kUpRSnqQ4gKs2srEWi1TwFKgj8F10DZfNI6lMtfpNkSgUi3jBhq5fqRMpcaxic9sVmVrgHTSSvkA
ntctcNxsxS3hgYABJMTwHHXpB+IMEQJRzPiU6Zo5Hq1G3IqcEB6OfW48y7/TJCe8hLRpe4hkFwDC
D9ClOe4XJ8PU3Tlw0vgINs2tepC0oAEm+GDScDxvu80tko09Txump4ZS9MfED1zwcjUS23yRbFgf
BdP5nKZUFPQKCZd60UqYH7CfruuzRbVpd93qai2EQga58KwBX7vsTiRH/jLxlwLm1rX94CiuiDq/
SIl3J/YYYBXjTN5++zL3PWUXycq1YHCSRj5kFQhRwky62pXK3BE3PocVx9kxhUF9jtGPoutIUVJh
nALtdnxjIx/KXfqQI2tYRLwxvrGrmMBc8s5lcsOy7zPfiNs+RI6qrND0rg5nRyQpt0LSlmG0C7yT
OxwHPGoRcQjluvj1rb1tx17/ERwbS7KCuNGWl6nSzDCuPUelbZTdC+BEoCv6rCiFKIUJ5Yn3QVJ/
98U4F4zy/Mopcp3onROVcW7kqGaWYtb5sooFItlcg1B/MMLEFSnUpVWLnRb6W49LLO4TOKH9ksaD
FhtHlxYQbEnh/TMWXjIvEB6KbH2thSDzoBEzPA136XSo6r4bluPnZjW6Rc6yFdTWrCS7o9ODlqmg
U7TfgICSx3Y6HZ6cjNih6eGC2FZF/oKb1YBzwVyTgkJsdVCS9zwV8C8g6B1J6dyZDOTij23RLKPO
qDzfK5Bqbi/Opkt/+J1sGCgLTw1aGl1Unvokbs5Ko7VbukMR8sFH73EPV+gum0I/kq31obpuFMGB
647jugEHwCzUOLiuLde1FCFt5PxSMYGyOBfx/axQ4huxLWfhM90s9jE0LQ//tNq293Z3EpWW9oxS
pEp3I3nYONJnyzohrAhlMlu1PN/jY1/uslcG0y/V3MheB9Qvw7b7+YqBUrkd9XMOUY+BI+uWuDzW
zxiKPvfc3SPNd9fOFNPX6K1iN6cljcSlVZTtUcrq+7IgSebTPTOA7kjthoFwL7tYL7iFTY4n8igH
ryrKtsSEmsHgxpSe2hor9cdLraFVAGUP1YVkp5DFXuypoyN+X0mDihj18sIqpppsOBQL50fAvI5S
5wgeJU/8CsfY/Nwc3DMYtpZPgI3jz5ebieguEtT+OG1bzl9kUmbV6vUw4P0fOSn0E5/qhiPMSL3y
tA6gFRlYr1xVixpsj9tdhfYUEhjGCdrtJi2Op47SPm56p7k2LpG+ERQYBIvuIpbRPot7FUgxvBBT
72rQ9OYegLUVxT7BSz7MVV1u3lvJ4HVOrmMHDF1xN0f2cGpmj1lAXz1E/cG0EykPf/MNqf6iyCF6
Fw3dLIbcOgLQA/eoyeLOAYmepFAioQPZkHI+kcjuy0nBJHKDoocbv/ICzIcgnf6rtx11x40p+Qw/
58stMK/OVQMiA7OSAz7N5LLLbHcIrDraKok9ZzUEum5+IIyxHfQLA8e4VNVyU+r2cHYPri2b8Kc4
N98MDnzpKxqPdsGg/iqcR1e2PE8qumEvMFTQW797dUTcRvf85e4wbX8sGbD0hw3+8SJewbuqgzdq
C9iJC6TbIlpXp8XSXl2rFs/2R8AmWj3OY3DZgnfQeTLmVP8l8WGq7wBRi5TA7i4THat0D3EdxRTq
RDZE+MpybfodNAuIH89OYyGywX/D/bA/aq+9k2n2BKtNqnjr5stXLDjk2SUYXoLTFZ9TdBq9fxAZ
HloFfmANpU5lwvRU6D5+bBZGxoUCluI+WEU0/ZfL75bsanwHSf7YWPPv9hYArbg36IRmYY/Doz91
CPWDjA1uggdzdtoCYKn1MFk+s7veyyrbA3/D2GNesKRZZbp8XHQTixBymWeIL/WjND5DjSkH9xC0
hZtjGbkBJD+0BK+f0HPFv0OcVbPSdyBQqRUpwVndAky3DCQRgnEFTEvRfbAXjZ8wLXCIsbhpJypo
ew5Day1JUpawqGc+5Ejk5BI+qFAfwKHkFooi252En7ks/RVxIx2vI4e1yrugy1G0Xf61Ic/Scbe5
4xf4m/gb5VoELl6NYJlaPvdzOqs+l1WJAVYNUs8Om0H4CQFvJsBASSSXMdbb4FzFNnBQyMCAEB8A
85vyDFMfZFq+5YTQOx52Ww2/u9jRau8qlgTxiyPGdmnGshMxZ42a5bYTvAo9Ic1vN9yxe6DhOV7b
1zgmG4KucPaZEhfrTcK+9V2QKUKfmGDZ5RndKOcWsZEHfINDWYkNpBFyMqV00TeSgMjS7xe403Eg
j2FOjZZiF8c/OlfoL2cPoIAPXa63am8C75sgUXLSXfyomoOFc2DTLQe1Oqy+QTxf/PDabInh6f+k
dt5+PuL92TmocgBorBEih/hC/rQbBy7aLRWhq2kjXLInvJcoLRWn/05vjFaCVa4xhFO5s/RnHWYC
ZcEl2bZIDNuk7ifuH455U+Aozt8zq4iqxK6v57jCFMKhl2phJh8H/otlFVyK4qSIXTeGEbb3HEam
qxyiUMD2/P9Owj+BKfTPvM4JtcTijBFge7ZvWIlCeV2KWmGGt/seq3gUoJL1wqER+BLwLvhIZIcT
ZWCbO6jkhyA41ahbowE3AxLK5LsPg2zmKoKkYF7Ho08Cm8RW4YFciAJsT0aCbNsE4lVFS7UWl76g
cYAXaB6ZhBtB3uWhbng1oGw1a7Vov93unKx9kaMHRM9h517Dw/EYR2TyxpJ6mLfbRm0rlzEnS/ig
siUzBUMJ0JtLtSrj7punem087+xNHnDw8bhMA+Jyv+rMtDeIISfd1LrNmUDreskXAQwBn3jeLWly
7NwW6T5cb47h+dzCK965a9VeknsgUw6JF4lJCy2O5Z6i2wg8kr347b4crzZzegwAN91weVfkKFmp
M9tZbEnzkVYzRMSzJtSZkL1Ff/v2E1HExOspiSMPEnExEtF7VJIa12ui8pY125sIJDnItclU4Cls
Jp6JqUJ/c0LjKVcKYite2zlEIoVafYgzdaMBIv1fM5IjSAKfrfOCJlm5pXCfqiUUnh9Dtxk9ebNw
/8x9pybROTy3wMkoJsC5zoR35JYyoiSgva140AJ68WN68w24cZaGX6mN9wjeAIZvGE4b4qbPqYpF
oEbUwnZwPeO1dmr1cQeNwGNyts9+8v82FomTUm2QUcg0erCpRCUVzeP1eVEpMFFKyf8EMKViQwVj
8qwjqU6/pnV3xkIW9o8AGgfTcD/Sd2m2kuteFYVfNlesDFSD5YiF0hf0ZmzzpUDuO9S/yCe9YPev
QgU6GFiRF5PlDbp9Sec3D2eYYmuC1jiB5m+Mf3FTAbRqXJ/K83VaRL10Jj3MtoCw2OvVnzC0ADlJ
b4y3fkLtEw5uiB5f7Y5TiEPhoRqlxlLV072cpG7cBRQA5qQ4amfmy64we0gzaTq8PORw8buNL1DD
nK03gtNC44Pg3TZQdlNFeQXuTem/Z06eLNczunQ5JvsPnBHemz8Gx73AMmRpnGv3Khzo1K70gp1d
F4xKwDM1SGjWyNZiUp4gteSRsRKxpH8KwczeHl8LIDDbe/WLn0bG+vNHyhTUpNWZgSQEv6TsP3nT
VOLvc1p04iLfWrx6W9sHSK1afMAP26bu+MRR/y/H+Xi/PsIW/AgaH1/MzMwMQb3xQ4FI32eodaac
ZOrr7L29WO8mXCU+Jd3dsKqxr20n7TK6mNI6b5sjvXPWl1yjdqXnUw+dX7u7YABzBctOrQXN1yfl
PeFCZSKerX6EE72+c4gQSHzL/4Dp9WUAumGcSofHXbvj//Qw2agxptmq5fzW04bSDss0tbCVXcg5
ZglG/wKtzboQZthxH7H7m+CbGiDdkXZd1EnH66rtQ6KX7fAnG0WvS3pQ7w9mH+EYe/GcRcQ4GUYW
8sWG9v0M/G4RpU0ZIFx+iSvEEy+3rUQ1igTYPr28J7GPHZC3A/UXdy2bu7HdS4BGr8RuglLczM5w
GL22hMprrlxeyGeQgg1IOx9iy83LwYuweKnicBprnLpJyDCj0RUgPk99/yY99+a73MSPjDCVG8FN
3KZLkUIxtHHlXhYy7z3DUMAVJVnyZnmWMS7KFOG/mq/KYgq5zvFMkVRa07aTpU6e8ujdfemiZu+9
Z0K49LPapLc3517M6sKtI22C/u6mi4ECMY+nMhammoIuLHxZxEQLqQxLYhOU0vjUt+3D9Yyuq2nw
x5TlUM7v+Tm3qmf9K8b8zoS/xldAjIXXVbWbKAB9NYwq3kjx+PpuS6L0Din8A/6DihLXh5L5A80t
ZX/i7V/h5cw/P9nkPNvPo/h1owLmyXJG/3CAJ05aUGJ5tLAUBVzJbTPOuFRdvofHZmpwcJjFTDXV
mweozSI9Ji8UxdjdA+3y6o/WhlRag0fblAiZxEPVdqSV+xoAst5/JSGuD/3KQ1XatcKzVwYyjee3
S8JiPQlL33pB7N9Clv9ykPl0NuByFIXv3P9b7yC0A7JaFSlhjDBmFI8CuzqRwb6exO9EiQq/QY+Z
sJ9BXZxBAcG+M55k0sZqsdHfrig0GPxvHzv7R+Dp5xyJGIwP9qLIjEUgvG1hBLSC/JqG5dyY8Xg6
bvtzZbMu7eNf846rMMrOPTS3hHk0JAmAWhR/9RnL83y1kgaixLzxCHbbdLUVQNFP1N9JdvUt0MJl
GRZUwBzcqI87dSP2m3U762+jGPmLWEVRujD40rYv9xGBKKyAwMZqKKk2ZjUy8kqjc8Wn+ox8CWQi
Ruk2Yg66Nl1sOnWMAWhrWYSZv+G3n/39ZwoCTQs2Z66blzqbLiKIPP6xro+K+2JZ2S/FdbAgVxcT
ZyWKEsiCUdUVbr+pOqjMNddHy0yOw5syIS0CqV7AfIUZHxZg2oywmrTDjv55kna+JpMVSuzX3tMX
9Gzfu04eByrYThoJTDitR6U3LeLEOpewddrC9e23YZi6gfbRwrjtH57jDJoLrRp+ht+G/d1bLVKb
HqeGuzqVVade4VVmyg/6/Haz7KzkPVl6V5qrlEQCxHkkdpJpEN743tIoTj/Ppw97g0kkYP8JLfME
N8z2yVf+Lg70H39ymF1+AxEOXHC4EBudTnF61YSHt48HYgusUV6JfTN66eBCfOt1s7EnOV07lX+o
yM+s72rXIL8OaiV96aAYLdC6tYvz/itHT8QwvXgaNXY1vGbLvA+VGvWC5gLDnN6SHMofcFFkzOT8
eYk8c+vggFwB5r1bnyG+cSmBzx2VUVT2encAyovTdyI7Yo4xrpyCEyWcFL+G4GGedfGb2JGvdKu7
5GrD9PeB3+p9g7DD61P+F3xdLkwEmsB/MjlWn8YSDAN0gbswLJzl2nms1t0nSTlQhLeB1GWsGsbq
SYk6TwDddXYxKeWxWx5crA48R/jXFn0g0v/XihzeNc13WM9wnKl2xC4Xo8O9I8sX12vtjHkPVVUX
zBsFl/PV1oV8wR+npW40oWE0FVFOyLC8J0OoorUC09TUuchuCfSYjpcVU7R9WjW8KDH8PhDxImx6
vZJmxKEoWsyMk8rQVN/FKv9wvz3a70htc3xdgYs+kINJZ1oYa6YmaScGTL65rxpPw1ad+DlsTbg/
DBR6Dk/3DIbSyDowppe2uP6VCtgMeCFhVYlnpIiTdD1yq7g4KKtnoM+Z7cJiAoi2IszCZKDq6Tmp
xrDIobp/+2HhDdrTOxNwr/+d/eAB2UyigyXHUk9oVU1OsVnKJTkf3vMimNcHjDf06hIlBzv4G5Y0
V1Ydw6eFciWBDesiH9Y8njfw+ZgaAd1lyagOY1luDg86sJvP92AMHTBHxFJROyzOvpKaykP189E4
lNkD5K1HSYxzwIq1qgstyGh/9tufj8uCYJOD5wTn+Cy1G15AzgcJN4obtEaVgYExxo3D3qPcT7IQ
QtE1WpSgR7cN5TaP2tQ1ATfSd2xrTNDpRfh9huZeBLErcQcTJM0Reke1amKXIrJ4ZZvUoThZGXDS
TpmkA48FagnvYGv7rWTPivlY/Wb2OJXJ7pf2/WKG7Gr3ZikHKVB0UIwhIMljexKxexWUNbkEzg7N
GCOjjsltbEiehBSGLg1gJ6TXwonBtKrYkZ4ig9OCTw0GBcAbxzQ90Qgt/88J8AF1+XS+IXYfyjh6
dT1cf9VYEcIODsBFaXOW8B6BkbBXbUGaS+yVAn6rcEQKBluOKVXGBSfoFOVeK8WFD03uwBRru5So
sznKTD1Sv/aI0cuwUs50ebldSCFUKnTiZ8KrEq8coglKCS7mZaAmFRh5zjLlJOhuXV6Na4yfFYcG
alpY/BAOhwAaAv4V+5VnSQRRHWRQOmnJnINCe+UgnQwfC6vLsABTPvsOg1Gvsd2JixDIMyrMDb05
bUJAv0if4Ed8psLdxuqSb85gEzEP5sDVjrKF+MJIffFz54qss5j38wuXSJNm/3uaxRx87BmiSdaq
AkqNwvdxtgmx4QJY07hvh8bJ71qq9xQKFMGfe8x7+Zonek67cMLxOsomG5W1MhensF/Rmt35NL7c
eTbwTUGFL4tuHUpwcjcOy96SDCZUmoa1fX/3+3oo8IL+vm1WVoZBdhwL+L8okcF/DEkuJFrXvhUE
dl138F2951vbXs545Wd+r0eooktYhLqm0jd7vR9Zvq6/bXkySCuUUupUBBm/mU6nyHpaYb1yol7P
YbjdRaMdZgeviAH+zillPUPJAD0elXA9OxX/tDNAaYDMvbi3XeCNuvor9D+Ee3NqOb1uRyU2+j3A
NnaM/w6Vk9wre90aBBprKhVvaEUNB9rGbodObaU6iUlfZPiSx45z7ENwalAAZEMrBqy3E7Mc0PJh
lRLinoIkRLPlnQiq7VgnYIVesXjxj5ZPxoEJ66qLKEAeGoMxptTqxpqH9DjRfR/X5L3J0pShCUhN
qAv2uaRtwxQ0bqN16AhvuVbe6PltLGABDBo1IERplWkjs/CraRyFSuDwtUX4hVQApx5nn/cu5MET
b1bMfK8zqgSvBHMqk64Y7mt2TRE6Bb8tn8AdtH13dtFtGc3u2OoUn/Giouaheo2XhV9YpazpFsT3
BuXqLJp5MSYvlRNKr5Wv/3or1GXW6HCiMBhhWFmw92K4+9B4LHMoKDxSjNhNJHpbHCByQww01k/y
/UV8pZcCb54yO2r26xZRf6LqLRbE43gtgezoXJmiNestRdNTZNrLj4/6QcRwirlipYIxGqRfiOcn
MBgWBgFuVjd6tC0T6xhP6XNU98Ow1IQMgsjXk5VGPCBW4E9DjymECAeY1Gvz8SqZ+vBc4ODvjg4K
KvGcsSgHhda2mraoWzEteSU7AQ3qqKr7MxjkRP5nUVbgFsDuP3jnrE7CcjQFpV0yzIuRZHj/z5AA
N1wrOsldU0+CGf8NXvvqiChxum/RnbdQoWopEqR/11qi8nAsqi5Azqk6m+ItL1gEscQMd0vesbhf
HtxHbyL+4oISmPOtEPbStaD+lHiqlvxYuwTZkMhmMk4llAW+2QVk/wZWFrV3M/RQ/lTlRAr9b4oc
6A8Tfj6bOVTJ+w5YFbJlGe/J4A/uqZEOqSiL1gka+7dyUlypytxSzBU6GwNy6zbeUJKmXYn5cpHF
EddbCauKe1kaOjH0UqLPGA+YT2CwUosCRhZvomyfDeJYytavVwzldNvWTT4RSVvtZsAGvAHt6M8V
Tw33bYEbrYWfW7iw5iGKIvWZeV2ZC9tx+M2ylKz3KXPhGPGOaB6sLt/la74fGOrf9xTgYOj0KSt8
GqLjGLywDfTQxu1NrU6Yh8Z+wuPGj/PCHTdzxrFpiJjucjT5y8UcrDfg4DE0O1xaV32Uu98SwXKE
jv/diQRlxTULdUdVyLCVzeQiasEh6X0cAMoXqrZNfi4jBKM53Elvw2yJ5GSLJF5uk0HmcN/95kl+
tFEilDlmJhrxI3H1NsRR2QQl6W5xjLW4K7BtmA9V96xivXT6FdOOjQihutkbBJR9nz122AxtPIsK
2WHJIQARdn6k0nO3oE93Ho7icAnQzC/es+QRNorzN3SCkQlm9LHNHtUtmsabOA4oT/h0eu9Np9wF
Iz2DSqY5IiILMkrwQfraWF2MalgCnGi/EB6rRH9E/4N3uF6cJf88QLQpvyXUsAvrlR4cKiDi2mOT
fAFgYN8Cvr7YeFOEpzv1y6waKI89kAXPTMioGiQH0afe1JagKxNrqwagtufAD2NHzrZWp0ZXFBQc
nufAZG3eSWDpcJ12gRDl6xCjjeRuUof2aremXhtWRhf2sIpBDuhgwtntRjYoerDAzV4ICX4MfhCU
5kmaZTYBawN8Z8ZgBCeAucCQdtKUqUWRnVI5mjDJvwJXA/CbNL0OTcHNIcDQkWfhRskWnP7O0I7Q
ku6AJFIhG/l71Uf1seGsRsIxcMonLzytsTgtL9L/wpoeUiljM9trdeGOS8T0mWKQ7Oh1Fox3cmLn
njuedOhoVE4aGI0nW2t+cqmEeqZftW2QRNLcQGs6jc1t0yKIeAz31Q8lJjeJRvLVd4aExugLIMbX
hDYM0YtciwPCW5l0rdJv9gtNIYaY61m6jl0NdEnpE6LZELHmCJY5z0frfDu/CbEuRuFC7KvnImPl
D9ZQopOM7ev8F7Kk1k/zxFDZsdnAmlRkHkqUf9+irnW5/tE0IceR8PvhiOSxF39w2mKpARjA2fY2
0K00hVsNKlIVWoyZpwA+e1MpGnOPd3XhrFB0OMrTWwb9L6wkUieFXDWlo+0adB4lUsJ4P059pOH9
iUb+fHjmmq1kBT21uz2Fn3fzK0ePX+v6m4EBhcfcavopnE6TQ7uh1Q/kmPymuBxrUjx5cqlFfehD
2bq+9g9WuZFK9/olTvsoGHTmC2dlhs3bzcwlZO4vdq/PLjxL+TWqRWfvCEzvNzuYjrhxOsUqLgcm
7p0kqQSd9J5RJN6b7zONKpLiPNTcCNrztFUIiRISxpIuTh/cFF7Dxiaw4e5tVaX6BVbnhY/FYe4M
Y+27wBpctrkjl3BGO8cITYV+/YaB4U73lLzccmMh8F3bCOoMqhzwNDOR1WZAbhfRQFq7TgYCQbgh
lPJo/JB0GjtAQx8UKX0/xppnWzbIyejg2L46Aw3SO9hIbyYJyOtlFbJjFi4VvXU9JJZc4HFOAgfq
4HlCXvzKrHi/3LDA2wLuFmV4xWeFThacJHqxSd1kqA0Y6L5NVm9VonP+FnQ4hXRZC8jMbqxUWH07
pf6FLPULjny8VmllOAyuab6NRrt6MK+1OEmYgFgOMDc7TGQPQy4KzOW3OPGsu4fTNcfsqDuyTJJH
cWbV0Hym89XXqwORBc7HwqNv9HE8q1DIB+FRPzK0xr4+ixJjVwaRcs6hmmUv8tujs2t6w2Hh+nPr
C9W2TlSimQKxTn1b6Aaeqh4aA9yhIJvJzZOtF2eai+14lEn6FYkQ7w3Id9M+Mb3ZRzXs6s48Ie/1
M7RomR/5ZccMscVNPu3SuL26J3Hq0K6pXRGV8WvjjJC8Pnq0sFaBQRcj1Oz5sfajWbs4Lon+ax2o
N46+GoXIWLWMmg7HVs1PbIAt0nea+6un8eKSJb6B4Fvcknez+238a6d0hFOVBzXne70VWTsiSPlZ
nrCDmjHt89qqBSJj+c7+20ECh6zWNIAhauU4m+0YRSKeDXBwXpaiWAu3UMHofGoWvkTmWAIPiYGp
583Mx84O8tswNpDganxssvsaedM87VoXGpLEI89ZRJIUip6EG5izOr73Mb6RcWwYVL2MRRbyLlhF
jQkJOQN7rOhQ7k/AIQFYFQZeEurKM71gQVbrIwc2bcoMhFGuwa1pvKksRPCtYKmU58npKydLL3du
SAOkecOis9xmR+r7jIm4N5qz6YnJViuLgeRhLqCbHe55D2JP1/NFqVfdIh+4wA/jnXjePf4Olgow
radmuf0tJqKGqzXixpC8l6TMaDCjljBg9vfThO1qDCE8G7W2kgG3HepwT6Ar44ZEjFy9b4ubT1qe
QYEtKjeUqXgVP78qX8CdgdA2QevMTKuhoyOpdpbLHEXmWqbINZBwdu4Udkf2ailWp/b2jEL6fLAD
k3SUes4m1umTDUeJ8cdfHY0OgrV/isfV3jpYZ6of3hHlmWozXUUem6OcVTgz3vlF5dN8mUHtQkBo
adCbxBC/izuZSXDszNwG0731YAcN7qveDnn5Eh5yHoy/41tfL51TsdAqPDz+KjCrdFJPONGnWtxW
X7xnpOYHudXVP/F7CwQC/mGzn/cIl5zmvYBNWMk/HgsjJoii5z23DW+OUYExpAmG1yamDfj4lt7I
yROkZnpIi6buC42+WWbbSTrpXUA8MhjGa8RKzcTEAqga2kgnnwULoPceOCR8FxhIBHzV4HoBeiFp
iecjhzsFWNPHBjw5QErrCA5mOQNxfxDMHZFGN/BYxIyVNxzXrGWMyeKQA1JiWR4PpQ1FL0JkuhAp
oiSJh8J0O6nvEf9VTjNkFofpMOy8alA1uoVIRJ5XR3M57q59CFG0qVGwaMVjqkI3sA0XNYIoO4gF
Swdt3UZWJpSfWiit+26Gpl/BHA9YjEpaD/xa9ITgt8FW7FhPk8bIeLIr4J3N24zliR0OZWbVM95A
ZICPuPHvd2pQG+yvUX2l0Vz23kQ/+rldv1KmZ1tCxSaBJ1MVv0b1SxM5tdTqDs3R5f5cbs5J0vgO
RHqzvSg0JeGCw1LY+tTx8ivl9v+rF5EusfEeAfc7Ne28gCDTj9pMJ6hwqeLTS6Z5p6PMluOZeYXe
zwhLhgX3BmkNh+lUa0QXW9z6J8R5ljYhhWQoWWMHyY2faDpGvgizGEw7AitAWf4cS/jet5/bzMCW
1iMpJ9/fFTTUU/foXLJNkW/lfuZKaxkTAiuvsbTO/ia1qerelMWUIS5wHm94XWoL7LMvxpf3AG7d
uUiG1bqFwiossqJ8dsT9NRvbMM3jCkxf9Rwi9GDKnZWFXtGldIFbfKLR2vut4qEnG1fH9WXBQXua
Qh2id9a6ZlQvwJjRPJAOsBUEXUcsgcZTqYd/Hqc6+hVVrN9qKvlLHHysdii749knjbLjwTPg4jdC
O0GoVApKM6OgMvDLl5Mthfa+q/0Pp6DVv8qeKMTQp/2yffqzdnOMxwPaeZA71VdT2RTNwBlXHvX6
aU5XpBLimfrnUqrNmhtUlJBfYkk3DlEdszhD6Y/vWMOF/p5Lvfa7UmcuIOI2sPM4LfPNbluz8Mz6
ZqpdGZ2z+9UzpNUehCVYuFcm/sVEMEjd7KGdnc5mwwhQ/2pi1/eOASVf6mNSXQ2tfRS9a/iihpsv
coCVyngcnU6D1pYcoKUMoo7sieOKC9WUwv2RBsmerT4UHCfRTu4f01tbzk3fdVXLwZ+ZPy076vSv
C/MfzR4klNRywIYiXMnf/3hwrvL4P7LiOqufPTGepj2flwRxxMN9DVI1t9GWvJudlq4An8ryGWST
9OqycHW8h2tq29soDBJlRUG4FrQF2SEkgmcm6rUrbBlrk6yrHGyTaT7aeFCSwOCskZGfqSPRNd2I
jKQ1iRFOXObd6HWu/8M78OhQXW0JY5VkEttUXWbMLtWA2HTcGIxmxUhdO94nuxamYUy6ajRpwE8K
GFpHD35JcMKZbKiUYBZVOMhATmjotICMvxlH5V6JN6y00VeYYbSFAKbBoXDzvLc+nfueoI3MZR9E
AFAuhnFyvOo7UGsK/Oz/368fKf/Nj4j4aATZuKcGeMO2QjDwsiBKBilZzoCmmortrXpdNN/Vjh5f
6q7QTghH1qVcnJiJjyau4iwdjc65W+fOhn76XvJ5yCjzXvQnvGhbao2Fud+Woq9BiFd8XJT4qo0r
lmWTvOipAr7IVt9YZWLz314S0ZMqEedbBlBcdyLyFODJi9iakeF+BNifZTc+imfGqEwL4EkL2uaB
6JMTLvwzji4WxrFekrKYXG0EO0HvKM1hQigPhQhlcMET1BTkFryw08bS73LBdqA9NqDdjYBRlR8F
Op00Dh+34d2S82CecY6CiiemswrwTjeXNWzoDUSqLBup1ruyuzOtb/qq9mRzX5fZLRq5ZVX9Sswf
8mC9qNK8hyqPjnzAmsWImTVQtxMHwT/s8e5s9NwpUHIsR6BRhXSD37fLRhsYkI2VA+5r477yi0WC
AXrf8IsfN+aGaRBXzEokCl1PL1yfVM2Sx+n8uTdS8AjhvhYjKu+dtXPPPi+BUxIjQ5KbuaQV6KP2
Jsc5PpoTWOuIrqPAxQpzKOOwZD28SC35I4A65bu8qFbzuPEb4ZW/XrIhSJ0xD4Xd9pNjf30TjOqf
+A+NuGZ4LQguxCpmzzozczhS6ZpLf1VLL84mGsgGtwG5hxOu/RfI1j2Ib3hvrXD+pmF/FteUAgFy
8vI1/w7UpFlG2mfZ6YMFIXB7yffdzFk8L8UZwmh54OcFIu2n+Ex2xSOJQcMZ9koiZ5XSO4xUVTrb
7389PDUPMh7eFQTmMIsU9XLqyjcQp0sUnIL8qzt2s0L1fWO607mSS2gmYI8LgocCQ4eaeV+f3n9R
tjM+mDuR1GRl465oHhy/cy1GLHf8rGoW8Ec5HdzNY1EHxOEQRz7ddvz3cIReLz+xTNQ/NYclj3Uo
UB9rQKtDd/16XFWzOiHYUxTVYvVb8UXkbjJBvY/cMutipq5EqbbMJvniZodnigVcuiLUWPiDnzPe
8XwGO1ClOrYOwmERMVTKo81WE4ihPWAZyp6lto54l70iGjbSq8vsHGLhm/R3LtbIDRSq8hrNCFoP
+Y2swnUQOQyx4h4tsJnT3gG8pzO+cMQ5mUuQPiLHbOpU0hJ9FRKAVpDd0iMYZ4HZHWKDB5QOj6zh
Y1vQtmr032ZQdOP8lwkTJWuxVAc3iZF1JevJ0+GAp97bs0IHVP2XND17+K9Gd+8+daRMJuxROx12
M9LgH/b4D8UufvmfGRMN/uePkEnhdZqv20lwk+SnJB9ZeiBQ4DS0jSrqXcx/n0t354IE5wx4m7Iy
WLzkii+WyP/n07AHWr5iCJvW3BqDguAnmOo8GwEGDfUa0DKYoD0kJyC+eDzO7C0hR/HgEuQ+hw1w
r2M4deWGe8ibfd1TvUgrgzeTqUsAoHZ42bxiEeMROtvOqF3YF+NU2jzQtlEKEWch1XB//YQ3jAuX
GTtLhZb9mFPrMFp0XwTe2LHrx8v0fKovL0b9TbwLlINX3X5DAXA4BwsCaFMHiFq8WPHi6+VzIQLs
kjm7c10FV/A5yjvRgZqRrIpp74Ueodyx8nBmQd1+Ez48O/bpqjy+rwOA8jzhNtFcnZ+5lhKqIuig
XXwBaJDLROBNQk58o2EZDb/DKEw3HtwPQjojDn5KYU50GiL4RoaU3RNByZq8yZs10/dSOsU9RFSD
MA006UwyH8bSLxxf7hOdWItFJKgdbMNRdMAnyWlqqw9Hl86L
`protect end_protected


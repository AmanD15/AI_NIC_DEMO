

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
AbrLtZEWaMZ9QRIEqn+KbGJaY9tnAHwhbFbsPC7WH49ehpa1EbqXv+qkeNRGupFwZ63XKanLVUyO
My0fDcdlyQ==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
jBjvZpZ5ZMxrEO8+CEfz6CEl8aMhkYM5vXXCdl+QFohneB/4ao6UdzksCSxNPxkQX54YmGSOciXP
wgiPEkvihckzTQ7V+IwmdcU3758CZsJi1jYV4WKld6YxfbWBrziJy4pEooel9pwm0aG1jMx1yNUM
erFXjNZfwKELIgXdp9g=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
bNlKYiiGIQP+R/ChMF9YxWObkJMdPWBzZKUDypAuNCvFSKj2ODeFkzLXYHokfw+rz7RZe5YojYmq
4UkICxShbV1k/N1YYli9QKFi7npsW0xHaRa8L0tSoNNqAKETg1msjVmjBV5kKgQ78l19v/4te7qL
zUqdthBriU3NcZYre5k=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
0gJe90X6qrVRqoGU7iK/i5s05zq/0GlJ22Kt2H/04aXbES5oZ4I0aGRfiLSYUCL8istn1JleJ/n3
1/LRSIHwjesRoSy/6j9iedPDLLSSnKq+N+ZcvCJl8gg/L6B9ChU+h5YNE7HqJVfqJzqKWKPqsHB4
WVtjQ/Uh+QwxJp4Q/GXnPw1qlnDs2s6lJ8EK8000R7Any16QZ06T5S1IW5s5v9bKhWJj2Oj7lmWo
6QSr9mTUFxCIV/m+pXzsIOsSgFWqsBmD8jksQw5AorgxI1HaqEa3+sl/imtv2p//6lwEVtz8coiR
PUlfIUpZ3ecBYh1Zuc/GrakwiRgEs/Yjfe+jCA==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
ux0aTH3zrSOSGrjxNBhNJ8nXWhxNzkLj/DcKiIgChJ1nxm8i4YMzp0L+VdbHtn6L3ZPNF7NTEh1P
v7Gcx16JuF2FM4sw/t6m+FCjX3oHl0zUFDs/HfDB1IEXz+2hsgoR9SYF+bXbSth9Ql5SVw6WlbpS
yFwlhS2eW7RGdfH7yFg8yRwWXcYySMv+L+udV6VzSwe0SODgbmC4o26VRMdm0RBQjLnYxl3eT+4N
Qf9DbWnbFLLU2LtQWORMV3hNidJEmt4J99c08slF3izsh110Cv87/wiU6Xuvi2AB6jI3wVkno8/h
1xSxQBnRHm/fJHMh/8PrydoVk8qMhMXs9UM3dA==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
A3eq7CQ1ZEC2Oz4Co0wE9eavdVVL5N2w7vnxu/t08WjNVvgkDcorbVB3GWcUKigHFQo0FHxElw0D
PA15/K+npi+dagAdVUmv5cfV+KYrdhCLG+Kvl0Tcm6fhXM4RH49frRlov9a41BctZWlMEXzlO2Ei
69nxF8+cDN/RPLjSUoKp8oVTX2g6+udi83fdCBYaBZQYCaaDSNeGqephcoL2zlXyK7vU9KpsDUWJ
oZshHV12Yw5hL+4YuSmKv1aODQadN1UJ8qyFc0vRYTAqwP+hcDUwxiR48olGBo7U7czJnFk4AkkD
qULDB9rPKRIK3YJacz6Pp3GAHUDGm2JO78Eg8A==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 74224)
`protect data_block
vSBjX61Nvft2xWAWTntJB+TclME1vfx/tU+V1Zgqe5qhWRwd0LNUEMw857X+yosHNPPKQuZsnEPN
F1lLrbG1Z+OWylFciacRqPPE301a96BcytjzskGChguOZF8urBEhbfPCoO2gIeYimAV/sK5AAM3P
1p0zlt+5IJrRYGa3XpekP8u14rHpaN3LQwKbfl5rOGtjEBL62jqzQ+HArRKakMHsSfhvK/mE1e+V
BPBbBXnpPNb5ycDzGvk+m0UySo5FOLKlIcqLQ6jb24a76GhOAVrcPG2fRWMotdrG5V4yOx/iqrd5
s/a663QizWztKiHdtwemBc7ap2TT7zjpWpeAfVUnDAtrP9C6TmPWgotI4ZvXHyqApOphpXrwKK3Y
MO+zUYdsykM4+rPCD+YQy0vQ8NlMtDPGP2jV0PCHTAy+WkLl8r7HKbg3nx1ndlyxCADXYa8DcrF2
hKInaKAtJUWYTWUdqy8kY7EpEuEa+tK87ft3ZCJfOxp6tRAlHFO51uGtZiq8uRKv0zZW1wbIbGFk
OtAq8U1g08cRyGzau2baWBf5lgI3L+ZhN2/r9pfBBkAGoOFDip2bOLMDZzg1c0hFlE16WWjfndCi
SrwkGXVHLM1nRJkYF/iDeWsW1Sskgc+pvshsqTCrsQoKFhvr/wY5ZYcdJ7K0DA5x3N45jwBGTlan
xxaa9Xb5HubwAYpiQYv9rinEOeydrQ2QpdWb81X35KwtQu+y9/tVuKAKCgVZCmD8UfAbEO4qWZq7
/d9RpFrxwHq55cnwJSUHBGbzpyB+AfkkROZChmpwbxQNbcpLzvDqCJFYsJd7oarNRoKhZQ1P2wwj
ZbdlVaPgcusnZRmwAsm1xLwH4gBUOBVX7NmVGx0lKz5RQUJ/InnablmIztakbeJ9RGyV7Z2oLFhB
/Ij8qdA45lwg1ts0i+8XN5b9biRyLcCqvUOAHKXlCjxntP2uBeSWrPfGH39Jc3Q1JWpxZD4BVwi6
gxDlGqn4CYowLzJYSzD2vG63yNFJYFUG6zCnz/QkP2T2+HvBB+eJp7JvIfFv2irw4ey5rqh4ViMg
SDdkPabXMYxxY6cJiSwJIjFhWwFoTl/sN0z9+Wyc5mgtBeBAgRQPydkwca67S5o6IAQ+TvDJfkUh
cGpxae4e+Ursf38KsB8m1ZZc36DNnzgQvnxPRWs9nXN1hZqt8Vq3UieWkoP9E1SCF+Qe1KWGlhF7
1vCRI0MRpZiriaPQWbES+Xm5hkAtFLutfU1VyBvcwsGky0ZbTmxc26V/qHl+0tcZ/fUKQ4OumcVg
pMzZYg4oQdlavsjvT6k98XZXVVnCm0RZR0Keebp33exEDwTYciZPDrqvtyVPbhmrzLi3W6Gs9eiU
0BtXlkXxDvtr6Ee/85MihIZSguPvHkJ8cD1ET2ZjoPWwxhmdmYijqJlfjizI4BbSjlQksKoJpbE1
XaT56fynNGshxaYgXcvxVzdvQvM9MQjnkWW4Ta1qgAAF0vajqwku83taUMmjWq8ih49FSvycxHFm
vnwcqcmUAPtyiEELufvJ7LIEnuot0NncAj90lUG8fqBJvC2qCREILoT6B39ymQaWyqn9gQfsJ8/f
lXHO02Y38MLp7YBORZV6Txh9KDxTbN18pgS4Z2eSQWtVbJ1OiSlykrPcStQ26AqPFaARKzyP0z7K
fAQkvHGUyGe54SRadB8cqCrungr04fG0MntQTqNRbfHSX0bTEAUbedbP2+p4WtBVddy+E/WgH7WP
xLP7gbxb/EQsaE4dyar+Ih32WLZr5PsJ9A2jfJz7MyuPRkm2TqU6sGkyso+JNqRI/MnntYSQKXsQ
YUHph/4HqgJ+jZ1U5aklJA7+1Y2sN/QC9gp5iDbn3wtZquGZZ1MEb5kXkvVmg1blAbQcYJdFmzsg
XyJyKG47NiopX8T1YXfO+/z0i1CpaqspPwEu7WU40hZlH1qFY2wOytyT991pjfurOy8/IaSpcZXY
gcnScnr0NbDre6sZv5Mfj0gRHstQGo9dXHdEyteywE442DfMU7mIlDSNetAmY6Jpq8/MwkK4uI19
gkMVij0HxjcAogJ2813GrI877EgwxEP/RPx7YwZmeSi145EMQTushXf0aeES2mXJsSxnZl9Nz3+p
rjT8JQ9ClRYS3KmXfQaoQ3rlcwnHZhy83eLDKE49bb4vnF/kaHeqSZtnahzRkJWjHwa6v/re7ckG
QOJ6fjrFXtD2a3SVp39Dq52R44O3GCMLe8ExUnSMXP/5BXPineJ/jZ5QeTS+UglLws8Sky02svfK
n+9kA/xUHTc8khQETADKOP7rj6cgD2U83JStdoKUtlJS6m/SfenbubgyK6aZwqQbArO2pfWYYNEX
+M6s8q05MMYayHIG1D9tbSeTB6haTPhWcsKTjfjW4YfvLyapX9QsgdxXgXFTdjGneKLFg+XrO7Ur
xsA8kgbnkMKRhrhlSfh9NkpoRGQFO/6rMHXCB1D+mHO3zg281OVq5I6Ssuszee4eNws3CYFoFGrc
UZxplmYcNNucRocpYawTr1j/FDBeNQWbdQMOSz50NxNLQXlKk47GC0WG8MrU2arScBbmdEvdSJwj
zhx9FFcggWSntg25uF+6fmrmesYjZ7BugHVqqbyYzhzEVZbt+7Aa7bqmGol3joh9OF6blIa264SZ
/s6e+Xu1iHARSUQUMeLYr4lHZdOpazysHQfv08fSeucp6q8F/fCT+zh7AEHgPDjIW823GqT9lfcD
tN7Y5UpIm7oDVLSOVLItzt3hflU7Q4btE6b/w7HDByDa3EAMXlanomzrbutncb5t/XXkkqrNH1DQ
/iGNK1Qa+SXjxdiDr78cs2Hqj1GMqxGCyeyL776Mc4pMRTDLSUfgd8L9VwUw/Myp/A898Ef62EHz
Hlj3IIldppvqhg+2XxZwUef9JpKvBEbDQFTgZ0rUP/KCJeabicz8072pgkvyT8bLdYuoORPEGMO8
Q1csggM279gGZtEy5667FnlzT1fADsjA7FXpAuMjBCanMTbHOfBi5AcKWFT5qMSMmhsz+PFqBb6r
mFi0T/FLViyWvVyHHrkikjRX+ZQJa36tpBs2NQMS/DgXWViIiLzuEfnB12K2zft03Sq2EK7H2aGj
pFUDkCh+y6n6i4EKydaoelz5L0yahhOqWHAEezU4DlTA4DXSrlGB0jifUaOr6MyrRUOMLw/dc2Th
okbvZzw1a1Y2R58gYRPWBdKDcXxQrnZZMimvDuFNSfI3sQEVoWI2TD/TRiP4gyK6BKaorFILVLRK
JiTmmqfg5zSS01shrNGpixgXypaZWdmspAIWonVG3Sviim5R97Au+is+2+zGziKzizy7HA7RbfDn
UMSPQXeDUNFD4xRPHDybs1K9VllERnsrLC7dAkDIQWmj7YtW6dT+qx1EAEQQ0p0sCmh8fmtlRfMO
2bqFabqGiRRT8nXqhZ8qVvw3bwPF9eq3Cy0sa8+FO2Kzsb4ZsYNxS9afwAuh7w4krpkWSIjOy1Uw
vd9BV0ECrjyYjwme4KjzsJ7L86qvF6BXhg0j+JAKt33n/IL1FwNuvf4MumvWe/VpBxJfUUyr2qO5
F6ovzyTIGhG4dXR2QV2MzNFlDzJQQ4QZ9raIWOewRAxXC4+MBloOnlfuJKwJr6Amqgp01LsAyJ8a
rJigtZK8if5coyh0/cXsBjfQy3bxk2/9n6KQ2PsiBl4GsWu68tU+CuRtsQ3i8+T5qll8k41B4gOu
oP0WeyTHKgQkA9dlgB4tFbNuRScx6BLuRNfh2BbsUSVN9RVqanE6oazHWt9FQujXETts4Cd7m7g9
mWb8EmvCNG08QvGPGvY1rJaiR0nwOjbE7uo92pEhFnS417IZSh+OdK4WtZ1XuqVCTCt/wBf5/iE6
XwfE5TCDVDxpfmqEuW1m2gekVBexohWnKcLKb+QKqpZswJ+Ap6XpQ2ZSmoRYS1q7Q2M8gN2xUHQ1
9j7gPmviHxqLE1lqlafkyZP8gEd2JNxDP5KZeB2NVjj128l9VqghzPHL8YgO6bnr2MhsL8o3e4qS
Ev9649f6A9Ka1NeMDZBL1fvEQQwWRDJPn8PvOca9mnNjoe3TrIb55aJNaCIzf+U1IPXePXy3eT9b
HI5LlR9feBSplx4aTrwakZexGfwFpFeE48x+EDEB1hhEq8H25Fth5Uaa4/woT/pNjtbearUni01Y
FL+zHUBrvUCDOp72A0OiN8Erjho6YprHBNDSdaJdwBoEGmeQeJshFn62vlE4EIjJIMnU5dWV76fr
bsXV677Wa5HN3h3Oqf6+nHD7HzN+R9dsWB6Qyz+YmvJA/7Yq7yFIeFxZVqqwgcVdJvv51mZubSTf
wEgd95J9gH2ubGBNcPOwJwNY856B8rccrVE/qwAxgppq5Sdxz5do1s5y/A/2+nftXu6SBv4CwIcq
nVT7B37ObdJru81zva+TaMuhKFxaQe4aH/pwav1sPgKtqd4InEQXW1YdI3E/62PGxQXZWICfjIBI
Jo2451zL2jf43pWGB8bLYytvE5n8HVQvrpBwwo68xDYbC8eFD3sT0uJYRroO/0qgkFoa1EY5rn0d
WsBEVw+qEc5HzIowFWBnGbu85DEPFQpQ00iI1NXa/24dgmPyV5hazEg/xKGAZpwCgBF8LhNXheEh
vDHrycZgdZyuqrqLDEuh0E/inrg07zpaB3NdoTVLe9GsjK7U3f8JXR71HXdDK6ElAE0IgMNPRoLZ
CkP2fpMuUL2wim3RbPbZvIqxsFvfSSItW80j5QgZ3mWhGCV61WOP10QJm53f/7r85aXsX4QBuVyS
StJKQO1mcMhVWyraIC7lB4eElwm/BHOBMOK5l+JFS2JFj/Srmtw9Gzr4kURR1cSxU+MY01hGZ59m
FGblBjnVuSdikYcUj3LavfJCPuO+AE4zaAimOC0R165kfXrASaTlTUpkX62ct7Muit4JV8ktpn9u
dIsIlsdixqHpAiAyRfQESVS+gRtq5mx4grtQ0x4UPhJSQapSZUEe38Gzmp/UTXk/aLC3fBlL+OUB
hKOnKhiQ7RZ+5qnx79/0/i8/5SgeS0hHjCuQV3N1DjgZ/5S94UidIfk/aAcoYH754bn1jw/HSTzr
5zSpE6/xkeohbqakQHKsj/2XL3QnGF4dsGqW4CCrJ1IEdjs/aeJP1r4mL7oWPq0y6NA15EA0CCvG
mJwKNRbeJVEWTBU0Bx28asM2J36+0CEepCGOo0/EW3nYw0bqSS4XVnrQAI979qpvtLk+2DcApM1s
Nt8vx/eAnH5ttFgfVZ4ozQqTCx3gRdYo/fWKzRJ8ksb4uFq8RUwXg71R6rfdOWcqNUv8QrijUR38
V6zxH9w+4aDHQluGAExIHR+OvmAALUNLa8IejDUYp66gsa7s4dlhV1Vzz/7BkV+O+jh62W+Mh0og
Uwcs9CGqg0MIqZC2pwaGN7oxQpzG3R//twOKmzU5/F637zteWzGItX7v7sYEL7Usv+yOgb/Fh7OU
uUNgno/868RipfGccZZsMcXgyWv620QkcfUy6ke8KuKDgpOAaqMpQ1eYQZJYQfLUwQGrm/naezrD
lJ4e4wXiXspT/3gEFgHXiTdIAcvNcwgi2OzRP3cWx7HiqZx6ITs0NCk3sGMFuXHkaEtjeYppZ6uU
QeLGNe8NjQp1tsG8j5XmxCTJRts8NFB4FWWWvANlhSKxkyJABFyeDq+ynYVEHwZ9waYF5Bwf7kyO
coMzt5EILYwvVRjlJwuPC2MWZATXWxVdNd5PSqKDXVSm4NXRGlBFZ5iWOWgvKULJ/y6sthyaLRSu
iCnJmiEFAUgkyy6BYKyKeaClmVmEI4yRXGz7hxKwB7aCk2YFkSSOLFVGSbmA9V0gPcW2w30T1733
u6sTEse/DJTeJAoFmVjSCCf+NBttp31p5l4bJBmUBXo0vQOjHdgsqZYuAOdYEOI1vR76AjWeq5vT
wUaU252xz0hGFcVFcpAPDAtKpdDgmRoy2thUQyolJuD5GRFnt0uNAe1sypZGLYTXbCdenQr5MZj7
zrlUboP7C6JkRKfJSgVFQQSk5x1Y6+KBhvH1Ohi2AkLznIyVnyC6gyBxaUxK9j0shFgJKhrjhIsG
q5AHHdQM2YtmnH3D5JYnMYhamFc7E03gFV3MkQF6i0zA6rLrNk0SsWty35Y4gytdMPqZ2YLv4D7h
Zz9nMDAImXy6ZGG1Kbny8iqAqcMh3o4dERpOUhy6w4GIJZmE+8oQq9bPIJ7JdhJ+YiF4yXu2DNi9
XYqKbXIeLEzJ/HMBTuwt337YUHzigy6TIdqYVugIroWTGWUD/Kv53YwPe7TcHVI/KKO5BocuB0X8
CZ7lHzi7PCOVp9xMKyHPmYRz5pi3y3Bewmd1Nh5v3Ex48zUAmPTb3TZ2TOIYbvOqXqHFCjKR3vC+
oE0YTPMTLXU93qo2cEJNfuHFfjLAhoePgXYkLIEsKSzolSfyPFDFc0WSKu7h2OEXsJeO/OT6FE2M
FbrYq76UG97ieDfqZQpzPu826GdZBbUzufQ7HOpCbxvQahi2Ezs60k9CrvIb73QOZxOettfHyScn
0//owyzgHTTsKFmmaeEsTWGYD8FyyBvGs94qgILUfi/vAd1m4eY0q4/U9xWyn5k+JqpgeR8L0jQ4
TY3lSwuHU6xL/qaK8MCyYj6gke3lJIA1ogW8peb27KUhmVhz2Q9FB1aykxBzgU1OYPoiA5SqF/BM
RbLHtgcr7oW2NbCZ7+o+W23ah9NoFzqpBGktM5yF8ZoZNH2DKEY0MVJFuBSLR2D6OlfCXe3BI9Z7
lLv9fo/vXkbN6y7Lbja8rbPPwGg+IPtklSNIz0PoBytJd+KKZrfM0jxnYDPdP0Er2FQYnLP8yRtf
wW1u6dkkYMp+qKW7UtJ7b+WI81Plwlf9PbTxoH38X72RDSXHjLYQ097y/YMVxviYYwVAwGYWiiex
A1MsLLvTvqBeg13fJhzfdjBLwahbNEnXPfIMBVnYLWJ+xE7NxlQ8FZan3D5Fl1lQcDuMIdkSmTZb
8nXNre9JbxdX7CbAse9XahY2RTVlrJt/3zt8bI1P+vwjVB8RS2iFjMPqwDxgbMHjzMpOk+lDTgfb
XbP76DxHBN1zn+tjnmPpNVBmUQQqTfR2EKGvzn96ZUeS7hKFMIqitZLfCQk1OX6dvw+WuJ9ZV/F9
2vrQ7o6bKXjQWWI1DT2CTHGsGZgDUt3x6IPv+00iOOGhDQ+xca3H41svNg9mVhFcqz3sBtDKj2H/
6fBCGFCbFIn8pghTLb4IqxE8I+4rxoGSrV2Gl+M1xy5LYh9maFOx5KYybk9OEC3mpgrD27RSHoKB
nkYLbDrNDE2Rc7ubdrDqgYFMzrYX73ZfsiVhTmgeQfu0vP8DPrtVFp01LyNiWNlQQCav0pcQie8Z
hJWwhcoqZmyGhB3sM7cJMDsaRMkishc+N6MCGE/PpGiI2oO3slK87BGDBq+bDtAU8RRQLGy/xSAo
A5BLlUyKxo0NghrlmciWDw4HxMRYv0Hqx/SeHJ7vu6Q2qW5i5qyFf0rCDjhvP4jayldJoTLV6CpE
LbbXjyXwVw0E1j1CmDy7QsjntexgCsud01V7LS12t29mNMcuamuM4p3tbv1K38x7U4znRODwr6wP
SXeswhsRHfuFBBe4kVmuhh7omi1HTrTTFj57jtv1ZQ8bzwHwOR7V+8MycWu7yO6JHUkCB5Lv3xOu
laJxnWEHu/w8tRAF4bTVe87AWpwg8lYr5Jf7pr9YB/xo/pI8CE/Ns7KNmj8pJLT8LtiDG1IFqdBG
7nOI3v4k+I6/kZvep55SN/sLsWNioO6wxNPOX7+joWZPOA1yw3zraCsUb80Sak4XUBFS5STb+1f0
ik7J294UK1jjGOEJjzmaR//4KnFTsHpx+sH+XBF0aksZW0aMPQTjWvScQr1uUL9PrP7nhf1Cni+P
qwNiyeWRcOf86ZclRtDiaaglPmq/N+vuTZS3u2FnK54Vr25pa0L58JRtjPEjqsYx28F6NgmCiqdV
xYcxGyrjWkXj7S+fwmpd6+eLPLuCFGNqqBZVO0hZMITD6p48XgaACC1+du2vmJwxPmbXgagBCMc+
iyKxTAlUx7cRukCzqFaqR9boUFSqIP78fukWWr/ng9PJNsbp0BYh4Xlf5n6UjbROPtYDaJod8tgO
+PwY9mY6c6JggNDHLjAtCBaVkgvhuWl36fTCkjt5/riXuJBPzsgPx2HZG2KTxXbqrz8MRBYsyhJr
v6CdGgElAyXLXhrOWXYdi+cSi0+ZcnIY+j/K/SxFP4nfLK691GV1NoQIqEdBFjx2bhNlbUs2pUFx
aMHCrDzEx91etRCwc95Fch4hRY5Kn/SnVgEEpoSdA6vU9Aix61LNShDIOvdyWBpuMuvBKs+zCEBk
lGQI90F8BXoHVmKm0ngGuybyumCkMGnIl5YyFz4mNqwffcJNTEGD1QzE/p2PzUEpM5vDb3cBVCME
LTFik+1CpJvmO0Wpwuof+xsIZ/eaonlP5ZD+zPpfVaZfCfkEROoQmPl64175McYRVQ9iFeANjM6K
/zqoMszA101KZuDKgMdwv5Bz0EjnHukl8RUpWH673FpDq2KX90uuIsjPIaRxlibosMlm21LQbcxk
mD8tmtas3+SD5tKSaEkM4i4HhtSAoH318yAltwi5cv0uoAdESmw7SXhUCkx0PgzAp93Qpm97lu6z
mx20qNTW7HIXOPH1XATHXQqjnIyqrni3u8KnZbOV+Urr7ZeU90GTRBRO5HwiLEJP/0brHXH5UiaH
TSgG4zwSQU2evNPCpqPsZ7bAlf7dyQVxDvThzvJ4v31vpDdLQoiS9pF9ymlE124n5BWNm5atEAo7
4SRuRfxRY49BCveKMvdoVi+U1TPFZ+aPVU5psCVCy+3Jpv7CCjCojdgSMggi3g1bD6QtSit5IjgH
VHYC3KBYiWvTnOl7D+5AvyRn0TGU2cqpTDjgM5cki2dD4btjIwHquN1vrtUb0CUi9DLQ/ieP7nYb
2M+7QYfihdiAm8b92sgr+l+BXhPw22Kz2JmNjXKH3PZ7U5Phf80YQeCuJOmJTCclZ+936UREkPGD
isgCfMIpvKOM7YjNeamIp1JqCT393SlOk4zJGlAJ9MKBvCccb0LLnb+3+6salDK2x9iIYhecaqT7
y4PrBP8bYvyTxSrFst2ZDVe9iW8cKtkVkhVcbRnrAai5SlckQLJu0w6JnwM8R2fR4LiE8Tml2gRV
rsr5oAxUuA/VFiizXULbTdbnLK2dtBnXIYytj2rY7hT0vC8syad1kplpRT9MMbVBXNSbulmFOyMu
Xlm1V2saSaTj32kL5ZWMt6GhJ3T+pYo8v+Ee4TfgA1dt2z25YZnukgxXiYG4oYeTDeaSluYWkAZa
rLWXgJ3CaDrNbDL+W3dkezbgl0WFIckwavFYJIZ0c0VUzGNz9lokHRrqGKuuUmQfCzYgWNvojggr
buqqLi/9UnsdGUpp5NRnWmwvw1gbE6t0dCwSRmF9UUrHVfl0fVLM82CJdi+boU+4ic4ILjxyvAM5
nWgJrKy9mx3LWEMsvbvnXzLPxEAA+39d+JiNvPH/MH9BqQyM8Z/7ySu5Bh1jHliKS7VX+owMPRub
2uumsvuudVDseednSUnPyWQZkd/pNpzYqjR794Hw/gbHW2VpILljX12ZhzSNx9rVUNqE9OhRLC0p
fvB1whIGSm0kOLEJ5gM1goyzEDOIoI6IVzfBiNAt0qSO8QXNouKGY4lne4NGhF17QjjwH2FLGlYx
RJmWedlzfk3ha0JbthOoqySWkuyAFyBdVUHjZtY8CyPDANOYiwkVcg2/YHhjCKKRCiASTNWh4jOD
phZAZyn3YFh+Bp9Mq/zzRuI3/Vk1S+k8QWLwGjOdO21+59MFWYl6LJt5spIlmprXSsnUadtbE5ji
w/NVTq5pyXvEFe45I6rz/flGcLBdU557K110UFP/asIsg6DRjT+RGUO255k5i+wCs8vtw+/D1Yek
29DbMYoKnM1wsaMajpA8vvX7H0S/bLhDt5o8yHl9ya9kQugnnouWtAYKv7etSkh/P/J+exTxN/1B
+cjGybYvbNvzpW2C8naYZ2pW9gxINphqBl7oQaBgAsY5XrCA2hwNfqY9XyE9Xor5OOZupH119Mhq
md7D+zu/6ChGAvsT30jfqWtqOZ3K4l1zFx4CyJxxqHkCAkcn673UOjmBTnL9TW0uBIp+CD4joG3R
93XbIx/T7+K6Om5xiR+7GltX6JEb8KXqdSLb3hDUvzG2wIT1NFz9NvilZhjgGlN5lROU5LhRgO5B
R4ENw3RFn6LNu0HwHae21wS5Ar4/kVuc8qp8NWVyCFe97XatFGkFt9ez4nNxFSL/ayULwnkeQnZp
oO3I7jfNcCXm2fjYvECKD8SWdZQsd2DJz03chRD78HDNx8i0GTqYpcKyvbq1VMM6Wrt4zOFh237C
emjKPH4IS9aVmyxHv/ut01bqU0llU7oZ2qgSRfSwfF/oH5dSEMskdq4FhEvwmNHlsHysnXhKZ+3r
gYV6vMoN8FaTd4hutbF2DsCwQ3EQtI6KpFtP+HTKwS63Im8xoTkEW3HiCGxFxjI1NnkBIr9x8aNf
M2auynrb/gUVb8PmbM0/UP0QL8M9zRr7uJ13Gpt2DzKVZK3Vv9SMSe7g2FF3rXISpcLsVowyx5r2
nKC1TePIjTu0phAgsx+HKgAWyPUgwM7toDZzHPwytNs0Bct5B9VXNUl3WOMvPIiF6KoonNFiDHvA
6WqzYC/kTvT4eAcdMHSOHNGgcqDUHo8ei3lzGtZF4qFNOUgxkPC3JzTIaTX8NAmoWCS4mrPWpHPK
x/Fq9NoSfYoqUZXYO0g/1nf7S+1EvIJqLqavY67Z0mzvUNpPk6h4GU45Jf0lsjdmSiGW/keM3adZ
nIhAGWYJWV4vhTsFGx0oxdn8/hxxv5ce/bpPSMj3ZeTK2R83lXnkCUyhU/J99jEn0Uj519QX4e6K
jCpr5GEKFDAmomMQQ3OoBN/4s1jUkaujic8gNXsv0OCb34zY7IYJ08L9DQVDGKG+cLXZ7ph1IUCG
nDV6WJvp1CL8qDlTPwLOO+/DTCzqGkWaGT+YcWzoxq3/N9/WJrFpU63yYnJMUPlMJbW53auf2PuR
uv5FxWE51cPI+0beQQoLd5v+g04nbwN8yjLjTa8dWfe3oZ4MIf2uoGfW6tg5F2G1sEWRrq9/y1KU
TChsE9SN6gwBiCD9N/ygryJvrMXdDzdRMAi2TRXFkSVfcTjBnjWkNVZZp/A6HlGqtdVNR5e3E27B
2xmiqv16QXGkdJBUz6Y/bJXOjogOBlFA058WkLNXs7zOPE5en/uy7D/qtRYm00uXtOnlNZyf8S8C
3hIaqGbIHXtu6wp9HpBDOmNrFFZ1rO/OxdKpZE/Ks4xBcEuVDtA5zC5GLx71MSMtTD3pjDeKQusa
Rl3zgw2Rbpxg5faSWoE/rqZjdYcIVh/uQbsJSrrGPXM0HQo3uwO1XVKMkDtvP9qGxnnwxuXq/7bj
ds7tDSxpJzD734Nai0QdTviiDqDxdJja8Mpo9RgwHUXhrvoswTUJrwgoecfrdEK33XDAg7ihoxxL
BaNYSlac0pGmz80P3KSi1jeCR0LjPzqZfEU1C6lvpd1jTKgAKpC6MQaPIfDB0ZRPdEiNixcg8/4l
xVQ1ErKspkbsnwEtXJpuBQy/RnoloQMAB15OYZdjOqlcpcGBFYOr3cRmHBk5pRQLQXPkvEvtdY3n
eNOU72RLdiFgQTsn0GLgwQjKG1QoXTNqgXLAZr/N3X7SC4FG0f3iwYNjRNwIuYbV7Qa0CjXQ3Dei
LK8EHP8ELsb72ReUzyVVZdnfYzIznNnlwruMCXZ70evA+1yYxrfRiJcJIm3F/er2tDrxx0hmCxRC
ZD6M8/boKS/dkFKM6Fhv48dI0O6bxufKThb5UgKgesCU46qvSWM6gToNHvlKLZquH03Yzk10pVed
/lR/sbF/z26Pk1LF+NVa1RUaguqNTk8S+XXjVUMgpL/KCV5sDa06qAHXLKVhmL/mCKpeyFKwrGnX
v10Ehr4STQndkXAKMtnn829nJWGBWXTgUOSlcI8e0D6CPOWimbaoQpkQ4LczS29ihgP47Dpd4dMm
QIkOVv+OuMOy6AERRsUFH/0ILwe+Q7f1CJmdlfJdaSL2R/SsGU36ZQgljDMgOjRwRK/MMsqPYIOc
01n9J3AgmYLuz9yoUCrSzdM94I5HzN2JSqF6nIoR3Szk3vexnBCPaVOnDwT6T6jB2zZj/iY5n22o
RqKAK7t3SkoTrLVckjylZM9oGEvh3EL6eE+oSugVzJiI6vIWyoPDjIDgM3HcGN7UcF44Po2RBKP+
tm31/qXqrozyqMMN5NK1YKJ7UcPdvpLHPoErs7eaE0vq2Vv9Qsw0L+rBesQ4NZkWouyXsEJSbcJ8
P9zG2HLVjyFEg0kdKj58HnhbYqJopuHhZr13RmPvX+gBRamuRyfn5LPk5UDGMYOkfq2k8qmxYXJR
wq1ZtBr/1q1mv7hSQp46Se2AIf1I7lj2DE3ia/abR5ew1A+XfMVtzPjDT4mLY301Ym07iuFaJp7E
fR+kVYL3dRDxOtiXdJCKO9agUd60pAALPWKcdGh8fxNaNwl33dsuJ2a4Cg8vKWhmoigiDtoW/IEq
MIE68bSi6MjwXQ4BDaA1TiJbI83bpEMXuiVqHkMNlSWKRMkJabiRtaD3icKydq1K8G/vUPE2Suj6
ka0U5oCDt5BoD64K65AbICtynD8vuwXKmdxMrqCto3OWJY+kyjcsDLAVxRCGtCIbipDgG2pJHuru
wOucGGYI9qTfUbXpx8vzEjkTRRoKWlI8JyRh1hftLYC8yWj9R+OO88Pi0RbDBqxmx1zYuJKZMk/f
/BDrvPpH1hHGnh/fJjBWoPKKLHjECZRYz0tVxZKCuVJQRUtfkFVvdn32P1fIqp0I1JgstEfW4PHh
NkHXjU9rXMypmS6+5pgfNLptdv+i/xbVkT1Dr0/8ucVfDVOpEhkZWMcK9msGbynuCWYgfYECHLzI
B2Bp45KABmWCo/rfKHPfqygUpIxyuJjhSuQfRNG0hKLAcvxBzwGvPRVNXBLLnhu8n9NoEQ6DAUZ6
eEfIUk1HYJO924RQkOq7yJ2juwA0Kwq62T7BTtyoZfmi9FL/3Z1LxLQzCxFrxyk/JjmDR8o5P9Kb
OYzg4w0rvcdtWH/0+TxtiPpKBj2ycgR3laoid5yjOFIJpK4Ezml7ep17aMoHy/I+11Bkmx0VDqNW
yn/ra8IIIBtEIHT/hHLPLwG2Ty2k8XhrHmpsdhPH/Ov+l5maSCwPAf1Wf1difm3KNjpgZzM9l9Jj
s3HT1crkbuKemRVT3+5PMqQLlVuK0TvhQsU12QqZ/Sn2nRVwcPM84smgBBcNrhQ4EFCZGEn0OR46
MOBwFNj+3xn5ciOrcL7R0AODNuxCZ5r8L14EIw/Bh+dLWXVvkG1bB3Lw3PSJCsTzdlbicejnhpcp
kKyDDhmUlo+7wEOugdstkTPz9kIx2jKUogg89819p8akU4HPm0cndMJmrwsIsrk2tvpP0TPEA1Bq
WO3dJzLpQJnFKSMrK4ykvS10yl8XqdBlUk/X3IpfA35zEwn4wBRbhNEWSmyUT9ZOhUxDksXoQBh3
K6s3MFoDLQT8Omk2woZJJTnCz+teeb5OuhCkGPy0+yeQmDlAyBAnrKbErqKu2iyqiSGrx0pz/k/7
+bsg1TUkqn0E3RmzBy3v+kN3BsA9pMuRU3+h6OXKQVmYbZCaiEut3frJAE17qjjdAMac5vMP2n6P
fhxzPM2Q3iUjDKhrNdCk2JwLM2/DNmjivA4b1VxOk30Umpe3cF50BptmbWk8gAIUPmIBOhBM4rVZ
Jp0Sm8s5JstumexMemX+YnTpCTHOmZ+HdQ4xXNwxO0pt33dpVhAxbGh9Xg+fpJGvvhrlb7Yc5nEE
hHYQtlXmS7eIDgSVQanxPdGREcGs/kzu3GQzQBXy1Pv9VlwHWDgBzDmcyV1QK9eLYNpeRd/+9hh+
3CzPsOhDWFbIDG55YtmWop5HCtif3fyIoe31BpSMWx31zSDg0KpV1Qbj3rRUpM5fJ0XQlvPZiW5K
f1YDqh1Em3jKhsAb9SPxN1lnpmc3O5Z49PxTBKAnn1/Oj39JVoajF7eEriF43k1mU8ttBKYf5GC0
110lgcWcYnrwpEVvKtqEGsZ8n2g96MnGepxihYoraL9rlIL7n7yRdi7XXPbRFGwpoL6Gw37tj5a5
7Q39cei3Zm+CYbMQ3ChD6/nG8vtUI/HxPwfRJJx/+DtauhFX6rgs+bnwfrLweBtHY91B0s2Y0CaP
BPd5ZxCjq6agyWuRn86nRuC5+5SPg4YeKtojdIxgT+l7U2T496AtQe4fKqhEplBUg1nImK9n21/U
2LdodJr/ozYQsshq6DD5v84tmRAlcUN7uvG8lC14EasM1wbO0LSwXJqma4kEZsU4h0e18aKQsTjY
UzZFCx0yEpPhGsqTK6hrwYI++84SJR/449lwpb6LuEKpmB/9AnvyjD8opMZFwOjj99scqNwyFAUg
4dMV/eIZ6vKpvjjyU94T2ZSS7eGI4wd5Qi5/ds7B8cn7eXUAoAwFHmQJYsvC9Dmzvw6q8hjlUJAC
JyDwVpcXqc0kCEYMC5CJq0XqtsTxvC1yFDSDdMViG+HAJ6mOYl+TPHTImpLcl7f4hjvILeq3iK5k
Quv9Y5U+uw2nR9+FhfuHibe5bcloi1wWkmJ/4qf0+fevr8VrIMeksYn9h1lUu29p+gt3RiEPAeg8
+5aBHefAz/ECvJamppxhujsil44pP+dSymAPtQZK+ffolABfiKFiWrnRBphO0lpp9cUGMcTRWSLr
noE+nG5TVxbw3yjDjf5vmrPNZ/4WBBTBKwbrnh7VeggTJZljdJJLzyi+cxR3iF34wB6mibm3VOPv
o9CGVUpFkRDCrbzlU6kfm5aewmvGZSq1xOuJ87q7t+cs/tbTdUnh7M0i1hMnUid+XOySwO4eCgkx
BRLCN9Fc03XVt8hqbfepN0HSYB48Xwj/Fjv8K/lz0LEz/ZUlb2Mbz+TLX2UZbj2lG9XO4QSZJSy4
W/C4LXjqqJr0q4NQ5iTjVQJAuOoPPRkPKz9AthhcbfCWgC59T/VMpwGpaAYQnAuPj0ocKtFOrXVu
+gu/1jmOKB9JMwoypX6rHv78VTdyrBGB1QwUQrqyzr2pU4bje7B6OpZdE1SqCUhL8Kt+2/z7TIMd
IhJ5YfBn5mwLqsTej/IJvprz5W9Ko7miwKQeHjlX/mDNs0vysBnT5qpci4Jf2yjfHkYUQPvNxk1V
ATZ7mAEwU2DZwvG3De/wdA27IXBqLdv7a9cyo1YXJLG2tFDBic26Wjz2POxw6CUSPbwcg2DuGzft
vOj4eYgyxu7tHFjnZqZng/zKbNnFy3YlW7nTGxHRk441fuAkSXkG1iU5W29uGBN4gmqcr9Sb5Sc1
Dn8hv7cvMpWsuGlKi1MBTjYBQVMLBOutOizo6LJ5ReEeKOFeTFAVl2u7tBxOww2avM0aRa7JY+rP
pbxuiwbaQcpobYQ0ObnHICAjN7vEmpr+ti8FfuMTve4HYw4Wqtn+gk/oXztqvxgu/gnntHRVJSKf
6QMxpTbQ3Y39+xdRZk8+Gtdxfj9oebaRnX6SdNKvI7JBV3lZSwdQr2vcfeuZs98GUn6mCFBCx9pM
IoVEOdEoitH24dagKodZEjvV4iBISHkn93p+g+vd8fYJheBpxSpqvHHy5bOMssuaxnIGrtFoKtgx
Vc/wRzlcU6Po3bEdmEEqk1H5bvzIdg1D2Q7ulvDr9OAOuhl5GV/YUf0bO2Jfzp0ppAGEUpBESFij
TKVDtbPpKxepNCrdGNP//MAU0TWHAlrT6FVvW1LiQOySGdo94DGRdIL5g1o2PEhgsde7SOUib9Lu
oLu2vEm/GoSHiWcUxS2Ls08DU06w9HoCUdAqUwOv9PKYjmvJ2xD1ZTCsxnHwy5gJkvO+F5IDaou5
HjD3Wg3vVasaS6SLyEXTB3qiyWkWql0LEICGZ4PV7JAXe7zNqfQrXA+4mV8nxpjpG7Ia8Mo8z/ke
u2/KHHc+DZL6Ga6HYheg3N67Rn4jwi9KArSHEGqobrBfdN6+TXe2W63bQTGtLcolfQHwnTHikPZh
SMKF4GH7WPZmFEjtPayi2vZaYvrS87qCW4EgbCY4sDi2KR5BEK4yeP3NbgYJ2pY4CWR0Axx8rOPh
oIzdu/8rW44XAOqif4U6xWnznk2ck6iPFv3WfRI3LGemWNWOROUOZintY/VWF+dtzvRRoQOl/fW8
EWRndhSBqnxAnaUkAoeI+QZph0gw0LnPICN/MXLB3rrJOBeNCRhUCrdzetJc7Tgk3/FWM99n3d9m
+2eFYVIg1tjOVsy1K4WX0/JL1n/ew8dm5myvMAq61IBFPFcYgul47lCSJHWb3QenfwK57urH/t/R
jatYDEZ0CL+QhYmQmyOrVfHReE0SvHvehwM+iO829+gWVQCM3VjOL53CzAF182VOElPmE+BdG//s
mg/+D7b3P/L/1zPYgQgGzM8NIjcdasLPpmJoB0NVTLTQGekclpYG/82RDzdQqoEzF85B2v5MWxuQ
HB8iNx3fyxiuci8Xf4+lIwC7MtiPRmIqOm/Jw/h3R61Uo9x9QWRr6AWVq/XJXZbKENELwRDN8uhh
JJzlcsu1G6wRlygFmQ/C23U5/KPqDMLRCPVk0tfh0MFEGZTUZEWUhOwMCTn34aeyy+XdzkV1bTja
xr/7C54X7rZwdgruSJh+NM4lKjdF9CKnqecEPGeY+0Nfa43RSUOcjDBvTeINKMoNROJDyHb3J0hg
FQkkWuKtCPfE5CFe66J4ma7VJ1/rrCsvJycGFtHg5ruNkBmnPUvohb7DzfBzfYcaY7yq52zfd9KC
dzp7OF9ew26e1O/rN0At4fD9UHOifYGVqFkdiYtzxYP7RcQ6zLi/28oj691MEK36UiODJX0GMzGP
/NeZWXtJ/i1rsm8Bz0KVu8JEbOf6og+C7ftkxqsSWze1DNWJ0OQFXT8l89MKotBq8eObARkUF2Qb
nf6OKTI89G4/wR+DYc3mEyhSEi6jKDFTc+1yDdALKjZWZGFRe3WcIggnSebgncVv70928P/pJ3fO
jJFm2RixPoI7QpKkQ7kf9q/n6trzF0QTBUwmuwQfDJL5H7k2aSiuf50hQRkiJrRSid0kFweeaSJX
NEbGz/0TBQHx7NpdCZC5nlHDpZ97PSNfwzwHTOkRaF8jG6Kwb90o3rURMUjv5+Vdtdtju8MLTwiK
qhs9TIZg3VUvuDdsibnqi8Exn9O1igq3c2RiGAdzbFAuRNS5DluJRu2J6Fr3cNRk5MuZCjuU9QBQ
yIph5pG6NCIyRNkpYs5LqDRo61K7xgJxTrjeLjCo+sk4Oty88C8RfhWAbny3KUS2LDcLEqgUJJKL
NrneGzG7tANgLJkKh2Ptl4rpDpy2KTH6DanKm++KwLp914wXweYHkkv+RdSbPn7KUbKMYIzaCN6D
FcHNgSAAcY3LCk/oCigPrZuuiKIfo48zxF9P7MKoWZpSekUoGjyDEkxSeZmqJ5rTy1K7RrwvzHVh
+JcGbjI7a3HLSZWeK3e7j+psA0ZBb/LGSggJIs7QhQaZBXwDtR8ZPokuY7hc6Rw6s+PnTIIxl5/v
Eii7hjY7JOxem/SQFrw2J9o8iNGXfFQAnV36rr6yIalM/GO1ejy7TorrAStV6bExeDw9V6q5357+
gDKdc3s86KupLFadPyNFjOialgEVOasvHH5uQKJIsB+mnz/deI6Hd4ABP8cTegWRZlU9jeKFGYVm
EFfqOU3wvIHNPexnOH+Vn6ImghyGEVF6Y1X3QSF0gTPoBnNVPMSJAOeU3Huvkx8jw5/r7qAswxK4
OnrRZoVp1ow6kFpHL1pzogH5J9cCG3xSFcRWmqGLU/NcAWQB/Z9he5zRZPxj1o9uWm+9pzJmrI6d
7VvB86qTbM+K1/t7RNCWKcLpP5oHVAVL/QrUEalekyARJb1X1HoqNa1tlFCMt/7EIWhAt88nkx9P
rsslcULjRTwJytJHcS+iJi8HP34Eyw5LsXgpPaYJhHwhEBsikOVxAbCGm+gvCvyWn4uzt5w8Tc5X
n10a9lXUUSQMn88AYWWlp/Ns9ynE/r2SyC/vA22/Bz3Xst11aL/nfubaVF/CX5PNaCnAg6zsNJfT
rmrrNzHwCHYsOW0x5fKFBqI3ugV1lkSi12Jer+zSY6YVdyZRqgSo4Q+9M6Cjp93WUHyA3Aqrck82
OKJjT9yVlbKnZWGcV2q/eg7LPaUFwqe5bLoNSYZiFonE0jvgc3QIhmf37zYil4DHCv7zAVHIOSOX
DeBhvHCPQw1zCSczDYH4J0CZeeDnaettvuntOsZR1ioapzB9d+ytmzFiNjxo8Qsf5FDKfxPCrUwG
OIm5JWrdVLRLPszxbk+igU84VRBEaLCx0RmeJhBTfVh22a25vTk54rqyxAwsroz73cnDDeR/tmu0
g1DOFrLQGvKNBA5nGWS0tctmF6vCeJQKShgN1dVfq9TsgkK4a0u7Z7k+oF1v84ssmHEUg76YQOqg
0wGHUAy2PKLRJJJlVmyjPZu2vZubrc/HZDIOED02vyeRWKd+VzoFNEXhDsYmFUWeo2ozGMe2c6ku
vtIre+Ifp1DXRdwLTJpOI7WhOSLmM059Naekpy5LoggnlKmhuTSwlboouPEafCRDTY/WdvaKKbKn
hOmDYfvcyOcjXDEVYOoCcSGtXvpE86gbMd9xiKJyaVOeRL5xXATk1WcxbxDxxa3Dbu/Ev4JHiifQ
Xj1mRNKRYidArv/PN8okPVZR1z2Qfkrjyp4nWhtIBIIbR713seIzEXwfpOnDE5XsOYcsKGfHlLCX
UiFCyjK9mxPgVvZbIo+JkTuoZOPKMxTAuitqofrnrESI7/hnSJDAMowCcwhhQCVvCDx7ohEsTKt6
zdMb0ilfcqkXNvSggqvJbGoaBsvFDNIZEhOIEHTsThymXgjHE+52eZi6V7HVbc1n80xAyqf/Ltfl
E0hW5+nUezYV3GSQ45sYsXk2OuUko0waA56eXk4NCfa3VCfhKzwOKyzZ21eHAFuezJo3Z667qy4x
YwQH8p4fXKHS6m5FLxs22hRzSZuUCx23rJkvsfVXsIS/UB8r6mBQrYyF3PJ8miUrV2jQ51pUuA2+
wXsgbF+TA1CbVAc3ga/95CcSZVdSAo5jfX6VqRNQGTo4ivfWAA9X6UWez/4bAiVbEn76BSkO0vti
vHFZQHhAqXeIrtJwvpKJkdADkEdVraDxYsS9wyBR1hJsnX1/XbR9X0LzBGWm8CwqLvxeRNqpjQxK
etw0Dp6Y3Wm9Eu/Csyu1NVFN6zZMTT45Bbaw/7dC38sQOcHqIlxt0TVaVNDy9EowpysRChTMyDfi
PhVaNl7gCcEe9JaZEizMAGJg4q/oONiETj+EqfQ5asYERJEfKH5dd9yEWAXG9m8eITplVkF0KQW3
s7CXgnTqrRivrNz+ZCgGvKSomTJK7lpt9B40/qesvAVeg/xrJeGaW52NsXR1txG2GfVmzmG9AN0e
bpjD+TSj2Lfxqc9ZlElt+0spcjFIjhv6aiG4SWrBuK6iaYTIBlarqvta+wuFXMzm1GAGTKKzqBEd
DO7PaCXYb9vRZ3tKFl9IwK22J3vQ28L0e1ijbdlCh37vNO1Ckt02pzoPnWcZ18zO2H3ncDXHcaKV
FAdMzdQPJFBsyY96LIGdIYrunMLLftORmTEISBJ2qGkCh0LWnuDGygEC729vYyhM7735Y+Rlf3cc
v8lQA/Yq3pF+F2uG3Bsyd6lS+3+18afpKTl0CVWAssE7w+iw7LSdbgXRnfLdy/ZLZaPJDtCrjSpt
u3L+Bn0nunmFQQxQwgBp0IKj2IMI4m5AC2BrojXizKFGtS6eYkZfqla/rrp6y8iQqHqErv4qH1C7
xCpOavzEKNZtKuMka4Ftk5UxNMyPXAt8s/UpMf0eCzFaul3XjSV27sF/ZHVKlMqltB5enhiuKwXH
wtZqhUb5+Fs9NCl1zRnTykes/JCuZuvv3jX0GMDoMKfrqfQfD/bJZ0Nu62FjoFU2nZb8beJli+m7
+FY+aMcqyny7qTCxr0kjekvGYPggqmt86YNOOiC0W8X0w4LSLzZICHya3NnQsuvwZe/EB9KJTtKd
0CjpUqMpSTDhTDjY0HqQYGacR7WID9fprmySxyiyp9iTwTfNvdyg8eNao+xOQSlz/0ItuIchDubi
oJjwXjIfg67rPa2z4zuO70CwCNtolnBvKzOK+FWo1F4oSV7rG0h7S0SwN91brnPCNbsLp1zPx1l8
d//vxn3j+F39dZxcA81w8jWJrOBSQf70zEt18CO+9uAvQ090LJALKhoYIvTZkIp3kXuHDyYlN4jn
GrsYV/2NCXRsj3xPOFmbG15RyjqE0uOTKAo48yD3MWp2YJNq4oJX5p9GINqFuaUtN8vb34WIvr0K
CGUtf2KyS/jb8uXW0zrmkQL0/emg3RPmcJl/cye/MRoNxBKXjBojxE7Uy27ZJ+z9gsJnSiNDdYDR
PoU7fhM5lbDi4SdIzRmvTnAbiF/MnSUYEhfRN/7Pt7qZjoyhqh2edvKB87FbVbJ7SsoOIGGiOU9A
Gj7K/RA53DRg2cHUiJc9eLxHk26pxsAMzAUoaL8F2/6P/w7srQgXtixgExSRtOhGnvZx+9dGe7b0
PRoXjcmaJ+XsA/2rQu5JuO3xn26p1F4ZaqWOEgnsiyKxsgSUEZ2UrAvF8hxrfcDtZQLDAeYgwbJ9
58p1xJS45IhtqNsuJZDbCJqpDZG9vT+Td87a1uvXPUgEh3tgz1Zk076t3wvMH/oyxj7kigaFtjx9
7IERYq+Yes2Ij+A2A7nbKCyVlWt+zFT5sDpqMlZp4WLTsYTbETTluRjCXR9r/Fepu7TfGigrNug7
dBYa7XiynuTJkHmJzEW3BMhBTWm1CdxoqnAzjGvJMiqvFLHSCX0LvdRhCuR+AVNNpFkUFeTUVsK3
4nf0Y34A/h4NoNwdSEo3TqS+ARETOUwu+LY10y/78xx9yh6uqqQvtGL/0WQ3xZMklFZJv07a1j/7
S/H6CQHn4LqTBn+mOXeT7qMRfKswO1A0YSpu3ctL4cs2kprIgYQoiUBd7rvO9OXCax84wYI1jwGS
BZ94l8hI1wBG0ikEpVNT2+W/8uT9UZkpH7deHwTwq8LF0laedCGNgkRlZzHnJh/1oA64/Q4wRejL
603FyZNDJPZQe8vna4OC440Q6jbTxZa5yE2PfoRD72JxVa9CEhl2dR5qCfuHuroIjng2b4aAuU2k
TIZA1CeFZJJrOErVNPd6FDK920a+NxfV+AE8OxWAfr6Dp0dsowPTYn6b8zbIbT/xbziKSxdlGzzF
2/rOVdVEhdCUbgxiVAkqQUwU44K0xlj7ieNiaj1WUXIza1h1Ep1ePeIQyzrQmhsvrGSFCpeQF5u2
likeO5grUu/roJKbcE0akGD51mDTnT/Y3rsPF1S5BqXU8n1hZgaGfAPI66cGAvFoGwkZkXVXivUs
Yisl10mlIb1QrxRS7C6oaLl22xqWNzNC9hZVcKt4MDoAhg5cz3m4pO1Ce/5iXSZTiIOic57viSdJ
gP6LlBrQ+qt+w3hiRB/XyHAs1TcAEJDCVXl5Cnl8r77PPMOuj95QRU77Cql6sbjMn0779JW8QVU6
ZFmBVkZ059FhmD6Su1llDxDsz8fkHWBhQKdjaCggcDNmzc555zEKHV5XEYKAwwiv07S79970eD6m
6Gz+e89onjstSHK1GWPIkKmw95MzjeDGGDKDVh2lfcvmhfjtZMegwOSmIK0kwKHNVHz6dSMjNkds
jdoSeZheWwLVtK+xGfIjQEnvsyPKwiuUw7mhlj5Q67jQHAmB1ZW/anfbBkq+6nnZjSB++MZPUhoY
KKK01DRrlM0s30a1Qd68Hzxk0zrtdL/D22fLMi39m4RqJcxSdicVrm84qTeDYYae5/IqguuOz+63
N6hvBA0Pyh2u/4Rnecogy9yKkQN3GLGBD7xCfGEOi6vfTKcBlKNVLOxKGHhStRVT4D59T64wBBAR
bceWoh7SkuG1J0fnbn2mjzgq52Bs84hUjSiUSyfqiQDsg1ZTXHe+qeKvLV01JuqYCGI2EzsTU5uC
qm2FxWAFEjsXOE4X7Cwq4P3jHrpxwP/SCT0X1BJQlX23SN+c7f5V8ujQyeP9UXUn1SdNADyG1kn6
yjoYtU98aXrBSGQXMIUO9a/eNRwAQ3WRJD0bPp6EdBeqCyEv+CBusN7MWPXRMKrgYErMHmv2prrL
fu/qHNzce8fpMn40MYjtBxytxb8p9IiOJPWQF2LkqgaDx5vdtiGbxtlNwx37pu9hsJ3pKCX8HtPe
adzk0pG1U0MkZDTU/BfQsRw7OM8vGotRnM7O5e90bmFB9TDRsjT9Dgj9elnfdSdU/Dbr0ZQqFMcI
Bjg42RCJPZxzjvrNmFfRs0rlGaHhe3xAjpK6vKZh+7ThBaaUGba7ZHV/F7uw6L0pdyooVo0YgRtX
Fmrume3FgW3OtW2RyMisqohcQXgw2y5A7k/upLmyUxro/p/p9YOmtlPejjvdDWZHtydeojKw/MXD
f1btLeUZnZuNcfmwMh29Kzpco2gfszI6OOqRbhQ1/aK0vM3cqpsyBwpf3r09kGH9pdneq3eZaKmQ
J6tT8cvAft2OyN/l+R3yVTvgwe0LPi4Jt09bABk44HFyhc3kaC+r5xBJizZ5hOwEhZBzpeDAgxtT
XBf0kNfyd5qmoJ8nTxKVZWz5LKjnYpOjU9ohUlWGgMA6WZMCGAu/M/BPA9nK0om/m8BmX9FyxMYS
4QGrfCiXMLARq7BfWduTb0UwHmD2xjnhcvlZeNLwVtXh13krbSeic85gvgtcdBNSBdiYRr5AAMIs
NosqA44Scwu3N+t59xNJUs6YUwL0PHHvKQieGur4lezr8DisRPUREzigSHMn43yXiYxYIVDtl/he
bFYWcB6xhSg69LZUZFoqpyq122TH2s5NNd11ZcLPD5NWZtCvdKmT/fl5k2UWLyVsUwSh/6z5Mor7
ZlJUFDPe6fwtt1ZVmxL4gHZ/J6xldi0aM886ebeYZuuGzHAbPIffXJILQj0GtmQXe+4o+cH6ivS1
i5LQH4H+ARjMCb6shwAP4sekxr0nt37TEECzd0Hec2H7MuV1jlE7e2v8j3fe/rW9ORTJqsOvHyxb
pu4GWwu8Igefute7sRZDb9rdJATkn1T5g1bXs5jR2vl3BmbhKO+BcuBERLA54kF95eWv9RhSt5Qo
4g2en/X+2aKXG9LKZEwKPEa7I4MgKFMHhbIzh3ZyexV/XNa8Z+AMO3TPDnbDLilY5ESbsQaPijJX
xSeAq5G/IkpR/1Rwahk++2O4VF5X+IjeMJpwoJHG9LtFxhnZrBn3d9ZKU98Z4RgA8gmgx01yrB+4
+ZocU5g5IpQ973lQd0HfAGhj6pBiv7Z/cQnnVijBEj0s8QyA7GIMt4PTqtb6srbv5s7puIM+ZR8C
vPismcUZhoHviF39gQhLNxsUQBGjHTkueA9XBo+l5PU9SSQKCgwbM/1G30pcG1tUFaFxMfQNh0uy
nvjPLxNhUjt9BZqLzBhW9mYuDZfakWoUMJUztx/exU+0UihNBRtccRFYIMg3EpK41MSMBIRYXz8S
Ai8/RF3wqhRDLP0maBZ6LRN9cvCbt0/PQfAfsqQFc+KcZpDD2z0PrNpVu2h+2uA0jiL9uVvnaduz
rcjmMB4tPNKuaGE0lu+au7jCfaAW4/ziOHFAtop6GG5LlVHi/Wa+kkrLlBrIbJFtJYpWC1hN3hZC
ydq0BgxjbJcTQSxWd9DcyzOI23riHrnGKRxoRD3l5OSJjXB6O/Yn1NCZrGUhgUoaSZWoJ+apn/RG
VtrITrNSLsItTQFzTvCfcXO4+9ReVfECOmhjvV2zreasdiUsgTkqW9bQbJAHrTu6zKVbRxboQ/AD
s4+hn3/BQFNw2EsbHQvRezngaT36n6FbHpt6bo4boGP2GR0crM7DCrWmCXZy/huXqmc4J+5Bfbm3
sAvoXnCv84a6laD1C+tQ2jsdxbZ+2jVQFvyN6RYBscPWc0Q5KIxumfznCHVPDOf5rS79JmeWIlpH
xyTn2drNQQuTFACrpXbG9JsTuqNZGnGzmj/O6mY25LLpnjrGYj9S2k0UEhK9N764hM7s8n4BRVg3
5Ezi1uruyBTVRRwur9KCiHjMGjvE6qs2U6DGEi3n8Wwq5I4FbRvl27UpBcK1xkrKUnBd7smgKrGj
bpwuFr+b16qysR3HkA32xk58zdJCQJdwLu1gc6m66L3jpIr3HABl0O9w7WegAxElMyNI1VwAInz4
0G+OwqC67MoY7g83Ro+2oZoUxT3iizt0WFXhd8RnCzW3eDvMY1mF991bK1MzvoGxaw1mKTe8M3Rv
4qBiCGwMfANhYrtj/vSO8SXSOIEuJxTQVwIKlnFVUlJfwUEQ+rie+7gjsixfDfunoWPnjmfoIUTx
pzEcT/ZaVRsja5xKklJepvpx3KBZhryxinQRPjblsPuwdIaEmcVr9/6YwK8tMIwFxd2P2Tk5WiZz
HVjm4XdbC3JWC6hpDxa6oCUQphLvEKGy8/CnYZ6V27LKC8qAgXhgpyB3PazkavEIkEoD+qbci7Xk
Vb7oo26qN6EKjce1nzltgm0gb/ZLJfwdgCIPfrEYtxudBQO7Yr+bY4OJA3EeUhsWUqgEAU8FjXmv
wQmKuAndLoI5k0gBTgoV+p80l7Ib+gl4eM1mgBEcxISTGoMToXgylXSv5dPE3WOD40rvEYeZLEjE
3hdg5r+kRFaVrdGWpej/UleYa2MqB0+jLOJrE6kplsD1kulRJiIcEC5aYIuXEVwqNTCLPwjppn2p
HbFa3l2OH/6DoMuQJG9l29ES+bipOLq5h/5rZyLX5OtRj/s/Dx3075DTjE6vAudgCXqCasu0hHJZ
95usfhQexBwEzDjn+BCIMgY8s9UWxoYAhkI8T8WVZO5YL7hn9x0I3KS8glNUA5keMi/tPzUhylk0
m9nA8meZAL+fPtmhAJZ/XOVysEZgk33xuTDzDzcdUeEAAUuLAtWp/xXZ3l/H22UAsvOBtmZi354+
xwpc1Py8P43kOqTPY3A9K/gJd6A0+8jUsq/DhTbETfYVm9DUqZspJJ5rTYVKJY6/zzAtJziwA5Gf
Dra858GutrxzFQ+mULn5JlBPHaiaXvcluPiBv39gX8POn3YZ8RfXCTJtlIpW/p2iQkrcTyPWYsn7
uO7NqxwD6ARgUBeOjUOt9zc0NwH593Nz9Q9CY6wo1y6Myknml0yxHXCVJZNgvJCNw/N7ET9ctb0u
iJ1WERF6YFKCcFhb753Fi/e95b79wBxBptBBYlhR0QHSwVyS7/U8kgIRPJLEO758I6HwPPa8mO7e
c7uc+06FQDKAn4WJUP7Q7FWrfxzDpZ4pYZfSFCpl4jPR6J6nNJPt7qPDvG/OXeqtlryR1DHLU/Cf
bkfb5ZLIXW8eCGDWtKKQM3FWsNDhcEafaqTIvGizTCC5RBidNT5nfiduSSkfQD6V4btWxOdIuBgO
bDXgL4Lz5O+WHsPjcJPljwlmlBrLxTAtK5uWJ68JsgJDtp72ymeGtxpqRpFACdrtz7qPSxKjX7Zj
0QF9u4fl142GYANJdVLfLUaoNevjJrVoRmolAPBZdadouv9itrcWdfK9Ia9MYjFpJRy43IARMZFr
lYs51Gw2iHXwHb/I64NbpAcTQo/T9HN3/L4CpNClgfzSsAWZNAXSLpp+mUMXNd0z8oyA1uYy2RB2
tzTkgg8jr3XsjzrbMlsbqMPX98SgdYkPeFYCWaINQqMGbOTVO6l0GFa/o/ZBEVU558aB30oJup1K
h0lsxtDgBMRirNvGdZWXveIzDemcnBedPKigxYQ/MH/WTVfe+GVLhV/shqNkXvG6CH2NMaoznfQ8
289mMI8pJp5yBT2fxtyQCB3JFHuWMz94KgG7XYJNqqPJDCNXPP0M3KVqYVqhH+QmRBHNiyOkAStE
oAW3GI5Wob83U5Uk8/rNLZRl7IofHmjezXXqxJ4rSfxwmfe7RAk0vftctSBnMAgb/d0IDTZMn1xo
bzRqI5rYG2/boeENiYthP30Svcus1h1GkQr+jQCQAjasWKx2+WYOYTeNmjV3zdXWtFtFO590AtIY
f92Q6oKsqdw2uqkn5mABxaSPJGuqs3hjhK3pEgbp1TrB/We03RbidDOK6bUZ0sdeu85W1/SOKe6c
9H/HigTREYDqgDeXFBoJp4Ae+2Pw84CcpGlMbJlI8cOicZpndmDqLC3Hd6dmnB9eSBVCjt64NIST
8i2rkiRrmAcO0xrpAx1ykkMUvHgLYgU2FWbBRBVxFVi4EyyWfGmJueTIkIW+SoXFZCjAxKP4xeu9
giqETOYv0SxesqO7yv87xea0gVxTJPAY5fIq4f7+ycigtRu2pQRcVDuWg08o85oncIBTSGvY0/24
RP5I3KBMg/CnWNTWsqg3f8KRIDrAx2qYSjrvNN+gDMq/aSK7BXQx9vERFp5yPI6PbiCBMoTDdOIe
B0qUzjCHNMmW8AnCuTq7BZaIxeB+xh0qzMB92MIzkKwUCw0OoI3sVwJDNrk+imv+mW/CQsFoO2ro
PRMYhRullQ0mQi7HC7E2gVOqFWiPVGvAEuT2p8X1NRlQunFP7BWc2oZ1kLOdQ2FUBkba2e/IborJ
sFVIK2wv+ro3py/aoTcekCXbOrU1xmcohHH75+RcXjFnE74QEueVhmbngK0MnWdEAXsw+n5pIQsm
eno8IsfTKmZjQhr4bdXZkx/iZU4QfX1IK+KdZNJzusPK2z9aGNeup7a/SisY5Y7mEAI5gRQzKS9Q
fAOYR1XsdmxltWZllwhhfKIA4VbrBIcMrCDcQzW79SVBWwcNcKZyWqlG7TVRwbyWU9S69MX3E+3m
JH7ng30typOvh2bmiWsZe277/WgyCGBGUFFLsTa6MeMjOEIM6Ast4Q0sdGffmS4HAuR0qyAC2gM/
OQ1AnM7yLuf1ksb0aTUdBlg90ROh0T+4yj39tNXWDT6glsNuuEVNvJ/wJYgPJXXphxUgMaDvroD0
R/Jv6imwNDaA8KJDhviEjQBPc4Tjjd8MKq1mKNXflMgDkhTOScGHBKh4NgzrOcJyiuDA/pgPcMdl
r0b1GzvqgqC3c1JUgPLsICe9bSfq95iuLcWzQN3EXhuCEDuZSSj6TZKQPiTG9/YWlGqspf1VJ5iB
4SlAFIhM4g8y854M6Au3sW9iHN67wBoFZUkPiYzKGVw7wMlDHJIoQ3QkLVHn2BRfc4eTrPS72Tgl
6EtSQwxB61xGw4vmJNaZ8XsXew6WhMVAG6PqRFR+x6OtXkvadJyXyp+DcbaTgff2cONznYx1HMWm
ssOb0HHF+tchczNlkidjtXl4YEew6/iHcI9LFf0Ii+rFsUmC/D63i7mjRlSOy19RsOZcdD6Z2eEL
v50yjzb4+YG7STo6WlRsscKNSi09Fvnf910oIqV3T4wOYLZMs6t/7PNY/dbew3SnmVyB507iCItC
8WkKT0CD/tiQSoatBrpkADYkuTMsEote+Nz3vbtNhw31KbAoZWIz5MTZwpWy2gIWZUtgtK/U6vDI
to4KAD0uEWyrmM7h1Fy1+2KlMPodGdJ0piKqo91kj0N8b7lyNtFSzDg17fHmz6kGBkguN4PmhsAE
GvQor9EicScipPMo82Yu9FDwaJj7TqoH3oBNtAB7o8r2HXwkZlzRaw0TQFvOKelIpU5vETUwRaG2
xUxoAln4o/PDjMUvdcOIu36xaMLnpy9CES5mOsW+bEsefiwElfBkzGcD63Qd0yNWi9S3cTzPGBU0
/VOb5Cae0z0dRdUs+uTTml4H0w5xddK5bgxFjAO7BTyEmHr3JGX1XN+jmkgsH0TbCukVnuFQmu3k
lLIxMIYT/E6IApkKQPz1WKlLFtpNmr/01GTAqc9HwLm8meP6zkO9W6JIXG+I1XAPDOLojsDcYCVK
eQtv4/BydeR9Zt+nVMilc/9KL77rNx/p1OCF1dhSrCqAj44I7+u99JDn47ViMQQG+nObZk7Fu2lO
9HQDwNUS4OKzGNmwkRZ/eWEqu83eG6cSbJvxgYLR8zhfGYRI3piiLIFN3WHK6obMqZCCiUpuX0UT
ob9+vNFxrzBzEO9arbGOENsQenmbC8NhBxn9p+eWK48Faru9J0yKMIC8EyqbBzxfly8EbM7H07Mt
5iRZDYMk3g0QeEbqgtsyJhjxF8P+sHwAqczqFSPse86dTzFs4DiYU/zrVHTXHXGf8+B+iOL4EXWu
QQ2MBGweWxyUDAcSOLweG6ye5k0Q6geC7aCX59IvQw8RH8I3Te34suAxQ0740HDKznaqHwvGej9T
jTAwQTFMgcYixRuuybBkPAyECMBz+Izuf+HV8ylQHkOILhYuWcRB+LGxCFuEWvgV1/FMgt7hiMUp
j1sg1eVhTuWxunF3xZcNkQpJmVroCJYh34jcb8w8OkLfuAZPj/XoM1iBy318WdjU3pkb7RkW5DXP
HMo5oJ2Rz0gZ+egf0ckPGsKcFVnq+atjDWBXOJD09Cr/nPNJwe+ppIoJFxb2/6nElokDn2UpO0tM
k1AoM5BPu0OqClvwDTPC5yPTNNFFo40VbbLSs9PyWZGL3C3oU8sSWmHxoBvIwPuicoq6dcS0FgK7
TlN1FJkviJCrCaTEAD6D5Fxx8enXZx7zDK0PwKvWEsgzRA5ldxgQgR9Sehhvt7PHVVWepO8mFUDN
WKdbGwItkJyXrI5ksEb9JizEVZr2UMHqIPTpVtWCY0lpAx1pXYq1U/QvV1mKWcz2UBgvNkVRyhYd
iPK08Xg7sEXnFfXz8p9uCO1iWPDSm3MDyPIj5NHrApgvhB6a829K9dotVwxXfdRW8AUi9qsaoNvc
c0rgiLqSNGHVyHetNQwD6L4r9rSdurvD6k7/VOvTLRnoeAgDa0PwQE5wMdmJbkZskjtNVxtmEe9m
TgqQF9odLXUhab765PHHFPQWxGUTuq0jJnnAJuHMIQJKCtAXBFUDEPbhX7W+mXMOnL1Pg4ayM3fb
F3B3SBcz8Ko/I3MZZhqYn8zSRGXF6HSaeB7CaP7WaaprUw0DZqsUPlXLnbTPgv8VA+qsJ7gpEmGY
GpnMWH9bjgM1CKe+OUJia0I5dgMq3D+fo0H/QC1K06b24fUosZRETFf2RdP+YNZaF0PdnyTWBFOB
TJhBV0gXcLuSsNhor/FldztnHNFyGOtEVbWSbDMDrzTdNYH/7c1Q5KXgAEy3zbCpq6VxHjsazZXx
4VBS4jwmG3+zIVgoD/0Md0SpoOXTSAKvwCoHRDNo1FWJSVHS3UcL40JHj30LA7zy1pLv9BAsebDE
9XGGJMp5HUcza3uqUAieTC3uynzkSIQ7QU2cJqoLfDdj3fsombTts/8Vfu0NiRuCPx5oYIN1GuM/
ZeyhPfTNMUxCnO7vQiqicOq2IZeNTfJlxu2tjQD2rxVevrlTEA9RnUciyrK64C/L1JWvKFr1EzVQ
O2hqgzJZZEhohw8iKssv/qBb3oQsxtX8791uCv0lduIDI7TJq7vZu/lWiY1dv07bMAuO22n8Yrjk
7SQNFPMvetqqjWmFwhTzdIwsTmh14H+T4Sm5cGnJlzqYhwf65aEk+mRQCK3l+vywhzpTXv321/jX
FCUPr7Sc9w51Hes5uKbAx2i3ldaeaWXCerPfxBimN7mQjN2rN5IY8ql1TaehaNe/bKp3f/VCC5cS
Wj4ovfSQ1FLJugdu4lDCkYva8v8XMvJ6V4uOyIIp9Uc/0euiUKLWWPUG+183hbmv7jMPYLZKkj9N
TvYipOkUfuij/CKlABo0AF51uKT6iCZaASIA+FWM84PJlhhTllgi+HE87Tt7rGoRdi6LfR4+tXV6
70wPoufFWGoEuXbuUbi+EfPeJB7awmB+fRsoqGoS8rUqbg8LrpCbkHVdBQkaehvZjnsgEXfrDhHt
6uixIuasPCj1wuiXmvs6fsS/cbrp656egVXbq4gX2iOzuZjXwjGgzk2WNbRDRe6LSy2aPXO2KJHe
ZdkT85ZyriC4tfW/QeJBWuvbcfOe3sCft83C1rdu9QhwP1038Mf4UNkPthYF9f9YeQKrw8/KWhmR
XI2dw4PjEYuXXrU1jc5n2C4wCQMBPV+zVmKQRtsjDzvrKM26w3oxHIJmXipFzLV7fFB7JWEPCsSo
xtKerzyELd+tL9gWYBA1D50jJQWGTLbo2/Z+HK4TsYIk1c+g7UfS6PTkUY6QPSyf6vtp6vr5aqf3
KDMQYlYdRhT42lNKP9isb8QdxIMcZxdSHGwFmRgBpM4sacFzSoKLLaNJSyi+0LGzQKMnNv7gjTIA
6gNsuwui0S7/SJvbHUW2pGIlOf0BC4UYFzOlTjK7AW4gE3VtU8RDCjYCVbdwRmkMmgRpytB9bgZU
6+tfD504BVLA19KPgoIxDJh0lqQXJ4L3VWOwX54dXUZQ56EUnfonHmb39nKrfVMWr02ZEdw2RA4b
LiDyWJUfKpPrPPyCqDyrWtA4iQlW/wuU7XVgXYHaJrnpQtWRk5U4/cEarNMvefn73vOKasx7AfRd
eWOEjuHTz1IjUbfFIoUeeo6XFsKijB8AFrVEfaSLvIlNJfR0QpMH/ecUsvv94hxGnQ8BIZT5hRcb
do8BHt6s7tzv0qQ6aDGGJYEECSzoKrivRKN/owgxtnPcurNENGZfrN8gQErfapHPBAj5vO8kEoJj
VGBnWFzcwG8Iis31dxFEbyYMOmg+mWIX6Z3oWSjjffacSN5W9EpACL1lprNUpRw4xoQGWNpt/DIZ
Mo4E0Q8mJNCwQzViTvmiVXJGBlWy+aL6OUQg5LT31xwiMa5DQlzRnLIlCKO/2lgdwEwn1fXiBZGx
0DK0ezyIIrSLR86jIxYSEzK9/b85pMz3PVS8lYngHtvw6Hxp0m2e+dme9xvC7mUEO6+LJ0ikAacP
ui28/OtO4Ls8GkjnCnEoaPyuTi3lT0brfthyuAo4QdDB8rlqvVO6HYarkkcgt2Dfmiurv7G0gPUx
5Efq6l3sd9FeY6miGWctVa9q/zLNqfDMcbHrFmHzLbNZhOFMY8SfZeUrEF4YJw7X3o+U6NFwfMWz
Ti8uV9M5ZEQ+YWMVzE2v/zR3GTLHJRv4vGiahvlbT7w43Hg1HHVIYXKqOuVjUL08KOtQRge9HT0L
UrIUcyjyjNLLsEMGEmeQETCWKikGzWg+lc8Fme6VOH5gkjvU2Dx7faK/4htbZt03Mn94mQFc1OYx
IN5FK9ZzHuDR17FyON/ZHDUiFBev8PSSUTTGnuinywYVNzG/+GLcQCbKPhfq+t0kqFIiZJEdbj7m
MWmNpkSuQhurs9DPZFGXVhu7BdCaolErl/itOQBv6Ye8EaJp5+k3tIjxMAIgBVs24W3QR3oD0SUS
EGNVCBcwq3c82A2v88GzfWVycr4Cgs3vR+PkyWb1g+xr0ZOXzN2vZ91OreK1x9ajhAvBnjfenPSb
6MXf2BsIxkteLGsJH34OkGJYIscBEddl+NvMbZk4FVB+ULQaDYdRRm9kREhV7k1FdBIzFTUtdTtQ
mGP7c1BsyLs9mxZxAXZfoGCd7cDKtbFApoEUX3/NpDrTfNpU2dqCqtwOBj/Da/qgPbR7VX1GsM4F
oDaeePRySmKtgpqRxvX6TM4Hxf1ZkemoXirP4UUNa3l4ZIRF/blq0lOOK77hS6hRus2pAriO13Nl
YyY5hpzOkiGnwZjuaxm+KAFMcPbiazpZswQZLgmnc/iJh+LyCJrzCgRxwNMveUJq+YOj42h8/pN4
zUgOiaQyetHoIQCs5/lBvoWXAroxZDojgex3eCzYwGffg/JOzxvVMSnocYFPotWPoBb3fIvDbms/
pubjU/rid13qLxJ4ha9NzZ0E8m5t1qIMsxBCDhz49zw9OOW2sh2R884IXDictVp8CHyxyv6A6sFF
svRbUeOieLLo3XDJcknHmOtR0lk31ei1oeWtbXVNSNAqsPjq8ZIcePy+1IQ0pS5Y8hPMXCt9aPPO
oiVU0XLEhL0DakDwItiYs9PNr/KEmdY2M17KaC1nFGEgJihMvpVAwpjiFS/dyqqsFn88T+Ud4nee
boE2qLeOQm8+4AOXhKziZkcD1aVEigBh8uWkfw/r+rYcMSCS9H/Dn83hzA8bO20Uvr096om+b6SC
J5g+VgcK83RnNBNpG5mLjvlUz5gUmY6SWc1+9JSxJnBLjUobntPyyS3X2ntZnkKW1vOc7JM9Uy5v
yjrEtjBEvFkz16OK4Jks990BGWxy8XQJq7b2g7aR3h74VvKvF2uyY1m+/WL7W3XPS2khdNI12eRd
CWwKwVPamlRv3TqkyOCTbtlR1yBHxT+3xPLILN/2RD2WuTpWgkw5XqJ6aLGri0sdSRfquC8IhCce
6GeMTd2q1kqfybeq3BtU3QSgD1wCmPHqn0rPAoFyi0RKeAcYTslLMkxad7puSAZIJ2evsqer/KVV
HD0IJcWfLfUrRY2/iKn7+nXYl8w3MBi/77ZDcvzQR3sBjUjNZkPKMoV6S8/ZVmwn6nN38FiDeXN+
JstYFcYeffR7meJ54+7FV+RE3iPpla9J1cPGtykdVGHi7ZheOGLls+MDOev8QsUFg6uht9PBylwX
/MbjCy7SSbmraD2jg+AE4h6hvhSDfIVl3TONNrFu6mDLa8mYI2k/l5cLUr/qr5nDrPpi6nATsdQ8
srKG9lDZ9/MSwFD3zkW/aDdSVEubH6uUaj3HFRMS4gMTRshKwLoScLeKL7UtA2gOr/Y/45xggICt
ua23R9vUH4faZWU9W8KWeXfbCd00yU9Q38VmuUMM/qiXzA+tpyvYittb1Dn5CSd2S4EDXFRznYiP
pIMJkagDTrVgEsyVHTI7p0M1iiOQ2DrCto4FUsqQOSmXwVTtTjS/kehYm3SYNir/m1a/9sOxJ5Cu
MqcJD085ElYnXAMZl2RNoWp5nj0zMCkASQ0Cm4TMe9yTU87rXLBtu1DZwW3IZNsaJAZIwoKQ9KHq
9vH/BNx3DCkB3H9BhuWIhElZgfJhZM15vh7bJ0G2z4qjIkaqmQVX90syYIAYmauMbmmC5+pmS5uY
QV8JuamARp0uaFtE7RRvUTGjDBAq2Od5L6pTHSZeaNgW2F11LrwRi8DRbLEss0j0lTaHw9qVQFLg
TNBy3zw4zOWXt+pNCuh/PI/AKjoG4RQxc7ewgQW3OVPmPzb/Jf8l0br2Etvk+HNATgUNawWReZBy
7bjdkZiZRxLoTRh+/+EqHCEbioYbxbQUubp1zCAV4hiW/49RxKcW7uw5KCQGl8UeTrE4Be/X9w6w
6CeTIp0SfShfbilVJGEiZ11qvCY4GJNvgydueycpgL4HEZEyaMrMCC4VBIKjOVMR6P44twxJTEDQ
lc2E0aITUeAVEd/mC2842Xxt+j847zIVHNKiGMLTEFaIWOJqO4O8A159p57PvQl3VnqEKOQoIZOR
JBfY8xZEvA7dEkeD7qLgTfjq1yqZ7OEKMQTjMzRvF5Q++sPR/8IX6yhqGiFMzWeLWH5zUEBjqrV1
FSWnBy89x/4vtJILfpmeX+v1TF/ye5b0GvJqZSDHMTnI1U4GHSFEtQfWTNgWqOl4jmqWfAjin86x
adwYzkjOHyxJ+DHe1nG75u/4poX0A59Azyt45qa9Di9qW248GmwAiDEHfyp7x7fw465uPdeMyoB2
5k3X92R1BZ7dXv4pdOZcRhLgNWKz/Ea89M4Un1YHszlW4JOD+Qd+G7NRStFGvmUYB9/mdkEc0Mg7
XinkKEEDMlSzbZDjiCSi3rmnjDRj2D/lmps1EOMNCtYhIW8B6p6okjUNZtplTl4VcVDHzDG9PeJA
ahz6rxvynK/WSPc/nEXAoRbbGuNf010fVefYVr9E3ZHv0ZIb0CisrwMjZK60Sev+ymDcINDHGbMB
4NGjPRHyBX/8bhrWwoFzfk72EbZ6HQzYDDeGyzwMVkYzpvPe10G0qR3lA1InETP72LkHFHZB+vDf
bcXrl4RE1HJPXf37YMpWuUXrxe4KxagFB9XM0SCfKNNTyDAbgc7+KZ44LJdeAlQTU/a3wOmgb/7s
JB6Iyt0D+fJhMR+RppG0+DkjoP+WuS930z2wrpInhj1qTJZYB2niGmNo6puHKs0GJllK8cRO/5r4
RxUbsMT9wEEqUt8tUclsME8TWV+har1wBE6guVZbDyU4tijhRbr9oWzjjR0y9LApJXWj5z0DYI22
/w0dROGYM8MuBohbUiBO0N74hSg4lXNyWwhNHcxHspf7a3d/aWDpuSu/jYianQg8Sq9BLDvam0Nj
a2vpBA7E0MnmZdIWV5Ax+gPoKZFaS70G+u3Z9dnVyqGLrsIPh4D5BZU4UnSR+eAJ9JVTxYxcENoV
PZihLra2wHg7tsprrIqqNq0H4qHH+PtJwuCRE8982tTDRcxzx4yQrx4Pa8/4UPMvgXjjmyWkGCpk
VpdsItmJl0WcQvOWcCP4Dpps7IS92Mi4yegRaUNkjYNDpgIXUbu95LoO4Sk6wa//r3BiNjrXntDJ
JHLNmA5CnYQflWNzR/YeQbsh0U4meMZ+S1zvfshnD1es5wmnUz7k0zRXAkUlJNMfKpsIcwYHOjac
J/Bpb0JbsYmi6MfzrczEEflIEWdS0PRez1qGhvqnuep3iEv15dVh/2cYyci4ThRrI0rD7UbVscEU
U1JKZGc/OxsHVGioyLRr4PPBuMFAI6A46mBcE2N/+4BXUku6Y0p39oHiucqS7OBUEpuyP0Mi9li5
ZgZ5NOAWV4AptGHJesoHhzqcLOKqxaDAbfMUkZVUTgcaSBXfD0iU1kQy8qKCSSUfLQDn6Qtn59uS
lzSs8fLI4mCl6HJFHostnQ1668xwdIjDSJlG/2epbrQ1mDOyUYSAgoxTyhvRXQc+jOQXgj5KuObJ
uDovSTIV6B4xPtQUsbkGi2YLYulpXIfE3aNJF5Hj2H+eqbpauUF6C2TevwZUsEwGaYK/RryjaznY
ajH4ne00oBWUsoFRQvlIUezGjY3G6/BOD1sVgEnzpU3CJkeuL6WH6xMCSkRAXTmzjE+sy3qWn1hr
8rVH5aQUtsibEHjGlfn+UlojAYHDqjLus4mqlz0HOeIyRvIP+0aU3vdOVwigccxLXfwpT6fHinLX
kVaxV74SvjZ2ZDSg039paZWHf9zNKAxhedq7RIE5PY3KHTQ2ozhxAmQHbheRFeLcv71tbtgdfxgE
50DTdc2Rf9wQMmhW46EjJjmfVBdFqkIvXLlOqCwwiLTZw0wJb3GvRBdo+zSqI0H/luynLVD2eD/h
V7iS1S6uqYj5ofITeMj3vyt6NEIel9ppPAieLw47ksfzEsUrJBlhqZy10A0+F5/6PGEYcXOEUZGt
HfOxFxCjFDT+ZatQ4swaJvCxT+VtxgJzvtTeDWghe5GtWzlCsT58Z0D1qi4RV+eyesa17Ne+lKmN
FRQKq3CzgYzlncKT8iSM//7Eax0ktrTXDJ5d9JC2Xqy6lpeUbeZTMTr2bLAFS40ywcwM8QPO14ue
/v6sXp6ISeM3Wsd6yM4QQUBSdXtqGO1B8wuwRcSpAV4fL0l7UoFspzb3qZPrwWPL971VQv83aA3j
KylPlIQaZsa9ztdKhHpsM4tQBatOBe80XbOhAlMvuovLoDHNBPTgGf+h03zzODinsY9N+V/38xYU
fJM+EmLLH+T+m4WLRkrMz7KSyZSrQpb6Pt9jY6NSLJjQ7+sqS/IFhrNXvvmTQXxOsxLtB9f1E6H1
21VVB2ziKvXc6BrPwGRB0lGc9/EqQJ5K1qJ8WuGERubHfk0CcH2QdM3YWsnlAj95MaLeYps1kSfk
T0CmAChGHedB60jQVncTXrPafF1ds7V+yqy+BYDkfbLBDGfWI2hGSJA29q0KdVgGlYfAk3V3Moeo
Ct7GJ3re5P2dm9TruuRK6Et+RtqWAQL5CVPfH9fVr/4j5ZE05/uZzjrVY0zq0dEEp4isT6upeAm5
GO+yCHL2hY0vym5rotlnrbG1pUXfCaCaiSduUdq9ZEO7F/i1mRfbnXpRbM2OKYVpEE4LFyW/wol2
ha99oTMvZedIwVv/9Rl7SO3apsjtAZ3K8sN9213yWpFKu83Fvbb5GlN0SBcIxEflJgAEsIFB4CN4
pH9zdnIj9gH3D0IdK1EIzTadjTF+QPmowS+95dc0AJcH5tkAewwF6JYw3B/OVCEoiLvbxIDGj2Z+
FLf5IvELeNKzOZfUt7krUC6E9BIs6Khs9asiWn3v1/yzOSBKrrO3NKihhCvB2FRXWYbePTPkOoP/
CxLMlpLrHk4rohm79ocZsmoZvnU/EEhYcuPVjJNLVQFWya5S+t6ikFL9t7QPClN2bkUUXiwrb6V6
mEPK1rTO/yCqKNbPuWDW4Qqu+9cM421qqg0JmO6aD06V3GJSRJLLgO7rZXCs21MXXWcLGq6XEG+b
GYiIz1aT5BEUpZa0erUskw8/jfKaDY/SFRD/6Znl6fF1q86RamabQHJHkofqHI/PmSgoHNBWX0YO
e3KsDBwSxDfK0NhbP3qPMlQDGbd6eVufv5PAGdmyVhoVnybTX2/X24+ZxXOE+cxyw7FntrMtgWJY
4cZIgXEB70QhdtB08OuIMKXPKk/GHMyYbaZ/XhKUSadfWfUVTDantAEBuu/4+qDImz+J8QGXnmwZ
TR89rDu26PwdufgKFwlVjlisKVzR7ao+IgrZknLAhsCHl/AVkJbF9IUWLasoyxvqTkLm1+lGaLdF
v7dZOgOPMljC1D6GelAmB0fChqP80W/2EhuZaMEi2oyLIeFfRt4KUyiisEIvGxDBD0v6SjrQ/saU
+Ytyxvy8YBz3SjQcJ3f/xUSuvQiOY5qcc7lPsBNylVAJGPtIcFB+2Zo+tr7L9Kowx1W9w3/Vto7a
gHGQu8ls2gpkEDsADFM6K2jeEoUO/c9fSJ858nkyt5kJPYgAsFEt64XLB8EEiF3+XQYzkTVOcgBm
OiA3VZjmpqcj5f5O611cVTAdup096jA5U1VzJtvKpBSLzW4/HkpFH4q9ZH5UlaaKlsqQ9VVpAS93
iuY7B2iO8U4MXoQvKuBmW9XQqLpO2E5uLr0rSUm/ynVy9kQDVLT6oyK5E3skb7VslIcy4k493db+
Ozpuq+OFF9YbyM/RbKUljEyvBreenidGTBDOh63MszGE2hMM9+SViTJDqYJ4ptsHRcFQy9zN9b2v
HzfFnPvRys5SitFbE9mDecM1MMQQEQm5Xixz070dFv0DaqSvrN2VSeMkWHGl9/YPa7NAZ1zS3Wpp
D/RWNRMY00tHDbiJqlktaW6MRo/3nIByY0CfJzAypBjvHogzveMvNhkf8GO3IaQ+31kXWJcg0YzZ
TFDNrBAjQJryS/7EsMpaHdlQ68w/Snaf8ITma4d8GucEF5JNZkYUhB+IMg2mmdrTcFF31NjtDYSy
VbOPqqi/f4KQu4x5u3sZ45d1gE8DDZEMZGz/yoOi9TWTPhAvyYNkULgKXjKZFZNyJi5ijqasK5G4
tZ0ryFYYUVV7kis378os3CSghDIndI7JMvn2Ix1tqYH4b1wFuLyMeu+yuUNLSPZ9lugH5dGp64a8
kzc/Or0785w75dAtINLi2ZNeLjzfS7M0myDVSpamkeJ2mwVBEGOjgOgJ3NqiMdY2uFS+eqldsDyf
EIvfZeVxV+X0EwsEaNAZJ2ooFGM/zZK8up/nzR14bPCBEYe/iwn9TfDo2bRjs5m6Ieg3i0gRGCsp
Qa5RrCZA7NxzThiW3lOir611EkG4se297mkpbM0rI+p46hJpBOAzkTr+zqp74d7vDnM+Wo3tUUr9
BQNcjftZT1cxkZyElcFKMzPdrvnpV5NY896BRfiUYFu8oCTm32hOQPbRPtRsGwLoV3L9cF+untVF
YUC5TV8wA/zfnsEHqr4D+KiSPzE74riWn7DOXTDnnko04+emZcN/oP5LYXOgxbhokhJ2U99gQCr8
rkz6JybylY/vvL6ThhZcpP7957bfQsUTnI2E+lfwv+KVy6YjV2nbIXrWu97LSDJt5pfBObb0Lx2/
756WDdf4sqrlB0Hj34sZ4oQ6S6V7IAhEr6fIstcVGNuZQoKk+Q0yEFBw2XR43mJKizyVGQAjQSwb
7t3iRY0u6xoGanDCrCPYrbnBKiU/NaTamxEa4OC08/UXesLO/ulhZqPBoPK4UC+0J/lZonXI+Yo2
fm6M/ViemScseDs3ymUk1KZVQS3uF8EB5a7RPTIXBa67chj+8KIHKCQmydQHWtVHL4L48kd3rpj3
/jmLZ2Wi77zE9Q5bjA+u+0vOWxN8pBzA1BCGcuVBv+U0yIQW0gVLNjx8A9TZ46Wvr+xhSRjom+1d
Gye1V6L6Iz7Z2CbnLq6K2AQO8sI1u+bv0eYSBgjs6Hgxh/O++YnUZMeUOckiL0ZdTTpa4T8S1jIp
OZCOEHuFyu+nBBOmYawTReIGz31W6Vd3oO/wIo1blAQBZ8F4Zdz2hysF8mZ3Nk4DIfPzAznkDdnK
P2ka3S9ssX54GQfSMcOAzvfmhT/goatQg+DTjqwI843/3wWUnJSzGoTjPg38bH0OidQJfcIbwfwU
jZElFkpxdlO90FxG/xyKBAKpnfE6G6ewXdmh2ikv9wAvXSDa3/UPkJtNLaV95RbYmAxs2cRUkU7c
T/v7GVIOv5xl/v3LFqZE6AprwSvJq7vxn715sA+8PXANlnyrnj16PIGBntfYwVlPYmYEPtFx6qZx
Ob6G3BBGGmwCZ2OlZT1eCMY7c4GnLt/paM+rwJbv04yNBxNYHiQKWTdCFydF0yQpiAue9CmQLoky
d+okzDDvc/wncJI89Gp9NlGlzkMd2SswDQsacwC654ruhL6K7ZP+UUV3KfCa/cvrMzeW44UCW4/X
572BInlF0PsieTuhrRVTj+N5aAHd0AeALn8fArSkZxa6MSGy5nbDMpQsJEeWyen/27yrkNWiunT1
qku/niuer60QCGsr4zSLXlwdxu/0rmK0RgBjqqsiE8OEEzB+ZN88JL+oZAwETAe/SzVIxwOgzKVC
aANTJZtQ/x64BW7lUQkD5ITJuY9O77g++qHKpBOA8P3D7VeWgnP85N/uQCbN1vaQdy0KdRQIfCPE
zB6UJQY5h+eHd5BmWFAXsv125Ttmv0FLhp4UGEUINS/05tXiojOIYJLzPPPAYYjP+TYBG2/LN4GQ
zAVNmSxOEaIuqxZUJ7fxWHQ2uvbH/10tknDZe0UuDCNtOpjxxyoldmzIQC2gP3vK+DcO34ujNNdY
85822K6Yeos8/9i+ioqHF8hDcXKL32vNpTrmzV+jRIcRnCrmgBSaywCJM+8O8ZANRysVBmK5T6vx
/gV4rWHpwhfhbrZb9WgZqoDXoSmowxzG2uy7Bmqm96/HlLWf/ac0Dtz1JMBZel6f0DJJZgbWlREV
yLSrZwJzLoR1GZSHHc5aG6YbFnvKqa8mX+AZjXgJQvob3ab2nq43F3Xbk1fcEkqjsZprS/GP/3Bw
C6xc0kuc1zIh0dfQ/yFZEDPmb3jntL7CqsH2oTMz+bg8O648Vr4mH0d/1uqpBQyO7hYpWR2+AnO7
MTRLe8/gXZ7YwIg1jX7F7EzOsFIXuPWyAkkeh3T1HL5JsdPDmwm/2zZHfbGElt+a0amS7TJuOUWX
hXMEGeRvhXEUYTL+4faV/9olsBPTXnjSl8fQyDREB7z9MAzQJRFAcduObl1leotHbI239lW2wRii
VBDpE8R27+MlH9JZt28Ki3J0xDKMXFEHtQTX3nu6U4Et8znes86SDg6H4O8sSfnGYPn0ZPQHBLDE
i4WklhC8fQVjTcuRFU6sfbHUGsyGDbvN+WbD4YaRmo7So6WnQk3jXjDNqTSgfpHbK0qK3iPbzHwj
PGCVv2YfwmOnZLVFmFUyGgLuCvwHB8lmG2ah5a95C4DNrrpT2K4IdbO5pphTGREchgYo84/DhRvg
I2hkLdRYtVMXsJoJBjf9l79YDFvocGb9SwzvX6gny2y8uodDarw4Bq20BVRfDMv80PiHwrC3xQXg
uRSgip69olPXPn3O6i/OT8OWeBV5dlL8gjH+IO70RQMPxL8UfugahindXbaNqtYyoeACed+v/4+V
KTmOXilVIeakM2jEVkDTA7/WaMC7YMV9ZVN0NRTzjL+/GKV+/I1O9HB7XlQ0g7R3t/Ibog8PLzyo
ZwidW+1z1LEG6fvVzO0YvzFggBUsCZFG44wuc7253rJyNmgf9ww4hrB9dygR/FdjEmTVxTqA8M1Y
adFM+gCXt+RZlBB/8EVPIO8Gh3u9yZSayabVN9qcajSWbpKcKVeYtDvga9+i7PpVoXjbcu896IpR
huIPmiBXFE+boVNOwQZZVDVNaDtye9icAT+Plg1n+RTsx5mNyBY5OthTag3QXT4DVTG2FhpcY1i3
x8FY8sRmNg3dxwGMij18D6cuEGJTyCBb1cUH3roCHkxRIY5KA+gM1gqiUv4+y3/xTZm0jVnyAE9D
o6u6muABFjBAnmncI8AVjhnB4uSNKSTv/ft8pt1Qx3ms6p42NIVLERk3vL/TziNLOlYOeJolmDmx
Fv/VfofpbWDd8WhnlpahcSZFYiGL8rnP4SjUiYOlYOBMv+vHZjcgaty3Q5VTfam1IePIs4a3ogmt
+vjSM6Ksgnzexu1jnm82IO984CnH0dvvqQ+W8F++XEDE5FT9UVcmnloYO5PvYnH1GB4H4VVhsJwe
sBklDncuDokp45ujKaEZrjdZ8FWQOzVxm7jElO9GbCdqkAMIFLTSxFam/uXe5M7FFLLOp8mMBc8V
C2V1WO1kZHVYmEiFE7iaHrXsvd5NmS/XpDoBm1KWAwJFGctzqXAR8pgXjodfYo9TtuxNvZbYqh56
ZQIDIXxGv6F7VWEzoFZlQwK8Bn35ffd7sABRwBuJmRMuQmFU1MjodH/RumHdfc4Tm8MBweeBpIOb
jmVwGbBCpAIt4OL44vL4mHLI0rB7j9Hsz0y+pzNHqEowO4ynJsVV+EHaNMgsoMOIS+oxysDSHaWf
kajUObaqGzWdRxBRjToU/38mw3d/SGWKINrdc2n3D025Y5yGCMYglfudDpFbNVmr5A4zS//ig3oY
/6rGCA+7sHT6tr66ajHZwACwUwmDVDxHO2pyGawGetaRNSwvdRmL1eRxKyyEokmjv5Rhz2tpeeG8
pPf9bdAqaPNaudZuhe6uklsdJMQbUFd50JHVQ3gpq1VLyZ82rK8Xj4yVmcCnGjw3U0DXQgWM9V/Y
kFnGg+v6CC3WDf5OOMx7hRR0zr7/4HoBhd4ZGuJTggn5oI0CevouxkoCay3yv3QRaOyOE9Miv78K
KyE0gGJuJgVjjzF/EGeMGLgNLMXM3H8Vfu8dZ0/9Qf29pdUO6pRXVnbSI0RHch4aW0jSP3+K/l3U
sfzmeIhQw1SmNhbL8ztolLDfjQThgJ+pNg25ZRBUeexcirj1Lzk/WGagT33jX2LEBrlZm6Vct2sD
9NK6U1dHc4AZ2zHqt4oAlkh4+HFlne1j51y1P5AA7LwrV5fR4kQINA7af3x9kxjH5Abb8+57iaCU
41cRJJnXG3ATJv3Xlb5ORRbWoLFhQgVocfOscUdCYpu2I4UtWgj5wwFNdy7pBRWurtBMqsgQDlON
oZuMeyNFaBXgsvITnsUOgr/4e6Q/Z0/94yUInl33OX5AUA/c5MZM0zrO+3VPaAkIg9ZUcTZP6zeD
dDa01vi25djKkuVDzPKbJyQpwhIJXgAS2dtDOywayOoVld3ALG+Ht8uSfrz0bUzNw0OhDdgjLwgz
6yY2bYpIuV0FJW75Gq1EZBb0X5kxEHgvZkDMzHh4sYoj91ITq1dt3EY62QY01mpVHwlrJKULKfCE
MQcQuftc+ba8yWlSDb7kKuo8B0zoPmV2Gc8H85qrh+B04+cbHyYNPxiTS/jrdgM4qvwLiFLUQqX/
McSC8Kfkri2/yINZu2YiLk49Q0+1qQY6OQOen4u3SSLLjDzjl2jkn8MSaUorEJ6g/+WQTdwQ0jjK
YHf9XrZx+jUEbOso3nkPVeLPS+nx2JW/Mup2KS57F1cjEj3EWSkhqgkC04zCk46pLIWxzHXMNZyz
yMCEGR7mszo2/M0mApoOXBvVlqGObGaacBytRNmALS8daaKKzeCHnIKLhyB36zALd67YZWCN9Yrr
Ddq8J+Jjlx7l08f7doofRWyG7bTfSQeLjHWsrJdjwO0t2wlT5iS33Rk6qumWvwtuPQHh2Cb6ABnk
Z3XwOUypWSwLZu8NKbTLbXD4kPeSE2aPK4jP/jnhmqbKF8uXFbX8o33ZDvFRUICOEQr0I8owa3we
9IHC2h7tmkT08FJvaJayBPaISwL4LkZEOYINbmduU6qlApRLJ0izUfoyPgwYAkddYgRnUts1Hark
0O38TuNunD6OLkSJFj6dj66FZEe/QNVhFYuzp7cXi26RInnTZK85WvIL/yaGU+6AscLkuMr5OCgG
KV+EBw/5fJPmRvJvN8DFbMOQUltE/bYfK5mjLfUS5HduYTYEoQzvZoKktiUcnVhOsRkK/SnqVCE0
Si44WDyWXzWqcMXm7DVCoqD7h1CNU+6sTcm9a0QlrtSZdroUUlJiyoXQ5ggHz9CLTVSOU+5L8PNV
YznfnMr0jGRYX2xm9wrDzld4jIJPfh44oZRpseDtHm+pcLtjeKied+F1ny00HABqqvgagT9Qnm28
y6nokzLqR53APRnb06DFBDHnwVAHlGZSQBbtkFaJhXEaNdgV5ZqkZV64eyCvuxyaARjvPWpuKoBG
OUw4EFI19QcdOV+1ENEshM3CUfbt7y0s5MLXBMjo5wM82mgx1vQI5yWochpY00MZt4cy7+SZ50G4
Clr8pP80+3XCvlMbgeeN1LKBjnaDGhLED9NNXo2oSOASwzcstQOmFdCg02u+lIfytghBUrHrFrEB
PGKg0ApKzqLh8UK/c3BxZZpbuyq257aL2lBIaqgc05zJ3ELt9fLIhlqpZZPjM/O8NE9fSDrkf0ms
G7ahVLeAdK//rAZ2ACAyRF012UlxHp1fTsjLezqAqR4vVDaFjXmnf9HH9RqFt+YEyYPa6KL5zqJZ
EyhbkUPcdEZBerjRAiAv4mQHkApphqIm7JlbopO2Q/CRXpz+FjnkWGx2tDR6adtL9wGg81P/wPTL
QuRLbZNb6ayRjfZ+b3baAHk8bGWey7bSB/QsuBeSpdhpTHm/EhdzRcKuJWXMEw2vNmr6TOqe+PJk
NHOo8fczUvckOckmWoglixMdkPHFr9W8dNYoNpOD4lxRBg0gmvPcXAvGebyBYWD+U49gKFa0/cCm
XtnBQctYB9YUvk/BP0vftphv1UB+wLO2dVopN4HjKFWdIKygsiCdfTxmOUHUbtIboEOtsD+DcuAR
fQ0ymuCsaLDIqNe5RyUGUEX6LAdlUqDCTkegDZk/FnqleAKL1FBJ6+QtyJBVQ0aJGAWNxQQ93urA
1dLMgaeW5lOY5/C9HuNDSWUC1V/ggqNfLYz3tgEZ1w0P2PsYrK29/5Cy5AP5eIJWLnZHgWEulcfH
S1HYgd/Yj3TXWzBoFTCh30BqpiCFZ915+1D0L03ahXK09h/PFxIG8Lh+aY/DFF2UvqarW3GVVOOV
t00Ukjq465+5DOqINFFysJzvYByCy0M0ffAhcEKb26HifEiFk0WhyKKzB3bwKZjPhKLndReyb7rs
iI9Hq30x9z9hVzf0Ln7iw3QWmYtXFYoalDb8oVqJ81P8RqY0WDU1UYf549K9Be+VpPe7owterR16
QQ20kKuHAOeowenX+96a9ykOEvoF040oenQBSC2S9E8jvj41jSrNXhK1cAQKdVkuPenbFWMm/Cwk
uidiOua32CjUjmTBwoTVWy8i6kAgKE1DwWqEKt/qtukLjDrinhThJek4eCH+dVl1wvd1NLg2qoFL
yjtRZyINVIcTahygU+OI+8NOTO+Dhy4f9u4s7Y6SVGnnwaEb/sGVSxJ5BiAaKdjwiIvmfll7H8JV
MJ/3eIAdU0vprZJlG5lG/IdZFZ1k636Lra5tUCd9i9hlOusW9V/F35M23KntUyljSGyCcSRQ/JNj
0WJtaLB5LvzGqzGoN9zsvNl96lqRcuCNrI4H5UZC5jn7lUgKrfZcVppmbtA+jdBdgpSb2eQkv5GZ
CVrlfPm1R7lEfIvwafmDMsRatMCRSrCTOLtKeYVhlmMiUWyNKgV53Dy+hN7BSy2N7yurZOswehUA
QRLEElTGE6csEd6HN/nUoManBvBrWD9QZnWss29Ls/I8Y27SIpqDhIeLauygxE1fgoXrkb/44Cwd
gzecEIOfbxMzB2xgjUEmuLMV3P0nBgPAlnsRPHSCcpYO8eUf3+CqLGQokmPneXLQZEw82NstTkpf
4KXB9v7O2PMTLcggShJGPK4DU2mxuAAOzpx7X0fgEcS40xsT8V6GIIR8EPn4BOSCEUALgyTtGKDc
viuxWNKBaxOKeeylKfFdtYBopnz5Or1eWlRRgG0HGiywvoqY+yOVWj/hbRfzYbhe2XUC2nP21i/3
1aVQE3yYfYmod3e5eRaRtz6l0wuALU6pmB6etB5LzBe5madsAwZehbuvtL3GRMoP2K4mXz+ddut7
laW2rFer5nECkzSjMBeRDIX7CxwLbi8T2Pn+PIQ2iGHjF1U5JSi/jgTNDAog+drKVi6AOxRAg287
BxaYCG7D/Pg6N06WZLdMt5rWYcsmVeiuG80Z7uaF1FvY/nkplwCFM8HhgchnsQ/h6paTUORa7ywB
j0XQl9PtaRVpmwwgFmrcapaCwpCD2R5uikaTJrwAPWue7DjQ9hIBlTNjFNdW2tNEkZN64g1Q6QK9
xPTtp+jCgKtTCsim90Z8It67RTxQkfTG4OLfLip7R2yZkMW8Txq0BlcFBo5VZxVlFXNZF/Hy5vJM
RArlLb/Uvbb3HuWpTHjL/r9mT/6Tyzc0VHuVJez6UBdz9D2ntVRrEFsuElL8RKverUyfWldoeCWR
5Zj6QVNZiHI7nnS+iKzcNaOGBtCjHL/OIiaffXffNJd2GY1uFVDmNvcfiMmonfbFeztnn+XY5HOQ
s8sNaLBR3s5ZcpL/htyY4ih1Ixn7FhAc6P2x13ayBY+W+iDv8BZ2MYfExOU5EgF607AuLScBIwSq
wgKKClBU+8wIt+bBtIhXFQgcd5Zc82d6ktYVazGOw+OOblkQdhAGCtLN7eMFQNqd77qkKqYrbQLW
08MceaNUmopZZY7iXCJUQeDUY9ZLpoS1NRFF4668GTQAvEHbB6+yXPgn6xp4k/yj029fxe4nPjAI
TQWs+cyX8orJhQqItBONPBUyLF6v2JI88R13ge50q9Zoy8TGlfjtMLJA+fXSO5YsRJI55X6vPGTJ
MsyFleXjHBo/JorP2MPoKzlqtoud3k/4yG6xjqI3kkKIqm7BjeFUlEvFt93ErNp+O/rkt7aJ3h/A
woU0v733ityyWWsN3MeJof19xFIrvy/n1WvebnKsTReOWn77VCTvXV9WPUOPKMiNqy5nRpve4dnP
rJjUYaKzSCWB0wYp9qMRnb+cZ9l5tXClVXLA4aJNN9RcsGiwpjPTuqMlNL3Uvj4DFJC4/vLGjPii
lqwA28k8UetJhVLXMJpL87wlJuekaJgkKi8Wbxtod/fgo71zVrKzhcHU4uatv4c+OlleQ6da9Vtn
Tkbgc4LTfL/o+T2DYKhofykCIx1T/NjKuX4aSI2yLIrXNlp/Gmm/jzitpaISdh53c5rIiSXjT0O7
/LtGQ4dCPiynXphHsFA8J0AaneaRYFdm3iCpjw/DRezYrVzRoFES8JomqIm5xLv03clIolpbSt7M
O/M2VMKefo19FFXdufyqvOtc+Szy/fvqGpGo22yIn2LhPJFcXAEkoCgYYtEIzlTz5IeOA56HmF9x
0gA9DF2fdBgmvvAA9cVFXkCjvyxtGaJ6rIgBq0+8G7fZ7lUXQnbgznUri4lQRobE/WRsI538rD/C
cDOrSQQSI5EEOHcMADW0lPn3Nxj9jWrqjolb1HzLtIh6KF5A8FxBja2ZCL7ffAiie9ueLn/udfmd
dlFekYZKBq3ZJ2dXCFczwCYiEHyzL4J5xdGvqNot9Wtuhm+vzV5GppPuVk6zo52TgNm32NUXuN1f
XhI4ESzpIimj9nY17xf8mzc8rSdLkKClrKfxgCr3lagPsjaDNmf7wvqurbJdAE8P0HgvVL6BJ8/c
Tk2Kn1op8UvFF4ntDI0wmuz/1qYKRa3TGVUo8OvfK0cv3miJ1haVfvEQNpSvO3rM4UhoxlCV0U18
BqhTvnJAm5oQhfyv0ODeYWj8BWolvO5yoHD8IYc50NsUGVUSewIXoTucmEz3TuE8Bj+kCfOL6QgH
t4wgQKOXLckWxdfef6BIolw++5rU2VVM7l7JpHOIiQsplxQS6Pn+kznpglP0xO7fXT7Q3dF2mBDQ
BTtM6TgsRKvxu8BeCuqxo4dO6wdSbVaBeOwEOXkshyo/0JeXCoRY6+bcasO4lTnVhsPLwUwmNDUg
/Z3wkaBS53FyMkuW1Gnbp19Q2CmvQGVeR9zb8fw9sf8ryMxCcscSKIDvicBra9WpuFJVZ6qZZ0bf
XHl5bZ8sxlSemJNAPMKHWz6KQPh77CSB4Mkq8WHPcCJ6of93Uo+gF1g7Eh97AqWx6Qzb6UmKeLpw
bDlOuqIlpxD9N6DmqinxRS1bC7+l5BHf+/ZRzRQLbDQRIoF5Pflt5Jg0iSG8xDH8phYn9kOJtcVX
sMvFGvuSnJmcIBOnvspaPWdy9DcrpRFeAR4xz9iuwbpjd7+wIhq91RznSAWQwPYD/ABYfC9aPyTY
4B1WbA5dEipU3lZGpApgDHXeIu1HXSz/igGP9Ot6Rcnnzm/1epSFR9sqVGSy+VmwX9/e86Y+UVZd
f2a58Zzh9yygLXnGCRHNlEcufsNy0SgC8yEf7K0nVN1bzU+z0g2IFx9ifGvzkNUoANmkziawEU8x
c88B/ddPqDQD+9fiOXMf1p67UmvxHc93HFK/MEWJUcSmltHMllTozyqJEJ+AhI1b0RTPWeTxOOQ6
VkKZApRFUGepOzPFhWEkxhOLZ5/zs8OgXFcIbtcttg4g7OlzAW4rnygzlwKVimXaVdIiVf07d+40
RGcM368VxXce4dUfgDDmadBRl95bZhB4Q8p3PEKptJCAAwdf/Df+qJBLqR94pdI5Ax5u8tL9lYyO
kg4BZviYB5fPmIpFKOcClaYyeDMIz0RzJqXTnMcaU5FqGwpiALYeez/lbRVpWdVeEwgDDcsTLJm2
F9+3F0zgAtqNbfpp9rRKG2OhCZtcmwzsc5lYXvlGq00FiIbSWfy9FLM0TWwdiOHRfP8CK1Ghviv5
zhUJKPe7/UoWL7jrPuqX1Emvaug2k+jgTOhkV+GXscSWk9LbyOwrH7VJbrkHN8zoMhFcxoJ8rO40
kWydMnVfJyoGPmplrpZnV03g20Q/u6/rSLoThb9S+JuDH/rc5IoPREAEmvdwSyR5V2pVX+zjFYWm
JBPcsLrE0zk3YtR81wiPdnWEVBlXTo7wwj5vQw0P3cfB2rCyxOu1W9uGE7/auJH8KdpfatKqHiQj
nXVpCoJiQz3ja3oKOMoon6PehvW4qBEh6W8L+X5kDto/u00p57EgX2T0L0B71qPFRGhqow4oG3I5
nCRc+UmObc4clgSfE7u5JlQ2dI9RFaRvgTBUAjVu4YX42sHDEUzNqoj0dDsxgu3ubeeXW54vK7eV
rptd1Gqreozo/XMoTQrmLQKQDFgCnsm4juUMPdxoNh+ilAdu6d9ZEoNupcINqFfNJu/QWsZNSA5A
rP1hietIr28s5IsZxgE0WB8kpjLsqXzvlILciEIwNtvu/jr1Gr4+vSbwkXv8/Bd9o/Jwa9Vd2kjy
NrbNbbdxKTIm5gUoQivwoxZtdEEE/L4+HqDfkn/UA1X1G7Hrdf+navo+no0Hh279eyxtp/zSUbtB
CmEOmCVvA+kzHJs5cFCYJjvvmyYKbJuEtGiXa/KWNEQBgPQNnC4XWe4b2VojJ7/+Y0L0o5eLTmK4
cCkhcKScK5wwd55egwC3E8v6vuyU+NDV/w1GpG3qtPmSnNc341S83dROfsxU0z1e53bLf1tp9KJ1
17WVu5U17h8c01J+V0BwEP9/ywsS1JyaSuYzxmIf1eWpszHLOg0miGeQk1bQJtCfzwc/5APPJ2i5
WWfDKPML9fbUG9a/4pMACaBrnTLN7Ojm8O2Gl1bdLbSKhWbqKjuAcBccXsMJwmF18VWIkMd2TAJU
DLpcqfBPuxEImuYfx0MolWEJC4/PQOKPhPjnzyXVsPdyDn3PsLvY9BWxlUza92ihXBNsGWYuaxRm
IFPMpy0BKKwo9+UptBn+7v2oWW0dP0Dv82220+YLPSf3XOJOYabB23kwY/0qIjClQmhy0R29FSh2
3zLmlvAA8j7/Mi6HXAFw30zTe5lLdg5245KEuzgHMka691v0PKN8KUw5yv1Qon6hy+0NelBzYVWT
n+4+x1zaWNuzysyzTEG+krZJLyY/3FJDyYv+jkj6cOMEEmywuHbbJdkmte+5jlSX3Cfk3x7DRAw9
9MZk74GOHsaxcAOlQfrL6MK01sMT/UGySKoZ64E/aS0rRMaANliJenceAdRArdFVK8H4EKWoe98a
MQy2iJtoZ0Et1A8p4dbeJZi5NaggmQR0sBsM1F1AbH2IGeuYudJIm2jfRqePJnnzks/UyvJFN1vl
aTJYFNPbbwTbmpYYogK/EDloHUzAN77WDmPgPXfntvOw+Yti/Q7nI88HF10uCcmfvuBnXt0ItAJb
SypBCntJR9GyR7K3Z8IG4EnphEBgS13KMQyrI0MCKeyW/mX8OiFaiD5uT+0UrAoxKO89YtHGwqSc
xCJscCZ/VDhbz4tCaL4YDgYql4tuuFAMlhhsCi+NIwou5eBkGhbZng/HtduPVJ8Vd+xNdCCrdNl2
6PfCItEfHrW5wBCUx0xzQ0u4K7A7FbUMHI/or2VDJircGgmYYeq/KvHeEVNmoP+aKTAd63inwE3g
jCrZIPGsNjBatzQwnapDVNUQSsbn/87JiONaNo+kK2yBbjhWaB/iJ188fRyOeQlj7SocA6r+lGiS
TpvIsSSQu4U5XiXhdH10WuJ3n5KqLPxNFBOcqtA1ASbZ92rG+TzH0GzDn6Ckc4f2EzMu0byPWJ4R
iUVnTYpuOUnurYjEU2+QCOi0Nu2iZftXflYfJEU19cL3zZ8Sc3+6FKX2KMZ0hdZCE1ulYfwVdZ9A
FECP1l/xim1YSYad/zkUAXMqqcSQw3Qz4UDc7lDEyGAY6F3VxDxXk1Eref+2lXeIX9E3X1pUlhjR
2i5g8kgtNg/VzrpDO3HzeVQvghk/zOEZ9pVBUD8HLpvGWL7VmiVaVBFIFTYQOTbfCvQshtNK1iRj
CJPryBKN7u9p+1mc0RBntJusxa0N/XT5FPs87ITjPJfpE2YRVqfvBwEdDTbGxDTw1Q+H3mUQTnRL
nQ/ZpoM6gAkCLHNxgDiD21EZeTrjediL5WWtFRI8SRc0DrBmMB0niYc3rOgpIpjKzyFgeovo37R7
bp0FhIhlxzun/9SeKzXMobOqdPPizyUWCbFfeCnzVgtwga36PkWxdTSMh9cWfsa04Ab7kul4T4p+
555h7xo3w8KW/rOQeIpFrkjzKCwV8jyKncFFKmU4rPFmMwWds1WL6gbJghAyvlbwc3Vp4pChghI+
FxWOteGvipzqaKjszi++y5yxPNTCi1RQQ6+lO6s5EAqNpvNuTvgk7/YT3zy/795oyNuCoVeMfNPM
5d2nzeXj6WQM858LoMGmLLBthpzQPRFCAit6VSdmnXdXLebJ4uRo5csR0zXbpVjz1yJ2bsTb3v8p
WgiMeNLW7syiYDE3xWZS37x9SfR6HBO1uNspepM+GlFLnXCBA9wmbdIRuPFUI8iavrHahTBhbDdP
yGgnuK7mDc9cUgCixqyZv+AMvFnRgpZEOb7Wutu1C5j9v6GruDJhWaj2Ayvxa34/0xek66YN4wO7
msJKnWFMPEneImdh1Cr7+wfpeFCrHfXz1tQivFt0a9wQXKRdBkQl8fHEqbDq5ki/E5S4LjX/2+nX
m9jayyxgeDpQRFEJND4GgEtMq0LmH8Kadi0WJj7SQccobq5VoDu9bSZ3PXE337N52b3MQDENtebK
/GIDj1VKCK/yisBnfTAwLT/1l1ARcTXar2myBkoC1cb8lyB/hd9CMjgHtQDL9d4qCDi3ERAphr/Z
3Rl/baYmUUd7KEzkHC8dnyds3/u5u0CTHvrtgorKEfPrZFq83VlzWRTe4rd71ydEUsC8QLmFqden
HD7QuQNB29vnKIrBv52cxTl7HWgT/Fc+NEG6hVqTY/m5I4PORDdG8NnpqjJmVndznWVdMeVOiWxq
AtPsuWPrPT6f+EeFzzQoQ4PBSaWhZjysm7p9vSFaqOslUGIxMrIXBq0ijlnQQIW1wovCHYGE30HK
oL2LIwr5I46XCuN1i4w/xwAnD6cpStqe1EwpJ+bl+V2Cp/fV6DD6ai8SF4AWQgZItRpy/No0ovGD
duiwLNjDmAiDty7zBB5B9Kci5gs4k9NjDNAjBJf5g35qxFNn1918TbjdLmMazXwEmAVtiX5Uv/n/
1kUAIxZi86SBdTXI+xdJS5fEaSJQxanNm9KrXmHH3IrTIBNKVK3ceKJeXGkMQIYQxqqKl5iZLZyv
JUCUdu3y9mob6359HKOdCweASEDXfctDxlx2aeRnucdvwP7KyCZrmDsC+Beyt0gdooerynfFms8A
bN7qdSkqUYfvnICyWFnEF//51uPeYtPsZl4jMSf9J2Sk4lH6QuCAYvup8AqB9vC3iD0IOw+tZGvw
RvE4afxZIyBgyiHj/Tmo6hYPASlywx28ew72Dnu+RxoiZEEMLCGh3KIdZt1OkLpw52ziEaGhlT0n
pJux6uGSrtdkHYnks61moiLOLF5ydGyhayGTFuaPJ5ZJe0c1azTkSJYIjehlKuRflL74aR8QcTHQ
1T/hJVh1rc5b3ypQnKRAsc5dylYO4wucTkavqAHq1FQPtuvOijohQexonU2p7vHCYsIsCmwuAsnq
uAlv1MiI8f778BC/XOs+sLIcHVX4srvP51JzcOsni0B7t8oLh3UFRBUxOLTiZrCoWWBTXXHNGQYX
6Hnkv9HLKCtpAZqZA5Evc+awXfpq7De1QK4lXmtsUBf7gjuq8bLD9zQNqu5WQ1YWkQHD3gKGv4Ue
kcbpyMtDxUbfp7Q8UKV1LBEOcYmv+VmLqdewSE1DOu756tG27EoQeuO1/XU14RAeSgc+4ChDgqVl
iBQWMltTNKbQtIdrPdeKxvSlYyfwKHwLNrJYEa/TL6UgDPCnaV95z6CtvvRwOSludey4vJZuBRX8
0faWJ7AwzAck1L50xDiJLB4ZTKJDw74LpGkDKM8VqG315Gktc8S+A/opldY9JdG4D62TarHeo7yI
QHZp8tgnbLJ56livMhVRm4OF1TTj9+hu5aHwSxcX6EWo794ievedSUfFvJHFhOGi9r9iNOymBFxB
2sUrWmlOjB1wpwtpWu80kBJegBR9rheg4D4fJWqKrHsTrwhJj9PW3i0BHiRjdH4N227GTun5pT6L
FXMUy+FamdV9pinhdba3LbnA8VjIda0ul2lUJW2G/6bhS5LDBxLJZTYY6wtPJv9ZBCqOkasFEHJw
qaf52slud8yHgO5SkaJKKDDqR0zOIynuc7dTNm0hIQpJxOavoiVGzqzv64oAsyFqNWJ18hqo4KO/
II+EsYaDp4qtJIGYZORj6DgRJg9COGk9TGEw64VlFntcj0mtYMUrxRxRahVPsSwNSrXOrRa/WNZm
5yvdn1w9rwt+0bxMB2Ur7K6drVhUAo2iNFYyet3BAzD2qTbKM4pfr3EKkdAFluNHFa+wtAvMLCJ3
dcvAqCDVuy1roNSoINSOG7VXPi4XLi59kdNCiAydoF2NxJWWhoU8dXe0tXTAJIsHieJtqORxkW2O
6rZbO1ZCn2lHt8BWPbAX/ufmtYr91lSTHx44IkNdq4anON/X8QOv8vjc5xL497suZsA7acqYBXZo
0HRtFp0tSzZGHaxqXtgcaDQQujby4cawPq/pGdwp6RI4xzjcbl58+oBSksfuxk+xstHDGySZW4T9
+5p1yWRDZrF4wtyAiZVJUQCQktI4lVDKuiVtNWdetq7MCaYSGXJR9A67I5oVINFQ2mbapcku/T0E
48/ehnF0AUNrnEQVaEBrp713IVNtO8IkPODOa8gaitmsRn1zaZVsB6srVvl57nv+WD4YPteBmOpv
CZX1JnpgGhjQ2jxs492w0K51CbpE/f9Q6dS8DHz9qxXL1pYg7KUx4MXdrE6DtQwKo5fmqfh1soin
AButclOR94/pyjAIzyHRcAgrZSyXJVp7syz6Wy2vo/HP7vz4YAAm+TtamQlMTWISN2gGtdK3zh5Q
9PXQ0ioQ55LjWEUJtL3P5n9ynrg2BrzqFats7tdxwqo3/1+b/AfEp9H0nT2njJatpXzO2Sllq3+O
CXTe0zORZP/FzsH9WHBBx6BtW8Duh8cxbI/kFsTlbzTlFLTDeWalnY7p/53PvDGwV7MclgopXHcr
PD+7kxHaiDlmQ+SbIgN8Gwa6crN9XWgKyMbNuYBQx2/hICusPg+1fp2t/mEppNp0KhhnZrUOtiCO
fiCoS/vnKdXR3r3eMvkTB3AMYyfxc54BBbxxYLB3fMkUMaqI67i+HGqJxDp/7nPEz8tur4zxXs3M
q7cS0vCOpwCHAgXnRDkbQFbmVp65iAD0qaw2L20lBIwupL5fTPdkv3HpdNGOsoCdMgGEvcM1/zq5
W+Em4dXeYTubRXEiHJuXmz19sn6D838jX/kI9rGSpZrHcKNVF/3ROSC5Q8+IN8bqbTTTasD5rc1W
M5aFaMC3MWTX4ZduqfxLity47b3lgxFbb8zAlyvlZp98DR3TTqhabhF/Sh9wcfnApfQ/F738FVQ8
IiV6oKqqgsT1Y5cWIZNBaS91mT3yBD86N4isnK8geXW14QdyqrAih9d00+jF2LKzr1PM2GTxGuBg
1CDo4rLhzMtgJKIrrF+U2enwynzMemDdNhG8CJi5PgHNefyRhQZa3ZNbW3HkeZZtqmZskkfOyLvx
LiDVv2/5t0RlE92NpF6DxZ8EkVAUlx25yVSZw7jTI8T9++TqdBtAL8JOQ6qBETfKS2FrxIhibf0B
maOtQOAJ4YIRz7UWliHbDCDn2LnAMG8jOG+DWKox7lhKmQTBUnvOMbT9xOov4p9ncJZWT7MKdcQi
0xzTjaEZQp2TFheN39sBdOwRa0DiVGtXMh0YDcTWsSAz9uQ67cKHUy69FmCbWmBzC4HAEL8bdbxR
gn8FZrmwpUCzH1dW103tgJQ1vxi60N/fhIqFLFQRohXqSqp0KuF9qhEiHPJLWVmsW/yulVRYbVC5
HRsxAObEh3b6NURVG/QpuzxUNhuvPmfLLzct8CULyrxM4ZRyChs89gs92VarbV+nHKjgnPcVtK/u
wJ4OD7FApOnRZlfKwn8enIZnymfqttXuWDcXonI98gxFY1E5EW/kbfRaOjLfdjwwmmauiSsgBOj5
o/GzF/T/9/iT/oArhoSNHQebXkLpxBexfAd+ox44t8snv2BVL+Y8IxuGhfBQsbnf9iLMMD2Mu0Xx
BCqJIaD7qWx8Sbfk+bdaLVMKjnqihM73N0im6vX5WxkqniXyQ6GgDTsE/gruLVoFENmIx0f+oM8t
BX2EiJQgsepEG7oGksLH5lHRNpt1/MhAyWsvPmjDN4VJv+pK8ZsWjhkpGjWH32AGcIUP+hJhiywE
ZNvy8wwpa6FiJewjCd71DdXVRN/7kSuKk07GIZO7c8HzAJ+6AR3VJuTJF7ZbBozumdtOFt61q/hV
NCR7MBdKnQsjzwbCA1ANRuZ6Z4VdQyrXQKfQsZip6/v4kV6kJpxD/q84sKcWuwIVZnJtcdciKyxu
u8p5Pf3cpg8Wu5870i2KEOc/S8ZLJH0m3Y1YqkEwGiv1R5/vZNvPRwHGfgwqmVgI0qxS9Bp+fFvC
GOPIfJh7dhieFsJs0J6HEOXpI2G58UIBeLqHG+WMZ0+Wlglav+Vx9LBpjkOPlzEfF1oGrh1Wll5j
H472ISaXDU4S/c3c3kyQ/QLo2iH2A8GSpU7cnywwdnmoGCcmxgc1sctXvOCRkSE57m25Jz+6Ym2I
K9lXuSqm7cstdvaPs8fu9ZYolzLu7eP6WlpkyGJpbjlkbmUlB9mYWhSfWkI+vJBQSmMkGLrlzSn6
Ed+SF9KmCAKw16806RmmoN0FqWc8ZnL2JITZ0v/vriCndI7ElG1DPj5qlPv9HjkyjfZVZq1reOGA
IIPHHXULk+fCVQF5qzSqt3aYtx5SG4ksDQTjp8zFdMxXvc2E5hgLk07h6yeI8QXIvKTXoi3Fa7GV
M15O3J3LvJ1IiAceWHR/L7o/qKBtROn63s+EZCAYKL+FzUPIfsnbR6lN4qc6VQfysQv/B3pJoQi9
atj9ZsaPnSyIFQWQHw68Koo6KaMhCatxwec1Oew5WfwVC7mVt/+XZ46TRYQ1Hg02ZPXl1iAFrpAd
whf4DhtRy/sjIjzKaZoV2+eJ/OHlAZg2nv1vE5sN0PrJJz3xHh87foYJsHifsinnO0MhvWoivUKn
4xM9OS/fEeSb436dig8hKPSzkCRIEjzu+50oibO7ttVu28Iv1fcgcJ1kzrotmXgLpJAHg0Ezhrty
OYVtybSKQlhExEOdNqwqiE/FQRV+6pl9PMdRVxffJ7YtIRFTH1ttOXnetmzPl4wnvwXjVcneNFv4
p1OpR92cX4tTNMAxfOs/i5PUZ61I7JV4Y+G45pxMC7VIpZib9oqbV/AZaNIrZhBPndBtXfOs48hN
FC5AFZuEJzxF2akLTSqcqcIwxD5hiiWvH9ZD94FCDCkBLdvluR9j/9CUfImygZupFyG57EXIl/lR
ND0IWZ/hrVVA49PfdhmEKO40AerLxjH0e0GEQ0Y67FLEdus/9I9MLpHuxdv3JZt8SI/xQPIrpYAA
0y0LlgpUV3MHhzKbUnDh++4pCrBRiJAFC9GOh79uDUD/86Ka7QoNhta/sfHCLbDUCxtKuCK9NYKP
RGjTzFfpfidxkXRZy1ttjssqzylO39E+BoDd+YSuSaFY3UJ5ec6O3BJfXwX99TEheXSzkR9RCysJ
ReDYgiwCkW6rf4ijxLNjqJm8GYIGjSjai6L6vqrxa9LO33JlTqpjCLYiEUuQwK2Xb6YNZBlaq6I9
oN/n/QOcTbrc/iAmySva8OnA3k1zMskhMVGR36S101X2MiLYs4eE657sX6sOQXpz1kKCAmJYeK5i
6z/u5Ycb02D7isdfKu5BfY9bw7Q3pv71cdOoz1fbvRBlgWED99oruVu39MKwY5tUSzEifV4o4ygM
9+ef99CB7OjV1+feRW3ewVDyTyYodUwJ+Nwggt+56pD6SpLNiNOLEAyjCF+U0fltBE6O3b2XgjAm
VAfELHycysASfP9TONatMX6IIwD0IjRywxw3/kcKw9tFF449UFZCczEGuuplXIXh/Og/WEK+K3ru
bbgdVH4xyM9vtrItO5DANfQL/q6893/j61FToInDsmhbAPKtKvwRvH3kwkiJBJwB4d/1BNq7uP/7
VavtI42JknGXTanV8U4sKi/5nbFgp2XwDhntyQL9uqEHP30o5tdEu5Wu+04zwBweMW0D+IQALhR2
cudOvuSfZs/wE1bdDjLRkb3hJio8qQaVwlLMKYp7CIw545UBtlbEiqhVOg2mk+zYQrlkELMM8q0L
82A1cTZO5FlYR+8wODc5LbDh3fIqk1N80RPYQYtMBAGtySLw9bEclObQnbOLi1CdEAdxeDH93Top
v1xnvSgBnN/o+c2v/aoYzMjOnaWJSyo5BiTEio9mIQ5ylNxmKy4FUtCP484CZv/gFBxKKFrnHff7
TC+ZtjHdWmGgw+sPyDko920D3x2qH+hFjVK3ZkMejP26ByksIMCzhtjkwgRwypz14R+Bc8Vf404h
64Sb4l7kmWKDSaEmKYVWVe9jnytWbYyqDlJNiG5uRXB4BDHxRE57J6L8vHbih9lpWttLUpZ/PST1
mzjCdnFqMUMK9/qwZqZJRzyeotcrrhzeHGKBnFEkmA3qapi+u6GhOEAtaiT0gzEnhmR6WQxblZN9
Jk5QJ8RfWSdR+pRIxShEdWwGDTRdtTlpcosCBlZEF2ZvIye0qdnhzsKUgPqyASevDqpeKjVoiC5P
uB//W8qcTmTfAd6PqWlwtCNqyDn427cMehdoU/FvGPwS6f5VE3RKpkww5dCjUghzbKdOJ/WBeFtW
RFrtCshepPN3P3+d8nD1zGBr/mybPl33+w1WC8WdtcVvjyMYsxGus3AgN0Ta4OaSSfV8EOwsTIn1
i5r9HyiCrIDE1R53WkiSYRHe810ixGkKwRJq5hD9WUf0IBCz0u1imQrQ4K2P8eV1LUKMOUCjsRi1
VDdSVsHuEf1sm4YRSEVDcD+Jx97Zz+XzZdElTcjC4rZ1uB0/OWAJFU+VA8mP7f6ZGO4T3g2+5N2G
xAQxm+zVEgzDeB5sShhd+IFwNHFala7Ic31DfrtBy7RNlX9tMpQClbz0dncEQDc7OVsmIv/Q/kbg
zorTsRxTc1dJs9e4C56mAQ+vbXFNHEg786RU5zibvMJtzFPXtdV05JV5/8dHXK2luBnC2lJnQbXR
shjx15U9FR8+LIZi37vXrgpn7zqC4DkAXRvjmvOYS6JCru+1kB0m4UkmiwCZQh4tHqu6QWGF4KS6
Zs6c1E1VwijuShuPrDMnLw0m++4iFtPJkj/gJEX6hiVSLXEJjba/j+KG6cOzqFqMGRSXssJVW/dk
kyu9WJLxnRCk6hRcgXIxOYW1QO6JGv9rnyvbG2LcOv3uC2rVLwAqDz9G1l2BJO3c0BMOT6MIj/eB
P1GodGLW/u4c76s6Zgo8xLMCiT5isK5KJBEzuOVk3gUE2RPLxshl8QmeKkq0OUDu/aYbY/fvfQSw
IrVPmIw51XLgO2y6Mx8912PBkbPyGJMYSIqxhgVaaaro2/vGvTLkIV+Z9tg6/WUxcHhj2oVfJeXx
tbmDiBN12K8GP7mUT6U4+ChFKlenWBNf4by/D+bzK17WEFuv0BioRj0bPqk5DmmEXtVKK6DDLwdb
seL2QgL0+iU79wqyP6dVJQS4k2i1VYo8XjFH26zR+s4gYOrpEAOu1AM/PNmwn9OjxTus3RwSvPgA
ktVF+Qj6j8fTy4RCcQCq2Vn3p7RS5pTVam6egWZ8DiNKAaUfvyplkH9sEGK1nKTJYx1WeyUvKQgw
lVhLWjuMVQ9YVmMY4lX7f9sN+JksGRediSQ9Md5BthQL7GPv6OP2TDszndum6J84iTcR5pxA1/pg
TZlfvWxVlv2o3ojkONZxVI0/USpelZz4gBYYlL7BlZ0UgO12ElhyL80kVgvYsqTCSvPoEXWFfUuX
9plmCb6BqpgqSBBWB9tt2NDP55ZLvYNyaBpK/P8taubOnl6IoiPMYbbG3qY/lf83gnQVkwEqlJc5
YqlKXuYtjopKMIC1+GcnIS4tVNWQ6GVf2xWPOM7qgtQzUgBJjQPNGogt2E3p32Ws0QZHIVvsXHHz
VRogMUL0qo3lIBrcdM0ll5gLqKDPGXs/HOrSbLku+2ZalDYQTKUDNVLbYWIhwFNA2+euHObCP9Kr
msfGQfZnHr0E8p9lgfgTWVe9JO+iHOQsxIve1sb7ZZfJkH/uGRqbLF4k0RhYLBjMO6D9mkTRKWLG
Ppyz0kvjSRGA24Eyoo9nn6Wa1vrjMjyU5nKKt94pu1rPnK/PpAcb0PBU8xVyYRPQ4W0vDK4MY+4t
H8AW9HO88/KctLgJZh26kyhvfsw/iJJQw2YigDwatFd6n2V7NKTDVuCYo6zs+uka/Bf5I+kXjDg1
gpZgvDAleUxPE8KgtT8kiIxllHB3fxU5EONYhuPe84fgkO4VF7UzUYZFHbYhLdrZmAcqCGGRP4UD
elpOKL6qhr/2O3f3IbpPqKkgYAOFDvBb71nZ4WaRGQcLNjo/N8TlcwDzdGBlXy8X/c8MqfPRVlS+
QGnT89lqsvTwBLGsGI82b7n9QucWtTNXayPPkivd/ukkmiDxHZ6ZkJ/fZ/kxzuQeJbK+KGSR9PQ+
hm88vbNXfN19/rO6pEz/YulGk3ByH016ijwGlZNe7Qby45aJHp3ZmeNIo6YXN6rur8SU4t2exSI+
lbm6z+2ezfGfdcKebzcdLHVir0KedYiTtcLHdvyqWVFOnn0b5Bk6QTQXaGUpk4ASpKyzlH/FaKj6
GoJXxCeT10MgwivXFZMLgjWHbkCC/wxEOOeEau8h3p4WPxUvYqPY3X4nAB1FL/xBL77NXu40sU8s
vKhKgKdkk2C5DqF1R7Lww0Z48lyp+YO/lnZEGP6JuUht1L2aJacIZgkCZAlMsumz/avLCp5koFGH
YLSbUoKDefqs7Ts2fYZsp4NekgZSDDkr1v6tewjXmOM7lLAsOHOu8HSHsaU7sWbohtO5AcI24WYc
kKDu65dKCykV6JsBH1ebSIg4frdfbcKvIjcXxMhoedSIirAf71prMgzhnYv/PRSHlYtVASUfoOkh
FIElpJ16v7Ow36WbK57/MQ9BLQWS5PoSoPEqHEa1zBnOFTBoFuFuqJx0srUxH8VretIsjWtYFiun
AQL9KRwl/DzPJYpn4jaYITI9GCScOrFwVbEHV1HaqSJHhL1lGb6U593EuNpbMByr9r69AN+JiHwC
W+afrYrA4JE8cDZPNCNatufPi8BUzAEz+vUHbY2bBtixiuoOUvvZ9sQhMKpiIIJLXNSQgK+L0lY4
NLfP5mmkUj8Yuy4fEFDTQxf+uVQb0qmB2I4DrGBClgbvFGE3yNsDa+LnwfZfgdZxACXZi0F3mKyd
N3FrwUM4dAKC5+ksQoQ/J7cPLTwTsR7X6YP6H+ezDvkgn7FH5gC2f4ZG0Ffvz0cVdtXRIAdyw6pY
D2eKM9nqtg7U4xobKFf/41OOyXRtUMZEM61ZMhAkq3USuMTvt5PWCH3vxwvb+ChvSEXB/bVL86li
U4bYgLFSynRURxS9wnYarKnLd4l1MyHTscWPzgCFevmaA44Rmcb6rC/VHXGhxQozTnWPMriOAp92
6LgGFnHE79Lo+bpB5D5hgnigpU7Doqlc2D8YC3yByTvo/df9r6BaZ+vVisS3M+2tJRNIzLd13p6c
ctA8baTGximaxReU6oj5bXinV8voXYecNycSzfTWk3QOJ2YGNwwh4U8OSlL/rj6JGWqduo8alWSE
FkL8HfUX0xcfrDygFw2Jqah4k/YzHpekWcOhtdqsts2BgbejHUDrBjlhag8FiudqJMJHzTixhdJs
gyNH4hzwygsY80uIAFQR3K5uwiXM33G/KlLSdEwiwGND7VHraxlRnWoot2SL0a8Vy1XRlwJiGDcx
2xf/xqxr5ddlNkkfF0xCFcDkTSCdwxdWwAU4698PmUzIj4BviqQguIuiAe3HGW7umdx/UzSckQK1
km01Zj6frWJB7qv4FIrfJDLNgy9VHbFr+opUEOF6N71sS8bGPAs3Me/ThFTmLW3uvfgbQ1FfJZsQ
eVksA1WTVvcM5CKTpsVWLQxa5BKDoPhZVdP9UVJKcVhKR9xxJNVKQuD+0WO+uQak7udS+hosilZX
VSFOZ2wewOSFX23fqLSn3DIyzHv+pxGFC/Ue0cydTZPSPFm2V2b7S/sQ/9+F21zWxH1al2CnJrmL
RJYxjUH8pTegi3dAEfHLT7ByjVyq4iqm9ibJ+S9PzAYoenkz6fHxFLS9G6z2DZBlfD+g9TJkBcYn
8+CZtQTlCYM3GEMzvhNhhRL6Bdb7PknLe4++mn+QH3b0mA3Tpo+IY2wZKoo0FpVGQ/LPDbITKZGL
lXA5IoxOut3b0Ot4ZWRohgP0836ryl5c9bl7F7Xm5gbCK3qOTqHbdrkENgfNarg3s/VCPuhNUPFM
7OlA3Dk0nirW7I12WzITA+ZZ4YzlIlivsTxj39Op3hjwNwLut1hAM2j6Np53Z/5sd58UK/X9yhU+
l8AQvG3Puhd5PqUzzrN9rnAfDAbJstB+3efGjsbjMeUSNw+04mYpb57sUVKJA/7z00+249NUWouV
HLkYk16vdqe5qJ98L7QFxztDi9G+mBGJ4MnU1NCnUbOepSpbGUIvm7s5Dr2/glRdtmgYRPhMdTs/
yJpMMqMwLw7dhjufTUNmF+vgk5uqJuTbTSH3m03/3zPM4tzlQClZgtXRRMJ+B94epyS+J4aF/Hpw
k2a/Pt6CnNCQw0SF0N7nPqnylx4GtwDhno5oXJXPWfC9rJQL+ZS3sbobRuFX0La/ytoMCBIpMVIu
EqeOye29HRIEVKE48Y9Qq+LsNHwr6JZXNMzYe/fXbVP18QDzTYS1Z810aR/qBskX8YwUl6IS3ZL7
Z1Q61nSG51ibMuOt0Q2XhoEKb+RfASNzLTWVwXdbBvCLcFCO8wkd7zUON32Yk1oSJ/o+A+pXRsKm
xWY5lMs+U7taEa2E0DioeiHTL98MHVoAJGoXt4oDyvxiVUzeKEeWTcUU81cri/qfEoG8Z/SL/m13
i995ksR5GfrNk3Aar3VQh3XRPj8CSRYfNYVVZ2A22hgEuUBbZ5UuDPQBSozU0hjgTQMtmqhxUBln
NF+4mjjCVLBvy3+4SgnY7IcWa3pW2Cyedo9Z/Iq6OoDFnm6dpuepxAs8x/EMSi6Xb13zKvJIy0Fm
2ISMZZJBCmBQKJbUiiTEhrHCUdQ2MIidYdltzFcpvKKx157XSVPhlam4uHEHZl+yApU7r4HwcIEj
UVQaFY5c7quj8oPkyowAI+sg8UaSyIbTRXJx8VF9aePmxaS97qBNAh567AvGHfnw7DZg1fBkCDlD
228jq46bvgI0r9f5Qk4KCrKTVtlijDILcZ6nIi5WZtpmpZveWC5stTO871goS+KYFXEmkXdcHyHs
ri7515znRwmXHQWMh7MFet/IPFvSa87AFjVp+bD83WgxqOvKgTGHL29yIaNYVUPmMqht+i/vBXbD
WUp7PPfiX+uJbJbbVXKOEzTAZeASo/LhF02z+Te9rrfjEjR1nzk+HTi+ybaqUZwKw5SOx9nNNpcw
XcSZAj6bTu5EX2RdeCzACib+rOfeq9uXZlTRaYm+2Y9i9RTjHwokUFQ/E8v4uKBq95hyrUcW11Gd
wML+ujKGcCKPLkK5alzdUcCPXsJfkv855GoKJxj/Xb9zODsLrwGHhRETSRD47EcnbfFJ46hiuiV6
jNSNSQreEV7ubx5bmasQjAF9FUwDfsu3ScDdKL4Qlh1lsuM6j1EVKz4L3kFY2WgnXZzXI+QlexFh
1Xi81S8WRP9l/BIZO7bvGltNAjvRHRjLzurNpdiCokGst0qSM1QySocaPl021G8AZ0hOm6T+zV1Y
w2LGXd6Nch8DKcjutpZaybJkWW3LVXsfrmcRuodfKiq3+YrenLVX2rC97U8e1R1iz9th6IKQEXsB
89Y65q/yzzAYXoDU5SIwhjbhIme/MYOPoKvhp+mN3vnoVG3vTWuF9gC2uBMV/dHaMd7dc521LP6V
ABYxK9bTMI0iL/WGiRSkeHA0N56jaByoPyXiFXc7dWrmBbUMi/ABp5sq+IBEMETJJAFHlwQW8Xba
tmgvFdchvN0TQGIEeYzuwVPXRAmmpY0DFCGIQ5Rn7lRjvZYArhe5JchuBSSEWhqlX2WDFkgv8eCQ
Ge5pXydoMzRcXQdtN6u79mNlkBAej0kc52LkydXLKu6P2jLsQTzuiKJT8Q5/IpqTrYHXbcxbFKq9
1iRC9R7Ai0QkEyY7qHe40isyvwhIPDjQFFxXEISqIECf8vI2eQxb5k0c6tRJ9EfiLGORVrIDZcXf
u3ltzkQLzvYjuotW1f5T7w+7o+p8MqW03RZaAjwPP/FxrxPU6UYBhnGh5Vpl+viG+9//HY2dQbxX
s2UGsHhedL/NE4Vp2GBmMHkpFjogNjc85J1j567edWL4sJwgbk2zVazpfEIa377Te+OOZ4iWW6sJ
hAJn4f5wbYa91OeEN4KAAO/6PvOItYPXcP5LGeBt1HlX2eG0ObKWELP8OLzaoc9QkK71C7QpnzOj
Y39VCU7PSMHpgmCSGs1W1MYiIl08X3x6uyn418MBE+y7Vis1j12Tyh5Lh9+GpCwJetdUqRGT3Evb
0EuoIbOpr2rLWD3YfqrfL2wzI2gaaHdY0/5UE9KuxSYkjanCJMIM6/TjhepwhEAVYNfss275L6K1
tQft88Fir6HYt6yjgeRCou0k84O0oLy5RPorECsaXe2q/JQNz0czGt3ly2ph2GsUei5GKfodcpdm
5fOhmjRzDV7Grw1v0hoR9lF9j3fqqcLNqqsfi+D0s/RO1wRDZYVX6G/UAtxdtfaYQo/Ky8D9WU0m
dsk5DFulUHxnlSYkAfssdVlbtUOwnGCMu3mrsZYxa8H3+4kb7qWf1R4Uybtv3xE+1gcgRZJuezVN
TK8I5xy/aZdXO5ffAfD0mufoYu7c+HU2u6z2nmytAq079vGjGc8ich22T3NXH/jriyDpz9y2a1rr
ddvBH/bgrjCCIdn3Pun1z4unPGaNTiFL2UkRdp+8bEYB/HGHfC74AU+wRrkTD0oGGSamODyess4A
2Cjxs0pxDw7osOfLwBXym48Yog+VsM2m8kLPpRhJoZ4uEtXGp58/aW8XF8GAwy+TRD9J4vVsqpsk
xb0RVm1OHSuftGZuf51jyQouY7Y1cFsQ0z/iGB9+mMjEOVMSkqb9H5CTWhaBv7Aju1tx4gPqJuyS
5TdtG3DLczSHzX5mwfTvgudBZPau5Xi+dn2/pNL5DRx6zfDLz1lyIDSJoqRw/Ft+t8vccBISW0xQ
UJ04Sxdkw9ef2FMbGDOOYeI5FpSJpK8Ur2tdJ/JZXDtKUuJ5FYDv4RSx52nke+NQsZ1Af2N6asMK
sjl1UhSE/Qzo6IBtPDbS0d85nTPUC6JezcRGuSbntuBngNNdsE8vaQ/I/s4hzn18CryFUHz9PuKp
6oHIbXkOw9bwMykuTMwv3JVeIPrxIzN/9sUtZ6uI5F6B+I3xFYFrQGpYkp+M26XR00NhVDCYvKYn
RitAPsd1+bSaY72knmbq50Nc8YT28AZeRRsLT1mu1tTspoRj9HLmtqyl2hp0sfN4Cv8fC8WcDp91
7bCUDIMGSSLSdI9j2OifZT7q0O2bwxgweCVWM4nTEb0OyGMZ3srx0h67y/DD0RWdGsjsB4T9WgNy
FNyCvJptRflDBOzR2a7suN21/R+7rKdPQi6J0oHpUVaVN3zOnSJ76g8nvjmIMhDgyQtN+9DZtvnr
/t5BIGmN2lthJFpPq/MJ9g6ULe9K6yETI928amyqTTDjY9sGBhYR5y/Xu2YTdqguQsRvvbZ5zrRy
r0nItVTviyJXsIsqu0cCuMhppbGQCt/s0t98Ilr/CErQLZao8xRSLA/6Pqp4v3SVV/GECO5oi9Iy
IkFyJnYm/8FPkRDsGKBjjmC4iR3ITYM0d5vLS0/Gril6FRj1838G5SFN6wS9ZLBqkQapIb5bzsak
Q1ZQClM9kYZntHC3mXIFQ1wZIENHEWdXuDoPQ1DAwNImGqVuYTW/XPElE5/ENqSce4rSZiXRFEeW
eRN0XsDyWoq7DvHC68+E2PUtw5DMWTafjJSmNdSxExzIMypTXVwX5tqPsCf5RKJOdVX5yPyEA9rD
FxDrlghvIFJ0SeffzuONAckiXqCv8XOmhnGtt3VbJsi6SPpf8CD0G8aE++TVVQ+OLo9tFIf/i6Kl
9V4jxa9cnDtjSifUXzf32NILo0fTHyypNcIaId1ebjYWyKH/Lwo9zHR3wxP+6mkOLVtevVVE7+Ue
LgX4KqUOdQ9oX+JCDKOuJUGAXOvYvy0++r1ddQAX171mOvFtvKGr8yXKGT4+beu5OOMOT6RhAByL
y7C1NBI0kZeszTtkWE8rPezrywGoRbSMAw4EV81v/0B/szlz4k4DJP+4w0xvAljnd9o0JrGpBkBA
cuG5AIgXOnE+yDd4vTp1Hg+Uuejar5HqFMAjmizWs5NReacTjus6XkTVFxY2vwjIzQ2IPiqAtRn4
lcoOBwgG8oCvTgzBFrG7JC5pv6gYw2wo5/PM6PK7y0SoKJRr+CBRNIzvl/eVk1D+zSuoOSXyZSAG
xzXG1fYcACw699yIojaKNhiniCuLwcIpVM8hPZkHYoEh3KeTecz/wXGcQC7Tob7Zl0m9ZikdPbi5
Qx98xKQCbz2Wo7qITJ54b9KSe0AjS47dVuQa4iEbaRvLLGh/fLDpXHYzLd4vfSZjiMJr9fU9JjGS
N3/GBbzL18t3t/iYnNmOHrDCQRbi5t0yFpmQE4hVWB8QXYxBL54/0wC5YQwE/dac4FEQE/M4v1XP
IXf/kAKZ9/MVhOgDniHel9MJGk/SsyH5lWCdKzYKWDt8YA67I6211ga2IpEx9h0OXt8IbRhZFhGv
9vFajnFD/L9Bb58jmY6Gks/cOLAZ+v9net15XkGNgVD5bTvwCL76p8kz0QSePVN9KadR44oh2pm1
fHV/Ck+GKtc8gDMLk5Hux1p977QVfmSyd/TZyeDv8gpe/5yFpR83x38/5ioWpCjSQIsDl60cpFTx
BX/6lcc4D9gHg7QkBZyfEAiDziJFKngdav4khNPqOmeER5v5QQmpzsqE4DhrBHz6I54sDLpCyA+5
5O6jU+8G63NadsFTO75J12BfXvJmrU1HRUmTw3pjEuRu8vFlmcmtTUhno6F9SmPs3wuFXhOZ4Z3c
lxSlK9l2XQ6KImS3ZG13bGeK8ADerFQDYN5ydu9rhgah1hkuqTZ/76sW7VtIjz7NDy/7Wm2bV62N
IZDi26gEbbDmCc5NVCPLO1U5Ylg3g9wYcqRVw2aqqdBbZ6TzjGSROo9OPXqpSGv8h/jx0I8zMLCr
2+/hhumwXrEhXN71x/vmOTMBS2rHpYNbDqHm50AKwvhwfSs1vN6JDzzQFtKEXjCc4lqr32syA6Qi
LaEtyjo0b8E6ExQqqQMdfFocqoXH5bDGG9NLZv3tb8I8ZuV32P1oRhfHl7WYxdD0LkMDZn/Z/JnE
cdcdDzoMKUyf3iwZx1zjuXPXmduddYW0hHnsBUJ9qfzM8wXwx5RdOBTJn9kZAHX2BR/6cBn4OIY6
37nMk5ZcUjjAc07y/ioAyGIsWcQ3LBE7qLic6AwwwlC6IqXXB2cvI+mUzC79UwR+TkVacrpJINvi
1Cwq0WUu+Ghcg06niLJrSCr34jJDicIXiXhA4BL09FsfeH6T7MpKgaOL0FLUuW7pwYL4d+1Mep5c
+GsMpE2FDn4VkiQ42Cobj3xL4/r0x1uUr/ueGcKZsU5YLaifFVkJw2fLIur9FkJgmg+jCKATsn4o
bkGZZoX70s6wzCeldGBud6T18O7jFp46TG+XrsxJe845GeIGWtXdvQXWfoNEoj9laKIANc03JLDn
6t3FO/o3Up06OfRtKjF4kLuR+CrctvF0xBoGln78TOnAcLMV7V0oJtDLI7k9AuIiYiH31X+Ki6Gv
zHM7yiwGhM09IDkPGqzk6dFTzET5FEDkNjv0paOC2UXi9eLIPFnNJwklURIbJ8ACcMvzuXRYR3b9
I0KQX9DQNbbqeLm/IdKqIlJ1wiYuX7XKZamvp+BoaTWInhEROyYImNss/St0J2qdoFX2s5sOwLMq
prTrZRMe9IsWM6Nyd6vscgZ/IZ9UNJtpZ+uybmF3JdGw5AVQbfRcH9Bht87ZsvfKAO45LLljNBR+
IcWh7WHjCQGCCaVcqZ6EFhUQ5d69frlt04XUUiwKyolXM1Kal3DtSmVWgLmWCik4CPZti4NZb8QM
QY0dE556lXKL6qg0yDOwk6MGzSZvXlkBblHPrnv8pNhuOuYAQe/06QwVuZ2jxeMOqI0w7qUMgeSA
f9p8kz/DiNQPOXGL+ep8Uq/jFZ7FQjmEK1jW09Ar2Nn+kAG/GRIQZIjOodXUvQzniSMVYldSPAzT
sGniwStWUhr4L/zSm3iNcsbvKsJGrFTzvACfZP56atP6NDCNScEE0CcVAeCaionSE1DOPdjTFwTI
bUvcxQlWfctwtnXTahGPMEC4mxhyCJY3uN5ZxvLvSLmqL5J7AyeITVZLLxAZtwocFciT8ZnarHXP
XwCr0uvMT4NIJWY2qNq86EPVoaWhPNygCe5yXPda+wIRwEyBJPGH27oZu7C741ccbWhjygcSfmdA
fLhqa9k/Li/youUDsBV0gWAWQxVd5WuDgDEHm/2q7/u19Kh0FeSkjuKsSJbBjy/XZeYrVYUbkYrS
wq658XNZVZQ94GHFtXtNJLGLIDpm0Fv+9kFwvScts/k78Qnr36A++baqyAXNmu6785Af+inPCrRP
I7GsBHpAezVgeXRY830C0Dm++U8scU4PXF5l0CrdshRZXRhS0JfUIh+Wx3uWuSXu7wXDd0bFFK09
x3M1KupfjiXxc2etDPOE3+tQla/L35mNU4T0a7C3PkRnZ2z2OL0gonsAA7FfchLd+vhIpYZwWXiz
H0esjdC6c/SZfvKOCAdU/sSAz6UE+W3JFQdrfMEfP60fnh8U/vkd0ZiX32ZJio+GAeQCevMUFk5x
dWegO/7Awq0LFlGy0odFE0V4tMmCKj96COlvZsL7YyT/RYRu0m6hYz5Ug79TbkKPyxSDbogTIUmD
fHc5rF3KDhEU3aAXJzbBCmQD7+LKUgR2LDX0vfJ7DXZg3B19fwU0Zn+jPRJmxdeUwHIM3V8c8cFT
eXX8czA3IpZYydC1K7tiM++6QtNwGuPIpTHNYQl4QdsBrY8TDslHfCk4gvg1psSQYrcJksXhGxl0
wmxIjBHu1HtgOJOP37d5OMiOUFo0EA46sUXfLFNEFr4zQGUG8BPxxae45c9yoZcio3W/FHR6R1jH
9qjVZub0wYCowGfgmVIUrOAsp1l1Lv0Miis43S581B1PwE2cOO7ER52jWTAjhx8o07aY4nqc4VYT
RBqLQiVgJrmStB4Djyk8aOrUe3I7WCmzueE4EE6woktZOjEOeGHy25u9UnYeoo/UC8M5oGI/B4YW
SM0HUxybFILoljjI4YJwUP7Zx5fYikX4Qzjp0ePwspY3vCuvJ2rMgEIl1+7usaHBFrEZSEyMQmZJ
rLvABaqTBPEAOnBXFgT5RCvFbduSTMn0zbE2bnSA2OY16gYM3KvV+sCoGNNSFXhO1Zw+NwYTX7R6
K9xut4deKwzqlp+zXtYmG/BWNtwCAc6XH/kQXmEt/iBwFg02ea8h0BFZ8rEJb6otX0gLNFQgoIXp
lcUmQ4yp6RPVDU4a+5EEUyLOhKBJupRCDt2tftA/wEvFBMG4UVynu+FhZ/228q9h44Q5/aSYgUcf
EoqooIWumklAogqMwoetEzf6dJ6Fr6zdNRnwglrYXdGBa9tEGUPMizbFnnaPSIC5FhGvZzvqKh7/
RGVFvFb0CkSeCzrg3CTs2+vdIIlRRXAK1XJkQdKswkwGdeZCSa8orN7qH5v5YlqVV8xrSrsPCB1U
Aq2S0g/E5Mu9a3TFckIc10Hyz28fyc+hO0UWE/X3/uqfCwt4BwROcSwXGYoT4tREw3f041UFGTZc
Onea5RSVL09QIXpXanGxeQhQtaos3R+No0hEaTqAzGPdiQcmYwhDiHrgWqwoprrELdeM7pPwPDQI
C68FkianEE5d4s7js0mYxunHi5j9QXpUdLhjSGXJWnLqhxbIX8wuTWnhOvrof9kr2CX924YZEj+3
AnNnO/H8EnTa9+Ddc9JnUJYFMlvIY4GYiBMyZlx9N4msSmlMSdvb7bIgLfQ4uViYOaQKoOzkhJlm
TcPNLb63iYCiEqKHQZ4d5Fks2rqZMqVUqn64aZiYcCp09RHx1IxGwsFUvrd3oPaQKE/vovISM9AR
YIp0NIoiixoq01f5qOLmXs3rFct6zYNd/NLONm6Welk/umgL/w4K/0paYtuvfrNrOUXj3L0/31Ht
yenQ9y86wyMQtomYKYyRZOM22rUeKfimxLGR1TWzkxvk3Kl7DgyoIHZbV5QFsZUjB0jzHPSYb4QJ
rKsnbqWe4JI/KcKJtawuQz3Czid/zaYH/cgAHAgQv8FudQrk4fcBGLEt2cUGXvMVLiYFb8rMzHhL
BBcXzt31ExaQklHX+90t8wkHGsC0TpvJNxk1MMH0JxbxI+0QKITd6i4BmF39puRUxqxP3geHzjWl
AvFiHLE8yng9qH3oDNSKHHfUiyYWBlN54JtISz9VWPZrctEdikyiF0JPja4mVVXYjHfadOERqGjN
Yanqx5B61aCDgD2VVJ1+JGyQTEs2Acn5rJWDV6DY1U5SjwVd78A6OS7PBvYV8fh4Mh5Dau/Vio81
k80P6NiEAU+qGI9ffErb4HxIynMw5T1NFUWaelLXFCCiMcwCtd6nlzan/lzXPkav4c8pUUMA30IT
3PrrJx+cr7LaeFNAtdnzOqUxuOuhWKEQ/kuShwLkKcIwLxqqQfN2zOGL6l1N1+e/5FN025uNgRll
LUZowcy/UxIGBTz62nFpBxD79Z2tXfC4WSLI8WWAB9NQeLkQ+/YQ6W/psZ+lMECZ3Cie1DjH9Ny8
JK3gbcoP9I/wRbya2rag0PGrPEH04rLCZH9WsNQmC6MOlfGAiuz0JWy8piML4zOYRAJzptp8HGXT
Njz9vZbMUeEXyvI8gBmLyk+ZfkaXQHR3VmFpX4E/MJVjuSxKJNUZ+tcHZnORdRt1+6z7UxMwp0Pj
2wO9dzNsRujzK0TZ5U6dYRAVJSbCsBXXpSLHjUterqqeMQ7s9OPmVuwk2gqzbUKjB0dXft4E4DRR
oyY9SXnx7icOF5dx/7qmKFTjiJwg5vLghiptqXrCxPPt+Um75w85h0Mj+6wCq7EqKnItKX+SUVfq
aBEjzC5rrOx8od1VUzN0+5buAKeremZpGMgVAafWzMNfYHpw9k8+kJnQnH0Koc+eVDOU4QNVz+3S
yJnboyicwphu05VNPnZN661wQ6Q8U0TrhYPy8XfELmUoQZ2WTgsy30BuLm4PakdKGccpgSU+6ie9
9yzi9U8p5LWznFIpPRm6zVzdIfY33loJhwICADOCyFb9+b883QaNUn0e9JCfRRYaTVacdk5i39Yk
lL1Pj7KbO4Ch4MmO6eWnAkX+xi9tsVKyBBbtLr95kH63mieKJgDxNbgbCOtiAiFDWRuZpaiBzZVa
BpVfUDieWlInSs6oJMCeNTuzooS2g6a/vABmCPJcuc5lozlLs1SVDF64Kk1hms74go82Kg1yS/kr
YhA1JWEVRFtR8qkeowz2WwUgCGqpC8FFR9aVTB5rtHLU1qfaWVk/mMna4Hadl4d68HpAb9F2EwLm
IhxxQP5bvB8EhwZ99NIZbEbzfmk5pVB9Mz8D6Laporarr507LzZagGwxXXqcFF6kcbKDpLva8lOQ
kTWqZyKzzM0F5yXIAFmA8RDRc2ytzU57MfNP4pnC3cO+TndqMAQRvyIYt8JkOhw7OXMBgmHKvVQQ
APaOqCnQ7AnpeMGBI42ugsfg/1kS38DLbcSxUzvDBQIWAdizgBWLgzxnXGa0guGodsVAc7oMpoGU
bsk4PzUC9jZFWT/nYgt8roeDUN8KMa8pJ3l6m17YG3HYYVVvVb7Z+39o6enX3q22ZNRPn0rBnHb4
FirB5PrGZRFiZDCLRYiED02RkiCttDnXuhG+cUUVzrK9UkCgnmWBwNz7ugoO4WlRohi2CosL1AcX
C6/noqqbOSSAwrVMWaV9SNFavK+rJGuGUPF27yLD5rOD4RxRggY1LErq5Y0bKPK2T5hvKzr9bZI1
BLu25X65yWTT6pD078Pkki+lO9tbqLSZ7QGRWX1HQ51553VUgp9kgpBCzWsgbrJDmuciWFDA89Cc
t/O46XdLVz+5498CiHOxzxjxD71jBb45J8wqZ6VNCo1GB8nkZSLcttxE2nPFwm2wv3b6EkHYC7Dn
/yLoTa/PK3CkrbM/VZL5kj0t3CcdrOb1XX83O3kC5e4kY8cMIhUsGmgUBZb7iDvkwaZjaPQNK/2W
Ip1yCy0kzg6GngPAHOV68czBDNbCGvcg6K8wm0t+bV6095ANFUejIpLo1og//1qmR7eSVs364cqw
aH90ObKYnWEnrbDMMxKfVXDutXOQ/AHjuQEN9nkD/yNJQ2QqekR/VKVS/PjVlXDfwrwrv6Xnqo9Y
XtTTn4uOvNuWh0tQkKQB+ozPnehTKc2B+mpcklvTCOPPGaSJqwEHQrUPFBh9uBR6gy/sGzKyRIUe
XfZ4zWXQC6a55jwcQ+K6+Er996rZp0wlhRycUPxTB0ZM7LXailY87IcuvS8eNZigtVKBjQ+c+Pyf
rOD1n/g7rrz8OLDqdEKzSS+TETrINpP4OWtxfKK5OZzoh7GmqnLXLHCYsofNGvynJTr9hPEcS4Xb
Wkdd3b3b61KPaOPb5RNluV9GmYghMeTJTsdaxWlTYxaKVU+wjFJ3apdeZMBml6D9oAjF9hAi3sz9
rapi96mMBr2qrrH8VOn2R9hPlHZeaCrSKol3cn9YasRtDPFrgkdtOIYO8igfKNwhlugPPgphgNuH
juWzfXUB9AbYbf9Ez1Sp/z9qExGt49ET7DXr53sMtzAaYe03shL2an0zRwJfYqHRmPmFxMAfeT7Z
gAJY6YnoSNL7mkr39xzLgCxlw0GVXr0Z4QS/S7E4gqzdN6Z2qRDh1hwZX1F9IdmcL7/zaTy7QzHz
kct0KnIH3kQ5KvevgtqIUDxUJaIfeiDNShHxERjTa59eEAuLHJeiD1h4BhxMBu/7sDYiBAs/inNN
BqKv7JAhiY1fOujSpRuIMIQckaNlmQTb/aYwNN2X55tXOgVj74NiUo2vdR46SWQ3LBbuDHDClTre
+YgTUaNQVlQPwEBt9Ru35ruVTcjAMcC5p+OSnFFiljoTVgAESLXsQm4R4smPM9GsbBjyeib12mjU
MTU04f7+ZKVJgxs9whCAL8x/ZwOy3uOm5LJyM0fNGFX3P1MG4rSk+aG1Zxj+moWyF2ordp42Dmf1
Ri8hWkpBzHv82kirqz9b5stjsr/L4wNWALHrv/D7Ve9ODluxQA1uHlmjPEj8asa7k3/OKakXB7cW
jvO8kPbLOywT6V/O5SLFXZtgt+1JBw8qykdYwz6RrOXrIO9CV2hB6QrrEuKBphM5zxONArceOJzh
ihyFJTbi0nAzK+qSNEHWO0Zpo/eLEI2lh6KDtlxFsh4FKGu8KLsxep5BuvA16pPcBkR0HkIeMvpA
+OCEApv0cpn4ORhfQDPg0Mi0OlCewN7ajJwYc74UWN58bt7adu/cXHAP/xwzeNNlyXYtJmZxUPsx
lv6KQZXqWjGU2vSYMVMZzJKYxGRRAVn1ekgbwieB28BIhI0MbyZ74XoNqg+3SBI96iDajh8WAm4T
wsJu1APyRJTsrCEnOVSH3pc1gbLxm4BDP2X7EHgHCk/nX76hO7ZTAogkFZfk0lmPoVk0MPKGpYsf
hV/UGMDnq6HA3kBXHgcfR3vX65mjwsWAoZUt6rBWR4xtViO31D3IyQY7D0YXxjxZsFQAD9s0DtIo
wFpBPek2+n6bqR0+rZzKMo5drfYyC0YRsbEt7o8/go1tuV7I90R05vneSnX/xyVZn09elx0mDf6U
W0HRsYY/NCuWIWI/VhZID3ZetwwcPM1JWPY4F3oEnmX4Nn1Lm+nOq/0GxApaQbF+uavN0+p67yWM
byHOSwGIROtENPrFTRejF5rzGFMErvd/369PKisKRbIR+kW+4T7dVN1ssVNoCf2yt2geE65sF6NW
P42hitPmay3m6iU63hHS4zNWCXNpZvftasBdzcIIV0SyFVHdN7jXG5QLM5NNLuMfr4eq0P3vpL8J
8lxu55jTOduobytZkqPBoMiSKy2oC9fDASjze4+cwMJ53rPXzOsmxUMynFc7rBjJgSnPv7r9yFBU
BhuvhNMDAoQi64a49ETE5yzQfYN+JPB8R5snIS9ROeLJw0XitfqKwK4PN+dqcb6YqcGPE9NcCxGC
XnzUKVFjQY7tfd7KlYNIuY1vOFsdUpvbPwIo2PzK1KXa6wqJVoKo4EnM9lTL8CZQuK8l4h+2E/nb
goso4rR4Zr8eyJjInJQObcFl7yKg4P/81wWHuzwMHE256KvI3SrzHN16KaiY3xKuijA+lJ/gBBFl
tvEqrNR3fnEMO7PzRRqPxwggwKNbt2cuabyPSTVfs/ySy2enmSe22OPoC7w+bFKsYek6AWVTjo6b
c5gfAHDj+PQ3xSCqTvoYqgGPoYbuKsuTFKVH1bntyKQ3c4KtkztRd4M1YOc4qWzMIxJT/JKNxHL3
ye99yk/Yl+rXioYm1snNMq6B08UwkbnD46XwtscGZKl+j+Y3NnSnia+ncXH2ebDXH2rQfzR0iC0t
0AP6lSKpzUvubeWtvKwng3+l9d7n8u1Tv9/a8M9h5CCOmjp9lvBaVQPt8dUsEU4q+/x5T3wt+qBZ
WA2nzqFFMVs2szerDeabCGJksQ0WjFSvZqAQWajD1PKb4WUq9bFTP31ky131x0++gqu/LhRaPO6W
BhOi0m3LGMJZdxrJ3XDNoybE4Vl7e4z1jpcEwwjJjT8YJeXngUxPatfQItE8eF6aXslACsKRqdoN
J0juuLUix0uAklGpNCktTdtRV/r5+4LXq5K5CKamguwmgEURvizXFEXeeENfUwmDg3xJoTfLgfpl
l7pzn96poqdt3Hu+PJ2BOWcv7LHNNH5xyg5xvPLLkJpnX8R7z2K0+wlT0HxMcpnMxitYlxKcFixM
T05xcl0vkd0ihwlVf4bItfdrrvCtZ9Q4JUQvnpsg0AhinXtODQzAQmXwgMv9PEiS+oyAePHjaQJ8
e+rn7vMWYoKTNNUupqOEgRgt6N1H8SeDACl8qzVOlFkYKSrV8+CZvfM7OvT9+1xr77bjKxxLx3z4
66v5RdeOGbCNL3SbC7ltPnXzAlAKiCdkNZ+I/Wb7MNnl1ak2s6I6fgoGecK3nPwmWW690SmNgadW
igMB1kKroLKwjhG44MW3uSy3HDyd1DPS3tCLn6CnVmLxxqxrbrVzvYoT4IMqnlGUzOazgfaXKRkP
wbZ0cfvUhDOdxFOnGsF0i9pIVhRnXk13GvYmWkjRP03j+oaWyLY6m6Gu5+y4Vs71hAxMhlIPhwQ/
6WnazDs7JzkiXdgosFPnwHMlBFlAQEqPFDYiVZoshjq4RLeTvxDEq8wlc24FcbOb8b6syNnFiwkK
79PNgA6JjahZOF4A1ce0WFnzEuUR93uln0aBxNGWR61UHY9h7ixk5IUib31fNQ/qM3TGlCjdOj1S
s4fuZG0gA5Bp6Jby2DwHARm148i1pkF0mlwLz3qlPtqWrVhp+coJS/LrxmsM6qL1kFj8EoiRex1C
YrSFR+HRAEFlQOsjUxfUDDI8SJBFO42+AA35EEoP5lNM8/sFNKjCOow15PeVofKofOOA5Q5lOLMk
8Ja5N8Ofg6aAuHsKlAaOb+5zn5Fld6ytVnuXfXiGvWQH12u5WFsYqlqh84VFiNiQmaBOxkqEkwO4
Ifp6hk16blh2mx6cXqGmLpHhsxzYmRxNDeglN/micAgiuiFfc2FFpcxldV2wEqdiWZFeOoW6/BMJ
xTWg6Xmr8t/tNv8hmWW/EFJqb0gEA5XtHVgGFd8m4yJhJYijHGNipZlsly05Ha45qxpurNmwpqzi
KwOwAp/jnvyWK3Cnu6qUIC8qviQTOcDtrCLwr9bLzF6vpApbYSyVNjeAHhsSLKLKHVbMfmQ55h1e
Ar9CE5P9TKc/7S6QETxmU8+F7VJCz0ObS5C9pQ21sn7znaB/bz6+0abNm9287FATvs9MAIZVOiKa
MdTNu+QWQnArPNP4Q67sk/obo6NeoOpKcbx32Zt1k5TZKh3bQr7VHfItTYmWnDfX2fa3y3/TVfpo
7UvEuUR7wlyiCWrdkDgYUzrU0No8leinrlsQMGxuXXwWghkEWSq0Y8L24Mxeb0kaRfdAwmG/pI3e
YmS2qZxq9Dg3kWSQUZgDMtlpHP3RefuuJxf8g9l3dnLWTEgEqB92nxwlatWYAP/1javz09bBwODB
PZ2azrFZzrNoR0rqgAw5NrMofS8lnf204WOJMiPt83tCXQy8QakBP+kSvaYnkcyb/W5v/MapkXqk
YFIotj8a6m/+VTiFv3KOU7BJ89ylTr90B4Xuov6bIObTFwECDtd+1bVh9ud22CpkKybsM2Liv+BC
yk35XobhaMHKOr/Pg5GSGaYJOhkvbwLuGx8N9XCPPc7rp2MGsfzF/HGK7G6u5BUbFXLzu330TYJx
QHSQhxE/sja8FTOk8/lvKY3/3wCW3vT3DUhOV5xkvy5Bfdt/6BT4Iv03AD1mMS+nhtVM45RFXIoE
hg4LYE6DLEBO0+c8AKHXWqxEU1jH84jdYe05KRWazRp2lpEaB8vaWQaRpf+YCtt6xyKdU5ueUMED
DckkbJKyJIk643+T97aTGSTMePwx9S5+ge1BY0jMcoBWQAeuMadaArzUq+uIwQLNsiG1IMHn68eT
qssLuC/c7H1AtnvGRX13A6BYRvM3Y/Qz2hnT3wtE+0RCaHWyOSpgFzu+vbX9Y34UmtLzOwibxAbJ
yFRshlKcg9FvlZgwTkMK3e9UFvwjHM4Gkl4/KZIrUPj2+27tGhc96dnQFvmxfhsYCBe5L5/QR+g3
PP37uFehw30XxJf6duC6UGhEshdCgfRZohigEmI1oFVK7ggzbHyde9Yl2Ib1GrOCvSbpih4Oiw8I
Awf4ee8YnJEowW6K2ZYOXE0A6B8AH4MtXKufC5wetNdA1yCLotzUHWQlQaCML29Kk9VjBsCYuT3M
rHrMjcbAltS7BsBWFDc1w+QkyMcl7b1yabbGj2flmG5/2XrDrXw9tbA6kfkBwMgsNOA8FwYensX1
EDgd1CXXvyvq2jsxPwqG116mr5OpNggJPYMt3wPthhtIXct6SIY1LYfm7SYfbRYEIPFzuuoSc1sV
zy0Hzt60+W84mX8HIXPGLTgZYf2hp46BliveLTzUIkjjLjgSxWBJZ5wu+dHt1cDZMSvpeV7YSLKx
SS3Y2PXRAZdrm/xWaqpkVwLGzvU8iQE8nriUx/e+bETdXH1crNzI1EYn1fyNt/Zrq5tZupTCL77t
5wd9OAdeiyPcmrLR1aUx+aC/+0CQfqH1glSbxS/TMsW0nJ7I8bRqdePKnrisOMjUuyzLD7Nfg9K2
HwRa2IBff3l2tQ9giCknDrsw54i2CJ+u6HJ8IGmWz8O01Nek/YLPIOBhheXRPdMn32caPjVkS+uK
nyr2Qf6Zmlwq8UTlKmW7ynyZ8TWRdepY8f19qlwKrUa5jnd2xNJ6FvMMwahwiI5iixNisW6/a2lG
vNuvdEmPKuTXZhgtDnB2xtsA8SX0ZtUOuEtY1FThukLUDCM4v9RLYnE2D3woBqQc+/+ZgYXnFDQn
wtutwu22kgK6ga3MfkBgoq984x7xEq4sA5/zlwJEOHnojhPOeiompSsEFwXO1hH1tr2mm7iY/ni6
0tFxIhyg2BqogzxnAb7O7qgHwZxwX0bN2GlpTzfd6yZuDWB31+ng+KqI3mJ4NRYFevvlDA1rkA5G
/Lk5ZWaIM10xdCy7knWVdaB1UFcmlbloYovdSMNhJjP42HjQakxj07vfDqnLg1e5H/NLbYKDckZO
9cuGdefkuJMOf1T8tFOSAO96tb/rYsP7nX+kfMfDbj9m2bucJeNsiqTMJfleBZG5it83w6V0YNg/
0Jcn+fqK6KFS6fjv5ngFrvdy6pMD3I7rbH7jeaaIV7Kd8Z3hqgj9IwQrT0q7Lx2R+mPfWWliSpLr
EY+rIHYvjQ4hPYQo4TnewRysDOON5CZviRG25nQBX/nH5ra9hX5AnrlmgIXFrwYGsVs7M0mbr7yN
ZxIjplSAcmQ+tWDCG64/o5ELgGqaaOENL6W6kPyAjrdp4TGX6drS62U/cqQraBMABb/xSAJ1yyIV
FuuT1+EJDoJWYSw4vTNEdNmZxtu6ZKfmOkOsZQ6RTTZQCyTL0Bq0iG38gaXBY9/FrfTpwzPSgkxF
qcPrLfqJccXb/eHf5UK+EySV/fsetVYyUafPzRencVo2iDUdEyJ7604kVh/S6B83ubG1LzGr2JhA
W4EzGX6nTgQgANIsiBIut96gWj3gy9C/Za6n8zJ78N4YctvDngMx0BuWjzrixmN8JsmuFNvzkd75
nLQ+xYEeJw19ITUDbTIrBwK2Oj3PGdLWy4T5A38J3oC1y8Sr6lCky4RSuxF8UpV1zMe5FgnSCKqc
H8m7UPTD1Dc1fWSKHuGHpGuhPEJlnkRvK4BsyklJHTZhWxTlK79EksllSV4pUSXEkvZszaCxY0r8
85iXK/XziSUHYyX0TqisdFgeixsAMJLzpfVEdipOXcxKrkiVr4qilQTemQ+PUH8587KGPnkpxZcw
u90VBNtqcmIjBcQuv/HApO/swKmUm0BB87ZNhZl7HNOQXJtCJUnQgifB3m5VPLp+1Z5YfBdGrVVU
NiqZpWn15EIIsJkEil3qIey23hDRXPnzy+WSZ+05ASEvINtctlwUPQfRzKC8rM800Qm66B0Z/bwZ
AMfq/arnidsjM5kGUo4zC41bISTid/owCgLgCY0Rb6YlZNrmvcWyFZDUOIIWAcG56aaYifNSWXzU
OOlOalEhFY6zPIBjQIz8Owa2WdoLaRX9yvo1bwZyEV0GBlCTzBJ6RT/zJ9YdlkP292BpTtbXdLPY
gAOLg6GgWLRCJYsuIOtbyfs6RMoij2+DKGoyOsucim50/qSmvfGsFFpJ5xaQ3Sr7n9Joyjn13q3W
KIRBljzKo9+bSnwtHSEh3PEfB2D3Z552BVT1cVzr8PYmmtasEKBSEA7g8aMXyK4S7cCcoUKspDbq
qmboqkxBTL/BG0/E7nt1XJ47J1zKGw7og68xUj/grLTkJePhw7xBPiuU3GjClPcTi0xLtoeqnwo2
hZfOGDaEnp0SEFysRxB4U3nOE6oah+L1fHYaqJGzZFclOXHO/T/88RJQIuAJpqusIBOy5koxq+Oz
75oxAIxa6UfyFZapTnNvWH0lUUdiFZdimRU3UnqRRDoSDPpjm24OfTud2KQdXTKjZLzZQiOKmAo8
Ght4TJMq156N7aaKNWubRMjR5z0IBmf2KYf6ib7zp8ooqhBQlwL06Sfd5qZ4t0qhgEaK0+0Y1EF2
7cBmDX/fZKGYBUmd+SRxYOtTqA44vSbrDPfDDp5coRaIz29r2H9ytfnuXaMyXb/Rf+gWEaf5AvHq
jPnTU7Y79MyqUJR59sgKF/o0/qNS0tRcdCV//PW0tFYLC3lLsbi9icaUhrwBIIP5Ktrb1VgIIxxz
fb3JbQbR0YoQ6DLXUWaEgG5eGLXNgOZAZKk3hUSqlaJyPXBTKgParOVFc2XHPO4/S3AAhzN9Fthh
8kDHY4kHqdObs/6VgiT7AfIYmvEL4+gYpLLSnRE07ArFq0ypYwfhQdbrDGRWLNt9nsFPxTpyz5h8
n0D7GyalLBuoKY5+BtRQ/cprrIGFkA/NLOuaDRPfGixxxHo5h3dH6C/8CuMR7psrvuJBl8lyOb5K
srgF0SEntEUqiDKWqjl/H9ckz6qYVcFkDoo25S8mTFPuTJlIi67yulQG2CE2AQkY7ZyWksrNMA0L
dvRXX+5pAj1+vBrvkQrFkDz/uas0EAAUCfUsVSbqMmLi2R+M4AFpZtJX3r9037EI8HpNeHu61rlb
K12TWZdR7vdMzjQBPY36j/Qo+QVL2yA0deji3CufsGQiosIaBgEJF4lpKxlke8eiktVSaQ/0H+RT
7jO/f/iJ1iXHrooziqp79q55IutmibEMY7IYOjy3YSp8M/PHzLXbr/z4vMSz547FE/ZcHjQxp1Un
YSt1FFgHUL7F+J1Mb5VYB+++8MucsEOXhu9i3jB8JTCieGktBAOJEW8FCdSmTbv0zIDBvIwGa5Ys
jkvOP92NkTcmXmYpliHvgQ+QxZMNOv8on5z9WmUUIfAAL/HrHe2EkF483EEQTN4CL2dnv8c30LDN
p2Akuabh3FLn19aRkE/BKzNyfu0CzU+oexbBFINgmND4xEaYH/Co0AJ4tiJFaGDW5DQ2baAZvShs
O6u2QOYgJQwWyy+aEaLsciP4AB4S7b4H+d+0npa6JOEjhhEvb7zhPzI3/qfx787jpMCvg3EuVG0E
hlhfujErZQ7BOBm4KngsH0IN9VbutpL6zpGTGds7ppPieauFs9Ga4zRNUC51WjDlBlutxMA8VF+l
wZO4bWtd76gQUoz+Zj1EI7quXiZrxs3eMzM2aqmhOA7dsdfOhhWntEoEb9lQev11jc7IJifB906c
oCAZjwtApZAJZJFYHrh+AuD+LnqKqZVqezWeymJH5Q5WdLLchCKAkgg1E5u9heZKiZpqdbpZ1XTY
qnGPwcw96aHQP9bSAx0IvAV6IIIfCPmC3zxl4BNh1Wl1SaqfIVqWjOyg4iy8hJD5uolerw82unrk
XPwbcIfEGBVgFZwBt6qXR0gRUk8aSSXJNXrCpFYZzkOIh4Gy5HwyF36c15ZTQvTtdXcnzprp7cRB
qxhG8kWw1GCD0MElH4lWOJIB/aKgyh2YFXJdB8mhWZ9st1totkoTQklzCN0iNR8Ff6Vg1z+/IXS7
qhyHTi3Uq1EMofAqa5mKeEPjacBQireRCBMPtQYn9JeXnxmZJwgbB25kajwwpz9icJzkYbw9pr39
LrcU9H46qVweAfvYIbNi98XGnxeh8KsP1pQDw2L+WYJ5Z4pCIAuTGr2PIj7UYRUIfbFQqqVYnoBT
IUj/3gTt17QFagMHsGv2aT+EkzFpqUznDnZozYvPCjY3MfFDPaPwRlljU1zK4LZW//WLBYkm5ubl
JwRv8laQ7QL6XcMq2mmpCBmDqY0j2/pKgOjlaCa0/Ww6aN7lXUo1UL3RbLdnXkNbB8meSCDQgzwm
sGdJHVc/ss/sMDa5hupwdF4ZiMpdw1+UmuIjYcp5gk0DlaG5VSnQ7HJjVih5mpj/KPee9Jm+gt5Z
4Xsq4VWaQXeGrEW/xeudVWjw5y1l9QgRx9a2cbix9AaW/cLBpBEUpaBkAwRybUgDBxLU9Lz+BNpk
h2PYj1nGu3WtGeCLDMiumMcZFb96MGcbWDatLhNcc/wgSGXNsjU4DZY6GXrq4FItBqq/IQgLuNTc
t+GJx3PN3H0ybZ25uF4vIDnJMjfdzR53Cf+bowCgriUib6NlLZXOvTJtxXIE7NGs7G5jCDe/8LCW
KYF102M9SCEJ+Vfx0/07Cfd+N8T01B/uqdruZUX5h+0e0GX7E6PTBOXKQgDI0krlZPpRuWhjklWO
hNC7op8SBScIE/Ex2UyJpB1UyQlKySuWdlYHTGrNKdfuU5ZOoDAotIxK5/4gy/NOuqV2wGEt2mja
MAefhzuQ3ePUi0TywkJIO3lLtuSFEKsMi4dFc/WbGjnMGjPzeUzsRfry1BiyLIgCU+EJhRyQ3EbQ
pDKlUO3sW7S2q3ngV7aMnlbCs9gXJfd0UzwcU8cpXNEu7IZi/xVPP1mAxApOOi8wVm95elQNNgxY
1GGb2RwlNtBKEdbKMbK7IoIuzwb1dSrzFnJaNokQbmmOys20VOoTVoVp4+6T1egvQuAhUmF/XCjA
PBPaz7HhA6RBzfJ6FYY1Dxrcku8HkV5OORUqF+HbnN32w5uPlzTu9fObKnDlhomyz096Bh9+CFvK
a+LZ/n5K3sNrpj9Rrx3o+3IEPuDlCtFleIa2xIcIC6gjG0qzCInDXdGegNPIVvHwfBT1knuUNxtd
S8KTbBg8zX76FvNA9hCVpoV1kj9sTDk1yPWh+EX41nwrno3/4j5EMlP0/TQYHP1QOgD6vmt93yN2
2sCBJd8dBgBKJYFC0QbeaC9TWRV7l7FBqzK/55Q/eVeaazxlTIcV8H5RZOiz3rXV/euNYVeLsc0q
AWXyBXKv3fTvk50d8Rk1VXqh/wUTKR9eVgtLbs66Y7zueR/NkPjjHGuNK8d0jaq+4QhkicPFVv0+
1Tg18VFsX3VTbJPfV8tTHiPLfBgg6zurnyg7pkg9S0rvHhAdOCvRApXa3q87MyNJMbJLxZ8QTGKa
bA29VlpgusxNX5Z78A1ZbmyLZu2Ya22wDTv6X6oiiOFxP9k1yoZI27ewFTFyP5956ejBP2gdm5GY
HdttmrU1Pq/fC2lRAXt3O/JTFTiwWNWO1fGPc/QJWcd95WB68yV8+0pU8S4I/0FYVyr6BDzwkLUE
NV/LFwgf3uyd0RYQkZSL1wtYsseE6SlyuiYPZfNFMqvFmfnsaib6Tw4t14Xc06wmel0a1zINgiUC
ztl7fC39YqR6hmhcLg0pxHbvp8G/9Tz3qhYQqr0jXc2Kpk0oTUcTw7JODvhHuZrRTBluoRUXNw6l
25xXUV6j8xaNe217Ox95MD8t038IHEVIX2dxAGPNRbwArBkoFfOlBV9c/P9qVs3TdIEnBYRCXjrZ
H1O09a0r4GbtdIMWWfYujDoQ5gD7UqNoxSyd18fdQH5n7PGCTHJDzMIwkIFVAYSVERMhjhxAxHwa
mhb4cpzaPbuvGjUzLJesTRjF/y7WoRWGGWY8/nFqjb3RA/PZK0IS1VSjUevhMJVr/JhGIljj7dC/
KC+YQcHiF/uIAqeiuhbXa80Xw+pVt2Lo8NRjqc+BdFX34SgdviIJhRTIC660dCFmtHStTg8syUbW
/tsDdW6WkAK8MdofjLeHXAYCkJCMO7UzZ5CbZMOePGHewRnTGTnuaTZpx4Uv4fRkgLUjtx9NvZa5
DYQ0VG8S1hvbS281L8CUHmB0/Fbqdb6DAXlDPTJb1h1fM9J6RPibdUMCgGY3MvaDBlJ32Y7Q/as5
Wklk7dIfbxiIsPvH1eW9gkPXStXjofMIkMTVFSD7rHeDjUN4/SHXq/GSeaFAQtJrsfxWynro+0TW
6otGDgddqXUO2pXpcXXMc3128oQkvA5HCDFkAhhEqc6GdjWcNvWa6tdIZPmPU7VLD5NoM8jthy+5
W4nSm/EjgO8/9uaYLkGQM4QW5eVC+QiavOn1mlfK3GIYxeKLYWE2miCVh6c/kISfBV6ByNiFXt5w
mi1EGo9+f3tQieFPFUCAtSBEEgE9R8RcI7k2Qq56+VmxOkZd7x0j1riAEOed6tNsyqxnP/ndNwk4
KQHK+pFrobH/61frsW/vl8zHdZcXYHfwSW1sDIrAda5J8tccBw+g6F3srVZWU7cR2a2RPTbcpElB
foosiwdDX3PMTS41mqy4yyGcwqkaJpvgQ4f6f6b9KYM3NvthHUX//tZSDFu8d/ye6PyBqodJXzMJ
KCicspB876GT6NhNWQQ2Hf/by+cC8pEaGbTOiLeIaCtbEHSskaUfOVtoPEbaZDnUvKP0AvBEvaGG
TJOLXrhDyo9BjPHq4Q8iqEZlXaEcKVX6ugE2acTyqXoGDWmLF22zA4/2h2mMGfeG4uVxN7TiYMjp
gywBoflMJv/oP9Wo7cZcnjY+QdsE8VudAlc8q/0nAtzqxBdIMyYXIY0jCoPj+bhRvQjrBsTjDioc
x49v9YmHWadvIdrLs6SD5SeMVXF6f0fP+N6BVdC+aQtuqiR7soX2E0O29dQkZxT0Gm7fxLQC6iI7
XQ9Q/sfoPCXmwfwhxG0ZvY3wkwCeZItc5sMyvrxvrIvRFzLMDuEX8b653ljMpLWQPjjXLj3SGOjZ
tBy0ybNAnHBr5/fo6OkeD7yUKt3NNwlH7uhxBpQosfhL/sYV6KL8NJWYhcLg7uoOn+B9xFxHvkwE
DScQ5YoMcUM9WT0PQEPAuoUs6QqcU/FrK3BnTDjy0z6OEH7cHK+1jFVvjyCPCmZNP2qjur0+gMQi
tPcQtslIYq5+thaR98UaRgoWCSfeeZlIqE11q+jkqpmZpNiEDhMkIMb0XWXm0f9Z4Q92r/Gf9u2O
2SYVV9EX5710DV6R/O611NNl7LOJ+7VWOY41YPtE7ASMujH0dfEiqwbOckVz1rAUiO3JrY8Nz5Nx
8ZUrYd1RW0WoBjXm1D32bIWonqnM7ziy3J/BTv9KD4M0iZkMvzElmqZC+plm0EA97MfHMsYLBkSr
7nfUPME2vUthAbr1M28QmNUkONatN++5BgnClF+qZacvPLzh2HPu+BhvcbQC3G0GVvlQy4iHwMm2
b3x5MrZjq8oHDR0cMO3RBMBhXOMktj8d2cY1uLUKnFypRKl+DE2AL2MFa1WL+6pYRQHn2kE1We0J
g/z/LYiiNdARm1OCB0a5ER/rj0dlpss85kv+bl2+FCu6NyjIPkCcwguow56vmPJlmUdn3NCSXfKG
HJQmalfH+7k2WX7JsB7UCcLe1IJlU3PvkSZPowvQ54jVJGFn2XQpkQV5RbrsnMLAhNpT+8phDeZs
5+OslQ/Fo0A7BtaflyTvtDjJ9bCUA0CqUNsBiGmRzcufHjz64f29XxxoCEBWFiEjXqt844bBLd57
GA/pCCLwVKU2w3TuErEYCTAF4ViA/TxjfkAoiFnrHV0LDSAvxi+Yq11Z2++qVfzQSBUhZc5MoQTl
HRRu11ZGmhgEagXXJinEBBAac0TqO2q5RvLTYbHv5U7AYgR1UJER5+bYYk3zRjgBjS3Mn9ybVdgo
yIH9FIpM/AjR4tsurgq1bSwCJ+ghwX1fk6o+iN4rq1L+ki/vPVqKvbqgKmPyz83Ds91OU4QQZbwA
6EH9e7tH14qZv3u8NrOO9NH5/XoKD6CXAQ0opQWTUR08Z/WrVwcNl2TrOE2ZwmY7PxKACy8jAhNq
Bb1QXjPE25cJFvYPyfNCsleWjgQLqMbMfGAI//UOA8rhhm4P4++WFpfzfwkpYzQRURTiyrHizYmA
Rc27xnwIauoIzCJM8m/WMTExXo3q2XddveNpjiu4SEFVHntdg3IasMBjkwmfkn1RNWn5FAxHGy4S
xskFufoCcwFFOqI2b3tNhHImqrninVFH1S8Ij/qH8uO6LTyhiWtws7bU8hzBeLzHbE/lNvT1iFhV
j3ABL68E3SjeHHww1FVd72QbUHA9kGsFl2GBAgaEPv1Pg+3FhEJERxAKYRR1A1R2ibf6wkt4nGtr
Mt2FfIqSALlrqGwRwIwaD0hWkuTubFubK3Lywm5Fr3dHiqSN2Q6Z4Bq4/7kxzLBdkimBoXecIrx4
xWM5Dmq1UsxDWIktvct5ZiRDh2X/kBVXGsmMbmZnhi27dZoqHzOb1AZm8HHRhIlTU7Nvovydf4kN
19cV6N0bqVwvi6aaSljnsoLeyhJFJ5YeiPjNtAK2N1R2Twf/irEthsuVimkqfZiJ05ALQGB620kO
w3hyLy4ScPmrlAE4iOp/aY6g4YKiV0q5KMwtIxYE/PYfJo5AZPLgj0nmY7vDv7MSnzLQGMXHftRi
W2wWyjpuTLYXYli1TMDzD1UyLUEXTkP/kA8fbs5PaQ9pkU1qxoIEjTF/gkloy+4NHq4JdtPnMtyC
H8hlQIW2C/i+c8pgHKh7OP0wDovgm6z80U3uK0e4uhK3xJ5pBDE50AFvhfmKp5DzYcPCX+q53FL7
e48U9k3bj5Ykn0dNisNpuiMXfe0/X95mxA4DW91bmiXshnTQpzhrEqYaxD7dZaHSFXJJIbrYhm/a
FlgZUj0Y3CC3Wft6Sx4kOJzDfVLHXGBczCyY6lNSD4KI1+zEWQWj3it+ymMlF4DQXXRGer5Iqggz
zNn3pOGMvpc1WVSU/HAWzMpCHxJb4gApQnM95imzpKlDaTa6wBzUbCz7Jdnt1uzsdVTMSX60Jih5
ROoPLGz9IgRpqDV/BUDaqNiDV0lq+2e9ByXRTXcjOpAGTlQVfJxhuJIPE5ZVibVloef4spJdj9Mx
q/pe3/pGbZZpSLP6JvYMKtVK6qhdBp2M7wXqWELhF6/CiAPBwroYWI/RIx6VSitP1JknbrG/FDbb
JO1qp5QHNFwvAMkdRWc5DcUaO7DDWLlzOywJRUGbDVb85gYO4ckLvUctsFOb8GGKSk++AhtC0nqS
Q4Jp9hApaEp/Cr5NDvVfuzY7UwfSI4R8hs9ZYELts9lxqdJKFr0MhIuPacwz57l/Ffg9No8eb5UA
n5kNi/0Z8HwhPkaY2p3RcT1wKsOtiwWOM/hTy52n+JjxWom1+7qn2h+HQsIwlcMp7IUDC/hv2gWm
Ir6JD+khZEhPz3sJR0y/85RFj+k7RMfeX1NIDrXDFWE73yXF9uLSv2br7oLTi+HcoV5KD9rhY6AL
t/zGBFCIq8+xciHJ4RfFaEtpRH3pgg6iYR5xYV+CNXrZHC/NokqBJdtCqUpWmE15O1pgGRMgTgQO
jwUVxC5hefc52qwQ+9NyTLO7Sb/6Fmj+yULa3QRPa0tA370Zx7DQ5PmWzUh89n2/7qQubtBeFNeJ
bjPk++O4od+enRcztx3bv3aKgCMXK4BOkylPKHcFaxTrhvpOIVfKjungI/n+6NqlEd5fT47kMq6a
mNGrz42VoyMKYgiCYm5Oit/parMBIVNIRfh6qAlJfYFsQVpXDz1WjTGPgV6Oqd8lKSecjUrX3ojC
T9Ogfcoq0HjfLeYirWhig6biUhIgMHoNVcPKxw80ffBRxhyRGAmhTiQHnI59ZljMmnnjkgA+APj7
SQ3gpdZM3s7F+6Cn7v5AwUjh8eHq6q+WA/WwhlOuvfGI3RBAoo54i4htNoJmBP+5g0ZXJ6kj4ZRs
uJ7yLWumusr7ePINzsTkpilnDfTMEpWn3zzlLJI4wCh6dtKk+s57nRIKBtZ05hYjuQs6YpNFmfP3
KIRcrvf2nEEHlBzHDonUuu+SDWpX2+jFaiafkw/slKEMnb3XAvJU6HTkSBckrccCRBBqcYgc5UZS
zGCdLEFssalxTGLz7YwsW6kgSSAXtRiUfFbeMURyhkvxV957PdLnNN8sO/q2z6ZHzEIz3jdxDT4P
Q/iHhcMIIM/5vX6frSqVNKbFwHGxIxOW0Upo9nSs81jiLr2A8kZqx6D08hIeG9PONTKwHswsl047
N+4uwPcf1oeio6mRUgazY4afFrFruZw/V8H+LcYtTTTylNJQ/AMPR80fGGyboTBAO3baIF3bE0Au
sLFHPTeByy9eQZK53mD2e5egkMrKzEsnUimoNsj8kjkg742LoGZbiXRazrf1+d1bFOOWh2K30MJa
yiLJh2n6fIlAb052iPXeIWpHASkuKlWQ3OfSnKuE+w3TzIfsOqyqOM7f/Bcgm7B0mtV/LWGSkb3J
bdssLq/hkhqBmWpFiHfwKSE+XQHRvGqwnZ3jrDxMe8T1brFW7bKUjH/H3vkJrOdYcHGJcKA7WiZp
uZNv5vFbODctdcwyFkOljJw39dZxEynclu2QiuoVeNT1TajS37DCCvSP0MJfjOpVknVG0GeDUmzJ
vC1MJ7BtatiGcYkShMGSLcuOJJlE2VFljoKD37dsjx7GFwboA0eZUZihmlHAbrulL10KeaUi0IpA
w9g566hMldUTtR4GYeTgPqdzfswPmgyPLH+7zDr/zHo01aoi9NMHh4XnreM1H68KV7/lS6MhcJSk
mCjgBwLfM0hl1I3Wb51pYGrtDYOSgIxXnLQtQH2ASd/XsyXKG54eOmrgENA80RZd4v20mMeXutxS
12NAxJ2kUqUgBb7J/zufe0VTD+/OQUHjdt4rElUW5ysUixfahPXjetvddoGXAXE0xLUh+ga490Z9
8aIMUHEgOcN2bLOVrdkA44E2PkP0jTSqb+p0F2rFo73oFygjMdMLmUpQ17DrxjGBrmAbHKF2z4gN
qm1axzHIbKAXl1rPj06UQ0AtQiUdNOuWcvhFl4rBjKUgKZyIuyFuIP35aRZmmCmhegVPtK6pb8DG
e4WwIvIvdv/NnVjOCx6etCzgVmXsHRttvN1+No5gJrTX7SRuc0OdnJhmuf3gqr0HeJN743nhHEXC
aaaZZyjr+aJK28yX0w3x9e3OGZgeD3LXAYQMTm5/Ob93p0FKvwZxUPq/B3kuIVQKPT0BiIdvidoX
N8dqKlFufO2rn99LApxcm3gljMSg6kLFy8v86tnSB+tY71s1FM6o/PwGMibccfFd5Gvg6JRTUHut
IFVyXBq76Fl45OOQIMdnhxab1Z+7rlRQpHmrFvpsXzK8h/zyr6cocLagXsXUqtjQsSaW3pFiIpdr
elbmoyIG4z1gXMZFHE1Z8Mnt3dkWSnqDM8wokqEQfu0K+lnwm6xHSwdTu5q3k+z62xau3S/x8s7k
pLGEUvNzi0gwo2GKF4pXZHPBiv5FIUtpEdf5PzFw6Ke1xJkVwucCnAs2rKZAbJ9xl28p+OY8ysii
dDw0PsNlR5I658ft/AVjssH8E9TiWcw3SvXQ3dJ0Y0YkytjPWiLlC7NdkqyKdYfjVrSwcrYSDdKV
4u614ngJgPV4gqu97K2mH7kZXkqUeMImv4Dk+GQI1+4O2Yh3kTMHe8lKaji7o26UbYP0TBXGsz1K
0PdTkFhkR9DFGuAdEk77HnKElYbKnYGjVbpfiiC6X8TFB2Ot4hGpNLyUN+Ne022wIycdi4MQiOJz
niu8dye6kyNWWwSMti5RQ0cxhwD8fwPdkSQ+BQM37/CL/oKSMT8YmlHZN1QciHa0WVcmI/PfLQgd
D9uk0wfFxydEZsBBrZoEKc4JQtcp+cdWkSvNyBhyqeAk4L/H10/Pz+G3QDIugGHEtWJozeYkXk2m
0e1H1bR5ppCyGigQquPkd41GhOZLDxF6nM1nMzsunueHQ/gY9SfMrcG3VZQg6wKk9j6EV+Oce2oG
/OwcxBMcNE9GeqIcZjMtO6b81RkEjREo/uJ3E/aUZA8EQTxB1X1UwrxMJ24iArYukuqpj7YAFlI1
iFCZuz1Nle7/It9LFfS4yuws1QFcplDBAvjC8ESouwJ3Akou2kuWIikavOmwndAoL1N54x2yTo+7
4vljMQOZu1nARj66wKgugkMNBlTsfrY8RJhOEuYjDEKRwhcUqWXgKl//CiXKUoOoHU6cshU6r3A1
S/ZieGhgwEV7q2vGYdKEnf9tBLSDQzLqxJlqPornxNOBWssm0qxw2iUoa4PIYezZmN5Q5k+U2Uzp
zwqh4RiDjruJDRdjLqcw3ryQE0aLHXgY58ENBCz+17JtMFAIVZ5dJeJWdsr5RUtWampfddT2tkFU
fFMSKICOt33qcrMyQ/Xphn/TUX7RRwlubMS1PG5TsR0WYEirNqSGfedkKumMKMbWPvcpn2KMuWfD
AnA9Fhm56/0r9mffK7LJEqil/4uw2dQJssOssxSPws0s9l8BXMZ8eoav9E6bUEEb/jnNZsWQg+LD
o0ZhoziIVnXVD0bou4+VRCgVEqPcFF4UYuT3jWM4LvMCM2QnInERY/dggDw5iXsYjynkNJ+pAYyH
7KZ5Yg9VWzAj2ifsCo/dxIOt8L6g8a2bO+5Db4H4Ck5RW+QsjQEdwXyyitDLxUHQKA6Xn/tCGgf9
IS4/mMDBp0bMuLRpCwl+Dg7qw6YMFAPoy1LEF1SImMfezDcyEnWrJ1oPD+pnAVUczxqiOU3OPVRm
jQePP+5BmJM7ekbOmYRquzHRza4dSn8edX4dQxNO/hHa0DXjVjwfbH+a+948htM8T7tnXdroCii8
y3NkGAJJLikFpq/R1inZysLQNYhl030UhiEI21d3NWUY6bgso2L4G/ID5V823RPfKy0wWEuAYUlr
DESKlhQDalkQxyoA3lexzc0THWYfJlawTlWip1Xr9pDhv66Jc/pDrEkWDz1nspBiT3mAXBEEbAsP
+5GSohaqHEeoJgWZF4IVtbziKNq1HQXpst7BWVTrv9DOK+ZCwpeBoOt/qwqaH5zLykCTxr8rjhXb
FnXef8mlLnxQcEwAyIK4r5NzeFJwv2gkP2LY3Xn/pfSzGiKH3/zh4Df7oqicr7tXFXkTpTczN9xC
ZbQj+WH0WXLKI1Rvmnh0/tRSKtDK5XuZwZxe+WdXVSGQuDZ1vAOKMzUr/Z7HnCcC2CJUz+OeoscJ
6BqjweIyNKhYjOAhioBMcuSktwRQR/oMpxEaqhER5AaVo7zx1Sk+baglFxsKv3VkCYKQv1pE7wXa
FGS97k1q62eJpa7RbIueBNzcRgKYAcWCcwmWwIYf5E3OWKIjSbTD8jx4XMKmJUt6sD+va3MxlrY3
Wr3/OHIx5FSvrNS7VJxTVclrhaEqm4lzfxPkcEkgmIMuhTTGcTQkvRuQZ4zeqpJABlXZ5Kbf4ynz
HGXk0uduwLijXrFKtubOqZNi+Y0lqFdfAImjJa8BQBA/3uloqI8y4l1MXZlTICRiPCcy/IxqeGup
UbooaKEIkoFdUBFpQMteVrHYKMTPLwJzki2q+TXoeSebiIhUfjjU82fcDjsImxZhTD4bUMKYou3u
CqjUfDO0trJl1zvs91tcs8vT5b9lx1Lz6WQNaQBjZQVj+mKAcnoPAYiFVESJcIhxaFfNQmFvfcpf
mL8jSAsIgd1KeiZr8BYarZdrQrbGMONOaaR9kbCu83AiTyQvumMmp2n8sbA9SuKgImqePxkSDhlU
GHC6v00nPJz8CXWSS6CqgW/VZoDsHbpUPRlwvjKn1qjDLkzslvOJUeHPhSK8Bf2yuwyuENjBvQ6v
tHRU6XWYmH//A3q5Pu5c1oAkvDbmdI8+j0wnTTwDk1ip6hCOqrv2+o5JsAp331PzSNtvtLp7co/8
3sKwSvI8lXg5MyB5LuXRxZCi28N49vfq10TijG3vAYLRK3sAgHQ4pURsMZGFQbCBzyQv8fxT+rwx
ZDkpBIRqU5C0HiOlNQHU9nyYAQTCKpy1OIj8CUlFf3D/tHn1TAlLS8LP7QuqaduntECE2StzFj1q
NXHgCipWGvEhsNLe3eO3XsMNscvDUyVn0YNjnKm9W8Tg4GDiAhzkU85jKmlI/87DBCehETPt9jD4
bht84ME+rXmR9Qk+Gr+rUaF/p3av7nyGKKX/7739NqVj6/zRJBusDeeJZrbeaQBh9dl/s9T/a7sk
gxg155QwrC/toXzjP1lce8/1/r08So9kHYnbHMIyjmPccCu4wwXXI7KKBPcBccrVqX7yE+aEkPJP
IZSomxeoC0AOa2dmTKDUO9fn07JxFJ5+k70oJ4j5zinHg8qPzZFbsS+hfQychmu0Sed8ZL+VF06X
+Cm95r6EEZ1ekbTG7QYtQi3fiI54TGC0yW7vQNWLB43I7TwNgryY5TvNpMqvr70haOInr4Nly7ff
5NLECmIIRhMaFzEW0ObAIixLUMV3KgE35Te8s8RJl6jsfP4zxfXg3DvvHUTy+SSHDuLO4lEYPxWU
rFE84WzSz6DspKETtbZonvGItGLZ4aGPwZV/UavxLb5GPPGIu1gWlwz+RslifxECdldr1XkPiqbW
inwbm96ay6cjmniycPK1sojED2quCIQcfD2pLh356hcgwmx7RqABQ5zFcFCqKvbAAlEsRUit1h1o
FpMr2KAwnQ2120defXhB4vG8n56m9BarVpePb3O1X6V4O7ZQTKRoJMFoxrO1Gn2pPnZaGTJcBjnl
m5R/n15FWxIiUcQrYbNbxlXo73RimVP3S12mD13/22BQSUdxOodRXlh7ZyIFdfQ3gCvHFTZ3KQqh
jH7m2LOXJPz8nB3vEMvbB8dwkmkmWho+sRY51oQInjPttk0g6WhD8VkGvyFsYVVYAfIy/dv10bY4
Vi96FR0q4cLIb5awmLPMnmKrj4C/fZlNwauvtZwgiBAkfe7MJBevLMKMA0cyBNgqbRKht2Yucd/r
I40hFLnfbK9tJkbTLnrugQyR3blnOaUmJYYfFd8fWpHMaTvwyQpAYgWT76EDu/XdNjrf3tasncbD
gb7dEE5MSQ/e+h819sqHnlEEGBRt10+lGgEfBdo9PY3526FUHo5OlNT5mIlTOKX7kFknhXVCia3d
JUiTdE9a6Fxk6wOBYk/lLkYFrGeG9qtFwxk50/vn4B6NgVDP8eS00RcG9vsPMxzKxzeZl7390Isw
qj976nGfTGGd28QY2G8my7Oox3sXP3VpTwoMOgXbqpwkA/QEkZ1DOocHj12ePtAtuvEt6fZQaXEJ
Gfp2dAdGsTstbTt4+MQZgB7dTRjY2jyGvfJWXCF/Jo9uFseqbcXUC5D77+XHt3ua61d2K2UUf2dI
nUc132W8pYEQcgugHy3OXeWOZJoOide92Td8b+BaHBPSkvWhOF3p7OSsoenubtjzqSMcQ1DQNoI1
sGD5dVwpxbsKouvaQnIrq0RlxaQ6683rXknW/uQEeG6NnzUiqkEY+KMISzcBhLnhF3I3bqw+WDhV
9nbVL+phJGHKvctxepkvQ/w/CBfRgtgUUCH61eXQ3HCElmjy7RiFpruuDAkrHcD0jmbDs1R4tRAK
haEaNpSETatPhK+E4YEQQAgF806g9FhoiWNijLAe2O8Ivmxh0yzFZVGsn2EOQb3ej7LtvdMimAOh
ja5b5Za32uVZon3pOHxzk7Ho4DHEtjIK7B0MHL5+Rp1lZadOAHkWLv6uOGOrVAtAtfEf/Br/KTfo
BYrryxAr01muUSbwwkZ3z8DSnO/pJ96uyhvSE5kPVi2IHPtmCFw7pMzs2otB6qHjN10aMB5/ND4t
Lc6tr3r/Y9pHrGLfuo2o5t0EX2Wk/rJPpSIE9CadJUER5Z1/zICyf77cCkTS1xXQIvsdUKxe97cF
ClXPKuIjlyjSyB23hPYc7Po1FuTOuUVIc+SnnKrFNJcrOsFlZP+BrMoALTbURDVmfkjRosM6FUem
e+VTrfdkBQkqVU3ggVfMmZ1vdYEMyLR10oyqy7BG+WCHmTZxzRVzBAIGXYgL2c5m0gN2To99lf5z
+nq5i1h2LKSe6bzfHUNjHVE2/RmAmrfw5McEnxu4OwWpSkgGWY1bVBfeRHGsUa3pUkF0Y8rK06Gd
lFf+Idt5oCJMNH5QtGKKODfqoAJ7Pr1Y1OUVRrd+xRmVt33kjsm8GZcVPj+uei74TyHP/afrY2ln
bpJHkv9ohXDajOHuo3fOWrEc4h4wArvvj1OKydhMPvYiEC95899Zw4Lpy9Iaer+8tp52Mok7zbZw
3QVNc1B7UWzJU2mdRKAvGfBXrskUxKG8NuQx1hdic6qokIHMMTkXBqM+ts94mRO933QMQI/Pu5TO
e81xXP10QSYqup1xMX5w0HsenazpEQYdKxQIOek2TBUEBCRF9YrWXqWr5S7+QBq29Hqwz5nXwmNE
XUi54ZO7XQE+ArvnFKRAxJRmFHFiy9mzdupcbAe795OuHf0XDbMtRACUT+I7NIsWd6XIU9FszIQU
ebBIVB5fG+d+ihRP1pWDLVRsUUwsrsgQRnmdodcGMkI8tAccMXto02/+w2nEVJq6joNVH5ND12R6
82sfZrFcqLusV91oWfnN1tPlf436x76aOxrUdSR5VH9CNYICh4N9FZdC6NmAxoywCmdtReYczvli
1xjMLjJ9RfpyF5CATnvisGkHGvB/K1KKhIEb4k/APrE6rXTnEfZGdCWDJsmbldc3IUwpy+swy4hO
FDMWy+1CJsvvKzQWPYOSnEqiCpcSdnf+qmBvCPZMcq2DfJwQrJw7Sq19XtP9y8PPSkdRtaPKWxXc
6U2Vy7dOUjzX2UBOm/AJDzThPMYA/BMszd8qZjoJnmecSMylptychqA2RIGqiJxldUn0F7oeYLMY
IClSPmfQYdjE2Q5/uzI1zXP+Ok+PeIGihjwa0+gzBUe77ZqjBv4ZlhGOdy9bjZRKWQTmE1fVa3NH
SqUYZ6MRFLXNRWficblio7VqV0KKqsUYWUvajMxp+1K4DfQ8fL6hy4e9wJUvTI62X8fxXq+oJxWE
7XkIBzyckFx480OrKYcP5gqMO3ocP9/EhBoeF+oR24Tv3epiATxUfwfWZvqAlyvbM9giW0mkelXD
UXKgni5Twsc+hSy9vQTUGNcXW2gqXYE4WKa+PljcpM/x/z1/V7wfuPHWNFygsi0ygqEUcQVBMmzf
LjI2u1EXJ3GveT4BkJi8fbifXOZCwb7Hhe3npaiJrjxUQtjyswJf9c5qZp2sNPdaVSkwy5CoZUat
f4qP8uTj8E+snkhsL9+A6GqElCCxU6LbIvvCd7H0ZXv4m5k/WDhljQGkMgB508F68DDJmWYNp9UC
OU/S6+xECi+cxn90xJwichi6Epgm7oB5XhhGYVSPcaCzcYYFBJeRVDLMACVHXD0vNnviD3o0I2YO
w3WYY0NhrFPEvPF5lRx2m+lcwK8c9opxQ02nuvkaO0mdDB2BYOVvM7Za0ripIyuzHeAyw8LnXJ1T
I7n1soI6ZHwke4gYfg9ossq3Y2KuFt1EOq8jfrQL+sFHjnk8kcyjVQLbxOpK2wRR88S1PFa8qGVK
4HVKYIA+3ajvDFMGhNK7z/LXcBvFtKP/vWxRNrBY3dwyKvqXIrNzBdOiH9saS58KORdupszvXAmj
JO8PSlPTfbQ74GrBvGImksDcs21O+c+qBo7WsmUfJ9/6Hyx1WEsa65HuU3DDYaGQHtrNfNFtrp+e
YiihOVFzSkmh6/XSQFxAKfqz6NGRHMRf57fQPmrqW2dAkjstO9X9jNBx8tKmQELOW15bza5reRCX
Y9B9BK82PNW0PtT7T5iIzpTGRVlLmNFkKCHhO/Vp/zCgPrSMcI2Rdowef/I4QZVaVp/jUyWt60f/
TA92mYSFip/yvVLjsvdylBrbFpW9S07bGeYr7KDmVUKRrzmV3q85zp2A/7Umk5254wTBad+5j8N8
AbJLW6v2ZEITKDjcC28LMqJl2fDQiPxwLvkE8lmmiUWfJZCPZHDoEnQ3DDGYnEyvildQsQFDzKh0
DFY5BQO0S9ciCQaacmqKF8L9VRTEXyxsHvP/gth7mvCPillMFcKhb9E38B6otdzIPsWEpYW9aRSW
A8aqthpwg/FbZTvvzudjywY85aI3cyKlogN0hX7FMgA2W5syPRUbrJZL19btcUf0/naZXGhuEy/F
Wv58AwskCV4u1Mjl4BJTfG+kvcGwH94QMINpQmlCOHIetuQRo44J9Tl/uPXhkz/ub36TAN/I07aT
Qdrv7DgoorCiIfLqfRlKHQOrZ0PiOudsETjJxBHrcFMNsTmd5KgH75yNVUDZHCbCmE+P2S+aBcsk
33yg+0hn/7ODnfAoXXTQUyvfKcVO9ha/ybgbWw3Y2B2X7LJroWwlRmYNY5mK2gTWPL2iPd8mpd1J
0nnHJsxu7eeDZRANUzeldpTqKQcNLN99+RroLBpOzM6SjVQVwkq81Brfao/n4jFUGRuKe+wT6OXx
/IxhO6ZILKnMguG+d5Awvp1efSwq6RUPssw2KCzyWdiIkWQuTyeRrt+htVzzNkG3UKf6dfNqSjEe
8rjih/GBu1+5iOZmAMlGSKZAKsHKleMb05d5lTK38WGIZeOSFvyclsBpWK/cUVQ5VBhvT5L2Y4d+
JCqZ/kM8po9X94v8VnOpi1zjq+amLHCD7X89J87HYVALwOSxUJ4SmhAlU91i3cJMuCa2fu6PIeiG
WKgnGk2Y7iPNKVoo56jtbGCr9XGlrVKRKPNQmAv72PRpO5EZmSEJr2tdRbjP60tmPMZSL8ddURI4
8Z0Dhl2P+45FbWFTja9CLckTe5JJ0mQkeWWDSeAJXpH8haJCzDy1Tf/5y5Aq2uEhBj9Mq6v/h/Y2
h0fgz3MUUXouxN6vlDG4oN/kfWplVUsD0aOS0ox5rGfRZ10r9iBmDnuv9pL1Gq1DlVgp+QX2HAYT
Gr4JoLRzDr+3uw2Vz7709T9Q/Q3HsOcR/p7UP4E/TlMQNchUtih+xuDbZ7cyg8nCpRk/Xcqoowgf
Pt6LYpKbPX6IzYS4rraGs4KVZ5er075t914o6yw4FQEkISzXXMrUnaxYL8tlLAKItOGZDBNycIbe
0oL/IXCQpKLW6c/RX52WM8cIhzqSNep3dUsNezghqxNu+bYTU8UXAVYMahGiiXIaJ3XN/TUaUwLP
siZ2pLTrxpm/BCFT+YfnJ8hlif0w/rjETCJDoeyxCZFzaZguZOJQ/hplP3Vb3MJfkocCjnEwZm8i
h0w9haKv8vn9M9ZtlM0YWDKQYP7RylB4WXrRvHXMi19Zk4k6/gRdlB35BHa2+kxwqFOMt1r3lws1
9u/Sn9vYhw/T7D8lKYFDfCh0y/XueiE2LNpSONtxVIr9z3UIhBgaOLGhPkDHaunMALNGy1FjzImM
aZWhXKGvTt7IPhMAinCHoQwichnwFrjluhFSqfdGsgcxNcSs+zMHBq6DHT7TKTYn9kEMHmypZECb
Rf/ri1pAUgZQvmJw8Y4SSNciRYJGfzThvAMzHf592MmSAJ9dzFdCAd/IJpHWxZ54z1YuFLhyDbwz
ruH2SYwuyzUfrj/4qyDgEcyI/xh8m0u3sFkYN3vDxJLD/pBdpSDIThStZDAkFGVpWT2Qshi56n9V
2qsRhFB7dgPMfR4LPfus5egNYs3qqFGwgOWFQJ8BWL6SEs+0jzvwGzlLWdtVcm4x7DRU9dehHUTB
5HOSAzjSRVSarvzaGaGonrRuLqE5OutgaA5OwotaI4XnZd3oDh7Uo+y32ekArHdA9InkpqXHEtKs
LNg4Pz3U5HTO68SSjKnn7kApELXYIlZvMqd/MxMbaGINRcHR+OT/spIbZ6n1Hzr/th40UtJmNAns
T+cWXpjc3Kx1CtPDvLQLv4PrmXuN7CMZMHkGyCy8oC4tpd+Tp0QTthgMr3XGJrcuTqzYUwTx4ep/
vjhWV/2MzKMOdmehNpTm0eSVjSJk6zbRnQYkKwUWuj3poxCfstb1EDQSVcrnC7gTIUN+l9XN0rs0
LJPTSIa/0FBPoaak/npJgWUMRsIwxE4mEbqut/XShoeQ6WOXSHgK5neXazBROr+Ia53FNPNrH0Mg
ro5UzWynGGWGCU0lGyvTE4z+pbTBkXyoGIw81iacqHpGHssUml6imx2sWWRPUgY4+TIQ7ziz842Q
tluMNa0zlRod746hAEN0MGWGGgNPCjVpgl5iHaJEPC2Iv668gYuwsv/tlnnH8KJ2mI5HPxDVqGa8
wz6gku+HnLHSzUgib0SSaoluSLqHHeIUca+XVidnAJNbnAA1JX6qqC+JC4HEJnvUJQ7WY6I5XoBf
KbIctsYA9WyLec6wQlVUyYQPX7h26GEvgZihor7qYwpHdM448aQCqjFM7Nx08u8/qL/Zh4ojGAMF
xukEzZr5mqocMTZAlxO7ZVDCPJMWX/gsPQk9akwlOJWuZnVYf70H6gfb0ADDLbfF8DA+NNbaI9Oy
nBEmyYPwrok0DTcFu5u+XdWJ9pnVMbDG144psgvgBcO4+berjXS5MgG8Ha+segOBPUr8sJJhKUjt
hXWngR9cD3LlVdz7WhwcizMz1x4mg5HLXfliMcGZuNS1CKRzrOhCpnoWpiKughThBSgQcMBl7X9M
ugnOqcFWdv5Imr97huSi468vtVP5giz0doiBcOmTR+wf83VlB0DJ8zJwGJsnMMGHhDfr88mxpNOW
elgv3yEIoKQCfimQlwNFhLMiGcKPdlbSN4PMEC7sjk0svf8qV7xEGOIXE8WPfwyI21M50ZN8KBo8
DkOnjpinFoYez1XwdAcnC8/DT1VPchIJj0ls1WQs9F1cgJKbyVgWGu3VSEjNXGoXumvFPmFf9Kg3
18HcqGNPFxUyUAwkpuuVRHEEWtfL1gj4USpEkIw6+Y1ziLU+Pv1TKvy6PvDE5U1bYW7wgfAYTXW4
9ZwH1g2RoBd6ywIyaS5AoBnHM7H4+AGE7a1VcZtjNdEs3twlZXc/xaMKODEM5BaehuuPoT8oEAmN
Kz6F/B8PSDSbWwvmoiXvylY3KvfvqCqi5ugYnP1wvbuKJi40iSmjF/ebP0Jzi2k75CcqjJjCbi+k
6mxaw3ynNXzBB54raja4FS1H+hIpB5mHCFmZk8gfijC2J0HlDlG6MrTmbQbiNKaAzaw/0LEUsBZN
4fZOZHz5Eb5QOyLmK/bCYeDG5UCEoRof0QOXgCpcwEAaUnhRVL/Mu+hQtTuqfrjdp8CGNUdFJe/l
QgtYPXTFp5WvupCKCwEoJ2oS3Q+sGN+FHnnV6UnrMp2aUXwIzQYX3mVjo6kiDq2EL4YQYm7nHYjZ
vDm4nkmyFSx/SL2pdSW/HWdqrj8EQGDeRtrYLmOh7t/XBDDmKOhwClI+znBSSe/jJTrSMH9zlq2+
1JpicwcdN38Ko72hN6KvOL6JcOi8ZjLkNZbuYTJ8q11JuKKay/AGBMstjzq5kxkd2Q1vScbOSEVg
ZzfN2MIqRaRKWsdOMqxT78WQo4l6A7NEwIIpmm3HDL8McQoaLEPN9XjrVTARvb4JCiVG3BxUrk8r
WSy/Z9Nu7JL4KON41OG3sRl/L8bhV+rk+SR1jGLUZxwgTD/MXUB6gwi49+K9zb4eWMwVWOTnSvK4
fslPCRirbfXHrk9OLy/j3cMcmnztOj6LeqKOY/f4dqqqSh5stQCGxwEWB/mA0LOFXqQOJxg49ehN
OvafAEvpZLMZ2yqvRWlEP328QvUQTs+o8Hbcyl3Em8eYovDjJ+RBz37k8vzuoflFSxH4hT8vBk25
xOi/iJ9Zm2a/S+Ljv6pOEyzBeHdLQPat8MomeOhOVJL+FWYk5xHeed/zc1Cr+a1wVjiJA34AetV3
+csBX+f8wO5HwlbEULZyCg6+3Um6pT3jq/FU12HM152RfNpJMyFWComDp71MvIp9Em18drLoRTBP
wURzs/OKe2vC7MbQRFU6agZcpzeW/X73B1VXd0m9t8ASCDtvY1pEVSnyDWOBcFv+Bc+rC7DGIUYJ
Mhz1AdDWCvZRMOIIAR4DrIUv01zqAF0suUO4elgRp+gWO56OSkL4a/12mJ4UlFVn2SSr7i48+/Eb
q9GSSsMb2b0oYsasl9wtzj6kyJtaOc99Hf3+QTUgtXe85X7JDKCwLAmWDQTLxisBNsBTPDnU99qT
kDLqsE+kyq8MKfTYjef0QCHIRyiYJNIwkFlStatG45ZFsfEdr1ar6OtfXjpa87RTi9ILwHfspDaw
WQrcDZVJ//4cAVYQ8E6lewLugxbWZRW8QU6HvJiTZGTD/Xe0JHG/V8ijuLObg0G/N/lhbhCbK5KL
7LoEEtTtBeiHd0PCXmYufLN7u+N+E1gaKZlbwUML9eGql4Xq++OwcyOBcDbO40+/e+trMgQCXhLD
VOAPQTr1ZubnVs5IVTXhHqfr/a/MtHGvSDj5FXd0uS+tgyzLjV8DSpFtoLSiPphZnpp0aM8mk0VN
CfrwPvDZsd8fW95vftkStlZccMaXnKqyllhcVNjFnzDKp6L99Kjo1i80GBOdcnahvEt72VBVN6C7
SE+VNE9AbY9HyEWXoWFJpzwNL7oKXhZlUyO2On8sLGKNdxSrOH5UGdFKbZnHHxgtvNmhnl17Q2JJ
ucFx6Qop7ONFpITjMHgTzDRZ8SwdDQQkagRORtRUyx7L8xGFjkQG6G4m7pQVifNPugObTz8jf6ME
/FEa1G05kFWo2etWZQoF8ldtVANWM+0D1baaraFeECWBtgNMZKEr9xobs15fKWFfgncrGdphrVq2
5BcweKXInUyEGDnnEXKrgpUSDFr9kK4zksUZ1VGUTwPylBnmPh5ffCqwP2mFAoaQKfjRxwl8ZA7x
oP+6d9+SCk94B8Xba7fUQ3FpTKAsRnpsd3nVrHUb4AR/isezm/FhnXrMWQB1K1rTTZxWlCor/k23
GgMGyToXIPw4EHi+dw6sMhoWOd/7ovvAkjrdo/9Nnl1hMhCwkqjvVMvQ8fXm0ktUACUyknIxO8M6
TfjIX1yzEE1SyTiFBY5q8wtj3aZh7r9Yn9ltjG/GrfI3TUjyESc8j+q1IXd01fFVrIxrLU9syeNQ
lP4j7cwqe+ju0dQgJ2lobXYSBUSGOSK785W7tD0GXUKyx1ZCdL9TqMtSYj4ttRypwzzLggpgDd8g
Fh8hkuTvUj0w/sj+OVmpiMclN+iumyxwte1degMuYRFnQswJbDzIg0f7QAOuoBtSYkXjcNmD5Gwh
Qh20nlx+ihCmabyf5pANaeQzkQ51DeeYnStf6jjShr8s5UyOl6wlB2+zAnWe5JoHp1nQUiX9lDZp
NNHHX+lJjPtkz0mrmbNRxbSfutVxBZHlh/Su0oNHq0wcGepmEDqRs28NWNCRm6vcIIYAofMRbDXz
JraS+UZstioNP0istgjvT22e09Ijv2XPOyA/DVB9D2n1WVeOXRuodpywotHayV6L+QXDGLkEjzKG
33KhT81CZAwPz2JWt1sxwywBTCNsWcnNIF15krdg+gU2Gc968xPFyroaeOYkPSZt4uWoITzoNnog
1j6SNE1IA63Dvw/geRs7EhIgRSW2++yJ7BDOs2L+AikFgTrlhhw8P7ulPcqTKltYiRgUePmVXdjt
Ld3qjTdP+cHn6yJw6bcVt7YKY7O94QlVT9ovbB7Qhuk+g0LJ5Pt2AJmpGZTQF6G8QqVb0n+8gfCl
snfVf6TBv5hMDITtM0dHFp/StTUL7k//RF4RqFqMZ+62l2sxNgL9mgZOgcN/hX4I5jEZz40LChMU
mWZqTzkPjEeswHxg29EM/pPw5mQ6nOHgqVZvYD5IacCjCgwy4sGHyYB0veB0CZKUha1VpUSDCJP9
GgQMzAy+WYzgduUueLbJylYSzK4x1pU8yFt5BdJe1YUCKG0tCYNMLEBi7GZebVm25YTOHfnoa5iE
KgFe4HfdJg71tQis7+Wnm3K6N7fcQlI5o8esKf89vKnqZsN5b1zhBALlBENpRuwDb/3RlQ8doqO3
AsXJdax70gZfC9g4Nt3Ld28kesGdriudJPCZZPZsJnLri/y5rvVhSYjj7+BCdHsWBDA1lA3iOV2+
mcZdH4hSOnkxnfwjDqe4+VoNAI8Tg0iEJ16RTypxmXMsXGpQuIfCGABwriubiSzaVKL2oV5n31hA
pcFxzwwIS+Pot4VEWbxVg9J9/ILJDkkIPIPHFHx6kVeYM61/D9cAISEtiK5rC56W+tA/GzZ/nNmI
0woWZYlBGjI7mpIb1D5wl7dFUNAG5xJHEA1oPcJ5qRhidQnsAK5beFbtmcVs5nENZuyLnn86gpq+
1QR/c227ln9Vetvl0NV5MAEly0bN0SQRkwTtDVVIAEF+fGYAt3XrQqLh09OZfrUFUGLg51vdB8Bf
TtG3IXWmz/n2X5w7nyG8zB57mInv57rM2So6AJ0lA5GpEU01gfcPqFrrJXAmsXNa1d31/cbN5zYg
5E3EXul23eVjCg==
`protect end_protected


library ieee;
use ieee.std_logic_1164.all;
package AjitCoreConfigurationPackage is
-- sleep time for ever-spinning modules.
  constant  CORE_SLEEP_TIME 	: integer :=     100 ;

-------------------------------------------- SPECIAL CONFIGURATION PARAMETERS --------------------------------
-- These are nominal values.  If modified, they should be modified as a group. See the HOWTO on processor builds.
--------------------------------------------------------------------------------------------------------------
  constant  TWO_THREADS_IN_CORE		: integer :=  0 ; -- two threads in core?
  constant  THREAD_IS_ISA_64		: integer :=  0 ; -- thread is 64-bit ISA?

  constant  DCACHE_BUFFER_REQUEST	: integer :=  0 ; -- buffer request inside DCACHE?  Adds one cycle to dcache hit latency!
  constant  ICACHE_BUFFER_REQUEST	: integer :=  0 ; -- buffer request inside ICACHE?  Adds one cycle to icache hit latency!

-- If buffering is used 
  constant  DCACHE_HIT_LATENCY       : integer :=     (2 + (TWO_THREADS_IN_CORE + DCACHE_BUFFER_REQUEST))	; -- DCACHE hit path latency (including buffering)
  constant  ICACHE_HIT_LATENCY       : integer :=     (2 + (TWO_THREADS_IN_CORE + ICACHE_BUFFER_REQUEST))    ; -- ICACHE hit path latency (including buffering)

  constant  LOG_DCACHE_SET_ASSOCIATIVITY : integer :=   2  ;   -- log of set associativity.
  constant  LOG_ICACHE_SET_ASSOCIATIVITY : integer :=   2  ;   -- log of set associativity.

  constant  DCACHE_ASSOCIATIVITY         : integer :=  (2 ** LOG_DCACHE_SET_ASSOCIATIVITY) ; -- dcache associativity
  constant  ICACHE_ASSOCIATIVITY         : integer :=  (2 ** LOG_ICACHE_SET_ASSOCIATIVITY) ; -- icache associativity

  constant  TREAT_NONCACHEABLE_AS_BYPASS  : integer :=  1 ; -- non-cacheables will be treated as bypasses...

--------------------------------------   CONFIGURABLE DCACHE PARAMETERS ---------------------------------
  constant  LOG_DCACHE_SIZE_IN_BLOCKS  : integer :=     9  	; -- Note: can be 7,8, or 9 (9 is 32KB)
  constant  DCACHE_SIZE_IN_BLOCKS      : integer :=     (2 ** LOG_DCACHE_SIZE_IN_BLOCKS)	;
  constant  DCACHE_WAY_SIZE            : integer :=     (DCACHE_SIZE_IN_BLOCKS - DCACHE_ASSOCIATIVITY) ;

--------------------------------------   CONFIGURABLE ICACHE PARAMETERS ---------------------------------
  constant  LOG_ICACHE_SIZE_IN_BLOCKS  : integer :=     9  ; -- Note: can be 7,8, or 9 (9 is 32KB)
  constant  ICACHE_SIZE_IN_BLOCKS      : integer :=     (2 ** LOG_ICACHE_SIZE_IN_BLOCKS)	;
  constant  ICACHE_WAY_SIZE            : integer :=     (ICACHE_SIZE_IN_BLOCKS - ICACHE_ASSOCIATIVITY) ;

--------------------------------------   CONFIGURABLE RAS  PARAMETERS ---------------------------------
  constant  LOG_RAS_DEPTH  : integer :=     4  ; -- small.
  constant  RAS_DEPTH      : integer :=     (2 ** LOG_RAS_DEPTH)	;

-------------------------------------------- CACHE PARAMETERS -------------------------------------------------
-- DO NOT MODIFY UNLESS YOU KNOW WHAT YOU ARE DOING!!
--------------------------------------------------------------------------------------------------------------
  constant  LOG_BYTES_PER_DWORD       : integer :=     3	;
  constant  LOG_DWORDS_PER_BLOCK      : integer :=     3	;
  constant  BYTES_PER_DWORD           : integer :=     (2 ** LOG_BYTES_PER_DWORD)	;
  constant  DCACHE_ADDR_WIDTH	      : integer :=     32	;
  constant  ICACHE_ADDR_WIDTH	      : integer :=     32	;
  constant  LOG_BASE_PAGE_SIZE	: integer := 	12 ;
  constant  BASE_PAGE_SIZE	: integer := 	(2 ** LOG_BASE_PAGE_SIZE) ;
  constant  PHYSICAL_ADDR_WIDTH  : integer := 	36 ;
  constant  VIRTUAL_ADDR_WIDTH   : integer := 	32 ;
  constant  LOG_CACHE_LINE_SIZE  : integer :=        6 ;
  constant  CACHE_LINE_SIZE      : integer :=       (2 ** LOG_CACHE_LINE_SIZE) ;   -- bytes.
  constant  CRITICAL_WAY_SIZE    : integer :=   (2**(LOG_BASE_PAGE_SIZE - LOG_CACHE_LINE_SIZE)) ; -- 64.

------------------------------------------------------------------------------------------------------

---------------------------------------------  DERIVED PARAMETERS ----------------------------------------
  constant  DWORDS_PER_BLOCK 	      : integer :=     (2 ** LOG_DWORDS_PER_BLOCK)	;
  constant  DCACHE_TAG_WIDTH           : integer :=     (32 - ((LOG_DWORDS_PER_BLOCK + LOG_BYTES_PER_DWORD) + LOG_DCACHE_SIZE_IN_BLOCKS))	;
  constant  DWORD_SIZE_IN_BITS         : integer :=     (BYTES_PER_DWORD * 8)	;
  constant  BLOCK_SIZE_IN_BITS         : integer :=     (DWORD_SIZE_IN_BITS * DWORDS_PER_BLOCK)	;
  constant  ICACHE_TAG_WIDTH           : integer :=     (32 - ((LOG_DWORDS_PER_BLOCK + LOG_BYTES_PER_DWORD) + LOG_ICACHE_SIZE_IN_BLOCKS))	;
------------------------------------------------------------------------------------------------------


----------------------------------------  FIXED MMU PARAMETERS ------------------------------------------------

  constant  DEFAULT_CACHEABLE_BIT				: integer :=     0 ;  -- keep it 0 if you dont know what it means
  constant  DWORDS_PER_LINE					: integer :=     8 ;


  constant  LOG_NUMBER_OF_L0_TLB_ENTRIES				: integer :=     1 ;  -- should be >= 0 and  at most 2
  constant  NUMBER_OF_L0_TLB_ENTRIES 				: integer :=     ( 2 ** LOG_NUMBER_OF_L0_TLB_ENTRIES ) ;
-- 8 bit context.
  constant  L0_TAG_WIDTH						: integer :=     ( 8 - LOG_NUMBER_OF_L0_TLB_ENTRIES) ;

  constant  LOG_NUMBER_OF_L1_TLB_ENTRIES				: integer :=     2  ; -- should be  >= 0 and at most 7
-- 16 MB pages, so 8 bits to identify page..
  constant  NUMBER_OF_L1_TLB_ENTRIES 				: integer :=     ( 2 ** LOG_NUMBER_OF_L1_TLB_ENTRIES ) ;
  constant  L1_TAG_WIDTH						: integer :=     ( 8 - LOG_NUMBER_OF_L1_TLB_ENTRIES)   ;

  constant  LOG_NUMBER_OF_L2_TLB_ENTRIES				: integer :=     4 ; -- should be  >= 0 and at most 6
  constant  NUMBER_OF_L2_TLB_ENTRIES 				: integer :=     ( 2 ** LOG_NUMBER_OF_L2_TLB_ENTRIES ) ;
-- 256kB pages, so 14 bits to identify page
  constant  L2_TAG_WIDTH						: integer :=     (14 - LOG_NUMBER_OF_L2_TLB_ENTRIES) ;

  constant  LOG_NUMBER_OF_L3_TLB_ENTRIES				: integer :=     6 ; -- should be  >= 0 and at most 8
  constant  NUMBER_OF_L3_TLB_ENTRIES 				: integer :=     ( 2 ** LOG_NUMBER_OF_L3_TLB_ENTRIES ) ;
-- 20-bit page id  (4kB-pages), of which bottom  LOG_L3 bits are rejected.
-- so 20-LOG_L3
  constant  L3_TAG_WIDTH						: integer :=     (20 - LOG_NUMBER_OF_L3_TLB_ENTRIES) ;


-- 2-entry tlb-0 (fully associative)
  constant  TLB_NEW_0_LOG_MEM_SIZE				: integer :=     1 ;
  constant  TLB_NEW_0_LOG_SET_SIZE				: integer :=     1 ;
  constant  TLB_NEW_0_LOG_NUMBER_OF_SETS				: integer :=     (TLB_NEW_0_LOG_MEM_SIZE - TLB_NEW_0_LOG_SET_SIZE) ;

-- 4-entry tlb-1 (fully associative)
  constant  TLB_NEW_1_LOG_MEM_SIZE				: integer :=     2 ;
  constant  TLB_NEW_1_LOG_SET_SIZE				: integer :=     2 ;
  constant  TLB_NEW_1_LOG_NUMBER_OF_SETS				: integer :=     (TLB_NEW_1_LOG_MEM_SIZE - TLB_NEW_1_LOG_SET_SIZE) ;

-- 16-entry tlb-2 (fully associative)
  constant  TLB_NEW_2_LOG_MEM_SIZE				: integer :=     4 ;
  constant  TLB_NEW_2_LOG_SET_SIZE				: integer :=     4 ;
  constant  TLB_NEW_2_LOG_NUMBER_OF_SETS				: integer :=     (TLB_NEW_2_LOG_MEM_SIZE - TLB_NEW_2_LOG_SET_SIZE) ;


-- 256-entry tlb-3 (4-way set associative)
  constant  TLB_NEW_3_LOG_MEM_SIZE				: integer :=     8 ;
  constant  TLB_NEW_3_LOG_SET_SIZE				: integer :=     2 ;
  constant  TLB_NEW_3_LOG_NUMBER_OF_SETS				: integer :=     (TLB_NEW_3_LOG_MEM_SIZE - TLB_NEW_3_LOG_SET_SIZE) ;

-- ICACHE RLUT.
  constant  ICACHE_RLUT_LOG_MEMORY_SIZE : integer :=   LOG_ICACHE_SIZE_IN_BLOCKS  ;
  constant  ICACHE_RLUT_MEMORY_SIZE      : integer :=   (2 ** ICACHE_RLUT_LOG_MEMORY_SIZE)  ;
  constant  ICACHE_RLUT_LOG_SET_SIZE    : integer :=   ((ICACHE_RLUT_LOG_MEMORY_SIZE  + LOG_CACHE_LINE_SIZE) - LOG_BASE_PAGE_SIZE)  ;
  constant  ICACHE_RLUT_SET_SIZE         : integer :=   (2 ** ICACHE_RLUT_LOG_SET_SIZE) ;
  constant  ICACHE_RLUT_LOG_N_SETS      : integer :=   (ICACHE_RLUT_LOG_MEMORY_SIZE - ICACHE_RLUT_LOG_SET_SIZE)  ;
  constant  ICACHE_RLUT_N_SETS           : integer :=   (2 ** ICACHE_RLUT_LOG_N_SETS)  ;
  constant  ICACHE_RLUT_DATA_WIDTH       : integer :=   (VIRTUAL_ADDR_WIDTH - LOG_CACHE_LINE_SIZE) ;
  constant  ICACHE_RLUT_REDUCED_DATA_WIDTH   : integer :=  ((LOG_ICACHE_SIZE_IN_BLOCKS + LOG_CACHE_LINE_SIZE) - LOG_BASE_PAGE_SIZE) ; --
  constant  ICACHE_RLUT_TAG_WIDTH        : integer :=   ((PHYSICAL_ADDR_WIDTH - LOG_CACHE_LINE_SIZE) - ICACHE_RLUT_LOG_N_SETS) ;



-- DCACHE RLUT.
  constant  DCACHE_RLUT_LOG_MEMORY_SIZE : integer :=   LOG_DCACHE_SIZE_IN_BLOCKS  ;
  constant  DCACHE_RLUT_MEMORY_SIZE      : integer :=   (2 ** DCACHE_RLUT_LOG_MEMORY_SIZE)  ;
  constant  DCACHE_RLUT_LOG_SET_SIZE    : integer :=   ((DCACHE_RLUT_LOG_MEMORY_SIZE  + LOG_CACHE_LINE_SIZE) - LOG_BASE_PAGE_SIZE)  ;
  constant  DCACHE_RLUT_SET_SIZE         : integer :=   (2 ** DCACHE_RLUT_LOG_SET_SIZE) ;
  constant  DCACHE_RLUT_LOG_N_SETS      : integer :=   (DCACHE_RLUT_LOG_MEMORY_SIZE - DCACHE_RLUT_LOG_SET_SIZE)  ;
  constant  DCACHE_RLUT_N_SETS           : integer :=   (2 ** DCACHE_RLUT_LOG_N_SETS)  ;
  constant  DCACHE_RLUT_DATA_WIDTH       : integer :=   (VIRTUAL_ADDR_WIDTH - LOG_CACHE_LINE_SIZE) ;
  constant  DCACHE_RLUT_REDUCED_DATA_WIDTH   : integer :=  ((LOG_DCACHE_SIZE_IN_BLOCKS + LOG_CACHE_LINE_SIZE) - LOG_BASE_PAGE_SIZE) ;
  constant  DCACHE_RLUT_TAG_WIDTH        : integer :=   ((PHYSICAL_ADDR_WIDTH - LOG_CACHE_LINE_SIZE) - DCACHE_RLUT_LOG_N_SETS) ;


-- invalidate cache.
--   8-entry fully associative cache.
  constant  SNOOP_CACHE_LOG_MEMORY_SIZE : integer :=  3 ;
  constant  SNOOP_CACHE_LOG_SET_SIZE    : integer :=  3 ;
  constant  SNOOP_CACHE_LOG_NUMBER_OF_SETS    : integer :=  (SNOOP_CACHE_LOG_MEMORY_SIZE - SNOOP_CACHE_LOG_SET_SIZE) ;
  constant  SNOOP_CACHE_TAG_WIDTH             : integer :=   ((PHYSICAL_ADDR_WIDTH - LOG_CACHE_LINE_SIZE) - 
							SNOOP_CACHE_LOG_NUMBER_OF_SETS) ;

-- coherent memory controller assumptions.
  constant   NUMBER_OF_INVALIDATE_SLOTS_PER_CORE	 : integer := 		12 ;

------------------------------------------------------------------------------------------------
-- FIXED parameters for the L2 Caches.
  constant  L2CACHE_LOG2_ASSOCIATIVITY 		: integer :=                3 ;
  constant  L2CACHE_ASSOCIATIVITY 		: integer :=  (2 ** L2CACHE_LOG2_ASSOCIATIVITY) ;
  constant  L2CACHE_LOG2_LINE_SIZE		: integer :=  6 ;
  constant  L2CACHE_LINE_SIZE  			: integer :=  (2 ** L2CACHE_LOG2_LINE_SIZE) ; 	        -- Bytes. 
  constant  L2CACHE_LOG2_LINE_SIZE_IN_DWORDS	: integer :=  3 ;
  constant  L2CACHE_LINE_SIZE_IN_DWORDS 		: integer :=  (2 ** L2CACHE_LOG2_LINE_SIZE_IN_DWORDS) ; -- double words.
------------------------------------------------------------------------------------------------


--
-- instruction buffer to be used in dual threaded CPU's.
--
  constant  ASI_FAKE_INSTRUCTION_BUFFER                : integer :=   127 ; -- whatever.
  constant  INSTRUCTION_BUFFER_LOG_MEMORY_SIZE         : integer :=   7   ; -- 128 entries.
  constant  INSTRUCTION_BUFFER_LOG_ASSOCIATIVITY       : integer :=   0   ; -- 1-way.. do not touch.
  constant  INSTRUCTION_BUFFER_LOG_N_SETS              : integer :=   7   ; -- 128
  constant  INSTRUCTION_BUFFER_TAG_WIDTH               : integer :=   (29 - INSTRUCTION_BUFFER_LOG_N_SETS) ; -- 28
  constant  INSTRUCTION_BUFFER_DATA_WIDTH              : integer :=   (64 + 3) ; -- ipair, acc

  constant  LOG_IBUF_CACHE_SIZE  : integer :=  6 ; -- instruction buffer cache in ifetch.
  constant  IBUF_CACHE_SIZE      : integer :=  ( 2 ** LOG_IBUF_CACHE_SIZE) ; -- nominally 64 entries.
  constant  IBUF_CACHE_TAG_WIDTH : integer :=  (29 - LOG_IBUF_CACHE_SIZE)  ; -- tag

-- for EE_1 processor
  constant  EE_1_INTERNAL_MEM_SIZE_IN_BYTES  : integer :=  (128 * 1024) ; -- EE_1 munit internal memory size.

end package;
package AjitGlobalConfigurationPackage is
	
	-- change the following to true for implementing
	-- the chip.
	constant use_tristates_flag: boolean := false;

	-- this should be at most 36. We need 22 for OS boot,
	-- 16 for running verification tests.
	constant sram_stub_address_width: integer := 20; -- for testing purposes.

        -- for simulations, truncate addresses.
        -- if false, an error will be signalled....
        constant sram_address_truncate_for_sims: boolean := true;

	-- can customize the number of lines in the ICACHE and DCACHE.
	-- For 180nm SCL, keep these at 8, In 65nm, 9.
	--   Superseded by entries in AjitCoreConfiguration.
	-- constant icache_log_number_of_lines: integer := 9; -- 512 lines, each line has 64 bytes.
	-- constant dcache_log_number_of_lines: integer := 9; -- 512 lines, each line has 64 bytes.

	-- MMU TLB entries... DO NOT TOUCH THESE, BECAUSE MMU TLB
	-- access code in AA has some hardwiring in it.  YOU WILL NEED
	-- TO CHANGE BOTH TOGETHER....
	constant mmu_log_tlb_level_0_entries : integer := 1; -- 2-entry  L0 TLB.
	constant mmu_log_tlb_level_1_entries : integer := 2; -- 4-entry  L1 TLB.
	constant mmu_log_tlb_level_2_entries : integer := 4; -- 16-entry  L2 TLB.
	constant mmu_log_tlb_level_3_entries : integer := 6; -- 64-entry L3 TLB.

	-- MMU TLB entries... DO NOT TOUCH THESE, BECAUSE MMU TLB
	-- access code in AA has some hardwiring in it.  YOU WILL NEED
	-- TO CHANGE BOTH TOGETHER....
	constant mmu_log_tlb_new_0_mem_size : integer := 1; -- 2-entry  L0 TLB.
	constant mmu_log_tlb_new_1_mem_size : integer := 2; -- 4-entry  L1 TLB.
	constant mmu_log_tlb_new_2_mem_size : integer := 4; -- 16-entry  L2 TLB.
	constant mmu_log_tlb_new_3_mem_size : integer := 8; -- 256-entry L3 TLB.
	constant mmu_log_tlb_new_3_set_size : integer := 2; -- 4-way set associative
	constant mmu_log_tlb_new_3_number_of_sets : integer := 6; -- 64-sets.

	constant DCACHE_BYPASS_RESPONSE_QUEUE_DEPTH: integer := 8;

end package;
library std;
use std.textio.all;

library ieee;
use ieee.std_logic_1164.all;

package MemmapPackage is
  type ByteArray is array (natural range <>) of std_logic_vector(7 downto 0);
  procedure read_memmap_file(file_name: in string; byte_array: out ByteArray; line_count: out integer);
  function construct_init_byte_array (file_name: in string; array_size: integer) return ByteArray;
  function Select_Byte_Init_Value_By_Position_In_Double_Word (byte_pos : integer; init_val: ByteArray)
    			return ByteArray;
  function to_std_logic_vector(x: bit_vector) return std_logic_vector;

  function insertByteIntoU64(orig_val: std_logic_vector; offset: integer; 
					insbyte: std_logic_vector) return std_logic_vector;
  function updateU64UsingByteMask
		(orig_val: std_logic_vector; byte_mask: std_logic_vector;
						insert_val: std_logic_vector)
			return std_logic_vector;
end package;

package body MemmapPackage is

  function to_std_logic_vector(x: bit_vector) return std_logic_vector is

	alias lx: bit_vector(1 to x'length) is x;
	variable ret_var: std_logic_vector(1 to x'length);
  begin
	for I in 1 to x'length loop
		if(lx(I) = '1') then
			ret_var(I) := '1';
		else
			ret_var(I) := '0';
		end if;
	end loop;
	return(ret_var);
  end function;

  procedure read_memmap_file(file_name: in string; byte_array: out ByteArray; line_count: out integer) is
    variable address_var: integer;
    variable data_var : bit_vector(7 downto 0);
    variable slv_data_var : std_logic_vector(7 downto 0);

    alias  r_var: ByteArray(0 to byte_array'length-1) is byte_array;

    File INFILE: text open read_mode is file_name;
    variable INPUT_LINE: Line;
    variable r_line_count: integer;
  begin
    r_line_count := 0;
    while not endfile(INFILE) loop 
	  readLine (INFILE, INPUT_LINE);
          read (INPUT_LINE, address_var);
          read (INPUT_LINE, data_var);
	  slv_data_var := to_std_logic_vector(data_var);
	 
  	  if((address_var >= 0) and (address_var < byte_array'length)) then
		r_var(address_var) := slv_data_var;
		--assert false report "mem[" & Convert_To_String(address_var) & "] = " & 
		 	--Convert_SLV_To_String (slv_data_var) severity note;
	  end if;

 	  r_line_count := r_line_count + 1;

    end loop;
    line_count := r_line_count;
  end procedure;

  function Select_Byte_Init_Value_By_Position_In_Double_Word (byte_pos : integer; init_val: ByteArray)
    return ByteArray
  is
    variable ret_val :  ByteArray(0 to (init_val'length/8)-1);
    variable addr : integer;
    variable slv_data_var : std_logic_vector(7 downto 0);
    alias r_init_val: ByteArray(0 to init_val'length-1) is init_val;
  begin
      for I in ret_val'low to ret_val'high loop 
        addr := (8*I) + byte_pos;
        if(addr < init_val'length) then
        	slv_data_var := r_init_val(addr);
        	ret_val(I) := slv_data_var;
		--assert false report "Select_Byte_Init_Value: byte_pos= " & Convert_To_String(byte_pos) &
                       --"  mem[" & Convert_To_String(I) & "] = " & 
				 --Convert_SLV_To_String (slv_data_var) severity note;
	end if;
      end loop;
    return (ret_val);    
  end function Select_Byte_Init_Value_By_Position_In_Double_Word;
  
  function construct_init_byte_array (file_name: in string; array_size: integer) return ByteArray is
	variable ret_array: ByteArray(0 to array_size-1);
	variable line_count: integer;
  begin
  	read_memmap_file(file_name => file_name,
				 byte_array => ret_array, 
					line_count => line_count);
	return ret_array;
  end function;

  function insertByteIntoU64(orig_val: std_logic_vector; offset: integer; 
					insbyte: std_logic_vector) return std_logic_vector is
     variable ret_val : std_logic_vector(0 to orig_val'length-1);
     alias lorig_val  : std_logic_vector(0 to orig_val'length-1) is orig_val;
  begin
     assert (orig_val'length = 64) report "wrong word-length in insertByteIntoU64 " severity failure;
     ret_val := orig_val;
     for I in 0 to 7 loop
         if(offset = I) then
             ret_val((8*I) to (8*I)+7) := insbyte;
         end if;
     end loop;
     return(ret_val);
  end function;

  function updateU64UsingByteMask
		(orig_val: std_logic_vector; byte_mask: std_logic_vector;
						insert_val: std_logic_vector)
			return std_logic_vector is
     variable ret_val : std_logic_vector(0 to orig_val'length-1);
     alias lorig_val  : std_logic_vector(0 to orig_val'length-1) is orig_val;
     alias linsert_val  : std_logic_vector(0 to insert_val'length-1) is insert_val;
     alias lbyte_mask    : std_logic_vector(0 to byte_mask'length-1) is byte_mask;
  begin
     assert (orig_val'length = 64) report "wrong word-length in updateU64UsingByteMask " severity failure;
     assert (byte_mask'length = 8) report "wrong byte-mask-length in updateU64UsingByteMask " severity failure;
     ret_val := lorig_val;
     for I in 0 to 7 loop
        if(lbyte_mask(I) = '1') then
             ret_val((8*I) to (8*I)+7) := linsert_val((8*I) to (8*I)+7);
	end if; 
     end loop;
     return(ret_val);
  end function;
   

end package body;
library ieee;
use ieee.std_logic_1164.all;
library AjitCustom;
use AjitCustom.MemmapPackage.all;

package AjitCustomComponents is

  component Simple4StageSynchronizer is
    port (clk, reset_asynch: in std_logic; reset_synch: out std_logic);
  end component Simple4StageSynchronizer;

  component  GenericCacheArray is -- 
    generic (name: string := "anon";
		log2_number_of_blocks: integer := 9; 
		log2_block_size_in_bytes: integer := 6; 
		address_width: integer := 32;
		log2_data_width_in_bytes: integer := 3);
    port ( -- 
      trigger: in std_logic;
      done: out std_logic;
      access_mae : in  std_logic;
      access_array_command : in  std_logic_vector(2 downto 0);
      access_byte_mask : in  std_logic_vector((2**log2_data_width_in_bytes)-1 downto 0);
      access_array_addr : in  std_logic_vector(address_width-1 downto 0);
      access_dword : in  std_logic_vector((8*(2**log2_data_width_in_bytes))-1 downto 0);
      dword_out : out  std_logic_vector((8*(2**log2_data_width_in_bytes))-1 downto 0);
      clk, reset: in std_logic
      -- 
    );
    -- 
  end component GenericCacheArray;
  component GenericIcacheArray is -- 
   generic (name: string := "anon";
		log2_number_of_blocks: integer := 9; 
		log2_block_size_in_bytes: integer := 6; 
		address_width: integer := 32;
		log2_data_width_in_bytes: integer := 3);
  port ( -- 
    trigger: in std_logic;
    done: out std_logic;
    access_mae : in  std_logic;
    access_array_command : in  std_logic_vector(2 downto 0);
    access_array_addr : in  std_logic_vector(address_width-1 downto 0);
    access_dword : in  std_logic_vector((8*(2**log2_data_width_in_bytes))-1 downto 0);
    dword_out : out  std_logic_vector((8*(2**log2_data_width_in_bytes))-1 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
  end component GenericIcacheArray;

  component GenericCacheTags is -- 
    generic (name: string := "anon";
		log2_number_of_blocks: integer := 9; 
		log2_block_size_in_bytes: integer := 6; 
		address_width: integer := 32;
		tag_length: integer := 1;
		log2_data_width_in_bytes: integer := 3);
    port ( -- 
      start_req: in std_logic;
      start_ack: out std_logic;
      fin_req: in std_logic;
      fin_ack: out std_logic;
      init_flag : in  std_logic;
      access_mae : in  std_logic;
      access_S : in  std_logic;
      access_is_read: in std_logic;
      access_is_ifetch: in std_logic;
      access_acc: in std_logic_vector(2 downto 0);
      access_tag_command : in  std_logic_vector(2 downto 0);
      access_tag_addr : in  std_logic_vector(address_width-1 downto 0);
      is_hit : out  std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0);
      permissions_ok : out  std_logic_vector(0 downto 0);
      clk, reset: in std_logic
      -- 
  );
  -- 
  end component GenericCacheTags;

  component GenericCacheTagsWithInvalidate is -- 
    generic (name: string := "anon";
		log2_number_of_blocks: integer := 9; 
		log2_block_size_in_bytes: integer := 6; 
		address_width: integer := 32;
		log2_data_width_in_bytes: integer := 3);
    port ( -- 
      trigger: in std_logic;
      done: out std_logic;
      init_flag : in  std_logic;
      access_mae : in  std_logic;
      access_S : in  std_logic;
      access_is_read: in std_logic;
      access_is_ifetch: in std_logic;
      access_acc: in std_logic_vector(2 downto 0);
      access_tag_command : in  std_logic_vector(2 downto 0);
      access_tag_addr : in  std_logic_vector(address_width-1 downto 0);
      -- invalidation channel for cache coherence and synonym avoidance.
      invalidate: in std_logic_vector(0 downto 0);
      invalidate_line_address: in std_logic_vector(((address_width-1) - log2_block_size_in_bytes) downto 0);
      is_hit : out  std_logic_vector(0 downto 0);
      permissions_ok : out  std_logic_vector(0 downto 0);
      lookup_acc : out  std_logic_vector(2 downto 0);
      clk, reset: in std_logic
  );
  end component GenericCacheTagsWithInvalidate;

  component GenericDcacheTagsArraysWithInvalidate is -- 
    generic (name: string := "anon";
		log2_number_of_blocks: integer := 9; 
		log2_block_size_in_bytes: integer := 6; 
		address_width: integer := 32;
		log2_data_width_in_bytes: integer := 3);
  port ( -- 
    trigger     : in std_logic;
    done        : out std_logic;
    init_flag : in  std_logic;
    access_mae : in  std_logic;
    access_S : in  std_logic;
    access_is_read: in std_logic;
    access_is_ifetch: in std_logic;
    access_acc: in std_logic_vector(2 downto 0);
    access_tag_command: in std_logic_vector(2 downto 0);
    access_tag_addr : in  std_logic_vector(address_width-1 downto 0);
    -- invalidation channel for cache coherence and synonym avoidance.
    invalidate: in std_logic_vector(0 downto 0);
    invalidate_line_address: in std_logic_vector(((address_width-1) - log2_block_size_in_bytes) downto 0);
    is_hit : out  std_logic_vector(0 downto 0);
    permissions_ok : out  std_logic_vector(0 downto 0);
    access_array_command : in  std_logic_vector(2 downto 0);
    access_byte_mask : in  std_logic_vector((2**log2_data_width_in_bytes)-1 downto 0);
    access_array_addr : in  std_logic_vector(address_width-1 downto 0);
    access_dword : in  std_logic_vector((8*(2**log2_data_width_in_bytes))-1 downto 0);
    dword_out : out  std_logic_vector((8*(2**log2_data_width_in_bytes))-1 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
  end component GenericDcacheTagsArraysWithInvalidate;

  component GenericIcacheTagsArraysWithInvalidate is -- 
   generic (name: string := "anon";
		log2_number_of_blocks: integer := 9; 
		log2_block_size_in_bytes: integer := 6; 
		address_width: integer := 32;
		log2_data_width_in_bytes: integer := 3);
  port ( -- 
    -- start it off
    trigger		     : in std_logic;
    -- is it done?  This will be asserted for
    -- exactly one clock cycle.
    done		     : out std_logic;
    
    init_flag : in  std_logic;
    access_mae : in  std_logic;
    access_S : in  std_logic;
    access_is_read: in std_logic;
    access_is_ifetch: in std_logic;
    access_acc: in std_logic_vector(2 downto 0);
    access_tag_command : in  std_logic_vector(2 downto 0);
    -- invalidation channel for cache coherence and synonym avoidance.
    invalidate: in std_logic_vector(0 downto 0);
    invalidate_line_address: in std_logic_vector(((address_width-1) - log2_block_size_in_bytes) downto 0);
    is_hit : out  std_logic_vector(0 downto 0);
    permissions_ok : out  std_logic_vector(0 downto 0);
    lookup_acc : out  std_logic_vector(2 downto 0);
    access_array_command : in  std_logic_vector(2 downto 0);
    access_addr : in  std_logic_vector(address_width-1 downto 0);
    access_dword : in  std_logic_vector((8*(2**log2_data_width_in_bytes))-1 downto 0);
    dword_out : out  std_logic_vector((8*(2**log2_data_width_in_bytes))-1 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
  end component GenericIcacheTagsArraysWithInvalidate;

  component VaToIndexInSetTlb is
	generic (number_of_entries: integer := 4; 
			set_id_width: integer := 8;
			index_in_set_width: integer := 1;
			va_tag_width: integer := 25   -- Va tag.
		);
	port (
		lookup_va_tag:    in std_logic_vector(va_tag_width-1 downto 0);
		lookup_set_id: 	  in std_logic_vector(set_id_width-1 downto 0);

		erase_va_tag: in std_logic_vector(va_tag_width-1 downto 0);
		erase_set_id: in std_logic_vector(set_id_width-1 downto 0);

		insert_va_tag: in std_logic_vector(va_tag_width-1 downto 0);
		insert_set_id: in std_logic_vector(set_id_width-1 downto 0);
		insert_index_in_set: in std_logic_vector(index_in_set_width-1 downto 0);
		insert_acc   : in std_logic_vector(2 downto 0);

		match: out std_logic;
		matched_index_in_set: out std_logic_vector(index_in_set_width-1 downto 0);
		matched_acc: 	  out std_logic_vector(2 downto 0);

		insert: in std_logic;
		lookup: in std_logic;
		erase : in std_logic;
		clear : in std_logic;
		clk, reset:  in std_logic
	);
  end component;

  component GenericSetAssociativeCacheArray is -- 
    generic (name: string := "anon";
		log2_number_of_blocks: integer := 9; 
		log2_block_size_in_bytes: integer := 6; 
		log2_associativity: integer := 1;
		address_width: integer := 32;
		log2_data_width_in_bytes: integer := 3;
		ignore_byte_mask: boolean := false);
    port ( -- 
     -- it is the responsibility of the one who triggers the activity
     -- to ensure that the match_index_in_set field is valid!
    trigger: in std_logic;
    done: out std_logic;
    matched_index_in_set: in std_logic_vector(log2_associativity-1 downto 0);
    access_mae : in  std_logic;
    access_array_command : in  std_logic_vector(2 downto 0);
    access_byte_mask : in  std_logic_vector((2**log2_data_width_in_bytes)-1 downto 0);
    access_array_addr : in  std_logic_vector(address_width-1 downto 0);
    access_array_write_dword : 
	in  std_logic_vector(8*((2**log2_data_width_in_bytes))-1 downto 0);
    access_array_read_dword_vector : 
	out  std_logic_vector(((2**log2_associativity)*8*(2**log2_data_width_in_bytes))-1 downto 0);
    bypassed_dword_out : 
	out  std_logic_vector((8*(2**log2_data_width_in_bytes))-1 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
  end component GenericSetAssociativeCacheArray;


  component GenericSetAssociativeCacheTagsWithInvalidate is -- 
    generic (name: string := "anon";
		log2_number_of_blocks: integer := 9; 
		log2_block_size_in_bytes: integer := 6; 
		address_width: integer := 32;
		log2_associativity: integer := 1;
		log2_data_width_in_bytes: integer := 3);
    port ( -- 
    trigger: in std_logic;
    done   : out std_logic;
    init_flag : in  std_logic;
    access_acc: in std_logic_vector(2 downto 0);
    access_tag_lookup : in  std_logic;
    access_tag_clear_line : in  std_logic;
    access_tag_clear_all : in  std_logic;
    access_tag_insert : in  std_logic;
    access_tag_addr : in  std_logic_vector(address_width-1 downto 0);
    -- invalidation channel for cache coherence and synonym avoidance.
    invalidate: in std_logic;
    invalidate_line_address: in std_logic_vector(((address_width-1) - log2_block_size_in_bytes) downto 0);
    -- valid tlb match info...
    valid_match: in std_logic;
    match_index_in_set: in std_logic_vector(log2_associativity-1 downto 0);
    -- outputs.
    lookup_is_valid : out  std_logic;
    access_index_in_set_valid: out std_logic;
    access_index_in_set: out std_logic_vector(log2_associativity-1 downto 0);
    access_acc_out: out std_logic_vector(2 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
  end component GenericSetAssociativeCacheTagsWithInvalidate;

  component GenericSetAssociativeCacheTagsArraysWithInvalidate is -- 
    generic (
		name: string := "anon";
		log2_number_of_blocks: integer := 9; 
		log2_block_size_in_bytes: integer := 6; 
		log2_associativity: integer := 1;
		address_width: integer := 32;
		log2_data_width_in_bytes: integer := 3;
		icache_flag: boolean := false
	  );
    port ( -- 
    -- start it off
    trigger		     : in std_logic;
    -- is it done?  This will be asserted for
    -- exactly one clock cycle.
    done		     : out std_logic;
    
    init_flag : in  std_logic;
    access_mae : in  std_logic;
    access_S : in  std_logic;
    access_is_read: in std_logic;
    access_is_ifetch: in std_logic;
    access_acc: in std_logic_vector(2 downto 0);
    access_tag_lookup : in  std_logic;
    access_tag_clear_line : in  std_logic;
    access_tag_clear_all : in  std_logic;
    access_tag_insert : in  std_logic;
    access_array_command : in  std_logic_vector(2 downto 0);
    access_addr : in  std_logic_vector(address_width-1 downto 0);
    access_byte_mask : in  std_logic_vector((2**log2_data_width_in_bytes)-1 downto 0);
    access_dword : in  std_logic_vector((8*(2**log2_data_width_in_bytes))-1 downto 0);
    -- invalidation channel for cache coherence and synonym avoidance.
    invalidate: in std_logic_vector(0 downto 0);
    invalidate_line_address: in std_logic_vector(((address_width-1) - log2_block_size_in_bytes) downto 0);
    is_hit : out  std_logic_vector(0 downto 0);
    permissions_ok : out  std_logic_vector(0 downto 0);
    lookup_acc : out  std_logic_vector(2 downto 0);
    dword_out : out  std_logic_vector((8*(2**log2_data_width_in_bytes))-1 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
  end component GenericSetAssociativeCacheTagsArraysWithInvalidate;

  component IcacheFrontendCoreDaemon is  -- system 
   generic (tag_length: integer := 1);
   port (-- 
    NOBLOCK_CPU_to_ICACHE_command_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_ICACHE_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_ICACHE_command_pipe_read_data : in   std_logic_vector(40 downto 0);
    NOBLOCK_CPU_to_ICACHE_reset_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_ICACHE_reset_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_ICACHE_reset_pipe_read_data : in   std_logic_vector(0 downto 0);
    noblock_icache_backend_to_frontend_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_icache_backend_to_frontend_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_icache_backend_to_frontend_pipe_read_data : in   std_logic_vector(101 downto 0);
    ICACHE_to_CPU_reset_ack_pipe_write_req : out  std_logic_vector(0 downto 0);
    ICACHE_to_CPU_reset_ack_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ICACHE_to_CPU_reset_ack_pipe_write_data : out  std_logic_vector(0 downto 0);
    ICACHE_to_CPU_response_pipe_write_req : out  std_logic_vector(0 downto 0);
    ICACHE_to_CPU_response_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ICACHE_to_CPU_response_pipe_write_data : out  std_logic_vector(89 downto 0);
    icache_frontend_to_backend_pipe_write_req : out  std_logic_vector(0 downto 0);
    icache_frontend_to_backend_pipe_write_ack : in   std_logic_vector(0 downto 0);
    icache_frontend_to_backend_pipe_write_data : out  std_logic_vector(41 downto 0);
    MMU_TO_ICACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_req: out std_logic_vector(0 downto 0);
    MMU_TO_ICACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_ack: in std_logic_vector(0 downto 0);
    MMU_TO_ICACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_data: in std_logic_vector(26 downto 0);
    NOBLOCK_MMU_TO_ICACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_req: out std_logic_vector(0 downto 0);
    NOBLOCK_MMU_TO_ICACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_ack: in std_logic_vector(0 downto 0);
    NOBLOCK_MMU_TO_ICACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_data: in std_logic_vector(26 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic);
  end component; 

  component IcacheFrontendDaemon is  -- system 
   generic (tag_length: integer := 1);
   port (-- 
    NOBLOCK_CPU_to_ICACHE_command_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_ICACHE_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_ICACHE_command_pipe_read_data : in   std_logic_vector(40 downto 0);
    NOBLOCK_CPU_to_ICACHE_reset_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_ICACHE_reset_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_ICACHE_reset_pipe_read_data : in   std_logic_vector(0 downto 0);
    noblock_icache_backend_to_frontend_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_icache_backend_to_frontend_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_icache_backend_to_frontend_pipe_read_data : in   std_logic_vector(101 downto 0);
    ICACHE_to_CPU_reset_ack_pipe_write_req : out  std_logic_vector(0 downto 0);
    ICACHE_to_CPU_reset_ack_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ICACHE_to_CPU_reset_ack_pipe_write_data : out  std_logic_vector(0 downto 0);
    ICACHE_to_CPU_response_pipe_write_req : out  std_logic_vector(0 downto 0);
    ICACHE_to_CPU_response_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ICACHE_to_CPU_response_pipe_write_data : out  std_logic_vector(89 downto 0);
    icache_frontend_to_backend_pipe_write_req : out  std_logic_vector(0 downto 0);
    icache_frontend_to_backend_pipe_write_ack : in   std_logic_vector(0 downto 0);
    icache_frontend_to_backend_pipe_write_data : out  std_logic_vector(41 downto 0);
    MMU_TO_ICACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_req: out std_logic_vector(0 downto 0);
    MMU_TO_ICACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_ack: in std_logic_vector(0 downto 0);
    MMU_TO_ICACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_data: in std_logic_vector(26 downto 0);
    NOBLOCK_MMU_TO_ICACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_req: out std_logic_vector(0 downto 0);
    NOBLOCK_MMU_TO_ICACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_ack: in std_logic_vector(0 downto 0);
    NOBLOCK_MMU_TO_ICACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_data: in std_logic_vector(26 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic);
  end component; 


  component IcacheFrontendWithRlutInvalidateDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
    	NOBLOCK_CPU_to_ICACHE_command_pipe_read_req : out  std_logic_vector(0 downto 0);
    	NOBLOCK_CPU_to_ICACHE_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
    	NOBLOCK_CPU_to_ICACHE_command_pipe_read_data : in   std_logic_vector(40 downto 0);
    	NOBLOCK_CPU_to_ICACHE_reset_pipe_read_req : out  std_logic_vector(0 downto 0);
    	NOBLOCK_CPU_to_ICACHE_reset_pipe_read_ack : in   std_logic_vector(0 downto 0);
    	NOBLOCK_CPU_to_ICACHE_reset_pipe_read_data : in   std_logic_vector(0 downto 0);
    	noblock_icache_backend_to_frontend_pipe_read_req : out  std_logic_vector(0 downto 0);
    	noblock_icache_backend_to_frontend_pipe_read_ack : in   std_logic_vector(0 downto 0);
    	noblock_icache_backend_to_frontend_pipe_read_data : in   std_logic_vector(101 downto 0);
    	ICACHE_to_CPU_reset_ack_pipe_write_req : out  std_logic_vector(0 downto 0);
    	ICACHE_to_CPU_reset_ack_pipe_write_ack : in   std_logic_vector(0 downto 0);
    	ICACHE_to_CPU_reset_ack_pipe_write_data : out  std_logic_vector(0 downto 0);
    	ICACHE_to_CPU_response_pipe_write_req : out  std_logic_vector(0 downto 0);
    	ICACHE_to_CPU_response_pipe_write_ack : in   std_logic_vector(0 downto 0);
    	ICACHE_to_CPU_response_pipe_write_data : out  std_logic_vector(89 downto 0);
    	icache_frontend_to_backend_pipe_write_req : out  std_logic_vector(0 downto 0);
    	icache_frontend_to_backend_pipe_write_ack : in   std_logic_vector(0 downto 0);
    	icache_frontend_to_backend_pipe_write_data : out  std_logic_vector(41 downto 0);
    	-- RLUT related.
    	NOBLOCK_RLUT_to_ICACHE_pipe_read_req : out  std_logic_vector(0 downto 0);
    	NOBLOCK_RLUT_to_ICACHE_pipe_read_ack : in   std_logic_vector(0 downto 0);
    	NOBLOCK_RLUT_to_ICACHE_pipe_read_data : in   std_logic_vector(31 downto 0);
    	ICACHE_to_RLUT_pipe_write_req : out  std_logic_vector(0 downto 0);
    	ICACHE_to_RLUT_pipe_write_ack : in   std_logic_vector(0 downto 0);
    	ICACHE_to_RLUT_pipe_write_data: out std_logic_vector(7 downto 0);
    	tag_in: in std_logic_vector(tag_length-1 downto 0);
    	tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    	clk : in std_logic;
    	reset : in std_logic;
    	start_req : in std_logic;
    	start_ack : out std_logic;
    	fin_req : in std_logic;
    	fin_ack   : out std_logic-- 
  	);
  	-- 
   end component IcacheFrontendWithRlutInvalidateDaemon;

  component DcacheFrontendDaemon is -- 
   generic (tag_length : integer); 
   port ( -- 
    NOBLOCK_CPU_to_DCACHE_command_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_command_pipe_read_data : in   std_logic_vector(142 downto 0);
    NOBLOCK_CPU_to_DCACHE_reset_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_reset_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_reset_pipe_read_data : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_data : in   std_logic_vector(120 downto 0);
    noblock_dcache_backend_to_frontend_command_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_dcache_backend_to_frontend_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_dcache_backend_to_frontend_command_pipe_read_data : in   std_logic_vector(83 downto 0);
    -----------------------------------------------------------------------------------------------
    NOBLOCK_DCACHE_TO_CPU_IU_BYPASS_pipe_write_req: out std_logic_vector(0 downto 0);
    NOBLOCK_DCACHE_TO_CPU_IU_BYPASS_pipe_write_ack: in std_logic_vector(0 downto 0);
    NOBLOCK_DCACHE_TO_CPU_IU_BYPASS_pipe_write_data: out std_logic_vector(92 downto 0);
    -----------------------------------------------------------------------------------------------
    NOBLOCK_DCACHE_TO_CPU_FU_BYPASS_pipe_write_req:  out std_logic_vector(0 downto 0);
    NOBLOCK_DCACHE_TO_CPU_FU_BYPASS_pipe_write_ack:  in std_logic_vector(0 downto 0);
    NOBLOCK_DCACHE_TO_CPU_FU_BYPASS_pipe_write_data: out std_logic_vector(92 downto 0);
    -----------------------------------------------------------------------------------------------
    DCACHE_to_CPU_reset_ack_pipe_write_req : out  std_logic_vector(0 downto 0);
    DCACHE_to_CPU_reset_ack_pipe_write_ack : in   std_logic_vector(0 downto 0);
    DCACHE_to_CPU_reset_ack_pipe_write_data : out  std_logic_vector(0 downto 0);
    DCACHE_to_CPU_response_pipe_write_req : out  std_logic_vector(0 downto 0);
    DCACHE_to_CPU_response_pipe_write_ack : in   std_logic_vector(0 downto 0);
    DCACHE_to_CPU_response_pipe_write_data : out  std_logic_vector(71 downto 0);
    DCACHE_to_CPU_slow_response_pipe_write_req : out  std_logic_vector(0 downto 0);
    DCACHE_to_CPU_slow_response_pipe_write_ack : in   std_logic_vector(0 downto 0);
    DCACHE_to_CPU_slow_response_pipe_write_data : out  std_logic_vector(71 downto 0);
    MMU_TO_DCACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_req: out std_logic_vector(0 downto 0);
    MMU_TO_DCACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_ack: in std_logic_vector(0 downto 0);
    MMU_TO_DCACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_data: in std_logic_vector(26 downto 0);
    NOBLOCK_MMU_TO_DCACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_req: out std_logic_vector(0 downto 0);
    NOBLOCK_MMU_TO_DCACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_ack: in std_logic_vector(0 downto 0);
    NOBLOCK_MMU_TO_DCACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_data: in std_logic_vector(26 downto 0);
    dcache_frontend_to_backend_pipe_write_req : out  std_logic_vector(0 downto 0);
    dcache_frontend_to_backend_pipe_write_ack : in   std_logic_vector(0 downto 0);
    dcache_frontend_to_backend_pipe_write_data : out  std_logic_vector(119 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
  end component DcacheFrontendDaemon;

  component DcacheFrontendWithStallCoreDaemon is -- 
   generic (tag_length : integer:= 1); 
   port ( -- 
    NOBLOCK_CPU_to_DCACHE_command_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_command_pipe_read_data : in   std_logic_vector(142 downto 0);
    NOBLOCK_CPU_to_DCACHE_reset_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_reset_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_reset_pipe_read_data : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_data : in   std_logic_vector(120 downto 0);
    noblock_dcache_backend_to_frontend_command_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_dcache_backend_to_frontend_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_dcache_backend_to_frontend_command_pipe_read_data : in   std_logic_vector(83 downto 0);
    -----------------------------------------------------------------------------------------------
    NOBLOCK_DCACHE_TO_CPU_IU_BYPASS_pipe_write_req: out std_logic_vector(0 downto 0);
    NOBLOCK_DCACHE_TO_CPU_IU_BYPASS_pipe_write_ack: in std_logic_vector(0 downto 0);
    NOBLOCK_DCACHE_TO_CPU_IU_BYPASS_pipe_write_data: out std_logic_vector(92 downto 0);
    -----------------------------------------------------------------------------------------------
    NOBLOCK_DCACHE_TO_CPU_FU_BYPASS_pipe_write_req:  out std_logic_vector(0 downto 0);
    NOBLOCK_DCACHE_TO_CPU_FU_BYPASS_pipe_write_ack:  in std_logic_vector(0 downto 0);
    NOBLOCK_DCACHE_TO_CPU_FU_BYPASS_pipe_write_data: out std_logic_vector(92 downto 0);
    -----------------------------------------------------------------------------------------------
    DCACHE_to_CPU_reset_ack_pipe_write_req : out  std_logic_vector(0 downto 0);
    DCACHE_to_CPU_reset_ack_pipe_write_ack : in   std_logic_vector(0 downto 0);
    DCACHE_to_CPU_reset_ack_pipe_write_data : out  std_logic_vector(0 downto 0);
    DCACHE_to_CPU_response_pipe_write_req : out  std_logic_vector(0 downto 0);
    DCACHE_to_CPU_response_pipe_write_ack : in   std_logic_vector(0 downto 0);
    DCACHE_to_CPU_response_pipe_write_data : out  std_logic_vector(71 downto 0);
    DCACHE_to_CPU_slow_response_pipe_write_req : out  std_logic_vector(0 downto 0);
    DCACHE_to_CPU_slow_response_pipe_write_ack : in   std_logic_vector(0 downto 0);
    DCACHE_to_CPU_slow_response_pipe_write_data : out  std_logic_vector(71 downto 0);
    MMU_TO_DCACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_req: out std_logic_vector(0 downto 0);
    MMU_TO_DCACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_ack: in std_logic_vector(0 downto 0);
    MMU_TO_DCACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_data: in std_logic_vector(26 downto 0);
    NOBLOCK_MMU_TO_DCACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_req: out std_logic_vector(0 downto 0);
    NOBLOCK_MMU_TO_DCACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_ack: in std_logic_vector(0 downto 0);
    NOBLOCK_MMU_TO_DCACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_data: in std_logic_vector(26 downto 0);
    CACHE_STALL_ENABLE: in std_logic_vector(0 downto 0);
    NOBLOCK_INVALIDATE_SLOT_RETURN_pipe_read_req : out std_logic_vector(0 downto 0);
    NOBLOCK_INVALIDATE_SLOT_RETURN_pipe_read_ack : in std_logic_vector(0 downto 0);
    NOBLOCK_INVALIDATE_SLOT_RETURN_pipe_read_data: in std_logic_vector(0 downto 0);
    dcache_frontend_to_backend_pipe_write_req : out  std_logic_vector(0 downto 0);
    dcache_frontend_to_backend_pipe_write_ack : in   std_logic_vector(0 downto 0);
    dcache_frontend_to_backend_pipe_write_data : out  std_logic_vector(119 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
  end component DcacheFrontendWithStallCoreDaemon;

  component DcacheFrontendWithStallDaemon is -- 
   generic (tag_length : integer := 1); 
   port ( -- 
    NOBLOCK_CPU_to_DCACHE_command_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_command_pipe_read_data : in   std_logic_vector(142 downto 0);
    NOBLOCK_CPU_to_DCACHE_reset_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_reset_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_reset_pipe_read_data : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_data : in   std_logic_vector(120 downto 0);
    noblock_dcache_backend_to_frontend_command_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_dcache_backend_to_frontend_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_dcache_backend_to_frontend_command_pipe_read_data : in   std_logic_vector(83 downto 0);
    -----------------------------------------------------------------------------------------------
    NOBLOCK_DCACHE_TO_CPU_IU_BYPASS_pipe_write_req: out std_logic_vector(0 downto 0);
    NOBLOCK_DCACHE_TO_CPU_IU_BYPASS_pipe_write_ack: in std_logic_vector(0 downto 0);
    NOBLOCK_DCACHE_TO_CPU_IU_BYPASS_pipe_write_data: out std_logic_vector(92 downto 0);
    -----------------------------------------------------------------------------------------------
    NOBLOCK_DCACHE_TO_CPU_FU_BYPASS_pipe_write_req:  out std_logic_vector(0 downto 0);
    NOBLOCK_DCACHE_TO_CPU_FU_BYPASS_pipe_write_ack:  in std_logic_vector(0 downto 0);
    NOBLOCK_DCACHE_TO_CPU_FU_BYPASS_pipe_write_data: out std_logic_vector(92 downto 0);
    -----------------------------------------------------------------------------------------------
    DCACHE_to_CPU_reset_ack_pipe_write_req : out  std_logic_vector(0 downto 0);
    DCACHE_to_CPU_reset_ack_pipe_write_ack : in   std_logic_vector(0 downto 0);
    DCACHE_to_CPU_reset_ack_pipe_write_data : out  std_logic_vector(0 downto 0);
    DCACHE_to_CPU_response_pipe_write_req : out  std_logic_vector(0 downto 0);
    DCACHE_to_CPU_response_pipe_write_ack : in   std_logic_vector(0 downto 0);
    DCACHE_to_CPU_response_pipe_write_data : out  std_logic_vector(71 downto 0);
    DCACHE_to_CPU_slow_response_pipe_write_req : out  std_logic_vector(0 downto 0);
    DCACHE_to_CPU_slow_response_pipe_write_ack : in   std_logic_vector(0 downto 0);
    DCACHE_to_CPU_slow_response_pipe_write_data : out  std_logic_vector(71 downto 0);
    MMU_TO_DCACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_req: out std_logic_vector(0 downto 0);
    MMU_TO_DCACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_ack: in std_logic_vector(0 downto 0);
    MMU_TO_DCACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_data: in std_logic_vector(26 downto 0);
    NOBLOCK_MMU_TO_DCACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_req: out std_logic_vector(0 downto 0);
    NOBLOCK_MMU_TO_DCACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_ack: in std_logic_vector(0 downto 0);
    NOBLOCK_MMU_TO_DCACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_data: in std_logic_vector(26 downto 0);
    CACHE_STALL_ENABLE: in std_logic_vector(0 downto 0);
    NOBLOCK_INVALIDATE_SLOT_RETURN_pipe_read_req : out std_logic_vector(0 downto 0);
    NOBLOCK_INVALIDATE_SLOT_RETURN_pipe_read_ack : in std_logic_vector(0 downto 0);
    NOBLOCK_INVALIDATE_SLOT_RETURN_pipe_read_data: in std_logic_vector(0 downto 0);
    dcache_frontend_to_backend_pipe_write_req : out  std_logic_vector(0 downto 0);
    dcache_frontend_to_backend_pipe_write_ack : in   std_logic_vector(0 downto 0);
    dcache_frontend_to_backend_pipe_write_data : out  std_logic_vector(119 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
  end component DcacheFrontendWithStallDaemon;

   
  component nonCacheablePageTlb is
	generic (number_of_entries: integer := 4);
	port (
		lookup_virtual_address: in std_logic_vector(31 downto 0);
		lookup_supervisor, lookup_read, lookup_ifetch: in std_logic;
		insert_virtual_address: in std_logic_vector(31 downto 0);
		insert_acc: in std_logic_vector (2 downto 0);

		match: out std_logic;
		insert: in std_logic;
		clear : in std_logic;
		clk, reset:  in std_logic
	);
  end component;
  component DcacheBypassController is -- 
    port ( -- 

    cpu_bypass_command_available: in  boolean; 
    cpu_bypass_command_accept   : out boolean;

    cpu_fast_valid		: in std_logic;
    cpu_slow_valid		: in std_logic;

    is_memory_write		: in std_logic;
    locked_access		: in std_logic;

    cpu_asi		        : in std_logic_vector(7 downto 0);
    cpu_byte_mask	        : in std_logic_vector(7 downto 0);
    cpu_address			: in std_logic_vector(31 downto 0);
    cpu_write_data		: in std_logic_vector(63 downto 0);

    cpu_slow_ready_for_bypass_response      : in boolean;
    write_to_cpu_slow		            : out boolean;

    cpu_fast_ready_for_bypass_response      : in boolean;
    write_to_cpu_fast		            : out boolean;

    response_to_cpu		: out std_logic_vector(71 downto 0);

    be_ready_for_request	: in boolean;
    be_write		       	: out boolean;
    to_be_from_bypass 		: out  std_logic_vector(119 downto 0);

    be_response_ready		: in boolean;
    be_read			: out boolean;
    be_dword			: in std_logic_vector(63 downto 0);

    bypass_response_pending : out boolean;

    clk : in std_logic;
    reset : in std_logic
  );
  -- 
  end component DcacheBypassController;

  component generic_single_port_memory_with_byte_mask is
   generic ( name: string; 
		g_addr_width: natural := 10; 
		g_data_width : natural := 16);
   port (
	   datain : in std_logic_vector(g_data_width-1 downto 0);
           dataout: out std_logic_vector(g_data_width-1 downto 0);
           addrin: in std_logic_vector(g_addr_width-1 downto 0);
	   bytemask: in std_logic_vector((g_data_width/8)-1 downto 0);
           enable: in std_logic;
           writebar : in std_logic;
           clk: in std_logic;
           reset : in std_logic);
   end component generic_single_port_memory_with_byte_mask;
   component protoBoardMemX2MB  is
	generic (tag_length: integer := 2);
	port ( 

		read_write_bar : in std_logic_vector (0 downto 0);
		byte_mask  : in std_logic_vector (7 downto 0);
		address    : in  std_logic_vector (18 downto 0);
		write_data : in std_logic_vector (63 downto 0);
		read_data  : out  std_logic_vector (63 downto 0);
 	   	tag_in: in std_logic_vector(tag_length-1 downto 0);
      	   	tag_out: out std_logic_vector(tag_length-1 downto 0);
		clk, reset: in std_logic;
		start_req: in std_logic;
		start_ack: out std_logic;
		fin_req: in std_logic;
		fin_ack: out std_logic
	     );
   end component protoBoardMemX2MB;

   component protoBoardMemX64KB  is
	generic (tag_length: integer := 2);
	port ( 

		read_write_bar : in std_logic_vector (0 downto 0);
		byte_mask  : in std_logic_vector (7 downto 0);
		address    : in  std_logic_vector (12 downto 0);
		write_data : in std_logic_vector (63 downto 0);
		read_data  : out  std_logic_vector (63 downto 0);
 	   	tag_in: in std_logic_vector(tag_length-1 downto 0);
      	   	tag_out: out std_logic_vector(tag_length-1 downto 0);
		clk, reset: in std_logic;
		start_req: in std_logic;
		start_ack: out std_logic;
		fin_req: in std_logic;
		fin_ack: out std_logic
	     );
   end component protoBoardMemX64KB;

   -- added for simulation purposes only.
   component generic_dual_port_memory_with_byte_mask is
     generic ( name: string; 
		g_addr_width: natural := 10; 
		g_data_width : natural := 16);
     port (
	   datain_0 : in std_logic_vector(g_data_width-1 downto 0);
           dataout_0: out std_logic_vector(g_data_width-1 downto 0);
           addrin_0: in std_logic_vector(g_addr_width-1 downto 0);
	   bytemask_0: in std_logic_vector((g_data_width/8)-1 downto 0);
           enable_0: in std_logic;
           writebar_0 : in std_logic;
	   datain_1 : in std_logic_vector(g_data_width-1 downto 0);
           dataout_1: out std_logic_vector(g_data_width-1 downto 0);
           addrin_1: in std_logic_vector(g_addr_width-1 downto 0);
	   bytemask_1: in std_logic_vector((g_data_width/8)-1 downto 0);
           enable_1: in std_logic;
           writebar_1 : in std_logic;
           clk: in std_logic;
           reset : in std_logic);
   end component generic_dual_port_memory_with_byte_mask;
   component generic_single_port_memory_with_byte_mask_and_init is
   generic ( init_file_name: string; 
		g_addr_width: natural := 10; 
		g_data_width : natural := 16);
   port (
	   datain : in std_logic_vector(g_data_width-1 downto 0);
           dataout: out std_logic_vector(g_data_width-1 downto 0);
           addrin: in std_logic_vector(g_addr_width-1 downto 0);
	   bytemask: in std_logic_vector((g_data_width/8)-1 downto 0);
           enable: in std_logic;
           writebar : in std_logic;
           clk: in std_logic;
           reset : in std_logic);
   end component generic_single_port_memory_with_byte_mask_and_init;

   component cpu_test_setup_memory  is
	generic (tag_length: integer := 2);
	port ( 

		read_write_bar_0 : in std_logic_vector (0 downto 0);
		enable_0 : in std_logic_vector (0 downto 0);
		byte_mask_0  : in std_logic_vector (7 downto 0);
		address_0    : in  std_logic_vector (11 downto 0); -- 8kwords.
		datain_0 : in std_logic_vector (63 downto 0);
		dataout_0  : out  std_logic_vector (63 downto 0);
		read_write_bar_1 : in std_logic_vector (0 downto 0);
		enable_1 : in std_logic_vector (0 downto 0);
		byte_mask_1  : in std_logic_vector (7 downto 0);
		address_1    : in  std_logic_vector (11 downto 0); -- 8kwords.
		datain_1 : in std_logic_vector (63 downto 0);
		dataout_1  : out  std_logic_vector (63 downto 0);
 	   	tag_in: in std_logic_vector(tag_length-1 downto 0);
      	   	tag_out: out std_logic_vector(tag_length-1 downto 0);
		clk, reset: in std_logic;
		start_req: in std_logic;
		start_ack: out std_logic;
		fin_req: in std_logic;
		fin_ack: out std_logic
	     );
   end component cpu_test_setup_memory;
   component cpu_test_setup_memory_dcache  is
	generic (tag_length: integer := 2);
	port ( 
		read_write_bar : in std_logic_vector (0 downto 0);
		enable : in std_logic_vector (0 downto 0);
		byte_mask  : in std_logic_vector (7 downto 0);
		address    : in  std_logic_vector (12 downto 0); -- 16kwords.
		datain : in std_logic_vector (63 downto 0);
		dataout  : out  std_logic_vector (63 downto 0);
 	   	tag_in: in std_logic_vector(tag_length-1 downto 0);
      	   	tag_out: out std_logic_vector(tag_length-1 downto 0);
		clk, reset: in std_logic;
		start_req: in std_logic;
		start_ack: out std_logic;
		fin_req: in std_logic;
		fin_ack: out std_logic
	     );
   end component  cpu_test_setup_memory_dcache;

   component cpu_test_setup_memory_icache  is
	generic (tag_length: integer := 2);
	port ( 
		read_write_bar : in std_logic_vector (0 downto 0);
		enable : in std_logic_vector (0 downto 0);
		byte_mask  : in std_logic_vector (7 downto 0);
		address    : in  std_logic_vector (12 downto 0); -- 16kwords.
		datain : in std_logic_vector (63 downto 0);
		dataout  : out  std_logic_vector (63 downto 0);
 	   	tag_in: in std_logic_vector(tag_length-1 downto 0);
      	   	tag_out: out std_logic_vector(tag_length-1 downto 0);
		clk, reset: in std_logic;
		start_req: in std_logic;
		start_ack: out std_logic;
		fin_req: in std_logic;
		fin_ack: out std_logic
	     );
   end component cpu_test_setup_memory_icache;

   component cpu_test_setup_memory_Operator  is
	port ( 

		read_write_bar_0 : in std_logic_vector (0 downto 0);
		enable_0 : in std_logic_vector (0 downto 0);
		byte_mask_0  : in std_logic_vector (7 downto 0);
		address_0    : in  std_logic_vector (11 downto 0); -- 8kwords.
		datain_0 : in std_logic_vector (63 downto 0);
		dataout_0  : out  std_logic_vector (63 downto 0);
		read_write_bar_1 : in std_logic_vector (0 downto 0);
		enable_1 : in std_logic_vector (0 downto 0);
		byte_mask_1  : in std_logic_vector (7 downto 0);
		address_1    : in  std_logic_vector (11 downto 0); -- 8kwords.
		datain_1 : in std_logic_vector (63 downto 0);
		dataout_1  : out  std_logic_vector (63 downto 0);
		clk, reset: in std_logic;
		sample_req: in boolean;
		sample_ack: out boolean;
		update_req: in boolean;
		update_ack: out boolean
	     );
   end component cpu_test_setup_memory_Operator;
   component cpu_test_setup_memory_dcache_Operator  is
	port ( 
		read_write_bar : in std_logic_vector (0 downto 0);
		enable : in std_logic_vector (0 downto 0);
		byte_mask  : in std_logic_vector (7 downto 0);
		address    : in  std_logic_vector (11 downto 0); -- 8kwords.
		datain : in std_logic_vector (63 downto 0);
		dataout  : out  std_logic_vector (63 downto 0);
		sample_req: in boolean;
		sample_ack: out boolean;
		update_req: in boolean;
		update_ack: out boolean;
		clk, reset:in std_logic
	     );
   end component cpu_test_setup_memory_dcache_Operator;
   component cpu_test_setup_memory_icache_Operator  is
	port ( 
		read_write_bar : in std_logic_vector (0 downto 0);
		enable : in std_logic_vector (0 downto 0);
		byte_mask  : in std_logic_vector (7 downto 0);
		address    : in  std_logic_vector (11 downto 0); -- 8kwords.
		datain : in std_logic_vector (63 downto 0);
		dataout  : out  std_logic_vector (63 downto 0);
		sample_req: in boolean;
		sample_ack: out boolean;
		update_req: in boolean;
		update_ack: out boolean;
		clk, reset:in std_logic
	     );
   end component cpu_test_setup_memory_icache_Operator;

   component single_port_16kX64_memory_Operator is -- 
     port ( -- 
        sample_req: in boolean;
        sample_ack: out boolean;
        update_req: in boolean;
        update_ack: out boolean;
        read : in  std_logic_vector(0 downto 0);
        -- 16K dwords..= 128KB
        addr : in  std_logic_vector(16 downto 0);
        byte_mask : in  std_logic_vector(7 downto 0);
        write_data : in  std_logic_vector(63 downto 0);
        read_data : out  std_logic_vector(63 downto 0);
        clk, reset: in std_logic);
   end component single_port_16kX64_memory_Operator;

   component mem_test_setup_memory  is
	generic (tag_length: integer := 2);
	port ( 

		read_write_bar : in std_logic_vector (0 downto 0);
		byte_mask  : in std_logic_vector (7 downto 0);
		-- 2048 x 64
		address    : in  std_logic_vector (10 downto 0);
		write_data : in std_logic_vector (63 downto 0);
		read_data  : out  std_logic_vector (63 downto 0);
 	   	tag_in: in std_logic_vector(tag_length-1 downto 0);
      	   	tag_out: out std_logic_vector(tag_length-1 downto 0);
		clk, reset: in std_logic;
		start_req: in std_logic;
		start_ack: out std_logic;
		fin_req: in std_logic;
		fin_ack: out std_logic
	     );
  end component mem_test_setup_memory;

  component icache_stub_daemon is -- 
      generic (tag_length : integer); 
  port ( -- 
    NOBLOCK_CPU_to_ICACHE_command_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_ICACHE_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_ICACHE_command_pipe_read_data : in   std_logic_vector(40 downto 0);
    ICACHE_to_CPU_response_pipe_write_req : out  std_logic_vector(0 downto 0);
    ICACHE_to_CPU_response_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ICACHE_to_CPU_response_pipe_write_data : out  std_logic_vector(89 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
  end component icache_stub_daemon;
  component dcache_stub_daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
    NOBLOCK_CPU_to_DCACHE_command_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_command_pipe_read_data : in   std_logic_vector(120 downto 0);
    NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_data : in   std_logic_vector(120 downto 0);
    DCACHE_to_CPU_response_pipe_write_req : out  std_logic_vector(0 downto 0);
    DCACHE_to_CPU_response_pipe_write_ack : in   std_logic_vector(0 downto 0);
    DCACHE_to_CPU_response_pipe_write_data : out  std_logic_vector(71 downto 0);
    DCACHE_to_CPU_slow_response_pipe_write_req : out  std_logic_vector(0 downto 0);
    DCACHE_to_CPU_slow_response_pipe_write_ack : in   std_logic_vector(0 downto 0);
    DCACHE_to_CPU_slow_response_pipe_write_data : out  std_logic_vector(71 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  end component dcache_stub_daemon;

  component dual_port_u64_mem_64KB_Operator is -- 
    port ( -- 
     sample_req: in boolean;
     sample_ack: out boolean;
     update_req: in boolean;
     update_ack: out boolean;
     read_0 : in  std_logic_vector(0 downto 0);
     addr_0 : in  std_logic_vector(12 downto 0);
     read_1 : in  std_logic_vector(0 downto 0);
     write_1 : in  std_logic_vector(0 downto 0);
     byte_mask : in  std_logic_vector(7 downto 0);
     addr_1 : in  std_logic_vector(12 downto 0);
     write_data_1 : in  std_logic_vector(63 downto 0);
     read_data_0 : out  std_logic_vector(63 downto 0);
     read_data_1 : out  std_logic_vector(63 downto 0);
     clk, reset: in std_logic
     -- 
   );
   -- 
 end component dual_port_u64_mem_64KB_Operator;
   

--------------------------------------------------------------------------------------------------
-- TLB's for MMU
--------------------------------------------------------------------------------------------------
  component accessTlbMemoryBase is -- 
  generic (address_width : integer := 8; data_width : integer := 32; use_mem_cuts: boolean := true);
  port ( -- 
    start_req: in std_logic;
    start_ack: out std_logic;
    fin_req: in std_logic;
    fin_ack: out std_logic;
    clear_flag : in  std_logic_vector(0 downto 0);
    wr_flag : in  std_logic_vector(0 downto 0);
    write_address : in  std_logic_vector(address_width-1 downto 0);
    write_entry : in  std_logic_vector(data_width-1 downto 0);
    lookup_address : in  std_logic_vector(address_width-1 downto 0);
    l_v : out  std_logic_vector(0 downto 0);
    lookup_entry : out  std_logic_vector(data_width-1 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
  end component accessTlbMemoryBase;

  component accessTlbMemoryBase_Operator is -- 
  generic (address_width : integer := 8; data_width : integer := 32; use_mem_cuts: boolean := true);
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    clear_flag : in  std_logic_vector(0 downto 0);
    wr_flag : in  std_logic_vector(0 downto 0);
    write_address : in  std_logic_vector(address_width-1 downto 0);
    write_entry : in  std_logic_vector(data_width-1 downto 0);
    lookup_address : in  std_logic_vector(address_width-1 downto 0);
    l_v : out  std_logic_vector(0 downto 0);
    lookup_entry : out  std_logic_vector(data_width-1 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
  end component accessTlbMemoryBase_Operator;

  component accessTlbMemory_0_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    clear_flag : in  std_logic_vector(0 downto 0);
    wr_flag : in  std_logic_vector(0 downto 0);
    write_address : in  std_logic_vector(0 downto 0);
    write_entry : in  std_logic_vector(46 downto 0);
    lookup_address : in  std_logic_vector(0 downto 0);
    l0_v : out  std_logic_vector(0 downto 0);
    lookup_entry : out  std_logic_vector(46 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
  end component accessTlbMemory_0_Operator;

  component accessTlbMemory_1_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    clear_flag : in  std_logic_vector(0 downto 0);
    wr_flag : in  std_logic_vector(0 downto 0);
    write_address : in  std_logic_vector(1 downto 0);
    write_entry : in  std_logic_vector(45 downto 0);
    lookup_address : in  std_logic_vector(1 downto 0);
    l1_v : out  std_logic_vector(0 downto 0);
    lookup_entry : out  std_logic_vector(45 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
  end component accessTlbMemory_1_Operator;


  component accessTlbMemory_2_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    clear_flag : in  std_logic_vector(0 downto 0);
    wr_flag : in  std_logic_vector(0 downto 0);
    write_address : in  std_logic_vector(3 downto 0);
    write_entry : in  std_logic_vector(49 downto 0);
    lookup_address : in  std_logic_vector(3 downto 0);
    l2_v : out  std_logic_vector(0 downto 0);
    lookup_entry : out  std_logic_vector(49 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
  end component accessTlbMemory_2_Operator;

  component accessTlbMemory_3_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    clear_flag : in  std_logic_vector(0 downto 0);
    wr_flag : in  std_logic_vector(0 downto 0);
    write_address : in  std_logic_vector(5 downto 0);
    write_entry : in  std_logic_vector(53 downto 0);
    lookup_address : in  std_logic_vector(5 downto 0);
    l3_v : out  std_logic_vector(0 downto 0);
    lookup_entry : out  std_logic_vector(53 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
  end component accessTlbMemory_3_Operator;

--------------------------------------------------------------------------------------------------
--  ram  for simulation
--------------------------------------------------------------------------------------------------

  component byte_ram_with_init is
   generic (name: string; g_addr_width: natural := 10);
   port (datain : in std_logic_vector(8-1 downto 0);
         dataout: out std_logic_vector(8-1 downto 0);
         addrin: in std_logic_vector(g_addr_width-1 downto 0);
         enable: in std_logic;
         writebar : in std_logic;
         clk: in std_logic;
         reset : in std_logic);
  end component byte_ram_with_init;
  component byte_ram_with_init_u64 is
   generic (name: string; g_addr_width: natural := 10);
   port (datain : in std_logic_vector(8-1 downto 0);
         dataout: out std_logic_vector(8-1 downto 0);
         addrin: in std_logic_vector(g_addr_width-1 downto 0);
         enable: in std_logic;
         writebar : in std_logic;
         clk: in std_logic;
         reset : in std_logic);
  end component byte_ram_with_init_u64;
  component dual_port_byte_ram_with_init is
   generic (byte_position: integer; g_addr_width: natural := 10; init_byte_array: ByteArray);
   port (
    	 datain_0 : in std_logic_vector(8-1 downto 0);
         dataout_0: out std_logic_vector(8-1 downto 0);
         addrin_0: in std_logic_vector(g_addr_width-1 downto 0);
         enable_0: in std_logic;
         writebar_0 : in std_logic;
    	 datain_1 : in std_logic_vector(8-1 downto 0);
         dataout_1: out std_logic_vector(8-1 downto 0);
         addrin_1: in std_logic_vector(g_addr_width-1 downto 0);
         enable_1: in std_logic;
         writebar_1 : in std_logic;
         clk: in std_logic;
         reset : in std_logic);
  end component dual_port_byte_ram_with_init;
  component single_port_byte_ram_with_init is
   generic (byte_position: integer; g_addr_width: natural := 10; init_byte_array: ByteArray);
   port (
    	 datain : in std_logic_vector(8-1 downto 0);
         dataout: out std_logic_vector(8-1 downto 0);
         addrin: in std_logic_vector(g_addr_width-1 downto 0);
         enable: in std_logic;
         writebar : in std_logic;
         clk: in std_logic;
         reset : in std_logic);
  end component single_port_byte_ram_with_init;

  component byte_ram_with_mmap_init is
   generic (mmap_file_name: string; g_addr_width: natural := 10);
   port (datain : in std_logic_vector(8-1 downto 0);
         dataout: out std_logic_vector(8-1 downto 0);
         addrin: in std_logic_vector(g_addr_width-1 downto 0);
         enable: in std_logic;
         writebar : in std_logic;
         clk: in std_logic;
         reset : in std_logic);
  end component byte_ram_with_mmap_init;

--------------------------------------------------------------------------------------------------
--  register file  
--------------------------------------------------------------------------------------------------

  component  window_update_daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      iunit_register_file_window_update_command_pipe_read_req : out  std_logic_vector(0 downto 0);
      iunit_register_file_window_update_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
      iunit_register_file_window_update_command_pipe_read_data : in   std_logic_vector(1090 downto 0);
      iunit_register_file_window_update_response_pipe_write_req : out  std_logic_vector(0 downto 0);
      iunit_register_file_window_update_response_pipe_write_ack : in   std_logic_vector(0 downto 0);
      iunit_register_file_window_update_response_pipe_write_data : out  std_logic_vector(1045 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
  end component window_update_daemon;

  component asr_daemon is -- 
    generic (tag_length : integer); 
    port ( 
      iunit_asr_access_command_pipe_read_req : out  std_logic_vector(0 downto 0);
      iunit_asr_access_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
      iunit_asr_access_command_pipe_read_data : in   std_logic_vector(43 downto 0);
      iunit_asr_access_response_pipe_write_req : out  std_logic_vector(0 downto 0);
      iunit_asr_access_response_pipe_write_ack : in   std_logic_vector(0 downto 0);
      iunit_asr_access_response_pipe_write_data : out  std_logic_vector(33 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
  end component asr_daemon;
 
			

--------------------------------------------------------------------------------------------------
--  iu operators
--------------------------------------------------------------------------------------------------
 component iu_umul32_Operator is -- 
    port ( -- 
      L : in  std_logic_vector(31 downto 0);
      R : in  std_logic_vector(31 downto 0);
      ret_val_x_x : out  std_logic_vector(63 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      sample_req : in Boolean;
      sample_ack : out Boolean;
      update_req : in Boolean;
      update_ack   : out Boolean
    );
 end component iu_umul32_Operator;

 component iu_umul32_Volatile is -- 
    port ( -- 
      L : in  std_logic_vector(31 downto 0);
      R : in  std_logic_vector(31 downto 0);
      ret_val_x_x : out  std_logic_vector(63 downto 0)
    );
 end component iu_umul32_Volatile;
 component iu_umul32 is -- 
    generic (tag_length : integer);
    port ( -- 
      L : in  std_logic_vector(31 downto 0);
      R : in  std_logic_vector(31 downto 0);
      RESULT : out  std_logic_vector(63 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
 end component iu_umul32;

 component fpunit_exec_pipe_merge_daemon is -- 
  generic (tag_length: integer);
  port ( -- 
    fpunit_exec_to_writeback_fast_pipe_read_req : out  std_logic_vector(0 downto 0);
    fpunit_exec_to_writeback_fast_pipe_read_ack : in   std_logic_vector(0 downto 0);
    fpunit_exec_to_writeback_fast_pipe_read_data : in   std_logic_vector(96-1 downto 0);
    fpunit_exec_to_writeback_slow_pipe_read_req : out  std_logic_vector(0 downto 0);
    fpunit_exec_to_writeback_slow_pipe_read_ack : in   std_logic_vector(0 downto 0);
    fpunit_exec_to_writeback_slow_pipe_read_data : in   std_logic_vector(96-1 downto 0);
    fpunit_exec_to_writeback_pipe_write_req : out  std_logic_vector(0 downto 0);
    fpunit_exec_to_writeback_pipe_write_ack : in   std_logic_vector(0 downto 0);
    fpunit_exec_to_writeback_pipe_write_data : out  std_logic_vector(96-1 downto 0);
    clk : in std_logic;
    reset : in std_logic;
    start_req: in std_logic;
    start_ack: out std_logic;
    fin_req: in std_logic;
    fin_ack: out std_logic;
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0)
  );
  -- 
  end component fpunit_exec_pipe_merge_daemon;

  component  fp_exec_in_args_mux_daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      fpunit_register_file_read_access_response_pipe_read_req : out  std_logic_vector(0 downto 0);
      fpunit_register_file_read_access_response_pipe_read_ack : in   std_logic_vector(0 downto 0);
      fpunit_register_file_read_access_response_pipe_read_data : in   std_logic_vector(172 downto 0);
      noblock_teu_idispatch_to_fpunit_exec_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_teu_idispatch_to_fpunit_exec_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_teu_idispatch_to_fpunit_exec_pipe_read_data : in   std_logic_vector(65 downto 0);
      noblock_fp_exec_in_args_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_fp_exec_in_args_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_fp_exec_in_args_pipe_write_data : out  std_logic_vector(238 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
  -- 
  end component fp_exec_in_args_mux_daemon;

  component mul53_Operator is -- 
   port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    L : in  std_logic_vector(52 downto 0);
    R : in  std_logic_vector(52 downto 0);
    RESULT : out  std_logic_vector(105 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
  end component mul53_Operator;
  component mul53 is -- 
    generic (tag_length : integer);
    port ( -- 
      L : in  std_logic_vector(52 downto 0);
      R : in  std_logic_vector(52 downto 0);
      RESULT : out  std_logic_vector(105 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
  end component mul53;

  component mul53_deterministic_pipeline_operator is -- 
    port ( -- 
      L : in  std_logic_vector(52 downto 0);
      R : in  std_logic_vector(52 downto 0);
      RESULT : out  std_logic_vector(105 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      enable : in std_logic;
      stall   : in std_logic_vector(1 to 1)
    );
  end component mul53_deterministic_pipeline_operator;

  component mul24_Operator is -- 
   port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    L : in  std_logic_vector(23 downto 0);
    R : in  std_logic_vector(23 downto 0);
    RESULT : out  std_logic_vector(47 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
  end component mul24_Operator;
  component mul24 is -- 
    generic (tag_length : integer);
    port ( -- 
      L : in  std_logic_vector(23 downto 0);
      R : in  std_logic_vector(23 downto 0);
      RESULT : out  std_logic_vector(47 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
  end component mul24;

  component mul24_deterministic_pipeline_operator is -- 
    port ( -- 
      L : in  std_logic_vector(23 downto 0);
      R : in  std_logic_vector(23 downto 0);
      RESULT : out  std_logic_vector(47 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      enable : in std_logic;
      stall   : in std_logic_vector(1 to 1)
    );
  end component mul24_deterministic_pipeline_operator;


  component fp_umul27_Volatile is -- 
    port ( -- 
      L : in  std_logic_vector(26 downto 0);
      R : in  std_logic_vector(26 downto 0);
      ret_val_x_x : out  std_logic_vector(53 downto 0)
    );
  end component fp_umul27_Volatile;

  component load_store_router_daemon is -- 
    generic (tag_length : integer := 1); 
   port ( -- 
    DCACHE_to_CPU_response_pipe_read_req : out  std_logic_vector(0 downto 0);
    DCACHE_to_CPU_response_pipe_read_ack : in   std_logic_vector(0 downto 0);
    DCACHE_to_CPU_response_pipe_read_data : in   std_logic_vector(71 downto 0);
    load_store_messy_to_router_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    load_store_messy_to_router_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    load_store_messy_to_router_pipe_pipe_read_data : in   std_logic_vector(97 downto 0);
    load_store_router_control_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    load_store_router_control_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    load_store_router_control_pipe_pipe_read_data : in   std_logic_vector(96 downto 0);
    teu_loadstore_to_fpunit_pipe_write_req : out  std_logic_vector(0 downto 0);
    teu_loadstore_to_fpunit_pipe_write_ack : in   std_logic_vector(0 downto 0);
    teu_loadstore_to_fpunit_pipe_write_data : out  std_logic_vector(77 downto 0);
    teu_loadstore_to_iretire_pipe_write_req : out  std_logic_vector(0 downto 0);
    teu_loadstore_to_iretire_pipe_write_ack : in   std_logic_vector(0 downto 0);
    teu_loadstore_to_iretire_pipe_write_data : out  std_logic_vector(53 downto 0);
    teu_loadstore_to_iunit_pipe_write_req : out  std_logic_vector(0 downto 0);
    teu_loadstore_to_iunit_pipe_write_ack : in   std_logic_vector(0 downto 0);
    teu_loadstore_to_iunit_pipe_write_data : out  std_logic_vector(77 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
  end component load_store_router_daemon;

  component load_store_router_reworked_daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      DCACHE_to_CPU_response_pipe_read_req : out  std_logic_vector(0 downto 0);
      DCACHE_to_CPU_response_pipe_read_ack : in   std_logic_vector(0 downto 0);
      DCACHE_to_CPU_response_pipe_read_data : in   std_logic_vector(71 downto 0);
      load_store_messy_to_router_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      load_store_messy_to_router_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      load_store_messy_to_router_pipe_pipe_read_data : in   std_logic_vector(97 downto 0);
      noblock_load_store_router_control_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_load_store_router_control_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_load_store_router_control_pipe_pipe_read_data : in   std_logic_vector(99 downto 0);
      teu_loadstore_to_fpunit_pipe_write_req : out  std_logic_vector(0 downto 0);
      teu_loadstore_to_fpunit_pipe_write_ack : in   std_logic_vector(0 downto 0);
      teu_loadstore_to_fpunit_pipe_write_data : out  std_logic_vector(77 downto 0);
      teu_loadstore_to_iretire_pipe_write_req : out  std_logic_vector(0 downto 0);
      teu_loadstore_to_iretire_pipe_write_ack : in   std_logic_vector(0 downto 0);
      teu_loadstore_to_iretire_pipe_write_data : out  std_logic_vector(53 downto 0);
      teu_loadstore_to_iunit_pipe_write_req : out  std_logic_vector(0 downto 0);
      teu_loadstore_to_iunit_pipe_write_ack : in   std_logic_vector(0 downto 0);
      teu_loadstore_to_iunit_pipe_write_data : out  std_logic_vector(77 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component load_store_router_reworked_daemon;

  component sc_iretire_join_daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      noblock_teu_stream_corrector_to_idispatch_pipe_read_req : out  std_logic_vector(0 downto 0);
      noblock_teu_stream_corrector_to_idispatch_pipe_read_ack : in   std_logic_vector(0 downto 0);
      noblock_teu_stream_corrector_to_idispatch_pipe_read_data : in   std_logic_vector(147 downto 0);
      teu_iretire_to_idispatch_pipe_read_req : out  std_logic_vector(0 downto 0);
      teu_iretire_to_idispatch_pipe_read_ack : in   std_logic_vector(0 downto 0);
      teu_iretire_to_idispatch_pipe_read_data : in   std_logic_vector(0 downto 0);
      noblock_joined_iretire_sc_to_idispatch_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_joined_iretire_sc_to_idispatch_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_joined_iretire_sc_to_idispatch_pipe_write_data : out  std_logic_vector(147 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
  -- 
  end component sc_iretire_join_daemon;
  
  component iunit_writeback_in_mux_daemon is -- 
    generic (tag_length : integer); 
  -- 
  port ( -- 
    iunit_exec_fast_alu_result_to_writeback_pipe_read_req : out  std_logic_vector(0 downto 0);
    iunit_exec_fast_alu_result_to_writeback_pipe_read_ack : in   std_logic_vector(0 downto 0);
    iunit_exec_fast_alu_result_to_writeback_pipe_read_data : in   std_logic_vector(108 downto 0);
    iunit_exec_to_writeback_pipe_read_req : out  std_logic_vector(0 downto 0);
    iunit_exec_to_writeback_pipe_read_ack : in   std_logic_vector(0 downto 0);
    iunit_exec_to_writeback_pipe_read_data : in   std_logic_vector(125 downto 0);
    noblock_teu_idispatch_to_iunit_writeback_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_teu_idispatch_to_iunit_writeback_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_teu_idispatch_to_iunit_writeback_pipe_read_data : in   std_logic_vector(83 downto 0);
    teu_fpunit_trap_to_iunit_pipe_read_req : out  std_logic_vector(0 downto 0);
    teu_fpunit_trap_to_iunit_pipe_read_ack : in   std_logic_vector(0 downto 0);
    teu_fpunit_trap_to_iunit_pipe_read_data : in   std_logic_vector(12 downto 0);
    teu_loadstore_to_iunit_pipe_read_req : out  std_logic_vector(0 downto 0);
    teu_loadstore_to_iunit_pipe_read_ack : in   std_logic_vector(0 downto 0);
    teu_loadstore_to_iunit_pipe_read_data : in   std_logic_vector(77 downto 0);
    teu_stream_corrector_to_iunit_pipe_read_req : out  std_logic_vector(0 downto 0);
    teu_stream_corrector_to_iunit_pipe_read_ack : in   std_logic_vector(0 downto 0);
    teu_stream_corrector_to_iunit_pipe_read_data : in   std_logic_vector(17 downto 0);
    noblock_iunit_writeback_in_args_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_iunit_writeback_in_args_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_iunit_writeback_in_args_pipe_pipe_write_data : out  std_logic_vector(372 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  end component iunit_writeback_in_mux_daemon;
 
  component iunit_writeback_in_mux_ajit_64_daemon is -- 
   generic (tag_length : integer); 
   port ( -- 
    iunit_64_exec_fast_alu_result_to_writeback_pipe_read_req : out  std_logic_vector(0 downto 0);
    iunit_64_exec_fast_alu_result_to_writeback_pipe_read_ack : in   std_logic_vector(0 downto 0);
    iunit_64_exec_fast_alu_result_to_writeback_pipe_read_data : in   std_logic_vector(140 downto 0);
    iunit_64_exec_to_writeback_pipe_read_req : out  std_logic_vector(0 downto 0);
    iunit_64_exec_to_writeback_pipe_read_ack : in   std_logic_vector(0 downto 0);
    iunit_64_exec_to_writeback_pipe_read_data : in   std_logic_vector(157 downto 0);
    noblock_teu_idispatch_to_iunit_writeback_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_teu_idispatch_to_iunit_writeback_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_teu_idispatch_to_iunit_writeback_pipe_read_data : in   std_logic_vector(83 downto 0);
    teu_fpunit_trap_to_iunit_pipe_read_req : out  std_logic_vector(0 downto 0);
    teu_fpunit_trap_to_iunit_pipe_read_ack : in   std_logic_vector(0 downto 0);
    teu_fpunit_trap_to_iunit_pipe_read_data : in   std_logic_vector(12 downto 0);
    teu_loadstore_to_iunit_pipe_read_req : out  std_logic_vector(0 downto 0);
    teu_loadstore_to_iunit_pipe_read_ack : in   std_logic_vector(0 downto 0);
    teu_loadstore_to_iunit_pipe_read_data : in   std_logic_vector(77 downto 0);
    teu_stream_corrector_to_iunit_pipe_read_req : out  std_logic_vector(0 downto 0);
    teu_stream_corrector_to_iunit_pipe_read_ack : in   std_logic_vector(0 downto 0);
    teu_stream_corrector_to_iunit_pipe_read_data : in   std_logic_vector(17 downto 0);
    noblock_iunit_64_writeback_in_args_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_iunit_64_writeback_in_args_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_iunit_64_writeback_in_args_pipe_pipe_write_data : out  std_logic_vector(436 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
   );
  end component iunit_writeback_in_mux_ajit_64_daemon;

  component interrupt_stub_daemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      INTR_LEVEL : in std_logic_vector(3 downto 0);
      ENV_to_CPU_irl_pipe_write_req : out  std_logic_vector(0 downto 0);
      ENV_to_CPU_irl_pipe_write_ack : in   std_logic_vector(0 downto 0);
      ENV_to_CPU_irl_pipe_write_data : out  std_logic_vector(7 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
  -- 
  end component interrupt_stub_daemon;

  component stream_corrector_in_mux_daemon is -- 
   generic (tag_length : integer := 1); 
   port ( -- 
    teu_idispatch_to_stream_corrector_pipe_read_req : out  std_logic_vector(0 downto 0);
    teu_idispatch_to_stream_corrector_pipe_read_ack : in   std_logic_vector(0 downto 0);
    teu_idispatch_to_stream_corrector_pipe_read_data : in   std_logic_vector(203 downto 0);
    teu_fpunit_cc_to_stream_corrector_pipe_read_req : out  std_logic_vector(0 downto 0);
    teu_fpunit_cc_to_stream_corrector_pipe_read_ack : in   std_logic_vector(0 downto 0);
    teu_fpunit_cc_to_stream_corrector_pipe_read_data : in   std_logic_vector(14 downto 0);
    teu_iunit_cc_to_stream_corrector_pipe_read_req : out  std_logic_vector(0 downto 0);
    teu_iunit_cc_to_stream_corrector_pipe_read_ack : in   std_logic_vector(0 downto 0);
    teu_iunit_cc_to_stream_corrector_pipe_read_data : in   std_logic_vector(16 downto 0);
    teu_iunit_to_stream_corrector_pipe_read_req : out  std_logic_vector(0 downto 0);
    teu_iunit_to_stream_corrector_pipe_read_ack : in   std_logic_vector(0 downto 0);
    teu_iunit_to_stream_corrector_pipe_read_data : in   std_logic_vector(89 downto 0);
    noblock_stream_corrector_in_args_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_stream_corrector_in_args_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_stream_corrector_in_args_pipe_write_data : out  std_logic_vector(326 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
  end component stream_corrector_in_mux_daemon;
  
  component stream_corrector_in_mux_daemon_v2 is -- 
    generic (tag_length : integer := 1); 
    port ( -- 
      teu_idispatch_to_stream_corrector_pipe_read_req : out  std_logic_vector(0 downto 0);
      teu_idispatch_to_stream_corrector_pipe_read_ack : in   std_logic_vector(0 downto 0);
      teu_idispatch_to_stream_corrector_pipe_read_data : in   std_logic_vector(204 downto 0);
      teu_fpunit_cc_to_stream_corrector_pipe_read_req : out  std_logic_vector(0 downto 0);
      teu_fpunit_cc_to_stream_corrector_pipe_read_ack : in   std_logic_vector(0 downto 0);
      teu_fpunit_cc_to_stream_corrector_pipe_read_data : in   std_logic_vector(14 downto 0);
      teu_iunit_cc_to_stream_corrector_pipe_read_req : out  std_logic_vector(0 downto 0);
      teu_iunit_cc_to_stream_corrector_pipe_read_ack : in   std_logic_vector(0 downto 0);
      teu_iunit_cc_to_stream_corrector_pipe_read_data : in   std_logic_vector(16 downto 0);
      teu_iunit_rs1_to_stream_corrector_pipe_read_req : out  std_logic_vector(0 downto 0);
      teu_iunit_rs1_to_stream_corrector_pipe_read_ack : in   std_logic_vector(0 downto 0);
      teu_iunit_rs1_to_stream_corrector_pipe_read_data : in   std_logic_vector(31 downto 0);
      teu_iunit_to_stream_corrector_pipe_read_req : out  std_logic_vector(0 downto 0);
      teu_iunit_to_stream_corrector_pipe_read_ack : in   std_logic_vector(0 downto 0);
      teu_iunit_to_stream_corrector_pipe_read_data : in   std_logic_vector(89 downto 0);
      noblock_stream_corrector_in_args_pipe_write_req : out  std_logic_vector(0 downto 0);
      noblock_stream_corrector_in_args_pipe_write_ack : in   std_logic_vector(0 downto 0);
      noblock_stream_corrector_in_args_pipe_write_data : out  std_logic_vector(359 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
  -- 
  end component stream_corrector_in_mux_daemon_v2;


  component bpbV2_Operator is
    port ( 
      sample_req: in boolean;
      sample_ack: out boolean;
      update_req: in boolean;
      update_ack: out boolean;
      bpb_init : in  std_logic_vector(0 downto 0);
      add_entry : in  std_logic_vector(0 downto 0);
      add_pc : in  std_logic_vector(31 downto 0);
      add_nnpc : in  std_logic_vector(31 downto 0);
      lookup_pc : in  std_logic_vector(31 downto 0);
      bpb_result : out  std_logic_vector(32 downto 0);
      clk, reset: in std_logic
  );
  end component bpbV2_Operator;

  component bpbV3_dual_port_mem_Operator is -- 
  port ( -- 
    init : in  std_logic_vector(0 downto 0);
    enable_0 : in  std_logic_vector(0 downto 0);
    addr_0 : in  std_logic_vector(7 downto 0);
    enable_1 : in  std_logic_vector(0 downto 0);
    write_bar_1 : in  std_logic_vector(0 downto 0);
    addr_1 : in  std_logic_vector(7 downto 0);
    write_data_1 : in  std_logic_vector(53 downto 0);
    read_data : out  std_logic_vector(109 downto 0);
    clk : in std_logic;
    reset : in std_logic;
    sample_req : in Boolean;
    sample_ack : out Boolean;
    update_req : in Boolean;
    update_ack   : out Boolean-- 
  );
  -- 
  end component bpbV3_dual_port_mem_Operator;

  component ibuf_cache_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    ibuf_cache_init : in  std_logic_vector(0 downto 0);
    add_entry : in  std_logic_vector(0 downto 0);
    add_pc : in  std_logic_vector(31 downto 0);
    add_acc : in  std_logic_vector(2 downto 0);
    add_ipair : in  std_logic_vector(63 downto 0);
    lookup_S : in  std_logic_vector(0 downto 0);
    lookup_pc : in  std_logic_vector(31 downto 0);
    ibuf_cache_result : out  std_logic_vector(64 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
  end component ibuf_cache_Operator;

  component ras_daemon is -- 
  generic (tag_length : integer := 1); 
  port ( -- 
    teu_ras_access_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    teu_ras_access_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    teu_ras_access_pipe_pipe_read_data : in   std_logic_vector(32 downto 0);
    teu_ras_top_of_stack_pipe_write_req : out  std_logic_vector(0 downto 0);
    teu_ras_top_of_stack_pipe_write_ack : in   std_logic_vector(0 downto 0);
    teu_ras_top_of_stack_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
  end component ras_daemon;
  
  component asr_update_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    core_id: in std_logic_vector(7 downto 0);
    thread_id: in std_logic_vector(7 downto 0);
    access_cmd : in  std_logic_vector(43 downto 0);
    read_val : out  std_logic_vector(31 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
 end component asr_update_Operator;

 component asr_update_64_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    core_id: in std_logic_vector(7 downto 0);
    thread_id: in std_logic_vector(7 downto 0);
    access_cmd : in  std_logic_vector(43 downto 0);
    read_val : out  std_logic_vector(31 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
 end component asr_update_64_Operator;

 component asr_update_core is -- 
  port ( -- 
    core_id: in std_logic_vector(7 downto 0);
    thread_id: in std_logic_vector(7 downto 0);
    access_cmd : in  std_logic_vector(43 downto 0);
    read_val : out  std_logic_vector(31 downto 0);
    clk, reset: in std_logic;
    trigger : in boolean
  );
  -- 
 end component asr_update_core;

 component window_update_core is -- 
  port ( -- 
    incoming_outs, incoming_locals, incoming_ins : in  std_logic_vector(255 downto 0);
    save, restore, write_psr: in std_logic;
    rd: in std_logic_vector(4 downto 0);
    rd_val: in std_logic_vector(31 downto 0);
    old_cwp, new_cwp : in std_logic_vector(4 downto 0);
    outgoing_outs, outgoing_locals, outgoing_ins : out  std_logic_vector(255 downto 0);
    outgoing_cwp : out std_logic_vector(4 downto 0);
    clk : in std_logic;                                
    reset : in std_logic;
    trigger : in boolean; 
    done    : out boolean;
    latch_locals, latch_outs, latch_ins, latch_outgoing_cwp: out boolean
  );
  -- 
 end component window_update_core; 

 component update_registers_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    next_registers : in  std_logic_vector(1023 downto 0);
    window_update_command : in  std_logic_vector(50 downto 0);
    new_cwp_and_updated_registers : out  std_logic_vector(1028 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
 end component update_registers_Operator;

  component window_address_calculator_Volatile is -- 
  port ( -- 
    cwp : in  std_logic_vector(4 downto 0);
    reg_id : in  std_logic_vector(4 downto 0);
    reg_address : out  std_logic_vector(5 downto 0)-- 
  );
  -- 
  end component window_address_calculator_Volatile;

  component window_registers_bank
	generic (name : string := "anon");
	port (trigger: in boolean; 
		write_enable_0: in std_logic;
		address_0, address_1: in std_logic_vector(5 downto 0);
		read_data_1 : out std_logic_vector(31 downto 0);
		write_data_0: in std_logic_vector(31 downto 0);
		clk, reset: in std_logic);
  end component window_registers_bank;

  component iu_registers_3r_1w_port_register_file_inner is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    rs1 : in  std_logic_vector(4 downto 0);
    rs2 : in  std_logic_vector(4 downto 0);
    read_rd : in  std_logic_vector(4 downto 0);
    read_cwp : in  std_logic_vector(4 downto 0);
    write_gpr_even : in  std_logic_vector(0 downto 0);
    write_gpr_odd : in  std_logic_vector(0 downto 0);
    write_rd : in  std_logic_vector(4 downto 0);
    write_gpr_value_even : in  std_logic_vector(31 downto 0);
    write_gpr_value_odd : in  std_logic_vector(31 downto 0);
    write_cwp : in  std_logic_vector(4 downto 0);
    reg_pair_values : out  std_logic_vector(191 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
  end component iu_registers_3r_1w_port_register_file_inner;

  component iu_registers_3r_1w_port_register_file_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    rs1 : in  std_logic_vector(4 downto 0);
    rs2 : in  std_logic_vector(4 downto 0);
    read_rd : in  std_logic_vector(4 downto 0);
    read_cwp : in  std_logic_vector(4 downto 0);
    write_gpr_even : in  std_logic_vector(0 downto 0);
    write_gpr_odd : in  std_logic_vector(0 downto 0);
    write_rd : in  std_logic_vector(4 downto 0);
    write_gpr_value_even : in  std_logic_vector(31 downto 0);
    write_gpr_value_odd : in  std_logic_vector(31 downto 0);
    write_cwp : in  std_logic_vector(4 downto 0);
    reg_pair_values : out  std_logic_vector(191 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
  end component iu_registers_3r_1w_port_register_file_Operator;

 -- NOTE: only for simulations.
 component dual_port_u64_mem_with_init_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    first_time : in  std_logic_vector(0 downto 0);
    read_0 : in  std_logic_vector(0 downto 0);
    addr_0 : in  std_logic_vector(28 downto 0);
    read_1 : in  std_logic_vector(0 downto 0);
    write_1 : in  std_logic_vector(0 downto 0);
    byte_mask : in  std_logic_vector(7 downto 0);
    addr_1 : in  std_logic_vector(28 downto 0);
    write_data_1 : in  std_logic_vector(63 downto 0);
    read_data_0 : out  std_logic_vector(63 downto 0);
    read_data_1 : out  std_logic_vector(63 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
  end component dual_port_u64_mem_with_init_Operator;

  component single_port_u64_mem_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    read : in  std_logic_vector(0 downto 0);
    -- 8K dwords..= 64KB
    addr : in  std_logic_vector(12 downto 0);
    byte_mask : in  std_logic_vector(7 downto 0);
    write_data : in  std_logic_vector(63 downto 0);
    read_data : out  std_logic_vector(63 downto 0);
    clk, reset: in std_logic
  );
  end component single_port_u64_mem_Operator;



  component mmuDcacheServiceDaemon is -- 
   generic (tag_length : integer); 
   port ( -- 
    DCACHE_to_MMU_request_pipe_read_req : out  std_logic_vector(0 downto 0);
    DCACHE_to_MMU_request_pipe_read_ack : in   std_logic_vector(0 downto 0);
    DCACHE_to_MMU_request_pipe_read_data : in   std_logic_vector(119 downto 0);
    NOBLOCK_DCACHE_TO_MMU_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_DCACHE_TO_MMU_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_DCACHE_TO_MMU_REQUEST_pipe_write_data : out  std_logic_vector(121 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
  end component;

  component mmuIcacheServiceDaemon is -- 
   generic (tag_length : integer); 
   port ( -- 
    ICACHE_to_MMU_request_pipe_read_req : out  std_logic_vector(0 downto 0);
    ICACHE_to_MMU_request_pipe_read_ack : in   std_logic_vector(0 downto 0);
    ICACHE_to_MMU_request_pipe_read_data : in   std_logic_vector(47 downto 0);
    NOBLOCK_ICACHE_TO_MMU_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_ICACHE_TO_MMU_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_ICACHE_TO_MMU_REQUEST_pipe_write_data : out  std_logic_vector(121 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  end component;

  component mmuMuxDaemon is -- 
   generic (tag_length : integer); 
   port ( -- 
    NOBLOCK_DCACHE_TO_MMU_REQUEST_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_DCACHE_TO_MMU_REQUEST_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_DCACHE_TO_MMU_REQUEST_pipe_read_data : in   std_logic_vector(121 downto 0);
    NOBLOCK_ICACHE_TO_MMU_REQUEST_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_ICACHE_TO_MMU_REQUEST_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_ICACHE_TO_MMU_REQUEST_pipe_read_data : in   std_logic_vector(121 downto 0);
    NOBLOCK_CACHE_TO_MMU_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_CACHE_TO_MMU_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_CACHE_TO_MMU_REQUEST_pipe_write_data : out  std_logic_vector(121 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
  end component mmuMuxDaemon;

  -- a generic fully associative memory for use in the MMU TLB.
  component genericFullyAssociativeMemory is
	generic (tag_width: integer := 8;
			data_width: integer := 32;
			log_number_of_entries: integer := 6;
			ignore_collisions: boolean := true;
			use_mem_cuts: boolean:= true);
	port (  start_req: in std_logic;
		start_ack: out std_logic;
		fin_req: in std_logic;
		fin_ack: out std_logic;

		-- clear all valids.
		clear_flag: in std_logic_vector(0 downto 0);

		-- add entry
		write_flag: in std_logic_vector(0 downto 0);
		write_data: in std_logic_vector(data_width-1 downto 0);
		write_tag : in std_logic_vector(tag_width-1 downto 0);

		-- lookup entry
		erase_flag: in std_logic_vector(0 downto 0);
		lookup_flag: in std_logic_vector(0 downto 0);
		lookup_tag : in std_logic_vector(tag_width-1 downto 0);
		lookup_valid: out std_logic_vector(0 downto 0);
		lookup_data: out std_logic_vector(data_width-1 downto 0);

		clk,reset: in std_logic);

  end component genericFullyAssociativeMemory;

	

  -- a generic fully associative memory for use in the MMU TLB.
  component genericFullyAssociativeMemory_Operator is
	generic (tag_width: integer := 8;
			data_width: integer := 32;
			log_number_of_entries: integer := 6;
			ignore_collisions: boolean := true;
			use_mem_cuts: boolean:= true);
	port (  sample_req: in boolean;
		sample_ack: out boolean;
		update_req: in boolean;
		update_ack: out boolean;

		-- clear all valids.
		clear_flag: in std_logic_vector(0 downto 0);

		-- add entry
		write_flag: in std_logic_vector(0 downto 0);
		write_data: in std_logic_vector(data_width-1 downto 0);
		write_tag : in std_logic_vector(tag_width-1 downto 0);

		-- lookup entry
		erase_flag: in std_logic_vector(0 downto 0);
		lookup_flag: in std_logic_vector(0 downto 0);
		lookup_tag : in std_logic_vector(tag_width-1 downto 0);
		lookup_valid: out std_logic_vector(0 downto 0);
		lookup_data: out std_logic_vector(data_width-1 downto 0);

		clk,reset: in std_logic);

   end component genericFullyAssociativeMemory_Operator;
   component genericFullyAssociativeMemoryNoData is
	generic (tag_width: integer := 8; log_number_of_entries: integer := 6; ignore_collisions: boolean := true);
	port (  start_req: in std_logic;
		start_ack: out std_logic;
		fin_req: in std_logic;
		fin_ack: out std_logic;

		-- clear all valids.
		clear_flag: in std_logic_vector(0 downto 0);

		-- add entry
		erase_flag: in std_logic_vector(0 downto 0);
		write_flag: in std_logic_vector(0 downto 0);
		write_tag : in std_logic_vector(tag_width-1 downto 0);

		-- lookup entry
		lookup_flag: in std_logic_vector(0 downto 0);
		lookup_tag : in std_logic_vector(tag_width-1 downto 0);
		lookup_valid: out std_logic_vector(0 downto 0);

		clk,reset: in std_logic);

    end component genericFullyAssociativeMemoryNoData;
    component genericFullyAssociativeMemoryNoData_Operator is
	generic (tag_width: integer := 8; log_number_of_entries: integer := 6; ignore_collisions: boolean := true);
	port (  sample_req: in boolean;
		sample_ack: out boolean;
		update_req: in boolean;
		update_ack: out boolean;

		-- clear all valids.
		clear_flag: in std_logic_vector(0 downto 0);

		-- add entry
		erase_flag: in std_logic_vector(0 downto 0);
		write_flag: in std_logic_vector(0 downto 0);
		write_tag : in std_logic_vector(tag_width-1 downto 0);

		-- lookup entry
		lookup_flag: in std_logic_vector(0 downto 0);
		lookup_tag : in std_logic_vector(tag_width-1 downto 0);
		lookup_valid: out std_logic_vector(0 downto 0);

		clk,reset: in std_logic);

    end component genericFullyAssociativeMemoryNoData_Operator;


  -- a generic set associative memory for potential use in the MMU TLB.
  --   This could probably be used in the caches as well..
  component genericSetAssociativeMemory is
	generic (
			-- width of tag.
			tag_width: integer := 8;
			-- width of data.
			data_width: integer := 32;
			-- size of the set associative memory is 2**log_number_of_entries
			log_number_of_entries: integer := 8;
			-- 0 means direct mapped.
			log_associativity: integer := 0;
			-- ignore write->lookup collisions
			ignore_collisions: boolean := true;
			-- use memory cuts or registers?
			use_mem_cuts: boolean:= true;
			-- ignore data
			g_ignore_data: boolean := false);
	port (  start_req: in std_logic;
		start_ack: out std_logic;
		fin_req: in std_logic;
		fin_ack: out std_logic;

		-- clear all valids.
		clear_flag: in std_logic_vector(0 downto 0);

		-- add/erase entry specified by write_* ports.
		erase_flag: in std_logic_vector(0 downto 0);
		write_flag: in std_logic_vector(0 downto 0);
		
		-- write data 
		write_data: in std_logic_vector(data_width-1 downto 0);
		-- write tag (computed by environment)
		write_tag : in std_logic_vector(tag_width-1 downto 0);
		-- write set id (specified by environment)
		write_set_id: in std_logic_vector((log_number_of_entries-log_associativity)-1 downto 0);

		-- lookup entry
		lookup_flag: in std_logic_vector(0 downto 0);
		-- lookup tag.
		lookup_tag : in std_logic_vector(tag_width-1 downto 0);
		-- lookup set id.
		lookup_set_id: in std_logic_vector((log_number_of_entries-log_associativity)-1 downto 0);
		-- lookup is valid.. hit.
		lookup_valid: out std_logic_vector(0 downto 0);
		-- lookup data.
		lookup_data: out std_logic_vector(data_width-1 downto 0);
		clk,reset: in std_logic);

  end component genericSetAssociativeMemory;

  -- operator form of generic set associative memory for potential use in the MMU TLB.
  --   This could probably be used in the caches as well..
  component genericSetAssociativeMemory_Operator is
	generic (
			-- width of tag.
			tag_width: integer := 8;
			-- width of data.
			data_width: integer := 32;
			-- size of the set associative memory is 2**log_number_of_entries
			log_number_of_entries: integer := 8;
			-- 0 means direct mapped.
			log_associativity: integer := 0;
			-- ignore write->lookup collisions
			ignore_collisions: boolean := true;
			-- use memory cuts or registers?
			use_mem_cuts: boolean:= true;
			-- ignore data, behave like a set and not a map.
			g_ignore_data: boolean := false);
	port (  sample_req: in boolean;
		sample_ack: out boolean;
		update_req: in boolean;
		update_ack: out boolean;

		-- clear all valids.
		clear_flag: in std_logic_vector(0 downto 0);

		-- add/erase entry specified by write_* ports.
		erase_flag: in std_logic_vector(0 downto 0);
		write_flag: in std_logic_vector(0 downto 0);
		
		-- write data 
		write_data: in std_logic_vector(data_width-1 downto 0);
		-- write tag (computed by environment)
		write_tag : in std_logic_vector(tag_width-1 downto 0);
		-- write set id (specified by environment)
		write_set_id: in std_logic_vector((log_number_of_entries-log_associativity)-1 downto 0);

		-- lookup entry
		lookup_flag: in std_logic_vector(0 downto 0);
		-- lookup tag.
		lookup_tag : in std_logic_vector(tag_width-1 downto 0);
		-- lookup set id.
		lookup_set_id: in std_logic_vector((log_number_of_entries-log_associativity)-1 downto 0);
		-- lookup is valid.. hit.
		lookup_valid: out std_logic_vector(0 downto 0);
		-- lookup data.
		lookup_data: out std_logic_vector(data_width-1 downto 0);
		clk,reset: in std_logic);

  end component genericSetAssociativeMemory_Operator;

 
  -- direct mapped, single cycle for write and read...
  component genericDirectMappedAssociativeMemory is -- 
  generic (tag_width: integer := 32;
		data_width: integer := 67;
		log2_number_of_entries : integer := 8);
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    init_flag : in  std_logic_vector(0 downto 0);
    insert_flag : in  std_logic_vector(0 downto 0);
    insert_tag : in  std_logic_vector(tag_width-1 downto 0);
    insert_data : in  std_logic_vector(data_width-1 downto 0);
    lookup_flag : in  std_logic_vector(0 downto 0);
    lookup_tag : in  std_logic_vector(tag_width-1 downto 0);
    lookup_match : out  std_logic_vector(0 downto 0);
    lookup_data : out  std_logic_vector(data_width-1 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
  end component genericDirectMappedAssociativeMemory;

  component accessTlbNewMemory_0_Operator is
    port ( -- 
    	sample_req: in boolean;
    	sample_ack: out boolean;
    	update_req: in boolean;
    	update_ack: out boolean;
	clear: in std_logic_vector(0 downto 0);
	write: in std_logic_vector(0 downto 0);
        write_tag:  in std_logic_vector(7 downto 0);
        write_data: in std_logic_vector(31 downto 0);
        lookup: in std_logic_vector(0 downto 0);
	lookup_tag: in std_logic_vector(7 downto 0);
        tlb_hit: out std_logic_vector(0 downto 0);
	pte: out std_logic_vector(31 downto 0);
        clk, reset: in std_logic);
  end component;

  component accessTlbNewMemory_1_Operator is
    port ( -- 
    	sample_req: in boolean;
    	sample_ack: out boolean;
    	update_req: in boolean;
    	update_ack: out boolean;
	clear: in std_logic_vector(0 downto 0);
	write: in std_logic_vector(0 downto 0);
        write_tag:  in std_logic_vector(15 downto 0);
        write_data: in std_logic_vector(31 downto 0);
        lookup: in std_logic_vector(0 downto 0);
	lookup_tag: in std_logic_vector(15 downto 0);
        tlb_hit: out std_logic_vector(0 downto 0);
	pte: out std_logic_vector(31 downto 0);
        clk, reset: in std_logic);
  end component;


  component accessTlbNewMemory_2_Operator is
    port ( -- 
    	sample_req: in boolean;
    	sample_ack: out boolean;
    	update_req: in boolean;
    	update_ack: out boolean;
	clear: in std_logic_vector(0 downto 0);
	write: in std_logic_vector(0 downto 0);
        write_tag:  in std_logic_vector(21 downto 0);
        write_data: in std_logic_vector(31 downto 0);
        lookup: in std_logic_vector(0 downto 0);
	lookup_tag: in std_logic_vector(21 downto 0);
        tlb_hit: out std_logic_vector(0 downto 0);
	pte: out std_logic_vector(31 downto 0);
        clk, reset: in std_logic);
  end component;

  component accessTlbNewMemory_3_Operator is
    port ( -- 
    	sample_req: in boolean;
    	sample_ack: out boolean;
    	update_req: in boolean;
    	update_ack: out boolean;
	clear: in std_logic_vector(0 downto 0);
	write: in std_logic_vector(0 downto 0);
        write_tag:  in std_logic_vector(27 downto 0);
        write_data: in std_logic_vector(31 downto 0);
        lookup: in std_logic_vector(0 downto 0);
	lookup_tag: in std_logic_vector(27 downto 0);
        tlb_hit: out std_logic_vector(0 downto 0);
	pte: out std_logic_vector(31 downto 0);
        clk, reset: in std_logic);
  end component;

  component memAccessRequestMergeDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      fast_mem_access_and_send_response_command_pipe_read_req : out  std_logic_vector(0 downto 0);
      fast_mem_access_and_send_response_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
      fast_mem_access_and_send_response_command_pipe_read_data : in   std_logic_vector(124 downto 0);
      slow_mem_access_and_send_response_command_pipe_read_req : out  std_logic_vector(0 downto 0);
      slow_mem_access_and_send_response_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
      slow_mem_access_and_send_response_command_pipe_read_data : in   std_logic_vector(209 downto 0);
      mem_access_and_send_response_command_pipe_write_req : out  std_logic_vector(0 downto 0);
      mem_access_and_send_response_command_pipe_write_ack : in   std_logic_vector(0 downto 0);
      mem_access_and_send_response_command_pipe_write_data : out  std_logic_vector(207 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
  end component;

  ----------------------------------------------------------------------------------------------------
  -- generic single and dual port memories.
  ----------------------------------------------------------------------------------------------------
  component genericSinglePortMemory_Operator

	generic ( data_width: integer := 32; address_width: integer := 32);
	port (sample_req: in boolean;
		sample_ack: out boolean;
		update_req: in boolean;
		update_ack: out boolean;

		enable: in std_logic_vector(0 downto 0);	
		write_bar: in std_logic_vector(0 downto 0);	
		write_data: in std_logic_vector(data_width-1 downto 0);
		read_data: out std_logic_vector(data_width-1 downto 0);
		address: in std_logic_vector(address_width-1 downto 0);

		clk,reset: in std_logic);

  end component genericSinglePortMemory_Operator;

  component genericDualPortMemory_Operator
	generic ( data_width: integer := 32; address_width: integer := 32);
	port (sample_req: in boolean;
		sample_ack: out boolean;
		update_req: in boolean;
		update_ack: out boolean;

		enable_0: in std_logic_vector(0 downto 0);	
		write_bar_0: in std_logic_vector(0 downto 0);	
		write_data_0: in std_logic_vector(data_width-1 downto 0);
		read_data_0: out std_logic_vector(data_width-1 downto 0);
		address_0: in std_logic_vector(address_width-1 downto 0);

		enable_1: in std_logic_vector(0 downto 0);	
		write_bar_1: in std_logic_vector(0 downto 0);	
		write_data_1: in std_logic_vector(data_width-1 downto 0);
		read_data_1: out std_logic_vector(data_width-1 downto 0);
		address_1: in std_logic_vector(address_width-1 downto 0);

		clk,reset: in std_logic);

  end component genericDualPortMemory_Operator;

  component accessRlutBase_Operator is -- 
    generic (
		g_LOG_BASE_PAGE_SIZE: integer;
		g_LOG_CACHE_LINE_SIZE: integer;
		g_CACHE_WAY_SIZE: integer;
		g_RLUT_TAG_WIDTH : integer;
		g_RLUT_REDUCED_DATA_WIDTH: integer;
		g_RLUT_LOG_N_SETS: integer;
		g_RLUT_LOG_MEMORY_SIZE: integer;
		g_RLUT_LOG_SET_SIZE: integer
	);
    port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    lookup : in  std_logic_vector(0 downto 0);
    update : in  std_logic_vector(0 downto 0);
    clear : in  std_logic_vector(0 downto 0);
    physical_addr_of_line : in  std_logic_vector(29 downto 0);
    virtual_addr_of_line : in  std_logic_vector(25 downto 0);
    syn_invalidate_word : out  std_logic_vector(26 downto 0);
    clk, reset: in std_logic
    -- 
  );
  end component accessRlutBase_Operator;
  
  component accessIcacheRlut_Operator is -- 
   port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    lookup : in  std_logic_vector(0 downto 0);
    update : in  std_logic_vector(0 downto 0);
    clear : in  std_logic_vector(0 downto 0);
    physical_addr_of_line : in  std_logic_vector(29 downto 0);
    virtual_addr_of_line : in  std_logic_vector(25 downto 0);
    syn_invalidate_word : out  std_logic_vector(26 downto 0);
    clk, reset: in std_logic
    -- 
  );
  end component;
  component accessDcacheRlut_Operator is -- 
   port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    lookup : in  std_logic_vector(0 downto 0);
    update : in  std_logic_vector(0 downto 0);
    clear : in  std_logic_vector(0 downto 0);
    physical_addr_of_line : in  std_logic_vector(29 downto 0);
    virtual_addr_of_line : in  std_logic_vector(25 downto 0);
    syn_invalidate_word : out  std_logic_vector(26 downto 0);
    clk, reset: in std_logic
    -- 
  );
  end component;

  component snoopFilter_Operator is
    port ( -- 
    	sample_req: in boolean;
    	sample_ack: out boolean;
    	update_req: in boolean;
    	update_ack: out boolean;
	rwbar: in std_logic_vector(0 downto 0);
	enable: in std_logic_vector(0 downto 0);
        pa_of_line:  in std_logic_vector(29 downto 0);
	send_inval: out std_logic_vector(0 downto 0);
        clk, reset: in std_logic);
  end component;
  component snoopFilter_1_Operator is
    port ( -- 
    	sample_req: in boolean;
    	sample_ack: out boolean;
    	update_req: in boolean;
    	update_ack: out boolean;
	rwbar: in std_logic_vector(0 downto 0);
	enable: in std_logic_vector(0 downto 0);
        pa_of_line:  in std_logic_vector(29 downto 0);
	send_inval: out std_logic_vector(0 downto 0);
        clk, reset: in std_logic);
  end component;
  component snoopFilter_2_Operator is
    port ( -- 
    	sample_req: in boolean;
    	sample_ack: out boolean;
    	update_req: in boolean;
    	update_ack: out boolean;
	rwbar: in std_logic_vector(0 downto 0);
	enable: in std_logic_vector(0 downto 0);
        pa_of_line:  in std_logic_vector(29 downto 0);
	send_inval: out std_logic_vector(0 downto 0);
        clk, reset: in std_logic);
  end component;
  component snoopFilter_4_Operator is
    port ( -- 
    	sample_req: in boolean;
    	sample_ack: out boolean;
    	update_req: in boolean;
    	update_ack: out boolean;
	rwbar: in std_logic_vector(0 downto 0);
	enable: in std_logic_vector(0 downto 0);
        pa_of_line:  in std_logic_vector(29 downto 0);
	send_inval: out std_logic_vector(0 downto 0);
        clk, reset: in std_logic);
  end component;

  component accessL2TagMemGeneric is -- 
  generic (
		LOG2_NUMBER_OF_LINES: integer := 12;
		LOG2_ASSOCIATIVITY: integer := 3;
		LOG2_DWORDS_PER_LINE: integer := 3;
		PA_ADDRESS_WIDTH: integer := 36
	  );
  port ( -- 
    start_req: in std_logic;
    start_ack: out std_logic;
    fin_req: in std_logic;
    fin_ack: out std_logic;
    init_flag : in  std_logic_vector(0 downto 0);
    tag_mem_read : in  std_logic_vector(0 downto 0);
    tag_mem_write : in  std_logic_vector(0 downto 0);
    read_set_id : in  std_logic_vector((LOG2_NUMBER_OF_LINES-LOG2_ASSOCIATIVITY)-1 downto 0);
    write_set_id : in  std_logic_vector((LOG2_NUMBER_OF_LINES-LOG2_ASSOCIATIVITY)-1 downto 0);
    tags_have_been_modified : in  std_logic_vector(0 downto 0);
    lwi_has_been_modified : in  std_logic_vector(0 downto 0);
    valids_have_been_modified : in  std_logic_vector(0 downto 0);
    dirty_bits_have_been_modified : in  std_logic_vector(0 downto 0);
    updated_set_tags : in  
	std_logic_vector(((2**LOG2_ASSOCIATIVITY)*(30-(LOG2_NUMBER_OF_LINES-LOG2_ASSOCIATIVITY)))-1 downto 0);
    updated_set_lwi : in  
	std_logic_vector(LOG2_ASSOCIATIVITY-1 downto 0);
    updated_set_valids : in  
	std_logic_vector((2**LOG2_ASSOCIATIVITY)-1 downto 0);
    updated_set_dirty_dword_masks : in  
	std_logic_vector(((2**LOG2_DWORDS_PER_LINE)*(2**LOG2_ASSOCIATIVITY))-1 downto 0);
    tag_mem_response : out  
	std_logic_vector(((2**LOG2_ASSOCIATIVITY)*(30-(LOG2_NUMBER_OF_LINES-LOG2_ASSOCIATIVITY))) +
			LOG2_ASSOCIATIVITY + (2**LOG2_ASSOCIATIVITY) + 
			((2**LOG2_DWORDS_PER_LINE)*(2**LOG2_ASSOCIATIVITY))-1  downto 0);
    clk, reset: in std_logic
  );
  end component accessL2TagMemGeneric;

   component accessL2TagMemX1024X8_Operator is -- 
   port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    init_flag : in  std_logic_vector(0 downto 0);
    tag_mem_read : in  std_logic_vector(0 downto 0);
    tag_mem_write : in  std_logic_vector(0 downto 0);
    read_set_id : in  std_logic_vector(6 downto 0);
    write_set_id : in  std_logic_vector(6 downto 0);
    tags_have_been_modified : in  std_logic_vector(0 downto 0);
    lwi_has_been_modified : in  std_logic_vector(0 downto 0);
    valids_have_been_modified : in  std_logic_vector(0 downto 0);
    dirty_bits_have_been_modified : in  std_logic_vector(0 downto 0);
    updated_set_tags : in  std_logic_vector(183 downto 0);
    updated_set_lwi : in  std_logic_vector(2 downto 0);
    updated_set_valids : in  std_logic_vector(7 downto 0);
    updated_set_dirty_dword_masks : in  std_logic_vector(63 downto 0);
    tag_mem_response : out  std_logic_vector(258 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
  end component accessL2TagMemX1024X8_Operator;

  component accessL2TagMemX2048X8_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    init_flag : in  std_logic_vector(0 downto 0);
    tag_mem_read : in  std_logic_vector(0 downto 0);
    tag_mem_write : in  std_logic_vector(0 downto 0);
    read_set_id : in  std_logic_vector(7 downto 0);
    write_set_id : in  std_logic_vector(7 downto 0);
    tags_have_been_modified : in  std_logic_vector(0 downto 0);
    lwi_has_been_modified : in  std_logic_vector(0 downto 0);
    valids_have_been_modified : in  std_logic_vector(0 downto 0);
    dirty_bits_have_been_modified : in  std_logic_vector(0 downto 0);
    updated_set_tags : in  std_logic_vector(175 downto 0);
    updated_set_lwi : in  std_logic_vector(2 downto 0);
    updated_set_valids : in  std_logic_vector(7 downto 0);
    updated_set_dirty_dword_masks : in  std_logic_vector(63 downto 0);
    tag_mem_response : out  std_logic_vector(250 downto 0);
    clk, reset: in std_logic
  );
  end component accessL2TagMemX2048X8_Operator;
  component accessL2TagMemX4096X8_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    init_flag : in  std_logic_vector(0 downto 0);
    tag_mem_read : in  std_logic_vector(0 downto 0);
    tag_mem_write : in  std_logic_vector(0 downto 0);
    read_set_id : in  std_logic_vector(8 downto 0);
    write_set_id : in  std_logic_vector(8 downto 0);
    tags_have_been_modified : in  std_logic_vector(0 downto 0);
    lwi_has_been_modified : in  std_logic_vector(0 downto 0);
    valids_have_been_modified : in  std_logic_vector(0 downto 0);
    dirty_bits_have_been_modified : in  std_logic_vector(0 downto 0);
    updated_set_tags : in  std_logic_vector(167 downto 0);
    updated_set_lwi : in  std_logic_vector(2 downto 0);
    updated_set_valids : in  std_logic_vector(7 downto 0);
    updated_set_dirty_dword_masks : in  std_logic_vector(63 downto 0);
    tag_mem_response : out  std_logic_vector(242 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
  end component accessL2TagMemX4096X8_Operator;

  component accessL2DataMemGeneric is -- 
    generic (LOG2_NUMBER_OF_LINES : integer := 11; 
		LINE_WIDTH_IN_BYTES: integer := 64);
  port ( -- 
    start_req: in std_logic;
    start_ack: out std_logic;
    fin_req: in std_logic;
    fin_ack: out std_logic;
    -- if true, read data line..
    read_data_line : in  std_logic_vector(0 downto 0);
    -- if true, write data word...
    data_write_dword : in  std_logic_vector(0 downto 0);
    -- if true, read data word (note: read_data_line will also be true in this case)
    data_read_dword : in  std_logic_vector(0 downto 0);
    -- write new line into data mem, (note: insert write dword if data_write_dword is true).
    data_write_new_line : in  std_logic_vector(0 downto 0);
    -- this is now redundant..  write_new_line is always the replaced line.
    do_write_replaced_line_to_mem : in  std_logic_vector(0 downto 0);
    -- byte mask for dword write.
    byte_mask : in  std_logic_vector(7 downto 0);
    -- address of line.
    line_id : in  std_logic_vector(LOG2_NUMBER_OF_LINES-1 downto 0);
    -- offset in line for write dword.
    pa_dword_id : in  std_logic_vector(2 downto 0);
    -- write dword.
    w_dword : in  std_logic_vector(63 downto 0);
    -- line to be written into memory..
    line_to_be_inserted : in  std_logic_vector((8*LINE_WIDTH_IN_BYTES)-1 downto 0);
    -- read data
    read_dword_from_data : out  std_logic_vector(63 downto 0);
    -- line that was read out of memory.. this line will be written eventually to main memory.
    writeback_line_from_data : out  std_logic_vector((8*LINE_WIDTH_IN_BYTES)-1 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
  end component accessL2DataMemGeneric;

  component accessL2DataMemGeneric_Operator is -- 
    generic (
		name: string;
		LOG2_NUMBER_OF_LINES: integer := 10;
		LINE_WIDTH_IN_BYTES: integer := 64
	);
    port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    -- if true, read data line..
    read_data_line : in  std_logic_vector(0 downto 0);
    -- if true, write data word...
    data_write_dword : in  std_logic_vector(0 downto 0);
    -- if true, read data word (note: read_data_line will also be true in this case)
    data_read_dword : in  std_logic_vector(0 downto 0);
    -- write new line into data mem, (note: insert write dword if data_write_dword is true).
    data_write_new_line : in  std_logic_vector(0 downto 0);
    -- this is now redundant..  write_new_line is always the replaced line.
    do_write_replaced_line_to_mem : in  std_logic_vector(0 downto 0);
    -- byte mask for dword write.
    byte_mask : in  std_logic_vector(7 downto 0);
    -- address of line.
    line_id : in  std_logic_vector(LOG2_NUMBER_OF_LINES-1 downto 0);
    -- offset in line for write dword.
    pa_dword_id : in  std_logic_vector(2 downto 0);
    -- write dword.
    w_dword : in  std_logic_vector(63 downto 0);
    -- line to be written into memory..
    line_to_be_inserted : in  std_logic_vector((8*LINE_WIDTH_IN_BYTES)-1 downto 0);
    -- read data
    read_dword_from_data : out  std_logic_vector(63 downto 0);
    -- line that was read out of memory.. this line will be written eventually to main memory.
    writeback_line_from_data : out  std_logic_vector((8*LINE_WIDTH_IN_BYTES)-1 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
  end component accessL2DataMemGeneric_Operator;

  component accessL2DataMemX1024X512_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    -- if true, read data line..
    read_data_line : in  std_logic_vector(0 downto 0);
    -- if true, write data word...
    data_write_dword : in  std_logic_vector(0 downto 0);
    -- if true, read data word (note: read_data_line will also be true in this case)
    data_read_dword : in  std_logic_vector(0 downto 0);
    -- write new line into data mem, (note: insert write dword if data_write_dword is true).
    data_write_new_line : in  std_logic_vector(0 downto 0);
    -- this is now redundant..  write_new_line is always the replaced line.
    do_write_replaced_line_to_mem : in  std_logic_vector(0 downto 0);
    -- byte mask for dword write.
    byte_mask : in  std_logic_vector(7 downto 0);
    -- address of line.
    line_id : in  std_logic_vector(9 downto 0);
    -- offset in line for write dword.
    pa_dword_id : in  std_logic_vector(2 downto 0);
    -- write dword.
    w_dword : in  std_logic_vector(63 downto 0);
    -- line to be written into memory..
    line_to_be_inserted : in  std_logic_vector((8*64)-1 downto 0);
    -- read data
    read_dword_from_data : out  std_logic_vector(63 downto 0);
    -- line that was read out of memory.. this line will be written eventually to main memory.
    writeback_line_from_data : out  std_logic_vector((8*64)-1 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
  end component accessL2DataMemX1024X512_Operator;

  component accessL2DataMemX2048X512_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    -- if true, read data line..
    read_data_line : in  std_logic_vector(0 downto 0);
    -- if true, write data word...
    data_write_dword : in  std_logic_vector(0 downto 0);
    -- if true, read data word (note: read_data_line will also be true in this case)
    data_read_dword : in  std_logic_vector(0 downto 0);
    -- write new line into data mem, (note: insert write dword if data_write_dword is true).
    data_write_new_line : in  std_logic_vector(0 downto 0);
    -- this is now redundant..  write_new_line is always the replaced line.
    do_write_replaced_line_to_mem : in  std_logic_vector(0 downto 0);
    -- byte mask for dword write.
    byte_mask : in  std_logic_vector(7 downto 0);
    -- address of line.
    line_id : in  std_logic_vector(10 downto 0);
    -- offset in line for write dword.
    pa_dword_id : in  std_logic_vector(2 downto 0);
    -- write dword.
    w_dword : in  std_logic_vector(63 downto 0);
    -- line to be written into memory..
    line_to_be_inserted : in  std_logic_vector((8*64)-1 downto 0);
    -- read data
    read_dword_from_data : out  std_logic_vector(63 downto 0);
    -- line that was read out of memory.. this line will be written eventually to main memory.
    writeback_line_from_data : out  std_logic_vector((8*64)-1 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
  end component accessL2DataMemX2048X512_Operator;

  component accessL2DataMemX4096X512_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    -- if true, read data line..
    read_data_line : in  std_logic_vector(0 downto 0);
    -- if true, write data word...
    data_write_dword : in  std_logic_vector(0 downto 0);
    -- if true, read data word (note: read_data_line will also be true in this case)
    data_read_dword : in  std_logic_vector(0 downto 0);
    -- write new line into data mem, (note: insert write dword if data_write_dword is true).
    data_write_new_line : in  std_logic_vector(0 downto 0);
    -- this is now redundant..  write_new_line is always the replaced line.
    do_write_replaced_line_to_mem : in  std_logic_vector(0 downto 0);
    -- byte mask for dword write.
    byte_mask : in  std_logic_vector(7 downto 0);
    -- address of line.
    line_id : in  std_logic_vector(11 downto 0);
    -- offset in line for write dword.
    pa_dword_id : in  std_logic_vector(2 downto 0);
    -- write dword.
    w_dword : in  std_logic_vector(63 downto 0);
    -- line to be written into memory..
    line_to_be_inserted : in  std_logic_vector((8*64)-1 downto 0);
    -- read data
    read_dword_from_data : out  std_logic_vector(63 downto 0);
    -- line that was read out of memory.. this line will be written eventually to main memory.
    writeback_line_from_data : out  std_logic_vector((8*64)-1 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
  end component accessL2DataMemX4096X512_Operator;

  component ajit_64kB_rom is
	    port (clk  : in std_logic;
	              en   : in std_logic;
	              addr : in std_logic_vector(15 downto 0);
	              data : out std_logic_vector(7 downto 0));
  end component ajit_64kB_rom;


  component rt_clock_counter is
	port (
			clk, reset: in std_logic;
			one_hz_rt_clock: in std_logic_vector(0 downto 0);
			count_value : out std_logic_vector(31 downto 0)
		);
  end component rt_clock_counter;

  component baud_control_calculator is  -- system 
   port (-- 
     clk : in std_logic;
     reset : in std_logic;
     BAUD_CONTROL_WORD_SIG: out std_logic_vector(31 downto 0);
     BAUD_CONTROL_WORD_VALID: out std_logic_vector(0 downto 0);
     BAUD_RATE_SIG: in std_logic_vector(31 downto 0);
     CLOCK_FREQUENCY_VALID: in std_logic_vector(0 downto 0); -- 
     CLK_FREQUENCY_SIG: in std_logic_vector(31 downto 0));  
  end component; 

  
  component uart_synchronizer is
		generic (baud_rate: integer := 115200);
		port (
				clk, reset: in std_logic;
				Rx_in: in std_logic;
				rt_clock : out std_logic
	     	);
  end component uart_synchronizer;

  component configurable_self_tuning_uart is
	port (clk, reset: in std_logic; 
		rt_1Hz: in std_logic_vector(0 downto 0); 

		BAUD_RATE: in std_logic_vector(31 downto 0);
		UART_RX: in std_logic_vector(0 downto 0); 
		UART_TX: out std_logic_vector(0 downto 0);

		TX_to_CONSOLE_pipe_write_data: in std_logic_vector(7 downto 0);
		TX_to_CONSOLE_pipe_write_req:  in std_logic_vector(0 downto 0);
		TX_to_CONSOLE_pipe_write_ack:  out std_logic_vector(0 downto 0);

		CONSOLE_to_RX_pipe_read_data : out std_logic_vector(7 downto 0);
		CONSOLE_to_RX_pipe_read_req :  in std_logic_vector(0 downto 0);
		CONSOLE_to_RX_pipe_read_ack :  out std_logic_vector(0 downto 0));
   end component configurable_self_tuning_uart;

   component configurable_self_tuning_uart_without_rt_clock is
	generic (BAUD_RATE: integer := 115200);
	port (clk, reset: in std_logic; 

		UART_RX: in std_logic_vector(0 downto 0); 
		UART_TX: out std_logic_vector(0 downto 0);

		TX_to_CONSOLE_pipe_write_data: in std_logic_vector(7 downto 0);
		TX_to_CONSOLE_pipe_write_req:  in std_logic_vector(0 downto 0);
		TX_to_CONSOLE_pipe_write_ack:  out std_logic_vector(0 downto 0);

		CONSOLE_to_RX_pipe_read_data : out std_logic_vector(7 downto 0);
		CONSOLE_to_RX_pipe_read_req :  in std_logic_vector(0 downto 0);
		CONSOLE_to_RX_pipe_read_ack :  out std_logic_vector(0 downto 0));
   end component configurable_self_tuning_uart_without_rt_clock;


  component afb_ahb_lite_master is -- 
  port( -- 
    AFB_BUS_REQUEST_pipe_write_data : in std_logic_vector(73 downto 0);
    AFB_BUS_REQUEST_pipe_write_req  : in std_logic_vector(0  downto 0);
    AFB_BUS_REQUEST_pipe_write_ack  : out std_logic_vector(0  downto 0);
    HRDATA : in std_logic_vector(31 downto 0);
    HREADY : in std_logic_vector(0 downto 0);
    HRESP : in std_logic_vector(1 downto 0);
    AFB_BUS_RESPONSE_pipe_read_data : out std_logic_vector(32 downto 0);
    AFB_BUS_RESPONSE_pipe_read_req  : in std_logic_vector(0  downto 0);
    AFB_BUS_RESPONSE_pipe_read_ack  : out std_logic_vector(0  downto 0);
    HADDR : out std_logic_vector(35 downto 0);
    HBURST : out std_logic_vector(2 downto 0);
    HMASTLOCK : out std_logic_vector(0 downto 0);
    HPROT : out std_logic_vector(3 downto 0);
    HSIZE : out std_logic_vector(2 downto 0);
    HTRANS : out std_logic_vector(1 downto 0);
    HWDATA : out std_logic_vector(31 downto 0);
    HWRITE : out std_logic_vector(0 downto 0);
    SYS_CLK : out std_logic_vector(0 downto 0);
    clk, reset: in std_logic 
    -- 
  );
  --
  end component afb_ahb_lite_master;
  component ahblite_controller is
	port (
		-- connections to AFB-AHB bridge
		AFB_TO_AHB_COMMAND_pipe_write_req: in  std_logic_vector(0 downto 0);
		AFB_TO_AHB_COMMAND_pipe_write_ack: out std_logic_vector(0 downto 0);
		AFB_TO_AHB_COMMAND_pipe_write_data: in std_logic_vector(72 downto 0);
		-- 
		AHB_TO_AFB_RESPONSE_pipe_read_req: in  std_logic_vector(0 downto 0);
		AHB_TO_AFB_RESPONSE_pipe_read_ack: out std_logic_vector(0 downto 0);
		AHB_TO_AFB_RESPONSE_pipe_read_data: out std_logic_vector(32 downto 0);
		-- AHB bus signals
		HADDR: out std_logic_vector(35 downto 0);
		HTRANS: out std_logic_vector(1 downto 0); -- non-sequential, sequential, idle, busy
		HWRITE: out std_logic_vector(0 downto 0); -- when '1' its a write.
		HSIZE: out std_logic_vector(2 downto 0); -- transfer size in bytes.
		HBURST: out std_logic_vector(2 downto 0); -- burst size.
		HMASTLOCK: out std_logic_vector(0 downto 0); -- locked transaction.. for swap etc.
		HPROT: out std_logic_vector(3 downto 0); -- protection bits..
		HWDATA: out std_logic_vector(31 downto 0); -- write data.
		HRDATA: in std_logic_vector(31 downto 0); -- read data.
		HREADY: in std_logic_vector(0 downto 0); -- slave ready.
		HRESP: in std_logic_vector(1 downto 0); -- okay, error, retry, split (slave responses).
		SYS_CLK: out std_logic_vector(0 downto 0);
		-- clock, reset.
		clk: in std_logic;
		reset: in std_logic 
	     );
   end component ahblite_controller;
   component afb_ahb_bridge is -- 
    port (-- 
      clk : in std_logic;
      reset : in std_logic;
      AFB_BUS_REQUEST_pipe_write_data: in std_logic_vector(73 downto 0);
      AFB_BUS_REQUEST_pipe_write_req : in std_logic_vector(0 downto 0);
      AFB_BUS_REQUEST_pipe_write_ack : out std_logic_vector(0 downto 0);
      AFB_BUS_RESPONSE_pipe_read_data: out std_logic_vector(32 downto 0);
      AFB_BUS_RESPONSE_pipe_read_req : in std_logic_vector(0 downto 0);
      AFB_BUS_RESPONSE_pipe_read_ack : out std_logic_vector(0 downto 0);
      AFB_TO_AHB_COMMAND_pipe_read_data: out std_logic_vector(72 downto 0);
      AFB_TO_AHB_COMMAND_pipe_read_req : in std_logic_vector(0 downto 0);
      AFB_TO_AHB_COMMAND_pipe_read_ack : out std_logic_vector(0 downto 0);
      AHB_TO_AFB_RESPONSE_pipe_write_data: in std_logic_vector(32 downto 0);
      AHB_TO_AFB_RESPONSE_pipe_write_req : in std_logic_vector(0 downto 0);
      AHB_TO_AFB_RESPONSE_pipe_write_ack : out std_logic_vector(0 downto 0)); -- 
    -- 
   end component;

   -- instruction buffer...
   component access_instruction_buffer_Operator is -- 
   port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    clear_flag : in  std_logic_vector(0 downto 0);
    insert_flag : in  std_logic_vector(0 downto 0);
    insert_addr : in  std_logic_vector(28 downto 0);
    insert_acc  : in  std_logic_vector(2 downto 0);
    insert_ipair : in  std_logic_vector(63 downto 0);
    lookup_flag : in  std_logic_vector(0 downto 0);
    lookup_addr : in  std_logic_vector(28 downto 0);
    lookup_match : out  std_logic_vector(0 downto 0);
    lookup_acc  : out  std_logic_vector(2 downto 0);
    lookup_ipair : out  std_logic_vector(63 downto 0);
    clk, reset: in std_logic
    -- 
   );
   -- 
  end component access_instruction_buffer_Operator;


  component instruction_buffer is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    icache_to_instruction_buffer_response_pipe_write_data: in std_logic_vector(89 downto 0);
    icache_to_instruction_buffer_response_pipe_write_req : in std_logic_vector(0 downto 0);
    icache_to_instruction_buffer_response_pipe_write_ack : out std_logic_vector(0 downto 0);
    instruction_buffer_to_cpu_response_pipe_read_data: out std_logic_vector(89 downto 0);
    instruction_buffer_to_cpu_response_pipe_read_req : in std_logic_vector(0 downto 0);
    instruction_buffer_to_cpu_response_pipe_read_ack : out std_logic_vector(0 downto 0);
    noblock_cpu_to_instruction_buffer_request_pipe_write_data: in std_logic_vector(40 downto 0);
    noblock_cpu_to_instruction_buffer_request_pipe_write_req : in std_logic_vector(0 downto 0);
    noblock_cpu_to_instruction_buffer_request_pipe_write_ack : out std_logic_vector(0 downto 0);
    noblock_instruction_buffer_to_icache_request_pipe_read_data: out std_logic_vector(40 downto 0);
    noblock_instruction_buffer_to_icache_request_pipe_read_req : in std_logic_vector(0 downto 0);
    noblock_instruction_buffer_to_icache_request_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
  end component; 

  component instruction_buffer_optimized is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    icache_to_instruction_buffer_response_pipe_write_data: in std_logic_vector(89 downto 0);
    icache_to_instruction_buffer_response_pipe_write_req : in std_logic_vector(0 downto 0);
    icache_to_instruction_buffer_response_pipe_write_ack : out std_logic_vector(0 downto 0);
    instruction_buffer_to_cpu_response_pipe_read_data: out std_logic_vector(89 downto 0);
    instruction_buffer_to_cpu_response_pipe_read_req : in std_logic_vector(0 downto 0);
    instruction_buffer_to_cpu_response_pipe_read_ack : out std_logic_vector(0 downto 0);
    noblock_cpu_to_instruction_buffer_request_pipe_write_data: in std_logic_vector(40 downto 0);
    noblock_cpu_to_instruction_buffer_request_pipe_write_req : in std_logic_vector(0 downto 0);
    noblock_cpu_to_instruction_buffer_request_pipe_write_ack : out std_logic_vector(0 downto 0);
    noblock_instruction_buffer_to_icache_request_pipe_read_data: out std_logic_vector(40 downto 0);
    noblock_instruction_buffer_to_icache_request_pipe_read_req : in std_logic_vector(0 downto 0);
    noblock_instruction_buffer_to_icache_request_pipe_read_ack : out std_logic_vector(0 downto 0);
    core_id: in std_logic_vector(3 downto 0);
    cpu_id: in std_logic_vector(3 downto 0)); -- 
  -- 
  end component; 
end package;
library ieee;
use ieee.std_logic_1164.all;

package RomPackage is
	type AJIT_ROM_TYPE is array (0 to 65535) of std_logic_vector(7 downto 0); -- 64kB
	-- for test purposes only..  Need to define based on rom contents.
	constant ROM_INITIAL_VALUE: AJIT_ROM_TYPE := (0 => X"00", 1 => X"01", 2 => X"02",
							3 => X"03", 4 => X"04", 5 => X"05",
							6 => X"06", 7 => X"07", 8 => X"08",
							9 => X"09", 10 => X"0A", 11 => X"0B",
							12 => X"0C", 13 => X"0D", 14 => X"0E",
							15 => X"0F", others => X"FF");
end package RomPackage;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

package UsefulFunctions is
	function accessPermissionsOk(S,ifetch,is_read: std_logic; 
					acc: std_logic_vector(2 downto 0))
		return std_logic;

	function InsertRdVal(offset: integer; save, restore : std_logic;
						rd: std_logic_vector(4 downto 0);
						rd_val: std_logic_vector(31 downto 0);
						reg_256: std_logic_vector(255 downto 0))
		return std_logic_vector;

end package UsefulFunctions;


package body UsefulFunctions is
	function accessPermissionsOk(S,ifetch,is_read: std_logic; 
					acc: std_logic_vector(2 downto 0))
		return std_logic is
		variable ret_val : std_logic;
	begin
		ret_val := '1';
		case acc is 
			when "000" => -- read:read
				ret_val := (not ifetch) and is_read;
			when "001" => -- read/write : read/write
				ret_val := not ifetch;
			when "010" => -- read/exec : read/exec
				ret_val := is_read;
			when "011" => -- read/write/exec : read/write/exec
				ret_val := '1';
			when "100" => -- exec: exec
				ret_val := ifetch;
			when "101" => -- read : read/write
				ret_val := (not ifetch) and ((not S) or is_read);
			when "110" => -- no-acc  : read/exec
				ret_val := S and is_read;
			when "111" => -- no-acc : read/write/exec
				ret_val := S;
			when others =>
				ret_val := '0';
		end case;		
		return (ret_val);
	end accessPermissionsOk;

	function InsertRdVal(offset: integer; save, restore : std_logic;
						rd: std_logic_vector(4 downto 0);
						rd_val: std_logic_vector(31 downto 0);
						reg_256: std_logic_vector(255 downto 0))
		return std_logic_vector is
		variable ret_val : std_logic_vector(255 downto 0);
		variable wr_val : std_logic_vector(31 downto 0);
		variable w0,w1,w2,w3,w4,w5,w6,w7: std_logic_vector(31 downto 0);

		variable reg_index : integer range 0 to 31;
	begin
		w7 := reg_256 (31 downto 0);
		w6 := reg_256 (63 downto 32);
		w5 := reg_256 (95 downto 64);
		w4 := reg_256 (127 downto 96);
		w3 := reg_256 (159 downto 128);
		w2 := reg_256 (191 downto 160);
		w1 := reg_256 (223 downto 192);
		w0 := reg_256 (255 downto 224);

		reg_index := to_integer(unsigned(rd));

		-- register 0 always contains 0.
		if(reg_index = 0) then
			wr_val := (others => '0');
		else
			wr_val := rd_val;
		end if;

		if(((save = '1')  or (restore = '1')) and (reg_index >= offset)) then
			
			reg_index := reg_index - offset;

			if(reg_index < 8) then

				
				if (reg_index = 0) then
					w0 := wr_val;
				elsif reg_index = 1 then
					w1 := wr_val;
				elsif reg_index = 2 then
					w2 := wr_val;
				elsif reg_index = 3 then
					w3 := wr_val;
				elsif reg_index = 4 then
					w4 := wr_val;
				elsif reg_index = 5 then
					w5 := wr_val;
				elsif reg_index = 6 then
					w6 := wr_val;
				elsif reg_index = 7 then
					w7 := wr_val;
				end if;
			end if;
		end if;

		ret_val := w0 & w1 & w2 & w3 & w4 & w5 & w6 & w7;
		return(ret_val);
	end function InsertRdVal;

end package body UsefulFunctions;
library ieee;
use ieee.std_logic_1164.all;

package CachePackage is

	constant CACHE_ARRAY_READ_DWORD  	: std_logic_vector(2 downto 0) := "001";
	constant CACHE_ARRAY_WRITE_DWORD  	: std_logic_vector(2 downto 0) := "010";
	constant CACHE_ARRAY_NOP	     	: std_logic_vector(2 downto 0) := "011";
	constant CACHE_ARRAY_PASS_THROUGH     	: std_logic_vector(2 downto 0) := "100";

	constant CACHE_TAG_LOOKUP	       : std_logic_vector(2 downto 0) := "001";
	constant CACHE_TAG_INSERT	       : std_logic_vector(2 downto 0) := "010";
	constant CACHE_TAG_CLEAR_LINE	       : std_logic_vector(2 downto 0) := "011";
	constant CACHE_TAG_CLEAR_ALL	       : std_logic_vector(2 downto 0) := "100";
	constant CACHE_TAG_NOP	       	       : std_logic_vector(2 downto 0) := "101";

	constant VA_INDEX_TLB_SIZE 		: integer := 2;

end package CachePackage;
library ieee;
use ieee.std_logic_1164.all;

-- Simple synchronizer... with 4-stage delay to simplify 
-- routing across the chip.
entity Simple4StageSynchronizer is
    port (clk, reset_asynch: in std_logic; reset_synch: out std_logic);
end entity Simple4StageSynchronizer;

architecture Obvious of Simple4StageSynchronizer is
   signal reset_synch_0, reset_synch_1, reset_synch_2: std_logic;
begin
  
 process(clk)
 begin
   if (clk'event and clk = '1') then
     reset_synch_0 <= reset_asynch;
     reset_synch_1 <= reset_synch_0;
     reset_synch_2 <= reset_synch_1;
     reset_synch   <= reset_synch_2;
   end if;
 end process;

end Obvious;

--
-- Written by Madhav Desai
--
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.BaseComponents.all;
use ahir.mem_component_pack.all;
use ahir.Types.all;
use ahir.Utilities.all;

entity GenericCacheArray is -- 
  generic (name: string := "anon";
		log2_number_of_blocks: integer := 9; 
		log2_block_size_in_bytes: integer := 6; 
		address_width: integer := 32;
		log2_data_width_in_bytes: integer := 3);
  port ( -- 
    trigger: in std_logic;
    done: out std_logic;
    access_mae : in  std_logic;
    access_array_command : in  std_logic_vector(2 downto 0);
    access_byte_mask : in  std_logic_vector((2**log2_data_width_in_bytes)-1 downto 0);
    access_array_addr : in  std_logic_vector(address_width-1 downto 0);
    access_dword : in  std_logic_vector((8*(2**log2_data_width_in_bytes))-1 downto 0);
    dword_out : out  std_logic_vector((8*(2**log2_data_width_in_bytes))-1 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity GenericCacheArray;
architecture Behave of GenericCacheArray is -- 

	-- dcache-array management commands
	constant CACHE_ARRAY_READ_DWORD  	: std_logic_vector(2 downto 0) := "001";
	constant CACHE_ARRAY_WRITE_DWORD  	: std_logic_vector(2 downto 0) := "010";
	constant CACHE_ARRAY_NOP	     	: std_logic_vector(2 downto 0) := "011";
	constant CACHE_ARRAY_PASS_THROUGH     	: std_logic_vector(2 downto 0) := "100";

	constant number_of_blocks : integer := (2**log2_number_of_blocks);
	constant bytes_per_block : integer := (2**log2_block_size_in_bytes);
	constant data_width_in_bytes : integer := (2**log2_data_width_in_bytes);
	constant dwords_per_block : integer := (2**(log2_block_size_in_bytes - log2_data_width_in_bytes));
	constant log2_dwords_per_block: integer := (log2_block_size_in_bytes - log2_data_width_in_bytes);

	--
	--  memory access signals.
	-- 
	signal  array_mem_address : std_logic_vector((log2_number_of_blocks + log2_dwords_per_block)-1 downto 0);
	signal  array_mem_write_data: std_logic_vector((8*data_width_in_bytes)-1 downto 0);
	signal  array_mem_read_data: std_logic_vector((8*data_width_in_bytes)-1 downto 0);
	signal  array_mem_byte_enable: std_logic_vector(data_width_in_bytes-1 downto 0);
	signal  array_mem_enable: std_logic;
	signal  array_mem_write_bar: std_logic;

	signal enable_sig: std_logic;
	signal dword_out_sig, access_dword_registered : std_logic_vector((8*(2**log2_data_width_in_bytes))-1 downto 0);

	signal  access_array_command_registered : std_logic_vector(2 downto 0);
	signal  access_mae_registered: std_logic;
	
begin --  

	----------------------------------------------------------------------------------
	-- state machine! Assuming that the memory is one-cycle.
	----------------------------------------------------------------------------------
	process(clk, reset, trigger)
	begin 
		if(clk'event and (clk = '1')) then
			if(reset = '1') then
				done <= '0';
			else
				done <= trigger;
			end if;
		end if;
	end process;
	enable_sig <= trigger;

	----------------------------------------------------------------------------------
	-- prepare inputs to memory.
	----------------------------------------------------------------------------------
	array_mem_address <= access_array_addr ((log2_number_of_blocks + log2_dwords_per_block + log2_data_width_in_bytes)-1
									downto log2_data_width_in_bytes);
	array_mem_enable <= (enable_sig and (not access_mae));
	array_mem_write_bar <= '0' when (access_array_command =  CACHE_ARRAY_WRITE_DWORD) else '1';

	-- enable bytes
	process(access_byte_mask, array_mem_enable)
	begin
		for B in data_width_in_bytes-1 downto 0 loop
			array_mem_byte_enable(B) <= array_mem_enable and access_byte_mask(B);
		end loop;
	end process;	
	array_mem_write_data <= access_dword;

	------------------------------------------------------------------------------------------------
	--  mux, register and forward to output stage
	------------------------------------------------------------------------------------------------
	process(clk, reset, access_dword, access_array_command, access_mae)
	begin
		if clk'event and clk = '1' then
			if(reset ='1')  then
				access_array_command_registered <= (others => '0');
				access_mae_registered <= '0';
			elsif	 (enable_sig = '1') then
				access_array_command_registered <= access_array_command;
				access_mae_registered <= access_mae;
				access_dword_registered <= access_dword;
			end if;
		end if;
	end process;
	------------------------------------------------------------------------------------------------
	------------------------------------------------------------------------------------------------
	-- line banks
	lineBankGen: for B in data_width_in_bytes-1 downto 0 generate
		lineBank: base_bank
				generic map (name => "linBank" & Convert_To_String(B),
						g_addr_width => log2_number_of_blocks + log2_dwords_per_block,
						g_data_width => 8)
				port map (
						datain => array_mem_write_data((8*(B+1))-1 downto 8*B),
						dataout => array_mem_read_data((8*(B+1))-1 downto 8*B),
						addrin => array_mem_address, 
						enable => array_mem_byte_enable(B),
						writebar => array_mem_write_bar,
						clk => clk, reset => reset);	
	end generate lineBankGen;
		
	------------------------------------------------------------------------------------------------
	--  output logic
	------------------------------------------------------------------------------------------------
	-- output
	dword_out <= (others => '0') when access_mae_registered = '1' 
			else array_mem_read_data when (access_array_command_registered = CACHE_ARRAY_READ_DWORD)
				else  access_dword_registered;
end Behave;
--
-- Written by Madhav Desai
--
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library AjitCustom;
use AjitCustom.UsefulFunctions.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

library ahir;
use ahir.BaseComponents.all;
use ahir.mem_component_pack.all;
use ahir.Types.all;
use ahir.Utilities.all;

entity GenericCacheTags is -- 
  generic (name: string := "anon";
		log2_number_of_blocks: integer := 9; 
		log2_block_size_in_bytes: integer := 6; 
		address_width: integer := 32;
		tag_length: integer := 1;
		log2_data_width_in_bytes: integer := 3);
  port ( -- 
    start_req: in std_logic;
    start_ack: out std_logic;
    fin_req: in std_logic;
    fin_ack: out std_logic;
    init_flag : in  std_logic;
    access_mae : in  std_logic;
    access_S : in  std_logic;
    access_is_read: in std_logic;
    access_is_ifetch: in std_logic;
    access_acc: in std_logic_vector(2 downto 0);
    access_tag_command : in  std_logic_vector(2 downto 0);
    access_tag_addr : in  std_logic_vector(address_width-1 downto 0);
    is_hit : out  std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0);
    permissions_ok : out  std_logic_vector(0 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity GenericCacheTags;
architecture Behave of GenericCacheTags is -- 

	-- dcache-tag management commands
	constant CACHE_TAG_LOOKUP	       : std_logic_vector(2 downto 0) := "001";
	constant CACHE_TAG_INSERT	       : std_logic_vector(2 downto 0) := "010";
	constant CACHE_TAG_CLEAR_LINE	       : std_logic_vector(2 downto 0) := "011";
	constant CACHE_TAG_CLEAR_ALL	       : std_logic_vector(2 downto 0) := "100";
	constant CACHE_TAG_NOP	       	       : std_logic_vector(2 downto 0) := "101";

	constant number_of_blocks : integer := (2**log2_number_of_blocks);
	constant bytes_per_block : integer := (2**log2_block_size_in_bytes);
	constant data_width_in_bytes : integer := (2**log2_data_width_in_bytes);
	constant dwords_per_block : integer := (2**(log2_block_size_in_bytes - log2_data_width_in_bytes));
	constant log2_dwords_per_block: integer := (log2_block_size_in_bytes - log2_data_width_in_bytes);


	--  tag width 
	constant tag_width : integer :=  address_width - (log2_number_of_blocks + log2_block_size_in_bytes);
	
	--
	--  memory access signals.
	-- 
	signal  tag_mem_address : std_logic_vector(log2_number_of_blocks-1 downto 0);
	signal  tag_mem_write_data: std_logic_vector(tag_width+2 downto 0);
	signal  tag_mem_read_data: std_logic_vector(tag_width+2 downto 0);
	signal  tag_mem_enable: std_logic;
	signal  tag_mem_write_bar: std_logic;
	
	--
	-- valid bits.. 
	-- 
	signal valid_bits: std_logic_vector (number_of_blocks-1 downto 0);
	
      	

	Type FsmState is (Idle, WaitForReceiveBuffer);
	signal fsm_state: FsmState;
	
	signal valid_bit_registered : std_logic;
	signal latch_request_info: Boolean;

	signal invalidate_missed_cache_line : Boolean;
	signal invalidate_missed_cache_line_block_id : integer range 0 to number_of_blocks-1;


	function blockId (x: std_logic_vector(address_width-1 downto 0)) 
		return integer is
		variable ret_var : integer range 0 to number_of_blocks -1;
		variable block_id_var : std_logic_vector(log2_number_of_blocks-1 downto 0);
	begin
		block_id_var := x ((log2_number_of_blocks + log2_block_size_in_bytes)-1 
							downto log2_block_size_in_bytes);
		ret_var := to_integer(unsigned(block_id_var));
		return(ret_var);

	end blockId;


	-- access-completed-registered.. indicates that
	-- an action has just completed.
	signal access_active, access_completed: Boolean;

	signal is_hit_sig : std_logic;
	signal permissions_ok_sig : std_logic;

	signal  tag_block_id : std_logic_vector(log2_number_of_blocks-1 downto 0);
	signal  tag_block_id_int : integer range 0 to number_of_blocks-1;
	signal  tag_addr_tag, tag_addr_tag_registered : std_logic_vector(tag_width-1 downto 0);

	signal rx_buf_read_req, rx_buf_read_ack: std_ulogic;

	-- for output stage.
    	signal access_tag_command_registered : std_logic_vector(2 downto 0);
    	signal access_S_registered : std_logic;
	signal access_mae_registered : std_logic;
	signal access_is_ifetch_registered : std_logic;
	signal access_is_read_registered : std_logic;
	signal fin_ack_sig, enable_sig: std_logic;
      
-- see comment above..
--##decl_synopsys_sync_set_reset##

begin --  

	----------------------------------------------------------------------------------
	-- state machine! Assuming that the memory is one-cycle.
	----------------------------------------------------------------------------------
	process(clk, reset, fin_req, start_req, fin_ack_sig, tag_in, enable_sig)
		variable next_fin_ack_sig: std_logic;
	begin 
		next_fin_ack_sig :=
			((not fin_ack_sig) and start_req)
				or
			(fin_ack_sig and (not fin_req))
				or
			(fin_ack_sig and fin_req and start_req);

		enable_sig <= 
			((not fin_ack_sig) and start_req) 
				or
			(fin_ack_sig and fin_req and start_req);

		if(clk'event and (clk = '1')) then
			if(reset = '1') then
				fin_ack_sig <= '0';
				tag_out <= (others => '0');
			else
				if (enable_sig = '1') then
					tag_out <= tag_in;
				end if;

				fin_ack_sig <= next_fin_ack_sig;
			end if;

		end if;
	end process;

	fin_ack <= fin_ack_sig;
	start_ack <= enable_sig;

	----------------------------------------------------------------------------------
	-- valid bit manipulation
	----------------------------------------------------------------------------------
	process(clk, access_tag_command, enable_sig, access_mae, tag_block_id_int, valid_bits, init_flag)
		variable next_valid_bits: std_logic_vector (number_of_blocks-1 downto 0);
		variable next_valid_bit_registered: std_logic;
		variable inserted_valid_bit: std_logic;
	begin
		next_valid_bits := valid_bits;
		inserted_valid_bit := valid_bits(tag_block_id_int);
		next_valid_bit_registered := '0';

		if(access_tag_command = CACHE_TAG_INSERT) then
			inserted_valid_bit := '1';
		elsif (access_tag_command = CACHE_TAG_CLEAR_LINE) then
			inserted_valid_bit := '0';
		end if; 

		if (access_tag_command = CACHE_TAG_CLEAR_LINE) or (access_tag_command = CACHE_TAG_INSERT) then
			next_valid_bits(tag_block_id_int) := inserted_valid_bit;
		elsif (access_tag_command = CACHE_TAG_CLEAR_ALL) then
			next_valid_bits := (others => '0');
		elsif (access_tag_command = CACHE_TAG_LOOKUP) then
			next_valid_bit_registered := inserted_valid_bit;
		end if;

		if(clk'event and clk = '1') then
			--
			-- note that init-flag is asynchronous and can appear at
			-- any time.
			--
			if ((init_flag = '1') or (reset = '1')) then
				valid_bits <= (others => '0');
				valid_bit_registered <= '0';
			elsif  (enable_sig = '1') then
				valid_bits <= next_valid_bits;
				valid_bit_registered <= next_valid_bit_registered;
			end if;	
		end if;
	end process;	
	
	tag_block_id_int <=  blockId(access_tag_addr);
	tag_addr_tag <= access_tag_addr(address_width-1 downto (address_width - tag_width));
	tag_mem_address   <=  access_tag_addr((log2_number_of_blocks + log2_block_size_in_bytes)-1 
						downto log2_block_size_in_bytes);
	tag_mem_enable <= (enable_sig and (not access_mae))
				when (access_tag_command = CACHE_TAG_INSERT) or 
					(access_tag_command = CACHE_TAG_LOOKUP) else '0';
	tag_mem_write_bar <= '0' when (access_tag_command = CACHE_TAG_INSERT) else '1';
	tag_mem_write_data <= (access_acc & tag_addr_tag);

	------------------------------------------------------------------------------------------------
	--  Registers
	------------------------------------------------------------------------------------------------
	process(clk, reset)
	begin
		if(clk'event and clk = '1') then
			if(reset = '1') then
				access_S_registered <= '0';
				access_mae_registered <= '0';
			
			elsif(enable_sig = '1') then
				access_tag_command_registered <= access_tag_command;	
			   	tag_addr_tag_registered <= tag_addr_tag;
				access_S_registered <= access_S;
				access_is_read_registered <= access_is_read;
				access_is_ifetch_registered <= access_is_ifetch;
			end if;
		end if;
	end process;

	------------------------------------------------------------------------------------------------
	--  Tag memory.
	------------------------------------------------------------------------------------------------
	tagInst: base_bank
		generic map		
			(name => "dcache_tag_memory",
					g_addr_width => log2_number_of_blocks,
					g_data_width => tag_width+3)
		port map (
				datain => tag_mem_write_data,
				dataout => tag_mem_read_data,
				addrin => tag_mem_address, 
				enable => tag_mem_enable,
				writebar => tag_mem_write_bar,
				clk => clk, reset => reset);	
		

	------------------------------------------------------------------------------------------------
	--  output logic
	------------------------------------------------------------------------------------------------
	-- is-hit?
	process(access_tag_command_registered, 
			access_S_registered,
			  access_is_ifetch_registered,
			     access_is_read_registered,
			   	   tag_addr_tag_registered,
					access_mae_registered,
						valid_bit_registered,
							tag_mem_read_data)
		variable hit_var : std_logic := '0';
		variable perms_ok_var : std_logic := '0';
		variable lookup_acc_var : std_logic_vector(2 downto 0);
	begin
		hit_var := '0';
		perms_ok_var := '1';
		lookup_acc_var := (others => '0');

		if((access_mae_registered = '0') and
				(valid_bit_registered = '1') and
				(access_tag_command_registered = CACHE_TAG_LOOKUP)) then
			if(tag_addr_tag_registered = tag_mem_read_data(tag_width-1 downto 0)) then
				lookup_acc_var := tag_mem_read_data (tag_width+2 downto tag_width);
				hit_var := '1';
				perms_ok_var := 
					accessPermissionsOk(access_S_registered,
								access_is_ifetch_registered,
								access_is_read_registered,
								lookup_acc_var);
			end if;
		end if;
		is_hit_sig <= hit_var;
		permissions_ok_sig <= perms_ok_var;
	end process;

	is_hit(0) <= is_hit_sig;
	permissions_ok(0) <= permissions_ok_sig;
			
end Behave;
--
-- Written by Madhav Desai
--
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library AjitCustom;
use AjitCustom.UsefulFunctions.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

library ahir;
use ahir.BaseComponents.all;
use ahir.mem_component_pack.all;
use ahir.Types.all;
use ahir.Utilities.all;

entity GenericCacheTagsWithInvalidate is -- 
  generic (name: string := "anon";
		log2_number_of_blocks: integer := 9; 
		log2_block_size_in_bytes: integer := 6; 
		address_width: integer := 32;
		log2_data_width_in_bytes: integer := 3);
  port ( -- 
    trigger: in std_logic;
    done   : out std_logic;
    init_flag : in  std_logic;
    access_mae : in  std_logic;
    access_S : in  std_logic;
    access_is_read: in std_logic;
    access_is_ifetch: in std_logic;
    access_acc: in std_logic_vector(2 downto 0);
    access_tag_command : in  std_logic_vector(2 downto 0);
    access_tag_addr : in  std_logic_vector(address_width-1 downto 0);
    -- invalidation channel for cache coherence and synonym avoidance.
    invalidate: in std_logic_vector(0 downto 0);
    invalidate_line_address: in std_logic_vector(((address_width-1) - log2_block_size_in_bytes) downto 0);
    is_hit : out  std_logic_vector(0 downto 0);
    permissions_ok : out  std_logic_vector(0 downto 0);
    lookup_acc: out std_logic_vector(2 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity GenericCacheTagsWithInvalidate;
architecture Behave of GenericCacheTagsWithInvalidate is -- 

	-- dcache-tag management commands
	constant CACHE_TAG_LOOKUP	       : std_logic_vector(2 downto 0) := "001";
	constant CACHE_TAG_INSERT	       : std_logic_vector(2 downto 0) := "010";
	constant CACHE_TAG_CLEAR_LINE	       : std_logic_vector(2 downto 0) := "011";
	constant CACHE_TAG_CLEAR_ALL	       : std_logic_vector(2 downto 0) := "100";
	constant CACHE_TAG_NOP	       	       : std_logic_vector(2 downto 0) := "101";

	constant number_of_blocks : integer := (2**log2_number_of_blocks);
	constant bytes_per_block : integer := (2**log2_block_size_in_bytes);
	constant data_width_in_bytes : integer := (2**log2_data_width_in_bytes);
	constant dwords_per_block : integer := (2**(log2_block_size_in_bytes - log2_data_width_in_bytes));
	constant log2_dwords_per_block: integer := (log2_block_size_in_bytes - log2_data_width_in_bytes);


	--  tag width 
	constant tag_width : integer :=  address_width - (log2_number_of_blocks + log2_block_size_in_bytes);
	
	--
	--  memory access signals.
	-- 
	signal  tag_mem_address : std_logic_vector(log2_number_of_blocks-1 downto 0);
	signal  tag_mem_write_data: std_logic_vector(tag_width+2 downto 0);
	signal  tag_mem_read_data: std_logic_vector(tag_width+2 downto 0);
	signal  tag_mem_enable: std_logic;
	signal  tag_mem_write_bar: std_logic;
	
	--
	-- valid bits.. 
	-- 
	signal valid_bits: std_logic_vector (number_of_blocks-1 downto 0);
	
      	

	Type FsmState is (Idle, WaitForReceiveBuffer);
	signal fsm_state: FsmState;
	
	signal valid_bit_registered : std_logic;
	signal latch_request_info: Boolean;

	signal invalidate_missed_cache_line : Boolean;
	signal invalidate_missed_cache_line_block_id : integer range 0 to number_of_blocks-1;


	function blockId (x: std_logic_vector(address_width-1 downto 0)) 
		return integer is
		variable ret_var : integer range 0 to number_of_blocks -1;
		variable block_id_var : std_logic_vector(log2_number_of_blocks-1 downto 0);
	begin
		block_id_var := x ((log2_number_of_blocks + log2_block_size_in_bytes)-1 
							downto log2_block_size_in_bytes);
		ret_var := to_integer(unsigned(block_id_var));
		return(ret_var);

	end blockId;


	-- access-completed-registered.. indicates that
	-- an action has just completed.
	signal access_active, access_completed: Boolean;

	signal is_hit_sig : std_logic;
	signal permissions_ok_sig : std_logic;

	signal  invalidate_block_id_int : integer range 0 to number_of_blocks-1;
	signal  invalidate_word_addr: std_logic_vector(address_width-1 downto 0);

	signal  tag_block_id : std_logic_vector(log2_number_of_blocks-1 downto 0);
	signal  tag_block_id_int : integer range 0 to number_of_blocks-1;
	signal  tag_addr_tag, tag_addr_tag_registered : std_logic_vector(tag_width-1 downto 0);

	signal rx_buf_read_req, rx_buf_read_ack: std_ulogic;

	-- for output stage.
    	signal access_tag_command_registered : std_logic_vector(2 downto 0);
    	signal access_S_registered : std_logic;
	signal access_mae_registered : std_logic;
	signal access_is_ifetch_registered : std_logic;
	signal access_is_read_registered : std_logic;
	signal enable_sig: std_logic;
      
-- see comment above..
--##decl_synopsys_sync_set_reset##

	constant ZZZ: std_logic_vector(log2_block_size_in_bytes-1 downto 0) := (others => '0');
	signal invalidate_word_address: std_logic_vector (address_width-1 downto 0);
begin --  

	invalidate_word_address <= invalidate_line_address & ZZZ;
	invalidate_block_id_int <=  blockId(invalidate_word_address);

	----------------------------------------------------------------------------------
	-- state machine! Assuming that the memory is one-cycle.
	----------------------------------------------------------------------------------
	process(clk, reset, trigger)
	begin 
		if(clk'event and (clk = '1')) then
			if(reset = '1') then
				done <= '0';
			else
				done <= trigger;
			end if;
		end if;
	end process;

	enable_sig <= trigger;

	----------------------------------------------------------------------------------
	-- valid bit manipulation
	----------------------------------------------------------------------------------
	process(clk, access_tag_command, enable_sig, access_mae, tag_block_id_int, valid_bits, init_flag)
		variable next_valid_bits: std_logic_vector (number_of_blocks-1 downto 0);
		variable next_valid_bit_registered: std_logic;
		variable inserted_valid_bit: std_logic;
		variable insert_index: integer range 0 to number_of_blocks-1;
	begin
		next_valid_bits := valid_bits;
		inserted_valid_bit := valid_bits(tag_block_id_int);
		next_valid_bit_registered := '0';

		insert_index := 0;

		if(access_tag_command = CACHE_TAG_INSERT) then
			inserted_valid_bit := '1';
		elsif ((invalidate(0) = '1') or (access_tag_command = CACHE_TAG_CLEAR_LINE)) then
			inserted_valid_bit := '0';
		end if; 

		
		if (access_tag_command = CACHE_TAG_CLEAR_LINE) or (access_tag_command = CACHE_TAG_INSERT) or 
						(invalidate(0) = '1') then

			if(invalidate(0)  = '1') then
				insert_index := invalidate_block_id_int;
			else
				insert_index := tag_block_id_int;
			end if;

			next_valid_bits(insert_index) := inserted_valid_bit;

		elsif (access_tag_command = CACHE_TAG_CLEAR_ALL) then
			next_valid_bits := (others => '0');
		elsif (access_tag_command = CACHE_TAG_LOOKUP) then
			next_valid_bit_registered := inserted_valid_bit;
		end if;

		if(clk'event and clk = '1') then
			--
			-- note that init-flag is asynchronous and can appear at
			-- any time.
			--
			if ((init_flag = '1') or (reset = '1')) then
				valid_bits <= (others => '0');
				valid_bit_registered <= '0';
			elsif  (enable_sig = '1') then
				valid_bits <= next_valid_bits;
				valid_bit_registered <= next_valid_bit_registered;
			end if;	
		end if;
	end process;	
	
	tag_block_id_int <=  blockId(access_tag_addr);
	tag_addr_tag <= access_tag_addr(address_width-1 downto (address_width - tag_width));
	tag_mem_address   <=  access_tag_addr((log2_number_of_blocks + log2_block_size_in_bytes)-1 
						downto log2_block_size_in_bytes);
	tag_mem_enable <= (enable_sig and (not access_mae))
				when (access_tag_command = CACHE_TAG_INSERT) or 
					(access_tag_command = CACHE_TAG_LOOKUP) else '0';
	tag_mem_write_bar <= '0' when (access_tag_command = CACHE_TAG_INSERT) else '1';
	tag_mem_write_data <= (access_acc & tag_addr_tag);

	------------------------------------------------------------------------------------------------
	--  Registers
	------------------------------------------------------------------------------------------------
	process(clk, reset)
	begin
		if(clk'event and clk = '1') then
			if(reset = '1') then
				access_S_registered <= '0';
				access_mae_registered <= '0';
			
			elsif(enable_sig = '1') then
				access_tag_command_registered <= access_tag_command;	
			   	tag_addr_tag_registered <= tag_addr_tag;
				access_S_registered <= access_S;
				access_is_read_registered <= access_is_read;
				access_is_ifetch_registered <= access_is_ifetch;
			end if;
		end if;
	end process;

	------------------------------------------------------------------------------------------------
	--  Tag memory.
	------------------------------------------------------------------------------------------------
	tagInst: base_bank
		generic map		
			(name => "dcache_tag_memory",
					g_addr_width => log2_number_of_blocks,
					g_data_width => tag_width+3)
		port map (
				datain => tag_mem_write_data,
				dataout => tag_mem_read_data,
				addrin => tag_mem_address, 
				enable => tag_mem_enable,
				writebar => tag_mem_write_bar,
				clk => clk, reset => reset);	
		

	------------------------------------------------------------------------------------------------
	--  output logic
	------------------------------------------------------------------------------------------------
	-- is-hit?
	process(access_tag_command_registered, 
			access_S_registered,
			  access_is_ifetch_registered,
			     access_is_read_registered,
			   	   tag_addr_tag_registered,
					access_mae_registered,
						valid_bit_registered,
							tag_mem_read_data)
		variable hit_var : std_logic := '0';
		variable perms_ok_var : std_logic := '0';
		variable lookup_acc_var : std_logic_vector(2 downto 0);
	begin
		hit_var := '0';
		perms_ok_var := '1';
		lookup_acc_var := (others => '0');

		if((access_mae_registered = '0') and
				(valid_bit_registered = '1') and
				(access_tag_command_registered = CACHE_TAG_LOOKUP)) then
			if(tag_addr_tag_registered = tag_mem_read_data(tag_width-1 downto 0)) then
				lookup_acc_var := tag_mem_read_data (tag_width+2 downto tag_width);
				hit_var := '1';
				perms_ok_var := 
					accessPermissionsOk(access_S_registered,
								access_is_ifetch_registered,
								access_is_read_registered,
								lookup_acc_var);
			end if;
		end if;
		lookup_acc <= lookup_acc_var;
		is_hit_sig <= hit_var;
		permissions_ok_sig <= perms_ok_var;
	end process;

	is_hit(0) <= is_hit_sig;
	permissions_ok(0) <= permissions_ok_sig;
			
end Behave;
--
-- Written by Madhav Desai
--
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library AjitCustom;
use AjitCustom.UsefulFunctions.all;
use AjitCustom.AjitCustomComponents.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

library ahir;
use ahir.BaseComponents.all;
use ahir.mem_component_pack.all;
use ahir.Types.all;
use ahir.Utilities.all;

entity GenericDcacheTagsArraysWithInvalidate is -- 
  generic (name: string := "anon";
		log2_number_of_blocks: integer := 9; 
		log2_block_size_in_bytes: integer := 6; 
		address_width: integer := 32;
		log2_data_width_in_bytes: integer := 3);
  port ( -- 
    -- start it off
    trigger		     : in std_logic;
    -- is it done?  This will be asserted for
    -- exactly one clock cycle.
    done		     : out std_logic;
    
    init_flag : in  std_logic;
    access_mae : in  std_logic;
    access_S : in  std_logic;
    access_is_read: in std_logic;
    access_is_ifetch: in std_logic;
    access_acc: in std_logic_vector(2 downto 0);
    access_tag_command : in  std_logic_vector(2 downto 0);
    access_tag_addr : in  std_logic_vector(address_width-1 downto 0);
    -- invalidation channel for cache coherence and synonym avoidance.
    invalidate: in std_logic_vector(0 downto 0);
    invalidate_line_address: in std_logic_vector(((address_width-1) - log2_block_size_in_bytes) downto 0);
    is_hit : out  std_logic_vector(0 downto 0);
    permissions_ok : out  std_logic_vector(0 downto 0);
    access_array_command : in  std_logic_vector(2 downto 0);
    access_byte_mask : in  std_logic_vector((2**log2_data_width_in_bytes)-1 downto 0);
    access_array_addr : in  std_logic_vector(address_width-1 downto 0);
    access_dword : in  std_logic_vector((8*(2**log2_data_width_in_bytes))-1 downto 0);
    dword_out : out  std_logic_vector((8*(2**log2_data_width_in_bytes))-1 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity GenericDcacheTagsArraysWithInvalidate;
architecture Structural of GenericDcacheTagsArraysWithInvalidate is -- 
	signal tags_done, arrays_done: std_logic;
	signal lookup_acc: std_logic_vector(2 downto 0);
begin --  
	done <= tags_done and arrays_done;

        tagsInst: GenericCacheTagsWithInvalidate
                        generic map (name => "dcache-tags",
                                        log2_number_of_blocks => log2_number_of_blocks, -- 9  
                                        log2_block_size_in_bytes => log2_block_size_in_bytes, -- 6
                                        address_width => address_width,
                                        log2_data_width_in_bytes => log2_data_width_in_bytes)
			port map (
					trigger => trigger,	
					done => tags_done,	
					init_flag => init_flag,
					access_mae => access_mae,
					access_S => access_S,
					access_is_read => access_is_read,
					access_is_ifetch => access_is_ifetch,
					access_acc => access_acc,
					access_tag_command => access_tag_command,
					access_tag_addr => access_tag_addr,
					invalidate => invalidate,
					invalidate_line_address => invalidate_line_address,
					is_hit => is_hit,
					permissions_ok => permissions_ok,
					lookup_acc => lookup_acc,
					clk => clk, reset => reset);

	   arrayInst: GenericCacheArray 
  			generic map (name => "dcache-array",
                                        log2_number_of_blocks => log2_number_of_blocks, -- 9  
                                        log2_block_size_in_bytes => log2_block_size_in_bytes, -- 6
                                        address_width => address_width,
					log2_data_width_in_bytes => log2_data_width_in_bytes)
			port map (
    					trigger => trigger,
    					done => arrays_done,
    					access_mae  => access_mae ,
    					access_array_command  => access_array_command ,
    					access_byte_mask  => access_byte_mask,
    					access_array_addr  => access_array_addr,
    					access_dword  => access_dword,
    					dword_out  => dword_out,
    					clk => clk,
					reset => reset
				);
	
end Structural;
--
-- Written by Madhav Desai
--   no byte-enables needed!
--
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.BaseComponents.all;
use ahir.mem_component_pack.all;
use ahir.Types.all;
use ahir.Utilities.all;

entity GenericIcacheArray is -- 
  generic (name: string := "anon";
		log2_number_of_blocks: integer := 9; 
		log2_block_size_in_bytes: integer := 6; 
		address_width: integer := 32;
		tag_length: integer := 1;
		log2_data_width_in_bytes: integer := 3);
  port ( -- 
    trigger: in std_logic;
    done: out std_logic;
    access_mae : in  std_logic;
    access_array_command : in  std_logic_vector(2 downto 0);
    access_array_addr : in  std_logic_vector(address_width-1 downto 0);
    access_dword : in  std_logic_vector((8*(2**log2_data_width_in_bytes))-1 downto 0);
    dword_out : out  std_logic_vector((8*(2**log2_data_width_in_bytes))-1 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity GenericIcacheArray;
architecture Behave of GenericIcacheArray is -- 

	-- dcache-array management commands
	constant CACHE_ARRAY_READ_DWORD  	: std_logic_vector(2 downto 0) := "001";
	constant CACHE_ARRAY_WRITE_DWORD  	: std_logic_vector(2 downto 0) := "010";
	constant CACHE_ARRAY_NOP	     	: std_logic_vector(2 downto 0) := "011";

	constant number_of_blocks : integer := (2**log2_number_of_blocks);
	constant bytes_per_block : integer := (2**log2_block_size_in_bytes);
	constant data_width_in_bytes : integer := (2**log2_data_width_in_bytes);
	constant dwords_per_block : integer := (2**(log2_block_size_in_bytes - log2_data_width_in_bytes));
	constant log2_dwords_per_block: integer := (log2_block_size_in_bytes - log2_data_width_in_bytes);


	--  tag width 
	constant tag_width : integer :=  address_width - (log2_number_of_blocks + log2_block_size_in_bytes);
	
	--
	--  memory access signals.
	-- 
	signal  array_mem_address : std_logic_vector((log2_number_of_blocks + log2_block_size_in_bytes - log2_data_width_in_bytes)-1 downto 0);
	signal  array_mem_write_data: std_logic_vector((8*data_width_in_bytes)-1 downto 0);
	signal  array_mem_read_data: std_logic_vector((8*data_width_in_bytes)-1 downto 0);
	signal  array_mem_enable: std_logic;
	signal  array_mem_write_bar: std_logic;

	signal fin_ack_sig, enable_sig: std_logic;
	signal dword_out_sig : std_logic_vector((8*(2**log2_data_width_in_bytes))-1 downto 0);
	signal selected_dword_from_access_cache_line : 
		std_logic_vector((8*(2**log2_data_width_in_bytes))-1 downto 0);
	signal selected_dword_from_mem_read_data : 
		std_logic_vector((8*(2**log2_data_width_in_bytes))-1 downto 0);

	signal  access_array_command_registered : std_logic_vector(2 downto 0);
	signal  array_mem_offset_in_line_registered: integer range 0 to dwords_per_block-1;
	signal  access_mae_registered: std_logic;
	signal  access_dword_registered : std_logic_vector(access_dword'length-1 downto 0);
begin --  

	----------------------------------------------------------------------------------
	-- Assuming that the memory is one-cycle.
	----------------------------------------------------------------------------------
	process(clk, reset, trigger)
	begin 
		enable_sig <= trigger;
		if(clk'event and (clk = '1')) then
			if(reset = '1') then
				done <= '0';
			else
				done <= trigger;
			end if;
		end if;
	end process;


	----------------------------------------------------------------------------------
	-- prepare inputs to memory.
	--    If the current address is A[31:0], then A[14:6] is the address of the line.
	--    index into array is A[14:3].
	----------------------------------------------------------------------------------
	-- (9 + 6 - 1) downto 3. OK.
	array_mem_address <= access_array_addr ((log2_number_of_blocks + log2_block_size_in_bytes)-1 downto log2_data_width_in_bytes);
	array_mem_enable <= (enable_sig and (not access_mae));
	array_mem_write_bar  <= '0' when (access_array_command =  CACHE_ARRAY_WRITE_DWORD) else '1';
	array_mem_write_data <= access_dword;

	bb: base_bank
			generic map 
			(name => "IcacheArrayBaseBank",
					-- address width is 9+3 = 12.
				g_addr_width => 
					(log2_number_of_blocks + log2_block_size_in_bytes 
								- log2_data_width_in_bytes),
					-- data width is 64 bits.
				g_data_width => 8*data_width_in_bytes)
			port map (
					datain => array_mem_write_data,
					dataout => array_mem_read_data,
					addrin => array_mem_address, 
					enable => array_mem_enable,
					writebar => array_mem_write_bar,
					clk => clk, reset => reset);	
		
	------------------------------------------------------------------------------------------------
	--  mux, register and forward to output stage
	------------------------------------------------------------------------------------------------
	process(clk, reset)
	begin
		if clk'event and clk = '1' then
			if(reset ='1')  then
				access_array_command_registered <= (others => '0');
				access_mae_registered <= '0';
			elsif (enable_sig = '1') then
				access_array_command_registered <= access_array_command;
				access_mae_registered <= access_mae;
				access_dword_registered <= access_dword;
			end if;
		end if;
	end process;

	------------------------------------------------------------------------------------------------
	--  output logic
	------------------------------------------------------------------------------------------------
	dword_out <= (others => '0') when access_mae_registered = '1' 
			else array_mem_read_data when (access_array_command_registered = CACHE_ARRAY_READ_DWORD)
				else  access_dword_registered;
end Behave;
--
-- Written by Madhav Desai
--
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library AjitCustom;
use AjitCustom.UsefulFunctions.all;
use AjitCustom.AjitCustomComponents.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

library ahir;
use ahir.BaseComponents.all;
use ahir.mem_component_pack.all;
use ahir.Types.all;
use ahir.Utilities.all;

entity GenericIcacheTagsArraysWithInvalidate is -- 
  generic (name: string := "anon";
		log2_number_of_blocks: integer := 9; 
		log2_block_size_in_bytes: integer := 6; 
		address_width: integer := 32;
		log2_data_width_in_bytes: integer := 3);
  port ( -- 
    -- start it off
    trigger		     : in std_logic;
    -- is it done?  This will be asserted for
    -- exactly one clock cycle.
    done		     : out std_logic;
    
    init_flag : in  std_logic;
    access_mae : in  std_logic;
    access_S : in  std_logic;
    access_is_read: in std_logic;
    access_is_ifetch: in std_logic;
    access_acc: in std_logic_vector(2 downto 0);
    access_tag_command : in  std_logic_vector(2 downto 0);
    -- invalidation channel for cache coherence and synonym avoidance.
    invalidate: in std_logic_vector(0 downto 0);
    invalidate_line_address: in std_logic_vector(((address_width-1) - log2_block_size_in_bytes) downto 0);
    is_hit : out  std_logic_vector(0 downto 0);
    permissions_ok : out  std_logic_vector(0 downto 0);
    lookup_acc: out std_logic_vector(2 downto 0);
    access_array_command : in  std_logic_vector(2 downto 0);
    access_addr : in  std_logic_vector(address_width-1 downto 0);
    access_dword : in  std_logic_vector((8*(2**log2_data_width_in_bytes))-1 downto 0);
    dword_out : out  std_logic_vector((8*(2**log2_data_width_in_bytes))-1 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity GenericIcacheTagsArraysWithInvalidate;
architecture Structural of GenericIcacheTagsArraysWithInvalidate is -- 
	signal tags_done, arrays_done: std_logic;
begin --  
	done <= tags_done and arrays_done;

        tagsInst: GenericCacheTagsWithInvalidate
                        generic map (name => "icache-tags",
                                        log2_number_of_blocks => log2_number_of_blocks, -- 9  
                                        log2_block_size_in_bytes => log2_block_size_in_bytes, -- 6
                                        address_width => address_width,
                                        log2_data_width_in_bytes => log2_data_width_in_bytes)
			port map (
					trigger => trigger,	
					done => tags_done,	
					init_flag => init_flag,
					access_mae => access_mae,
					access_S => access_S,
					access_is_read => access_is_read,
					access_is_ifetch => access_is_ifetch,
					access_acc => access_acc,
					access_tag_command => access_tag_command,
					access_tag_addr => access_addr,
					invalidate => invalidate,
					invalidate_line_address => invalidate_line_address,
					is_hit => is_hit,
					permissions_ok => permissions_ok,
					lookup_acc => lookup_acc,
					clk => clk, reset => reset);

	   arrayInst: GenericIcacheArray 
  			generic map (name => "dcache-array",
                                        log2_number_of_blocks => log2_number_of_blocks, -- 9  
                                        log2_block_size_in_bytes => log2_block_size_in_bytes, -- 6
                                        address_width => address_width,
					log2_data_width_in_bytes => log2_data_width_in_bytes)
			port map (
    					trigger => trigger,
    					done => arrays_done,
    					access_mae  => access_mae ,
    					access_array_command  => access_array_command ,
    					access_array_addr  => access_addr,
    					access_dword  => access_dword,
    					dword_out  => dword_out,
    					clk => clk,
					reset => reset
				);
	
end Structural;
--
-- Written by Madhav Desai
--
library std;
use std.standard.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.BaseComponents.all;
use ahir.mem_component_pack.all;
use ahir.Types.all;
use ahir.Utilities.all;

library AjitCustom;
use AjitCustom.CachePackage.all;


-- line data in Cache.  Organized into 
-- sets.  For example if associativity is 2 (i.e. log2_associativity = 1),
--
-- Address of a dword-pair  is
--       set-id   offset-in-line
--       [10:3]   [2:0]		
--       set_id offset_in_line  zero3
--  
--
-- with data width = 16 bytes..
--
-- There will be 2 banks, bank 0 keeps data with index-in-set=0,
-- bank1 keeps data with index-in-set=1.
--
--
entity GenericSetAssociativeCacheArray is -- 
  generic (name: string := "anon";
		log2_number_of_blocks: integer := 9; 
		log2_block_size_in_bytes: integer := 6; 
		log2_associativity: integer := 1;
		address_width: integer := 32;
		log2_data_width_in_bytes: integer := 3;
		ignore_byte_mask: boolean := false);
  port ( -- 
     -- it is the responsibility of the one who triggers the activity
     -- to ensure that the match_index_in_set field is valid!
    trigger: in std_logic;
    done: out std_logic;
    matched_index_in_set: in std_logic_vector(log2_associativity-1 downto 0);
    access_mae : in  std_logic;
    access_array_command : in  std_logic_vector(2 downto 0);
    access_byte_mask : in  std_logic_vector((2**log2_data_width_in_bytes)-1 downto 0);
    access_array_addr : in  std_logic_vector(address_width-1 downto 0);
    access_array_write_dword : 
	in  std_logic_vector(8*((2**log2_data_width_in_bytes))-1 downto 0);
    access_array_read_dword_vector : 
	out  std_logic_vector(((2**log2_associativity)*8*(2**log2_data_width_in_bytes))-1 downto 0);
    bypassed_dword_out : 
	out  std_logic_vector((8*(2**log2_data_width_in_bytes))-1 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity GenericSetAssociativeCacheArray;
architecture Behave of GenericSetAssociativeCacheArray is -- 
	constant associativity: integer := 2**log2_associativity;


	constant number_of_blocks : integer := (2**log2_number_of_blocks);
	constant bytes_per_block : integer := (2**log2_block_size_in_bytes);
	constant data_width_in_bytes : integer := (2**log2_data_width_in_bytes);
	constant dwords_per_block : integer := (2**(log2_block_size_in_bytes - log2_data_width_in_bytes));
	constant log2_dwords_per_block: integer := (log2_block_size_in_bytes - log2_data_width_in_bytes);

	--
	--  memory access signals... 
	-- 

	-- the number of distinct memory locations is number of dwords / associativity.
	signal  array_mem_address : 
		std_logic_vector((log2_number_of_blocks + log2_dwords_per_block - log2_associativity)-1 downto 0);
	
	type    MemDataWordArray is array (natural range <>) 
				of std_logic_vector((8*data_width_in_bytes)-1 downto 0);

	-- number of dword-width banks is = associativity.
	signal  array_mem_write_data: MemDataWordArray (associativity-1 downto 0);
	signal  array_mem_read_data: MemDataWordArray (associativity-1 downto 0);

	type    ByteEnableArray is array (natural range <>) 
				of std_logic_vector(data_width_in_bytes-1 downto 0);
	signal  array_mem_byte_enable: ByteEnableArray(associativity-1 downto 0);

	signal  array_mem_enable: std_logic;
	signal  array_mem_set_enable: std_logic_vector(associativity-1 downto 0);

	signal  array_mem_write_bar: std_logic;

	signal  enable_sig: std_logic;
	signal  access_dword_registered : 
			std_logic_vector((8*data_width_in_bytes)-1 downto 0);

		
	signal dbg_signal: std_logic;
	signal dbg_int_signal: integer range 0 to associativity-1;
begin --  
	process(clk, reset, trigger)
	begin
		if(clk'event and clk = '1') then
			if(reset = '1') then
				done <= '0';
			else
				done <= trigger;
			end if;
		end if;
	end process;
	enable_sig <= trigger;

	----------------------------------------------------------------------------------
	-- prepare inputs to memory.
	----------------------------------------------------------------------------------

	-- address is determined by set-id, dword-index-in-block.
	array_mem_address <= 
		access_array_addr ((log2_number_of_blocks + log2_dwords_per_block + log2_data_width_in_bytes - log2_associativity)-1
									downto log2_data_width_in_bytes);

	-- enable write only if matched index in set is valid 
	--   This is guaranteed by the one who triggers this module.
	array_mem_enable <= (enable_sig and (not access_mae));
	array_mem_write_bar <= '0' when (access_array_command =  CACHE_ARRAY_WRITE_DWORD) else '1';

	--------------------------------------------------------
	-- byte mask!
	--------------------------------------------------------
	dbg_int_signal <= to_integer(unsigned(matched_index_in_set));
	process(access_byte_mask, array_mem_enable, dbg_int_signal, access_array_command, access_array_write_dword)
		variable sel_var: std_logic;
		variable dbg_signal_var: std_logic;
		variable be_var: std_logic_vector(data_width_in_bytes-1 downto 0);
		variable  array_mem_write_data_var: MemDataWordArray (associativity-1 downto 0);
		variable  array_mem_byte_enable_var: ByteEnableArray(associativity-1 downto 0);
		variable  array_mem_set_enable_var: std_logic_vector(associativity-1 downto 0);
	begin
		sel_var := '0';
		dbg_signal_var := '0';
		be_var := (others => '0');

		array_mem_write_data_var  := (others => (others => '0'));
		array_mem_byte_enable_var := (others => (others => '0'));
		array_mem_set_enable_var  := (others => '0');

		for A in 0 to associativity-1 loop
			if(access_array_command = CACHE_ARRAY_READ_DWORD) then 

				array_mem_write_data_var(A)  := (others => '0');
				array_mem_byte_enable_var(A) := (others => '1');
				array_mem_set_enable_var(A) := array_mem_enable;

			elsif (A = dbg_int_signal) then

				sel_var := '1';
				dbg_signal_var := '1';
			
				if (access_array_command = CACHE_ARRAY_WRITE_DWORD) then
					array_mem_write_data_var(A) := access_array_write_dword;
					array_mem_set_enable_var(A) := array_mem_enable;

					for B in data_width_in_bytes-1 downto 0 loop
						array_mem_byte_enable_var(A)(B) := array_mem_enable and access_byte_mask(B);
					end loop;
				end if;
			end if;
		end loop;

		array_mem_write_data <= array_mem_write_data_var;
		array_mem_byte_enable <= array_mem_byte_enable_var;
		array_mem_set_enable <= array_mem_set_enable_var;

		dbg_signal <= dbg_signal_var;
	end process;	

	------------------------------------------------------------------------------------------------
	--  register and forward to output stage
	------------------------------------------------------------------------------------------------
	process(clk, reset, access_array_write_dword, access_array_command, access_mae)
	begin
		if clk'event and clk = '1' then
			if (enable_sig = '1') then
				access_dword_registered <= access_array_write_dword;
			end if;
		end if;
	end process;

	------------------------------------------------------------------------------------------------
	-- set + line banks
	------------------------------------------------------------------------------------------------
	SetBankGen: for A in associativity-1 downto 0 generate

	  withByteMask: if (not ignore_byte_mask) generate 
            lineBankGen: for B in data_width_in_bytes-1 downto 0 generate
	    
		lineBank: base_bank
				generic map (name => "linBank_" & Convert_To_String(B),
						g_addr_width => 
							log2_number_of_blocks + log2_dwords_per_block 
										- log2_associativity,
						g_data_width => 8)
				port map (
						datain => 
							array_mem_write_data(A)(((B+1)*8)-1 downto (B*8)),
						dataout => 
							array_mem_read_data(A)(((B+1)*8)-1 downto (B*8)),
						addrin => array_mem_address, 
						enable => array_mem_byte_enable(A)(B),
						writebar => array_mem_write_bar,
						clk => clk, reset => reset);	
            end generate LineBankGen;
          end generate withByteMask;

          ignoreByteMask: if ignore_byte_mask generate
             setBank: base_bank
				generic map (name => "setBank_" & Convert_To_String(A),
						g_addr_width => 
							log2_number_of_blocks + log2_dwords_per_block 
										- log2_associativity,
						g_data_width => 8*data_width_in_bytes)
				port map (
						datain => array_mem_write_data(A),
						dataout => array_mem_read_data(A),
						addrin => array_mem_address, 
						enable => array_mem_set_enable(A),
						writebar => array_mem_write_bar,
						clk => clk, reset => reset);	
	   end generate ignoreByteMask;

	end generate SetBankGen;
		
	------------------------------------------------------------------------------------------------
	--  output logic
	------------------------------------------------------------------------------------------------
	-- all entries in the set are presented to the output word.
	process(array_mem_read_data)
	begin
		for A in associativity-1 downto 0 loop
			access_array_read_dword_vector (((A+1)*8*data_width_in_bytes)-1  downto (A*8*data_width_in_bytes))
						 <= array_mem_read_data(A);
		end loop;
	end process;
	bypassed_dword_out <= access_dword_registered;

end Behave;
--
-- Written by Madhav Desai
--
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library AjitCustom;
use AjitCustom.UsefulFunctions.all;
use AjitCustom.AjitCustomComponents.all;
use AjitCustom.CachePackage.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

library ahir;
use ahir.BaseComponents.all;
use ahir.mem_component_pack.all;
use ahir.Types.all;
use ahir.Utilities.all;

--
--  tags and arrays..
--      For every triggering of this module, there
--      is a specified tag operation (lookup/insert/clear0
--      and a specified array operation (write/read).
--
--  To execute the array operation, we need to know the
--  location of the address in the set.   This is available
--  one cycle after the triggering.  For a naive implementation,
--  this would imply that the array operation is started one
--  cycle after the triggering.
--
--  Instead, we use a small TLB to store address -> index
--  translations which if there is a match imply that
--  the array write access can start simultaneously with
--  the tag lookup.
--
--  The Tlb is updated every time a tag lookup/insert
--  completes..
--
-- 
--  Pairs
--      tag 		array
--       lookup         read/write
--            On write, wait for tlb hit
--            or tag hit.  If hit, proceed
--            else nop.
--
--            On read, do array read and
--            tag read in parallel.
--
--       insert         write
--            For array, if va-tlb-miss,
--            wait on tag information.
--            start tag access immediately,
--            possibly using tlb match information.
--
--       Note: insert may create new entry or overwrite
--             existing entry in set and tlb..
--            
--       nop            write
--          (does this modify tlb structure?  No)
--             tlb must hit. if not write is a nop.
--
--       erase          nop
--          erase set (whole set) and tlb entry
--
--       clear          nop
--          clear all sets and entire tlb 
--
--       nop            nop
--
entity GenericSetAssociativeCacheTagsArraysWithInvalidate is -- 
  generic (
		name: string := "anon";
		log2_number_of_blocks: integer := 9; 
		log2_block_size_in_bytes: integer := 6; 
		log2_associativity: integer := 1;
		address_width: integer := 32;
		log2_data_width_in_bytes: integer := 3;
		icache_flag: boolean := false
	  );
  port ( -- 
    -- start it off
    trigger		     : in std_logic;
    -- is it done?  This will be asserted for
    -- exactly one clock cycle.
    done		     : out std_logic;
    
    init_flag : in  std_logic;
    access_mae : in  std_logic;
    access_S : in  std_logic;
    access_is_read: in std_logic;
    access_is_ifetch: in std_logic;
    access_acc: in std_logic_vector(2 downto 0);
    access_tag_lookup : in  std_logic;
    access_tag_clear_line : in  std_logic;
    access_tag_clear_all : in  std_logic;
    access_tag_insert : in  std_logic;
    access_array_command : in  std_logic_vector(2 downto 0);
    access_addr : in  std_logic_vector(address_width-1 downto 0);
    access_byte_mask : in  std_logic_vector((2**log2_data_width_in_bytes)-1 downto 0);
    access_dword : in  std_logic_vector((8*(2**log2_data_width_in_bytes))-1 downto 0);
    -- invalidation channel for cache coherence and synonym avoidance.
    invalidate: in std_logic_vector(0 downto 0);
    invalidate_line_address: in std_logic_vector(((address_width-1) - log2_block_size_in_bytes) downto 0);
    is_hit : out  std_logic_vector(0 downto 0);
    permissions_ok : out  std_logic_vector(0 downto 0);
    lookup_acc : out  std_logic_vector(2 downto 0);
    dword_out : out  std_logic_vector((8*(2**log2_data_width_in_bytes))-1 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity GenericSetAssociativeCacheTagsArraysWithInvalidate;

architecture Structural of GenericSetAssociativeCacheTagsArraysWithInvalidate is -- 
	constant associativity: integer := 2**log2_associativity;
	constant data_width_in_bytes: integer := 2**log2_data_width_in_bytes;
	constant log2_number_of_sets : integer := log2_number_of_blocks - log2_associativity;
	constant number_of_sets : integer := 2**log2_number_of_sets;

	signal tags_trigger, tags_done, arrays_trigger, arrays_done: std_logic;
	signal access_array_read_dword_vector: std_logic_vector((associativity*8*data_width_in_bytes)-1 downto 0);
    	signal bypassed_dword_out : std_logic_vector((8*data_width_in_bytes)-1 downto 0);
    	signal dword_out_pre_reg, dword_out_reg : std_logic_vector((8*(2**log2_data_width_in_bytes))-1 downto 0);

	signal tags_busy, tags_lookup_is_valid, tags_index_in_set_is_valid: std_logic;
	signal tags_index_in_set : std_logic_vector (log2_associativity-1 downto 0);
	signal tags_acc: std_logic_vector(2 downto 0);

    	signal tlb_to_tag_valid_match: std_logic;
    	signal tlb_to_tag_match_index_in_set: std_logic_vector(log2_associativity-1 downto 0);

	signal array_read_dword, array_write_dword: std_logic;
	signal array_read_dword_reg: std_logic;

    	signal access_array_command_qualified : std_logic_vector(2 downto 0);
    	signal access_addr_qualified : std_logic_vector(address_width-1 downto 0);
    	signal access_byte_mask_qualified : std_logic_vector((2**log2_data_width_in_bytes)-1 downto 0);
    	signal access_dword_qualified : std_logic_vector((8*(2**log2_data_width_in_bytes))-1 downto 0);

	type ArrayFsmState is (ARRAY_IDLE, ARRAY_WAIT_ON_TAGS);
	signal array_fsm_state : ArrayFsmState;

	type ToplevelFsmState is (IDLE_STATE, WAIT_STATE, TAGS_DONE_STATE, ARRAYS_DONE_STATE);
	signal fsm_state: ToplevelFsmState;

	constant line_address_width: integer := (address_width - log2_block_size_in_bytes);
	signal va_tlb_lookup, va_tlb_insert, va_tlb_erase, va_tlb_clear, va_tlb_match: std_logic;
	signal va_tlb_lookup_va_tag, va_tlb_insert_va_tag, va_tlb_erase_va_tag: 
					std_logic_vector((line_address_width-log2_number_of_sets)-1 downto 0);
	signal va_tlb_lookup_set_id, va_tlb_insert_set_id, va_tlb_erase_set_id: 
					std_logic_vector(log2_number_of_sets-1 downto 0);
	signal va_tlb_insert_index_in_set: std_logic_vector(log2_associativity-1 downto 0);
	signal va_tlb_insert_acc: std_logic_vector(3-1 downto 0);

	signal va_tlb_lookup_index_in_set, va_tlb_matched_index_in_set : std_logic_vector (log2_associativity-1 downto 0);
	signal va_tlb_lookup_acc, va_tlb_matched_acc : std_logic_vector (3-1 downto 0);
	
	signal arrays_matched_index_in_set:  std_logic_vector (log2_associativity-1 downto 0);
	signal arrays_matched_index_in_set_reg:  std_logic_vector (log2_associativity-1 downto 0);


	signal tags_hit, tags_miss, tags_insert_done: std_logic;
	signal tags_hit_reg, tags_miss_reg: std_logic;
	signal cpu_permissions_ok, cpu_permissions_ok_reg: std_logic;
	signal va_tlb_match_hit, va_tlb_match_miss, va_tlb_cpu_permissions_ok: std_logic;

    	signal access_mae_reg, access_mae_qualified : std_logic;
    	signal access_S_reg : std_logic;
    	signal access_is_read_reg:std_logic;
    	signal access_is_ifetch_reg:std_logic;
    	signal access_acc_reg:std_logic_vector(2 downto 0);
    	signal access_tag_lookup_reg, access_tag_insert_reg,
			access_tag_clear_line_reg, access_tag_clear_all_reg :std_logic;
    	signal access_array_command_reg :std_logic_vector(2 downto 0);
    	signal access_array_command_final :std_logic_vector(2 downto 0);
    	signal access_addr_reg :std_logic_vector(address_width-1 downto 0);
    	signal access_byte_mask_reg :std_logic_vector((2**log2_data_width_in_bytes)-1 downto 0);
    	signal access_dword_reg :std_logic_vector((8*(2**log2_data_width_in_bytes))-1 downto 0);
	
	signal debug_sig_0: std_logic;
begin --  
	-----------------------------------------------------------------------------------------------------
	-- permissions ok from tag lookup ....
	-----------------------------------------------------------------------------------------------------
	cpu_permissions_ok <= 
		accessPermissionsOk (access_S_reg, access_is_ifetch_reg, 
					access_is_read_reg, tags_acc) and access_tag_lookup_reg;
	lookup_acc <= tags_acc;
	tags_hit  <= cpu_permissions_ok and tags_done and tags_lookup_is_valid and access_tag_lookup_reg;
	tags_miss <= tags_done and ((not cpu_permissions_ok) or (not tags_lookup_is_valid)) and access_tag_lookup_reg;
	tags_insert_done <= tags_done and access_tag_insert_reg;

	process(tags_trigger, va_tlb_match, va_tlb_lookup_acc, 
			access_tag_lookup, access_tag_lookup_reg,
			access_tag_insert, access_tag_insert_reg,
			access_acc, access_S, access_is_ifetch, access_is_read,
			access_acc_reg, access_S_reg, access_is_ifetch_reg, access_is_read_reg) 
		variable S,ifetch,read, perms_ok: std_logic;	
		variable acc_var: std_logic_vector(2 downto 0);
		variable lookup_var : std_logic;

	begin
		S := access_S; ifetch := access_is_ifetch; read := access_is_read;

		-- acc-var by default allows only reads..
		lookup_var := '0';
		acc_var := va_tlb_lookup_acc;

		if(tags_trigger = '0') then
			S := access_S_reg; ifetch := access_is_ifetch_reg; read := access_is_read_reg;
			lookup_var := access_tag_lookup_reg;
		else
			lookup_var := access_tag_lookup;
		end if;

		-- permissions should be checked only in lookups!!
		perms_ok := (not lookup_var) or accessPermissionsOk(S, ifetch, read, acc_var);

		va_tlb_match_hit <= va_tlb_match and perms_ok;
		va_tlb_match_miss <= va_tlb_match and (not perms_ok);

	end process;


	-------------------------------------------------------------------------------------
	--  arrays control state machine...
	--          On trigger: 
	--             if read_dword/write_dword, wait until tlb match or tags done.. and then trigger
	--             arrays.
	-------------------------------------------------------------------------------------
	process(clk, reset, trigger, 
			access_mae, access_mae_reg,
			access_array_command, access_array_command_reg,
			access_dword,  access_dword_reg,
			access_addr, access_addr_reg, 
			va_tlb_lookup_index_in_set,
			tags_index_in_set,
			tags_trigger,
			tags_miss, va_tlb_match_miss, va_tlb_match_hit,
			tags_hit, tags_insert_done,
			array_fsm_state)
		variable next_array_fsm_state_var: ArrayFsmState;
		variable trigger_array_var : std_logic;

		variable command_var: std_logic_vector(2 downto 0);
		variable addr_var: std_logic_vector(address_width-1 downto 0);
    		variable access_dword_var : std_logic_vector((8*(2**log2_data_width_in_bytes))-1 downto 0);
    		variable access_byte_mask_var : std_logic_vector((2**log2_data_width_in_bytes)-1 downto 0);
		variable matched_index_var : std_logic_vector (log2_associativity-1 downto 0);
		variable access_mae_var: std_logic;
	begin
		next_array_fsm_state_var := array_fsm_state;
		matched_index_var := (others => '0');
		trigger_array_var := '0';
		command_var := CACHE_ARRAY_NOP;

		access_dword_var := (others => '0');
		access_byte_mask_var := (others => '0');
		access_mae_var := access_mae;

		case array_fsm_state is 

			when ARRAY_IDLE =>
				addr_var := access_addr;
				access_byte_mask_var := access_byte_mask;
				access_dword_var := access_dword;
				addr_var := access_addr;

				if(tags_trigger = '1') then

					--
					-- NOTE: the cache array write can proceed only after we
					--       know that there was a hit!
					--
					if(access_array_command  = CACHE_ARRAY_WRITE_DWORD) then
						if (va_tlb_match_hit = '1') then
							trigger_array_var := '1';	
							command_var := CACHE_ARRAY_WRITE_DWORD;
							matched_index_var := va_tlb_lookup_index_in_set;
						elsif (va_tlb_match_miss = '1') then
							trigger_array_var := '1';	
						else
							next_array_fsm_state_var := ARRAY_WAIT_ON_TAGS;
						end if;
					--
					-- NOTE: the cache array read can proceed even without a tlb 
					--       hit.
					else
						trigger_array_var := '1';	
						command_var := access_array_command;
					end if;
				end if;
			when ARRAY_WAIT_ON_TAGS => 
				-- Come here only on write dword....
				addr_var := access_addr_reg;
				access_byte_mask_var := access_byte_mask_reg;
				access_dword_var := access_dword_reg;
				access_mae_var := access_mae_reg;

				if (tags_miss = '1') then
					trigger_array_var := '1';	
					next_array_fsm_state_var := ARRAY_IDLE;

					command_var := CACHE_ARRAY_NOP;

				elsif ((tags_hit = '1') or (tags_insert_done = '1')) then

					trigger_array_var := '1';	
					command_var := access_array_command_reg;
					matched_index_var := tags_index_in_set;

					next_array_fsm_state_var := ARRAY_IDLE;
				end if;
		end case;

		arrays_trigger <= trigger_array_var;
		access_array_command_qualified <= command_var;
		access_byte_mask_qualified <= access_byte_mask_var;
		access_addr_qualified <= addr_var;
		access_dword_qualified <= access_dword_var;
		arrays_matched_index_in_set <= matched_index_var;
		access_mae_qualified <= access_mae_var;
			

		if(clk'event and (clk = '1')) then
			if(reset = '1') then
				array_fsm_state <= ARRAY_IDLE;
			else
				array_fsm_state <= next_array_fsm_state_var;
				if(trigger_array_var = '1') then
					arrays_matched_index_in_set_reg <= matched_index_var;
				end if;
			end if;
		end if;
	end process;
	
	-----------------------------------------------------------------------------
	--  top-level state machine.
	-----------------------------------------------------------------------------
	process(clk, reset, fsm_state, trigger,tags_done, arrays_done, array_read_dword)
		variable next_fsm_state_var: ToplevelFsmState;
		variable done_var: std_logic;
		variable register_args_var: boolean;
		variable tags_trigger_var : std_logic;
	begin
		next_fsm_state_var := fsm_state;
		done_var := '0';
		register_args_var := false;
		tags_trigger_var := '0';

		case fsm_state is
			when IDLE_STATE =>
				if (trigger = '1') then 
					next_fsm_state_var := WAIT_STATE;
					register_args_var := true;
					tags_trigger_var := '1';
				end if;
			when WAIT_STATE =>
				if((tags_done = '1') and (arrays_done = '1')) then
					done_var := '1';
					if(trigger = '1') then 
						register_args_var := true;
						tags_trigger_var := '1';
					else
						next_fsm_state_var := IDLE_STATE;
					end if;
				elsif (tags_done = '1') then
					next_fsm_state_var := TAGS_DONE_STATE;
				elsif (arrays_done = '1') then
					next_fsm_state_var := ARRAYS_DONE_STATE;
				end if;
			when TAGS_DONE_STATE => 
				if(arrays_done = '1') then
					done_var := '1';
					if(trigger = '1') then 
						next_fsm_state_var := WAIT_STATE;
						register_args_var := true;
						tags_trigger_var := '1';
					else 
						next_fsm_state_var := IDLE_STATE;
					end if;
				end if;
			when ARRAYS_DONE_STATE => 
				if(tags_done = '1') then
					done_var := '1';
					if(trigger = '1') then 
						next_fsm_state_var := WAIT_STATE;
						register_args_var := true;
						tags_trigger_var := '1';
					else 
						next_fsm_state_var := IDLE_STATE;
					end if;
				end if;
					
		end case;

		done <= done_var;
		tags_trigger <=	tags_trigger_var;

		if(clk'event and (clk = '1')) then
			if(reset = '1') then
				fsm_state <= IDLE_STATE;
			else
				fsm_state <= next_fsm_state_var;
				if(register_args_var) then
					access_addr_reg    <= access_addr;
					access_byte_mask_reg <= access_byte_mask;
					access_tag_lookup_reg <= access_tag_lookup;
					access_tag_insert_reg <= access_tag_insert;
					access_tag_clear_line_reg <= access_tag_clear_line;
					access_tag_clear_all_reg <= access_tag_clear_all;
					access_acc_reg <= access_acc;
					access_array_command_reg <= access_array_command;
					access_dword_reg <= access_dword;
					access_S_reg <= access_S;
					access_is_ifetch_reg <= access_is_ifetch;
					access_is_read_reg <= access_is_read;
					access_mae_reg <= access_mae;
					array_read_dword_reg <= array_read_dword;
				end if;
			end if;
		end if;
	end process;


	-------------------------------------------------------------------------------------
	--  TLB to keep translated VA -> index-in-set translations.
	-------------------------------------------------------------------------------------
        TrivTlb: if VA_INDEX_TLB_SIZE = 0 generate
		va_tlb_match <= '0';
		va_tlb_matched_index_in_set <= (others => '0');
		va_tlb_matched_acc <= (others => '0');
        end generate TrivTlb;

        nonTrivTlb: if VA_INDEX_TLB_SIZE > 0 generate
	  vaTlbBlock: block
	  begin

		-- lookup TLB.  Keep track of VA tag being used for lookup.. we are always lookup-ing!
		va_tlb_lookup_va_tag <= 
			access_addr(address_width-1 downto (log2_number_of_sets + log2_block_size_in_bytes));
		va_tlb_lookup_set_id <= 
			access_addr((log2_number_of_sets + log2_block_size_in_bytes)-1 downto 
							log2_block_size_in_bytes);
		-- always looking up, aren't we?
		va_tlb_lookup <= '1';

		-- lookup index in set.
		va_tlb_lookup_index_in_set <= va_tlb_matched_index_in_set;
		va_tlb_lookup_acc          <= va_tlb_matched_acc;
		
	
		-- insertion into TLB:
		--      On tags lookup, when the lookup is done, the tags block returns 
		--       a set index which will be used in the TLB.
		-- or
		--	On insert..
		va_tlb_insert      <=  tags_done and tags_index_in_set_is_valid;

		va_tlb_insert_va_tag  <= 
			access_addr_reg(address_width-1 downto (log2_number_of_sets + log2_block_size_in_bytes));
		va_tlb_insert_set_id  <= 
			access_addr_reg((log2_number_of_sets + log2_block_size_in_bytes)-1 downto 
									log2_block_size_in_bytes);
		va_tlb_insert_index_in_set <=  tags_index_in_set;
		va_tlb_insert_acc <= tags_acc;

		-- erase from TLB:
		va_tlb_erase <= '1' when (trigger = '1') and 
					((access_tag_clear_line = '1') or (invalidate(0) = '1')) else '0';
		va_tlb_erase_va_tag  <= access_addr(address_width-1 downto (log2_number_of_sets + log2_block_size_in_bytes)) when
					(invalidate(0) = '0') else invalidate_line_address(line_address_width-1 downto log2_number_of_sets);
		va_tlb_erase_set_id  <= access_addr(log2_number_of_sets + log2_block_size_in_bytes-1 downto log2_block_size_in_bytes) when
					(invalidate(0) = '0') else invalidate_line_address(log2_number_of_sets-1 downto 0);

		-- clear TLB
		va_tlb_clear <= '1' when (trigger = '1') and (access_tag_clear_all = '1') else '0';
	
		--
		-- the VA tlb lookup is in the critical path.  Keep the index tlb size=2
		--  (one per cpu thread!).
		--
		vaTlb: VaToIndexInSetTlb
			generic map (number_of_entries => VA_INDEX_TLB_SIZE,
					set_id_width => log2_number_of_sets,
					index_in_set_width => log2_associativity,
					va_tag_width => (line_address_width-log2_number_of_sets)
				    )
			port map (
					lookup_va_tag => va_tlb_lookup_va_tag,
					lookup_set_id => va_tlb_lookup_set_id,

					erase_va_tag => va_tlb_erase_va_tag,
					erase_set_id => va_tlb_erase_set_id,

					insert_va_tag => va_tlb_insert_va_tag,
					insert_set_id => va_tlb_insert_set_id,
					insert_index_in_set => va_tlb_insert_index_in_set,
					insert_acc => va_tlb_insert_acc,

					match => va_tlb_match,
					matched_index_in_set => va_tlb_matched_index_in_set,
					matched_acc => va_tlb_matched_acc,

					insert => va_tlb_insert,
					lookup => va_tlb_lookup,
					erase => va_tlb_erase,
					clear => va_tlb_clear,
					clk => clk,
					reset => reset);	
	   end block vaTlbBlock;
        end generate nonTrivTlb;

	-------------------------------------------------------------------------------------------------------------------------
	--         lookup/insert/clear-line/invalidate/clear-all.
	-------------------------------------------------------------------------------------------------------------------------
        tagsInst: GenericSetAssociativeCacheTagsWithInvalidate
                        generic map (name => "dcache-tags",
                                        log2_number_of_blocks => log2_number_of_blocks, -- 9  
                                        log2_block_size_in_bytes => log2_block_size_in_bytes, -- 6
					log2_associativity => log2_associativity,
                                        address_width => address_width,
                                        log2_data_width_in_bytes => log2_data_width_in_bytes)
			port map (
					trigger => tags_trigger,	
					done => tags_done,	
					init_flag => init_flag,
					access_acc => access_acc,
					access_tag_lookup => access_tag_lookup,
					access_tag_clear_line => access_tag_clear_line,
					access_tag_clear_all => access_tag_clear_all,
					access_tag_insert => access_tag_insert,
					access_tag_addr => access_addr,
					invalidate => invalidate(0),
					invalidate_line_address => invalidate_line_address,
					valid_match => va_tlb_match,
					match_index_in_set => va_tlb_matched_index_in_set,
					lookup_is_valid => tags_lookup_is_valid,
					access_index_in_set_valid => tags_index_in_set_is_valid,
					access_index_in_set => tags_index_in_set, 
					access_acc_out => tags_acc,
					clk => clk, reset => reset);

	-------------------------------------------------------------------------------------------------------------------------
	--         write/read dword or pass-through or nop.
	--		Note: on a miss, the array operation will be skipped..
	-------------------------------------------------------------------------------------------------------------------------
	array_read_dword     <= '1' when (trigger = '1') and 
					(access_array_command = CACHE_ARRAY_READ_DWORD) else '0';
	array_write_dword    <= '1' when (trigger = '1') and 
					(access_array_command = CACHE_ARRAY_WRITE_DWORD) and 
						(access_mae = '0') else '0';


	arrayInst: GenericSetAssociativeCacheArray 
  			generic map (name => "dcache-array",
                                        log2_number_of_blocks => log2_number_of_blocks, -- 9  
                                        log2_block_size_in_bytes => log2_block_size_in_bytes, -- 6
					log2_associativity => log2_associativity,
                                        address_width => address_width,
					log2_data_width_in_bytes => log2_data_width_in_bytes,
					ignore_byte_mask => icache_flag)
			port map (
    					trigger => arrays_trigger,
    					done => arrays_done,
					-- index in set valid
					matched_index_in_set => arrays_matched_index_in_set,
    					access_mae  => access_mae_qualified ,
    					access_array_command  => access_array_command_qualified ,
    					access_byte_mask  => access_byte_mask_qualified,
    					access_array_addr  => access_addr_qualified,
					access_array_write_dword => access_dword_qualified,
    					access_array_read_dword_vector  => access_array_read_dword_vector,
    					bypassed_dword_out  => bypassed_dword_out,
    					clk => clk,
					reset => reset
				);

	  -------------------------------------------------------------------------------------
	  -- select access_dword out of access_array_dword_vector..
	  -------------------------------------------------------------------------------------
	  process(access_array_read_dword_vector, 
			array_read_dword_reg,
			bypassed_dword_out, 
			tags_index_in_set,
			access_addr_reg, 
			access_array_command_reg)
		variable I: integer range 0 to associativity-1;
	  begin
		if(array_read_dword_reg = '1') then
			I := to_integer(unsigned(tags_index_in_set));
			dword_out <= 
				access_array_read_dword_vector(((I+1)*8*data_width_in_bytes)-1 
									downto (I*8*data_width_in_bytes));	
		else 
			dword_out <= bypassed_dword_out;	
		end if;
	  end process;	
	
	  -------------------------------------------------------------------------------------
	  -- permissions OK logic based on tags acc out and hit status.. 
	  --   Note tags_hit is a bit different...
	  -------------------------------------------------------------------------------------
	  is_hit(0) <= tags_lookup_is_valid and access_tag_lookup_reg;
	  permissions_ok(0) <= cpu_permissions_ok;

end Structural;
--
-- Written by Madhav Desai
--
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library AjitCustom;
use AjitCustom.CachePackage.all;


-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

library ahir;
use ahir.BaseComponents.all;
use ahir.Subprograms.all;

use ahir.mem_component_pack.all;
use ahir.Types.all;
use ahir.Utilities.all;

-- implementation of tags in associative memory.
-- will be done using single ported memory.
--
-- Two simultaneous activities may be requested
--    lookup/insert/clear-line/clear-all  AND invalidate-line
--
-- Now clear-line/invalidate will clear all lines in a set.
--    Note: if not, then the clear operation will take two
--          clock cycles which is not really affordable....
-- 
-- On insert, the tags for an entire set are updated
--    by a single write, using either
--       if there is no match in the valid index tlb,
--       then the next free index.
--	    (this corresponds to the first dword fill
--               on a line miss)
--          OR
--       the matched index from the TLB.
--	    (this corresponds to the remaining dword fills
--               on a line miss)
--
-- On lookup, the tags for an entire set are read out
--    from the tag memory, and the match information
--    is muxed out.
--
-- What about allocation of a set entry?   This will
--    be done at insert time..
--
entity GenericSetAssociativeCacheTagsWithInvalidate is -- 
  generic (name: string := "anon";
		log2_number_of_blocks: integer := 9; 
		log2_block_size_in_bytes: integer := 6; 
		address_width: integer := 32;
		log2_associativity: integer := 1;
		log2_data_width_in_bytes: integer := 3);
  port ( -- 
    trigger: in std_logic;
    done   : out std_logic;
    init_flag : in  std_logic;
    access_acc: in std_logic_vector(2 downto 0);
    -- tag commands.
    access_tag_lookup : in  std_logic;
    access_tag_clear_line : in  std_logic;
    access_tag_clear_all : in  std_logic;
    access_tag_insert : in  std_logic;
    --
    access_tag_addr : in  std_logic_vector(address_width-1 downto 0);
    -- invalidation channel for cache coherence and synonym avoidance.
    invalidate: in std_logic;
    invalidate_line_address: in std_logic_vector(((address_width-1) - log2_block_size_in_bytes) downto 0);
    -- valid tlb match info...
    valid_match: in std_logic;
    match_index_in_set: in std_logic_vector(log2_associativity-1 downto 0);
    -- outputs..
    lookup_is_valid : out  std_logic;
    access_index_in_set_valid: out std_logic;
    access_index_in_set: out std_logic_vector(log2_associativity-1 downto 0);
    access_acc_out: out std_logic_vector(2 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity GenericSetAssociativeCacheTagsWithInvalidate;
architecture Behave of GenericSetAssociativeCacheTagsWithInvalidate is -- 
	function isEqualSLV(x: std_logic_vector; y : std_logic_vector) return std_logic is
		variable ret_var : std_logic;
		variable t: std_logic_vector(1 to x'length);
		alias lx: std_logic_vector(1 to x'length) is x;
		alias ly: std_logic_vector(1 to y'length) is y;
	begin
		for I in 1 to x'length loop
			t(I) := not (lx(I) xor ly(I));
		end loop;
		ret_var := AndReduce(t);
		return(ret_var);
	end function;

	function OrReduceSLV(x: std_logic_vector; constant N: integer) return std_logic_vector is
		alias lx: std_logic_vector(x'length-1 downto 0) is x;
		variable tvar: std_logic_vector((x'length/N)-1 downto 0);
		variable result_var : std_logic_vector(N-1 downto 0);
	begin
		for I in 0 to N-1 loop
			for J in 0 to (x'length/N)-1 loop
				tvar(J) := lx(I + (J*N));
			end loop;
			result_var (I) := OrReduce(tvar);
		end loop;
		return result_var;
	end function;
		
	constant number_of_blocks : integer := (2**log2_number_of_blocks);
	constant bytes_per_block : integer := (2**log2_block_size_in_bytes);
	constant data_width_in_bytes : integer := (2**log2_data_width_in_bytes);
	constant dwords_per_block : integer := (2**(log2_block_size_in_bytes - log2_data_width_in_bytes));
	constant log2_dwords_per_block: integer := (log2_block_size_in_bytes - log2_data_width_in_bytes);

	constant associativity: integer := 2**log2_associativity;
	constant number_of_sets   : integer := number_of_blocks/associativity;
	constant log2_number_of_sets: integer := (log2_number_of_blocks - log2_associativity);

	constant line_address_width : integer := (address_width - log2_block_size_in_bytes);

	--  tag width 
	constant tag_width : integer :=  
		address_width - (log2_number_of_sets + log2_block_size_in_bytes);
	--  acc + tag.
	constant tag_mem_data_width : integer :=  tag_width + 3;
	
	--
	--  memory access signals.
	-- 
	type   TagMemDataArray is array (natural range <>) 
					of std_logic_vector(tag_mem_data_width-1 downto 0);

	signal  tag_mem_address :   std_logic_vector(log2_number_of_sets-1 downto 0);
	signal  tag_mem_write_data: TagMemDataArray(associativity-1 downto 0);
	signal  tag_mem_read_data:  TagMemDataArray(associativity-1 downto 0);
	signal  tag_mem_word_mask: std_logic_vector(associativity-1 downto 0);
	signal  tag_mem_enable:     std_logic;
	signal  tag_mem_read_write_bar:  std_logic;
	
    	signal access_lookup_acc_out: std_logic_vector(2 downto 0);
    	signal access_insert_acc_out: std_logic_vector(2 downto 0);
	--
	-- valid bits.. 
	-- 
	type   ValidBitArray is array (natural  range <>) of std_logic_vector(associativity-1 downto 0);
	signal valid_bits: ValidBitArray(number_of_sets-1 downto 0);

	type   LastWrittenIndexArray is array (natural  range <>) of std_logic_vector(log2_associativity-1 downto 0);
	signal most_recently_used_indices: LastWrittenIndexArray(number_of_sets-1 downto 0);

	-- No need for states... all operations complete in one cycle.
	signal valid_bit_registered : std_logic;

    	signal valid_match_reg: std_logic;
    	signal match_index_in_set_reg: std_logic_vector(log2_associativity-1 downto 0);
	
	signal lookup_valid_sig: std_logic;

    	signal access_acc_reg: std_logic_vector(2 downto 0);
    	signal access_tag_addr_reg : std_logic_vector(address_width-1 downto 0);

    	signal invalidate_reg: std_logic;
    	signal invalidate_line_address_reg: std_logic_vector(line_address_width-1 downto 0);
    

		
	function virtualAddressTag(va: std_logic_vector(address_width-1 downto 0)) 
		return std_logic_vector is
		variable ret_var : std_logic_vector(tag_width-1 downto 0);
	begin
		ret_var := va(address_width-1 downto (log2_number_of_sets  + log2_block_size_in_bytes));
		return(ret_var);
	end function virtualAddressTag;

	function setId (x: std_logic_vector(line_address_width-1 downto 0)) 
		return integer is
		variable ret_var : integer range 0 to number_of_sets -1;
		variable set_id_var : std_logic_vector(log2_number_of_sets-1 downto 0);
	begin
		set_id_var := x(log2_number_of_sets -1 downto 0);
		ret_var := to_integer(unsigned(set_id_var));
		return(ret_var);
	end setId;

	function computeNextValidBits (vbits: ValidBitArray;
					insert, clear_line, clear_all: std_logic;
					insert_line_addr, clear_line_addr: 
						std_logic_vector(line_address_width-1 downto 0);
					insert_index_in_set: integer range 0 to associativity-1)
	return ValidBitArray is
		variable ret_var : ValidBitArray(number_of_sets-1 downto 0);
		variable bit_val: std_logic;
		variable set_id : integer range 0 to number_of_sets-1;
		variable ins_bit: boolean;
	begin
		ret_var := vbits;
		bit_val := '0';
		ins_bit := false;
		set_id  := 0;

		if(clear_all = '1') then
			ret_var := (others => (others => '0'));
		elsif (clear_line = '1') then
			set_id := setId(clear_line_addr);	
			ins_bit := true;
		elsif (insert = '1') then
			set_id := setId(insert_line_addr);	
			ins_bit := true;
			bit_val := '1';
		end if;
	
		if(ins_bit) then
			if(clear_line = '1') then
				-- on clear line, we just clear the whole set.
				-- and there is no need to worry about matches.
				ret_var(set_id) := (others => '0');
			elsif (insert = '1') then
				ret_var(set_id)(insert_index_in_set) := '1';
			end if;
		end if;

		return(ret_var);
	end computeNextValidBits;

	function findNextFreeIndex(pre_val: integer range 0 to associativity-1;
					set_valids: std_logic_vector(associativity-1 downto 0))
	return integer is
		variable ret_var: integer range 0 to associativity-1;
	begin
		ret_var := pre_val;
		for I in 1 to associativity -1 loop
			if ret_var = associativity-1 then
				ret_var := 0;
			else
				ret_var := (ret_var + 1);
			end if;

			if(set_valids(ret_var) = '0') then
				exit;
			end if;
		end loop;

		return(ret_var);
	end findNextFreeIndex;
				
	procedure updateNextMostRecentlyUsedIndices
			(lwi: in LastWrittenIndexArray(number_of_sets-1 downto 0);
						set_id: in integer range 0 to number_of_sets-1;
						set_valids: in std_logic_vector(associativity-1 downto 0);
						vmatch: in std_logic;
						mindex: in std_logic_vector(log2_associativity-1 downto 0);
						insert: in std_logic;
						lookup: in std_logic;
						next_lwi: out LastWrittenIndexArray(number_of_sets-1 downto 0);
						most_recently_used_index : out integer range 0 to associativity-1
			) is
		variable curr_val, next_free_val: integer range 0 to associativity-1;
	begin
		-- return the index into which a new entry has to be created.
		-- Also, update the next free index for this set.
		next_lwi := lwi;
		curr_val := to_integer(unsigned(lwi(set_id)));

		next_free_val := curr_val;

		if (vmatch = '1') and ((lookup = '1') or (insert = '1')) then 


			-- move the free pointer to point to something other than mindex!
			next_free_val := findNextFreeIndex(to_integer(unsigned(mindex)), set_valids);
			
			-- the index which will be used by insert...
			curr_val   := to_integer(unsigned(mindex));

		elsif (insert = '1') then 
			-- if not, and if it is an insert, the free slot is incremented..
			if(curr_val < associativity-1) then
				next_free_val := (curr_val + 1);
			else
				next_free_val := 0;
			end if;
		end if;
			
		next_lwi(set_id) := std_logic_vector(to_unsigned(next_free_val, log2_associativity));

		-- this is OK.
		most_recently_used_index := curr_val;
	end updateNextMostRecentlyUsedIndices;
				    
	function incrementIndex (X: integer range 0 to associativity-1) return integer is
		variable ret_var:integer range 0 to associativity-1;
	begin
		ret_var := 0;
		if(X < associativity-1) then
			ret_var := (X + 1);
		end if;
		return(ret_var);	
	end incrementIndex;

				

      
-- see comment above..
--##decl_synopsys_sync_set_reset##

	signal active_lookup_index_in_set, active_insert_index_in_set_reg: 
					std_logic_vector(log2_associativity-1 downto 0);
	signal active_set_id_reg: integer range 0 to number_of_sets-1;
       		
	signal lookup, insert, clear_all, clear_line: std_logic;
	signal lookup_reg, insert_reg, clear_all_reg, clear_line_reg: std_logic;
begin --  
	

	insert <= '1' when (trigger = '1') and (access_tag_insert = '1') else '0';
	lookup <= '1' when (trigger = '1') and (access_tag_lookup = '1') else '0';
	clear_line <= '1' when (trigger = '1') and ((access_tag_clear_line = '1') or (invalidate = '1'))  else '0';
	clear_all  <= '1' when (trigger = '1') and (access_tag_clear_all = '1') else '0';

	----------------------------------------------------------------------------------
	-- register the inputs... etc.
	----------------------------------------------------------------------------------
	process(clk, trigger, reset) 
	begin
		if(clk'event and (clk = '1')) then
			if reset = '1' then
				done <= '0';
			else
				done <= trigger;
				if trigger = '1' then
    					access_acc_reg <= access_acc;
    					access_tag_addr_reg <= access_tag_addr;
    					invalidate_reg <= invalidate;
    					invalidate_line_address_reg <= invalidate_line_address;

					lookup_reg <= lookup;
					insert_reg <= insert;
					clear_line_reg <= clear_line;
					clear_all_reg <= clear_all;

					valid_match_reg <= valid_match;
					match_index_in_set_reg <= match_index_in_set;
				end if;
			end if;
		end if;
	end process;


	----------------------------------------------------------------------------------
	-- tag memory control process.
	----------------------------------------------------------------------------------
	tagMemCtrl: block
	begin
		
		process(clk, reset, 
				trigger, 
				lookup, 
				insert, 
				clear_all, 
				clear_line, 
				valid_match,
				valid_bits,
				match_index_in_set,
				most_recently_used_indices,
				access_tag_addr, 
				invalidate_line_address)
			variable next_valid_bits_var: ValidBitArray(number_of_sets-1 downto 0);
			variable next_most_recently_used_indices_var: LastWrittenIndexArray(number_of_sets-1 downto 0);
			variable access_tag_line_address_var, clear_line_address_var : std_logic_vector(line_address_width-1 downto 0);
			variable tag_mem_write_data_var: TagMemDataArray(associativity-1 downto 0);
			variable tag_mem_address_var :   std_logic_vector(log2_number_of_sets-1 downto 0);
			variable tag_mem_word_mask_var: std_logic_vector(associativity-1 downto 0);
			variable active_set_id_var: integer range 0 to number_of_sets-1;
			variable active_set_valids_var: std_logic_vector(associativity-1 downto 0);
			variable active_tag_var: std_logic_vector(tag_width-1 downto 0);
			variable most_recently_used_index_var: integer range 0 to associativity-1;
		begin
			tag_mem_word_mask_var := (others => '0');
			tag_mem_write_data_var := (others => (others => '0'));
			tag_mem_address_var := (others => '0');

			access_tag_line_address_var := access_tag_addr(address_width-1 downto log2_block_size_in_bytes);
			active_set_id_var := setId(access_tag_line_address_var);
			active_set_valids_var := valid_bits(active_set_id_var);

			active_tag_var := (others => '0');
			

			if(invalidate = '1') then 
				clear_line_address_var := invalidate_line_address;
			else
				clear_line_address_var := access_tag_addr(address_width-1 downto log2_block_size_in_bytes);
			end if;

			--
			-- update last written indices on insert (rotate to the right).
			--
			updateNextMostRecentlyUsedIndices(most_recently_used_indices,
								active_set_id_var,
								active_set_valids_var,
								valid_match,
								match_index_in_set,
								insert,
								lookup,
								next_most_recently_used_indices_var,
								most_recently_used_index_var
							  );
				
			next_valid_bits_var := computeNextValidBits (valid_bits,
									insert, 
									clear_line, 
									clear_all,
									access_tag_line_address_var, 
									clear_line_address_var,
									most_recently_used_index_var);
									
				
			tag_mem_address_var := access_tag_line_address_var(log2_number_of_sets-1 downto 0);
			active_tag_var := access_tag_line_address_var(line_address_width - 1 downto  log2_number_of_sets);
				

			-- tag mem is addressed by the set-id.
			if (insert  = '1') then
			    	tag_mem_word_mask_var(most_recently_used_index_var) := '1';	
				    -- write acc + tag into the specified index within the set.
				tag_mem_write_data_var(most_recently_used_index_var) :=  access_acc & active_tag_var;
			else
				tag_mem_word_mask_var := (others => '1');
			end if;

			tag_mem_address <= tag_mem_address_var;
			tag_mem_word_mask <= tag_mem_word_mask_var;
			tag_mem_write_data <= tag_mem_write_data_var;
			tag_mem_read_write_bar <= not insert;
			tag_mem_enable <= lookup or insert;

			if (clk'event and (clk = '1')) then
				if(reset = '1') then
					valid_bits <= (others => (others => '0'));
					most_recently_used_indices <= (others => (others => '0'));
				else
					valid_bits <= next_valid_bits_var;
					most_recently_used_indices <= next_most_recently_used_indices_var;

					if(lookup = '1') or (insert = '1') then
						active_set_id_reg <= active_set_id_var;
					end if;

					if(insert = '1') then
						active_insert_index_in_set_reg <= 
							std_logic_vector(to_unsigned(most_recently_used_index_var, log2_associativity));
					end if;
				end if;
			end if;
		end process;
	end block tagMemCtrl;

	------------------------------------------------------------------------------------------------
	--  Tag memory.
	------------------------------------------------------------------------------------------------
	bGen: for A in associativity-1 downto 0 generate
          tblk: block
              signal enable_sig: std_logic;
          begin
		enable_sig <= tag_mem_enable and tag_mem_word_mask(A);
		tagInst: base_bank
			generic map		
				(name => "dcache_tag_memory_" & Convert_To_String(A),
						g_addr_width => log2_number_of_sets,
						g_data_width => tag_mem_data_width)
			port map (
					datain => tag_mem_write_data(A),
					dataout => tag_mem_read_data(A),
					addrin => tag_mem_address, 
					enable => enable_sig,
					writebar => tag_mem_read_write_bar,
					clk => clk, reset => reset
			);	
           end block tblk;
	end generate bGen;

		

	------------------------------------------------------------------------------------------------
	--  output logic
	------------------------------------------------------------------------------------------------

	-- Some selection logic... needs to be fast
	matchBlock: block
		signal set_valids: std_logic_vector(associativity-1 downto 0);
		signal lookup_acc_aggregate: std_logic_vector((associativity*3)-1 downto 0);
		signal active_lookup_index_aggregate: std_logic_vector((associativity*log2_associativity)-1 downto 0);
		signal lookup_valid_aggregate: std_logic_vector(associativity-1 downto 0);
	begin
		set_valids <= valid_bits(active_set_id_reg);

		genPar: for T in associativity-1 downto 0 generate
			mb: block
				signal match_sig: std_logic;
				signal Zero3: std_logic_vector(2 downto 0);
				signal ZeroA: std_logic_vector(log2_associativity-1 downto 0);
			begin

				Zero3 <= (others => '0');
				ZeroA <= (others => '0');

				match_sig <= '1' when
						(set_valids(T) = '1') and 
						(isEqualSLV(tag_mem_read_data(T)(tag_width-1 downto 0), virtualAddressTag(access_tag_addr_reg)) = '1') and
						(lookup_reg = '1') else '0';
				lookup_valid_aggregate(T) <= match_sig;
				active_lookup_index_aggregate(((T+1)*log2_associativity)-1 downto (T*log2_associativity)) 
						<= std_logic_vector(to_unsigned(T, log2_associativity)) when match_sig  = '1' else ZeroA;
				lookup_acc_aggregate(((T+1)*3)-1 downto (T*3)) 
						<= tag_mem_read_data(T)(tag_mem_data_width-1 downto tag_width) when match_sig = '1'  else Zero3;
			end block mb;
		end generate genPar;

		lookup_valid_sig <= OrReduce(lookup_valid_aggregate);
		access_lookup_acc_out <= OrReduceSLV (lookup_acc_aggregate, 3);
		active_lookup_index_in_set <= OrReduceSLV (active_lookup_index_aggregate, log2_associativity);

	end block matchBlock;

	lookup_is_valid <= lookup_valid_sig;
	process(lookup, active_lookup_index_in_set, 
			lookup_valid_sig, valid_match_reg, match_index_in_set_reg)
	begin
		if(clk'event and clk='1') then 
		   if(lookup_reg = '1') and (lookup_valid_sig = '1') and (valid_match_reg = '1') then
			-- set entry must be valid if vmatch is indicated.
			assert (to_integer(unsigned(active_lookup_index_in_set))) = 
					(to_integer(unsigned(match_index_in_set_reg)))
				report "LOOKUP MISMATCH BETWEEN TLB AND SET!" severity FAILURE;
		   end if;
		end if;
	end process;

	-- index information.
	access_index_in_set_valid <= ((lookup_reg and lookup_valid_sig) or insert_reg);
	access_index_in_set <= active_lookup_index_in_set when (lookup_reg = '1') 
						else active_insert_index_in_set_reg when (insert_reg = '1') else (others => '0');
	access_acc_out <= access_lookup_acc_out when (lookup_reg = '1')
				else access_acc_reg when (insert_reg = '1') else (others => '0');

end Behave;
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;

entity VaToIndexInSetTlb is
	generic (number_of_entries: integer := 4; 
			set_id_width: integer := 8;
			index_in_set_width: integer := 1;
			va_tag_width: integer := 25   -- Va tag.
		);
	port (
		lookup_va_tag:    in std_logic_vector(va_tag_width-1 downto 0);
		lookup_set_id: 	  in std_logic_vector(set_id_width-1 downto 0);

		erase_va_tag: in std_logic_vector(va_tag_width-1 downto 0);
		erase_set_id: in std_logic_vector(set_id_width-1 downto 0);

		insert_va_tag: in std_logic_vector(va_tag_width-1 downto 0);
		insert_set_id: in std_logic_vector(set_id_width-1 downto 0);
		insert_index_in_set: in std_logic_vector(index_in_set_width-1 downto 0);
		insert_acc   : in std_logic_vector(2 downto 0);

		match: out std_logic;
		matched_index_in_set: out std_logic_vector(index_in_set_width-1 downto 0);
		matched_acc: 	  out std_logic_vector(2 downto 0);

		insert: in std_logic;
		lookup: in std_logic;
		erase : in std_logic;
		clear : in std_logic;
		clk, reset:  in std_logic
	);
end entity;

architecture Behavioural of VaToIndexInSetTlb is

	constant entry_width: integer := va_tag_width + set_id_width + index_in_set_width + 3;

	--
	-- each entry has the following fields.
	--      va_tag set_id index_in_set
	--
	-- On lookup, given up the lookup tag and set-id, return match if it exists.
	-- 
	-- On insert, create new entry, and also invalidate entries which 
	--   have the same set-id and index-in-set.
	--
	-- On erase, remove entry which matches tags.
	--
	-- 
	type TlbArray is array (natural range <>) of std_logic_vector(entry_width-1  downto 0);
	signal tlb_entries: TlbArray (number_of_entries-1 downto 0);
	signal valids: std_logic_vector(number_of_entries-1 downto 0);
	signal last_inserted_pointer, matched_insert_pointer: integer range 0 to number_of_entries-1;
	signal match_sig: std_logic;
	signal insert_match_sig:  boolean;
	signal erase_match_index_sig : integer range 0 to number_of_entries-1;

	function IncrementPointer(x: integer) return integer is
		variable ret_val: integer range 0 to number_of_entries-1;
	begin
		if(x = number_of_entries-1) then
			ret_val := 0;
		else
			ret_val := x + 1;
		end if;

		return(ret_val);
	end function;

		
	signal erase_match_indices : std_logic_vector(number_of_entries-1 downto 0);
begin
	-- match process
	process(tlb_entries, valids, lookup_va_tag, lookup_set_id, 
				insert_va_tag, insert_set_id, insert_index_in_set, insert_acc,
				erase_va_tag, insert, lookup, erase)
		variable match_var: std_logic;
		variable tlb_entry    : std_logic_vector(entry_width-1 downto 0);

		variable entry_va_tag    : std_logic_vector(va_tag_width-1 downto 0);
		variable entry_set_id: std_logic_vector(set_id_width-1 downto 0);
		variable entry_index_in_set: std_logic_vector(index_in_set_width-1 downto 0);
		variable entry_acc   : std_logic_vector(2 downto 0);

		variable insert_match, lookup_match, erase_match: boolean;
		variable erase_match_indices_var : std_logic_vector(number_of_entries-1 downto 0);
		variable matched_acc_var : std_logic_vector(2 downto 0);
		variable valid_var: std_logic;
		variable matched_index_in_set_var: std_logic_vector(index_in_set_width-1 downto 0);
		variable matched_insert_pointer_var: integer range 0 to number_of_entries-1;
	begin

		match_var := '0';

		insert_match := false;
		erase_match  := false;
		erase_match_indices_var := (others => '0');
		matched_acc_var := (others => '0');
		matched_index_in_set_var := (others => '0');
		matched_insert_pointer_var := 0;
		
		for I in 0 to number_of_entries-1 loop

			valid_var := valids(I);

			tlb_entry 	:= tlb_entries(I);

			entry_acc    := tlb_entry (2 downto 0);
			entry_index_in_set := tlb_entry (2+index_in_set_width downto 3);
			entry_set_id := tlb_entry (2+index_in_set_width+set_id_width downto 3+index_in_set_width);
			entry_va_tag    :=  tlb_entry(entry_width-1 downto 3+index_in_set_width+set_id_width);

			-- insert match
			if ((insert = '1') and (entry_va_tag = insert_va_tag) and 
						(entry_set_id = insert_set_id) and 
						(valid_var = '1')) then

				assert insert_match = false
					report "MULTIPLE INSERT MATCHES IN VA TLB." severity FAILURE;

				insert_match := true;
				matched_insert_pointer_var := I;
			end if;

			--
			-- erase if  
			--       erase = 1 and erase-setid matches 
			--		erase is applied to the entire set...
			--
			--       or  insert = 1 and not insert match and setid+indexinsetid matches.
			--
			erase_match     := 
				((erase = '1')  and  (valid_var = '1') and (entry_set_id = erase_set_id))
					 or
				-- if insert matches entries set and index ids... then the entry should be erased..
				   ((insert = '1') and (valid_var = '1') and
					(entry_set_id = insert_set_id) and (entry_index_in_set = insert_index_in_set));

			-- erase match? ....
			if erase_match then
				erase_match_indices_var(I) := '1';
			end if;

			-- lookup match if entry matches set and tag..
			lookup_match    :=  
					(lookup = '1') and (valid_var = '1') and 
						(entry_va_tag = lookup_va_tag) and (entry_set_id = lookup_set_id);
			if(lookup_match) then
				
				assert match_var = '0'
					report "MULTIPLE LOOKUP MATCHES IN VA TLB." severity FAILURE;

				match_var := '1';
				matched_acc_var := tlb_entry (2 downto 0);
				matched_index_in_set_var := tlb_entry (index_in_set_width+2 downto 3);
			end if;
		end loop;

		insert_match_sig <= insert_match;
		erase_match_indices <= erase_match_indices_var;

		match <= match_var;
		matched_index_in_set <= matched_index_in_set_var;

		matched_insert_pointer <= matched_insert_pointer_var;
		matched_acc <= matched_acc_var;

	end process;

	-- management process
	process(clk, reset, 
			valids, 
			insert_va_tag, insert_set_id, insert_index_in_set, insert_acc, insert_match_sig,
			erase_match_indices, 
			last_inserted_pointer,
			matched_insert_pointer,
			tlb_entries) 
		variable insert_pointer_var : integer range 0 to number_of_entries-1;
		variable next_valids_var: std_logic_vector(number_of_entries-1 downto 0);
	begin
		next_valids_var := valids;

		if(insert_match_sig) then
			insert_pointer_var := matched_insert_pointer;
		else
			insert_pointer_var := IncrementPointer (last_inserted_pointer);
		end if;


		for I in 0 to number_of_entries-1 loop
			if(erase_match_indices(I) = '1') then
				next_valids_var(I) := '0';
			end if;
		end loop;
				
		if  (insert = '1')  then
			next_valids_var(insert_pointer_var) := '1';
		end if;

		if(clk'event and clk = '1') then
			if((reset = '1') or (clear = '1')) then
				valids <= (others => '0');
				last_inserted_pointer <= 0;
			else
				valids <= next_valids_var;

				if  (insert = '1')  then
					tlb_entries(insert_pointer_var) <= 
						insert_va_tag & insert_set_id & insert_index_in_set & insert_acc;
					last_inserted_pointer <= insert_pointer_var;
				end if;
			end if;
		end if;
	end process;

end Behavioural;

library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library AjitCustom;
use AjitCustom.AjitGlobalConfigurationPackage.all;
use AjitCustom.AjitCustomComponents.all;

entity accessTlbMemory_0_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    clear_flag : in  std_logic_vector(0 downto 0);
    wr_flag : in  std_logic_vector(0 downto 0);
    write_address : in  std_logic_vector(0 downto 0);
    write_entry : in  std_logic_vector(46 downto 0);
    lookup_address : in  std_logic_vector(0 downto 0);
    l0_v : out  std_logic_vector(0 downto 0);
    lookup_entry : out  std_logic_vector(46 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity accessTlbMemory_0_Operator;

architecture SimpleTon of  accessTlbMemory_0_Operator is -- 
begin
	bmem: accessTlbMemoryBase_Operator 
		generic map (address_width => mmu_log_tlb_level_0_entries, data_width => 47, use_mem_cuts => false)
		port map (
    			sample_req => sample_req,
    			sample_ack => sample_ack,
    			update_req => update_req,
    			update_ack => update_ack,
    			clear_flag  => clear_flag ,
    			wr_flag  => wr_flag ,
    			write_address  => write_address ,
    			write_entry  => write_entry ,
    			lookup_address  => lookup_address ,
    			l_v  => l0_v ,
    			lookup_entry  => lookup_entry ,
    			clk  => clk,
			reset => reset);

end architecture SimpleTon;

library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library AjitCustom;
use AjitCustom.AjitGlobalConfigurationPackage.all;
use AjitCustom.AjitCustomComponents.all;

entity accessTlbMemory_1_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    clear_flag : in  std_logic_vector(0 downto 0);
    wr_flag : in  std_logic_vector(0 downto 0);
    write_address : in  std_logic_vector(1 downto 0);
    write_entry : in  std_logic_vector(45 downto 0);
    lookup_address : in  std_logic_vector(1 downto 0);
    l1_v : out  std_logic_vector(0 downto 0);
    lookup_entry : out  std_logic_vector(45 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity accessTlbMemory_1_Operator;


architecture SimpleTon of  accessTlbMemory_1_Operator is -- 
begin
	bmem: accessTlbMemoryBase_Operator 
		generic map (address_width => mmu_log_tlb_level_1_entries, data_width => 46, use_mem_cuts => false)
		port map (
    			sample_req => sample_req,
    			sample_ack => sample_ack,
    			update_req => update_req,
    			update_ack => update_ack,
    			clear_flag  => clear_flag ,
    			wr_flag  => wr_flag ,
    			write_address  => write_address ,
    			write_entry  => write_entry ,
    			lookup_address  => lookup_address ,
    			l_v  => l1_v ,
    			lookup_entry  => lookup_entry ,
    			clk  => clk,
			reset => reset);

end architecture SimpleTon;


library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library AjitCustom;
use AjitCustom.AjitGlobalConfigurationPackage.all;
use AjitCustom.AjitCustomComponents.all;

entity accessTlbMemory_2_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    clear_flag : in  std_logic_vector(0 downto 0);
    wr_flag : in  std_logic_vector(0 downto 0);
    write_address : in  std_logic_vector(3 downto 0);
    write_entry : in  std_logic_vector(49 downto 0);
    lookup_address : in  std_logic_vector(3 downto 0);
    l2_v : out  std_logic_vector(0 downto 0);
    lookup_entry : out  std_logic_vector(49 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity accessTlbMemory_2_Operator;


architecture SimpleTon of  accessTlbMemory_2_Operator is -- 
begin
	bmem: accessTlbMemoryBase_Operator 
		generic map (address_width => mmu_log_tlb_level_2_entries, data_width => 50)
		port map (
    			sample_req => sample_req,
    			sample_ack => sample_ack,
    			update_req => update_req,
    			update_ack => update_ack,
    			clear_flag  => clear_flag ,
    			wr_flag  => wr_flag ,
    			write_address  => write_address ,
    			write_entry  => write_entry ,
    			lookup_address  => lookup_address ,
    			l_v  => l2_v ,
    			lookup_entry  => lookup_entry ,
    			clk  => clk,
			reset => reset);

end architecture SimpleTon;



library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library AjitCustom;
use AjitCustom.AjitGlobalConfigurationPackage.all;
use AjitCustom.AjitCustomComponents.all;

entity accessTlbMemory_3_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    clear_flag : in  std_logic_vector(0 downto 0);
    wr_flag : in  std_logic_vector(0 downto 0);
    write_address : in  std_logic_vector(5 downto 0);
    write_entry : in  std_logic_vector(53 downto 0);
    lookup_address : in  std_logic_vector(5 downto 0);
    l3_v : out  std_logic_vector(0 downto 0);
    lookup_entry : out  std_logic_vector(53 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity accessTlbMemory_3_Operator;


architecture SimpleTon of  accessTlbMemory_3_Operator is -- 
begin
	bmem: accessTlbMemoryBase_Operator 
		generic map (address_width =>  mmu_log_tlb_level_3_entries, data_width => 54)
		port map (
    			sample_req => sample_req,
    			sample_ack => sample_ack,
    			update_req => update_req,
    			update_ack => update_ack,
    			clear_flag  => clear_flag ,
    			wr_flag  => wr_flag ,
    			write_address  => write_address ,
    			write_entry  => write_entry ,
    			lookup_address  => lookup_address ,
    			l_v  => l3_v ,
    			lookup_entry  => lookup_entry ,
    			clk  => clk,
			reset => reset);

end architecture SimpleTon;

library std;
use std.standard.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library AjitCustom;
use AjitCustom.AjitGlobalConfigurationPackage.all;
use AjitCustom.AjitCustomComponents.all;


entity accessTlbNewMemory_0_Operator is
  port ( -- 
    	sample_req: in boolean;
    	sample_ack: out boolean;
    	update_req: in boolean;
    	update_ack: out boolean;
	clear: in std_logic_vector(0 downto 0);
	write: in std_logic_vector(0 downto 0);
        write_tag:  in std_logic_vector(7 downto 0);
        write_data: in std_logic_vector(31 downto 0);
        lookup: in std_logic_vector(0 downto 0);
	lookup_tag: in std_logic_vector(7 downto 0);
        tlb_hit: out std_logic_vector(0 downto 0);
	pte: out std_logic_vector(31 downto 0);
        clk, reset: in std_logic);
end entity;


architecture Wrapper of accessTlbNewMemory_0_Operator is
	signal zero_sig: std_logic_vector(0 downto 0);
begin
	zero_sig(0)  <= '0';
	basemem:genericFullyAssociativeMemory_Operator
			generic map(tag_width => 8,
					data_width => 32,
					log_number_of_entries => mmu_log_tlb_new_0_mem_size,
					ignore_collisions => false,
					use_mem_cuts => false)
			port map(
					sample_req => sample_req,
					sample_ack => sample_ack,
					update_req => update_req,
					update_ack => update_ack,
					clear_flag => clear,
					erase_flag => zero_sig,
					write_flag => write,
					write_data => write_data,
					write_tag => write_tag,
					lookup_flag => lookup,
					lookup_tag => lookup_tag,
					lookup_valid => tlb_hit,
					lookup_data => pte,
					clk => clk, reset => reset);
end Wrapper;

library std;
use std.standard.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library AjitCustom;
use AjitCustom.AjitGlobalConfigurationPackage.all;
use AjitCustom.AjitCustomComponents.all;


entity accessTlbNewMemory_1_Operator is
  port ( -- 
    	sample_req: in boolean;
    	sample_ack: out boolean;
    	update_req: in boolean;
    	update_ack: out boolean;
	clear: in std_logic_vector(0 downto 0);
	write: in std_logic_vector(0 downto 0);
        write_tag:  in std_logic_vector(15 downto 0);
        write_data: in std_logic_vector(31 downto 0);
        lookup: in std_logic_vector(0 downto 0);
	lookup_tag: in std_logic_vector(15 downto 0);
        tlb_hit: out std_logic_vector(0 downto 0);
	pte: out std_logic_vector(31 downto 0);
        clk, reset: in std_logic);
end entity;


architecture Wrapper of accessTlbNewMemory_1_Operator is
	signal zero_sig: std_logic_vector(0 downto 0);
begin
	zero_sig(0)  <= '0';
	basemem:genericFullyAssociativeMemory_Operator
			generic map(tag_width => 16,
					data_width => 32,
					log_number_of_entries => mmu_log_tlb_new_1_mem_size,
					ignore_collisions => false,
					use_mem_cuts => false)
			port map(
					sample_req => sample_req,
					sample_ack => sample_ack,
					update_req => update_req,
					update_ack => update_ack,
					clear_flag => clear,
					erase_flag => zero_sig,
					write_flag => write,
					write_data => write_data,
					write_tag => write_tag,
					lookup_flag => lookup,
					lookup_tag => lookup_tag,
					lookup_valid => tlb_hit,
					lookup_data => pte,
					clk => clk, reset => reset);
end Wrapper;

library std;
use std.standard.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library AjitCustom;
use AjitCustom.AjitGlobalConfigurationPackage.all;
use AjitCustom.AjitCustomComponents.all;


entity accessTlbNewMemory_2_Operator is
  port ( -- 
    	sample_req: in boolean;
    	sample_ack: out boolean;
    	update_req: in boolean;
    	update_ack: out boolean;
	clear: in std_logic_vector(0 downto 0);
	write: in std_logic_vector(0 downto 0);
        write_tag:  in std_logic_vector(21 downto 0);
        write_data: in std_logic_vector(31 downto 0);
        lookup: in std_logic_vector(0 downto 0);
	lookup_tag: in std_logic_vector(21 downto 0);
        tlb_hit: out std_logic_vector(0 downto 0);
	pte: out std_logic_vector(31 downto 0);
        clk, reset: in std_logic);
end entity;


architecture Wrapper of accessTlbNewMemory_2_Operator is
	signal zero_sig: std_logic_vector(0 downto 0);
begin
	zero_sig(0)  <= '0';
	basemem:genericFullyAssociativeMemory_Operator
			generic map(tag_width => 22,
					data_width => 32,
					log_number_of_entries => mmu_log_tlb_new_2_mem_size,
					ignore_collisions => false,
					use_mem_cuts => false)
			port map(
					sample_req => sample_req,
					sample_ack => sample_ack,
					update_req => update_req,
					update_ack => update_ack,
					clear_flag => clear,
					erase_flag => zero_sig,
					write_flag => write,
					write_data => write_data,
					write_tag => write_tag,
					lookup_flag => lookup,
					lookup_tag => lookup_tag,
					lookup_valid => tlb_hit,
					lookup_data => pte,
					clk => clk, reset => reset);
end Wrapper;

library std;
use std.standard.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library AjitCustom;
use AjitCustom.AjitGlobalConfigurationPackage.all;
use AjitCustom.AjitCustomComponents.all;


entity accessTlbNewMemory_3_Operator is
  port ( -- 
    	sample_req: in boolean;
    	sample_ack: out boolean;
    	update_req: in boolean;
    	update_ack: out boolean;
	clear: in std_logic_vector(0 downto 0);
	write: in std_logic_vector(0 downto 0);
        write_tag:  in std_logic_vector(27 downto 0);
        write_data: in std_logic_vector(31 downto 0);
        lookup: in std_logic_vector(0 downto 0);
	lookup_tag: in std_logic_vector(27 downto 0);
        tlb_hit: out std_logic_vector(0 downto 0);
	pte: out std_logic_vector(31 downto 0);
        clk, reset: in std_logic);
end entity;


architecture Wrapper of accessTlbNewMemory_3_Operator is
	signal zero_sig: std_logic_vector(0 downto 0);
begin
	zero_sig(0)  <= '0';
	basemem:genericSetAssociativeMemory_Operator
			generic map(tag_width => 28-mmu_log_tlb_new_3_number_of_sets,
					data_width => 32,
					log_number_of_entries => mmu_log_tlb_new_3_mem_size,
					log_associativity     => mmu_log_tlb_new_3_set_size,
					ignore_collisions => false,
					use_mem_cuts => true)
			port map(
					sample_req => sample_req,
					sample_ack => sample_ack,
					update_req => update_req,
					update_ack => update_ack,
					clear_flag => clear,
					erase_flag => zero_sig,
					write_flag => write,
					write_data => write_data,
					write_tag => write_tag(27 downto mmu_log_tlb_new_3_number_of_sets),
					write_set_id => write_tag(mmu_log_tlb_new_3_number_of_sets-1 downto 0),
					lookup_flag => lookup,
					lookup_tag => lookup_tag(27 downto mmu_log_tlb_new_3_number_of_sets),
					lookup_set_id => lookup_tag(mmu_log_tlb_new_3_number_of_sets-1 downto 0),
					lookup_valid => tlb_hit,
					lookup_data => pte,
					clk => clk, reset => reset);
end Wrapper;

library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;

entity accessTlbMemoryBase_Operator is -- 
  generic (address_width : integer := 8; data_width : integer := 32; use_mem_cuts: boolean := true);
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    clear_flag : in  std_logic_vector(0 downto 0);
    wr_flag : in  std_logic_vector(0 downto 0);
    write_address : in  std_logic_vector(address_width-1 downto 0);
    write_entry : in  std_logic_vector(data_width-1 downto 0);
    lookup_address : in  std_logic_vector(address_width-1 downto 0);
    l_v : out  std_logic_vector(0 downto 0);
    lookup_entry : out  std_logic_vector(data_width-1 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity accessTlbMemoryBase_Operator;


architecture Mixed of accessTlbMemoryBase_Operator is

	signal start_req, start_ack: std_logic;

	signal ureg_write_data: std_logic_vector(data_width downto 0);
	signal ureg_write_entry: std_logic_vector(data_width-1 downto 0);
	signal ureg_write_valid: std_logic_vector(0 downto 0);
	signal ureg_write_req, ureg_write_ack: std_logic;

	signal ureg_read_data: std_logic_vector(data_width downto 0);
	signal ureg_unload_req, ureg_unload_ack: Boolean;

	
begin

   p2l: Sample_Pulse_To_Level_Translate_Entity
                generic map(name => "accessTlbMemoryBase-Operator-p2l")
                port map (rL => sample_req, rR => start_req,
                                aL => sample_ack, aR => start_ack,
                                        clk => clk, reset => reset);

   ureg: UnloadRegister 
		generic map (name => "genericAccessTlbMemoryBase_Operator:ureg",
				data_width => data_width + 1,
				  bypass_flag => true, nonblocking_read_flag => false)
		port map (write_data => ureg_write_data,
				write_req => ureg_write_req,
					write_ack => ureg_write_ack,
					    read_data => ureg_read_data,
						unload_req => ureg_unload_req,
						   unload_ack => ureg_unload_ack,
							clk => clk,
							  reset => reset);

   ureg_write_data <= ureg_write_valid & ureg_write_entry;
   ureg_unload_req <= update_req;
   update_ack <= ureg_unload_ack;


   l_v(0) <= ureg_read_data(data_width);
   lookup_entry <= ureg_read_data(data_width-1 downto 0);


   bmem: accessTlbMemoryBase 
		generic map (address_width => address_width,
				data_width => data_width, 
					use_mem_cuts => use_mem_cuts)
		port map (
				start_req => start_req,
				start_ack => start_ack,
				fin_req => ureg_write_ack,
				fin_ack => ureg_write_req,
    				clear_flag => clear_flag,
    				wr_flag => wr_flag,
    				write_address => write_address,
    				write_entry => write_entry,
    				lookup_address => lookup_address,
    				l_v => ureg_write_valid,
    				lookup_entry => ureg_write_entry,
    				clk => clk, reset => reset);
			
end Mixed;


library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.mem_component_pack.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
entity accessTlbMemoryBase is -- 
  generic (address_width : integer := 8; data_width : integer := 32; use_mem_cuts: boolean := true);
  port ( -- 
    start_req: in std_logic;
    start_ack: out std_logic;
    fin_req: in std_logic;
    fin_ack: out std_logic;
    clear_flag : in  std_logic_vector(0 downto 0);
    wr_flag : in  std_logic_vector(0 downto 0);
    write_address : in  std_logic_vector(address_width-1 downto 0);
    write_entry : in  std_logic_vector(data_width-1 downto 0);
    lookup_address : in  std_logic_vector(address_width-1 downto 0);
    l_v : out  std_logic_vector(0 downto 0);
    lookup_entry : out  std_logic_vector(data_width-1 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity accessTlbMemoryBase;


architecture Mixed of accessTlbMemoryBase is

	signal valids : std_logic_vector((2**address_width)-1 downto 0);
	signal base_bank_enable: std_logic;
	signal base_bank_address: std_logic_vector(address_width-1 downto 0);
	signal base_bank_write_data, base_bank_read_data, base_bank_read_data_reg: std_logic_vector(data_width-1 downto 0);
	signal base_bank_write_bar : std_logic;

	signal lookup_address_reg, write_address_reg: std_logic_vector(address_width-1 downto 0);
	signal write_entry_reg: std_logic_vector(data_width-1 downto 0);
    	signal wr_flag_reg, clear_flag_reg : std_logic_vector(0 downto 0);

	-- state machine: 
	--             curr-state  clear_flag wr_flag start_req fin_req   next-state action
	--           	 Idle        _          _       0          _       Idle      assert start-ack 
	--               Idle        1          _       1	   1       Idle      start-ack, write 0 to valids, send zero-response 
	--		 Idle        0          1       1          _       WriteState, start-ack start read. 
	--               Idle        0          0       1          _	   ResponseState,  start-ack, read valid, start read
	--               WriteState  _          _       _          _	   ResponseState, write valid, write modified read-data.
	--               RespState   _          _       _          0	   ResponseState, present data to output, assert fin_ack, wait.
	--               RespState                      1          1       Same transitions as Idle, assert fin_ack. 
	--               RespState                      0          1       Idle, assert fin_ack
	--               
        --
	type FsmState is (IdleState, WriteState, ResponseState);
	signal fsm_state: FsmState;

-- see comment above..
--##decl_synopsys_sync_set_reset##

begin


   process(clk, reset, start_req, fin_req, 
		valids,
		wr_flag, clear_flag, write_address, write_entry, lookup_address,
		wr_flag_reg, clear_flag_reg, write_address_reg, write_entry_reg,  lookup_address_reg,
		base_bank_read_data, base_bank_read_data_reg, fsm_state
	 )
   	variable next_fsm_state: FsmState;
	variable next_valids_var : std_logic_vector((2**address_width)-1 downto 0);
	variable start_ack_var, fin_ack_var: std_logic;
	variable base_bank_enable_var, base_bank_write_bar_var: std_logic;
	variable base_bank_address_var: std_logic_vector(address_width-1 downto 0);
	variable base_bank_write_data_var : std_logic_vector(data_width-1 downto 0);
	variable next_base_bank_read_data_reg_var : std_logic_vector(data_width-1 downto 0);
	variable l_v_var: std_logic;
	variable lookup_entry_var: std_logic_vector(data_width-1 downto 0);
	variable next_write_address_reg_var: std_logic_vector(address_width-1 downto 0);
	variable next_write_entry_reg_var: std_logic_vector(data_width-1 downto 0);
    	variable next_wr_flag_reg_var, next_clear_flag_reg_var : std_logic_vector(0 downto 0);
	variable next_lookup_address_reg_var: std_logic_vector(address_width-1 downto 0);
	variable lookup_index_var, write_index_var : integer range 0 to (2**address_width - 1);
   begin
	start_ack_var := '0';
	fin_ack_var := '0';
	base_bank_enable_var := '0';
	base_bank_write_bar_var := '0';
	base_bank_address_var := (others => '0');
	base_bank_write_data_var := (others => '0');

	next_fsm_state := fsm_state;
	next_valids_var := valids;
	next_wr_flag_reg_var(0) := '0';
	next_clear_flag_reg_var(0) := '0';
	next_write_address_reg_var := write_address_reg;
	next_write_entry_reg_var := write_entry_reg;
	next_base_bank_read_data_reg_var := base_bank_read_data_reg;
	next_lookup_address_reg_var := lookup_address_reg;


	-- returned values.
	l_v_var := '0';
	lookup_entry_var := (others => '0');

	case fsm_state is
		when IdleState =>
			start_ack_var := '1';
			if(start_req = '1') then
				if(clear_flag(0) = '1') then
					next_valids_var := (others => '0');
					next_fsm_state := ResponseState;
					next_clear_flag_reg_var(0) := '1';
				else
					-- schedule a read.
					base_bank_enable_var := '1';
					base_bank_write_bar_var := '1';
					base_bank_address_var := lookup_address;
		
					-- save write information.
					next_wr_flag_reg_var := wr_flag;
					next_write_address_reg_var := write_address;
					next_write_entry_reg_var := write_entry;
					next_lookup_address_reg_var := lookup_address;

					if(wr_flag(0) = '1') then
						-- write in the next-state
						next_fsm_state := WriteState;
					else
						next_fsm_state := ResponseState;
					end if;
				end if;
			end if;
		when WriteState =>
			-- schedule a write.
			base_bank_enable_var := '1';
			base_bank_address_var := write_address_reg;
			base_bank_write_data_var := write_entry_reg;
			write_index_var := to_integer (unsigned (write_address_reg));
			lookup_index_var := to_integer (unsigned (lookup_address_reg));

			-- write will validate write-index.
			next_valids_var(write_index_var) := '1';

			next_base_bank_read_data_reg_var := base_bank_read_data;

			next_wr_flag_reg_var(0) := '1';

			l_v_var := valids (lookup_index_var);
			if(write_address_reg = lookup_address_reg)  then
				-- if lookup and just written match, make it 1.
				l_v_var := '1';
				-- also bypass write-entry to lookup-entry.
				lookup_entry_var := write_entry_reg;
			else
				lookup_entry_var := base_bank_read_data;
			end if;

			-- ack it...
			fin_ack_var := '1';
			if(fin_req = '1') then
				next_fsm_state := IdleState;
			else
				next_fsm_state := ResponseState;
			end if;
		when ResponseState =>
			fin_ack_var := '1';

			write_index_var := to_integer (unsigned (write_address_reg));
			lookup_index_var := to_integer (unsigned(lookup_address_reg));

			l_v_var := valids (lookup_index_var);
			if(wr_flag_reg(0) = '1') then
				if(write_address_reg = lookup_address_reg)  then
					l_v_var := '1';
					lookup_entry_var := write_entry_reg;
				else
					lookup_entry_var := base_bank_read_data_reg;
				end if;
			elsif (clear_flag_reg(0) = '0') then
				lookup_entry_var := base_bank_read_data;
			else 
				l_v_var := '0';
			end if;
			
			-- lets not waste a cycle..
			if(fin_req = '1') then
				start_ack_var := '1';
				if(start_req = '1') then
					if(clear_flag(0) = '1') then
						next_valids_var := (others => '0');
						next_fsm_state := ResponseState;
						next_clear_flag_reg_var(0) := '1';
					else
						-- schedule a read.
						base_bank_enable_var := '1';
						base_bank_write_bar_var := '1';
						base_bank_address_var := lookup_address;
			
						-- save write information.
						next_wr_flag_reg_var := wr_flag;
						next_write_address_reg_var := write_address;
						next_write_entry_reg_var := write_entry;
						next_lookup_address_reg_var := lookup_address;

						if(wr_flag(0) = '1') then
							-- write in the next-state
							next_fsm_state := WriteState;
						else
							next_fsm_state := ResponseState;
						end if;
					end if;
				else
					next_fsm_state := IdleState;
				end if;
			end if;
	end case;
	
	
	start_ack <= start_ack_var;
	fin_ack <= fin_ack_var;
	base_bank_enable <= base_bank_enable_var;
	base_bank_write_bar <= base_bank_write_bar_var;
	base_bank_address <= base_bank_address_var;
	base_bank_write_data <= base_bank_write_data_var;

	l_v(0) <= l_v_var;
	lookup_entry <= lookup_entry_var;

	if(clk'event and clk = '1') then
		if(reset = '1') then
			fsm_state <= IdleState;
			valids <= (others => '0');
		else
			fsm_state <= next_fsm_state;
			valids <= next_valids_var;
			wr_flag_reg <= next_wr_flag_reg_var;
			clear_flag_reg <= next_clear_flag_reg_var;
			write_address_reg <= next_write_address_reg_var;
			write_entry_reg <= next_write_entry_reg_var;
			base_bank_read_data_reg <= next_base_bank_read_data_reg_var;
			lookup_address_reg <= next_lookup_address_reg_var;
		end if;
	end if;
   end process;

   memCutBB: if use_mem_cuts generate 
   	bb: base_bank 
		generic map  (name => "accessTlbTagPte:base_bank", g_addr_width => address_width,
						g_data_width => data_width)
		port map (
				datain => base_bank_write_data,
				addrin => base_bank_address,
				dataout => base_bank_read_data,
				enable => base_bank_enable,
				writebar => base_bank_write_bar,
				clk => clk, reset => reset
			);
   end generate memCutBB;
   regBB: if not use_mem_cuts generate 
   	bb: base_bank_with_registers
		generic map  (name => "accessTlbTagPte:base_bank", g_addr_width => address_width,
						g_data_width => data_width)
		port map (
				datain => base_bank_write_data,
				addrin => base_bank_address,
				dataout => base_bank_read_data,
				enable => base_bank_enable,
				writebar => base_bank_write_bar,
				clk => clk, reset => reset
			);
   end generate regBB;
 
	
end Mixed;
library std;
use std.standard.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library AjitCustom;
use AjitCustom.AjitCoreConfigurationPackage.all;
use AjitCustom.AjitCustomComponents.all;


entity snoopFilter_Operator is
  port ( -- 
    	sample_req: in boolean;
    	sample_ack: out boolean;
    	update_req: in boolean;
    	update_ack: out boolean;
	rwbar: in std_logic_vector(0 downto 0);
	enable: in std_logic_vector(0 downto 0);
        pa_of_line:  in std_logic_vector(29 downto 0);
	send_inval: out std_logic_vector(0 downto 0);
        clk, reset: in std_logic);
end entity;


architecture Wrapper of snoopFilter_Operator is
	signal zero_sig: std_logic_vector(0 downto 0);
	signal erase, lookup, update, tlb_hit, enable_reg, rwbar_reg: std_logic_vector(0 downto 0);
	signal sample_ack_sig: boolean;
begin
	zero_sig(0)  <= '0';
	sample_ack <= sample_ack_sig;

	erase(0)  <= (enable(0) and  rwbar(0));
	lookup(0) <= (enable(0) and  (not rwbar(0)));
	update(0) <= (enable(0) and  (not rwbar(0)));
        

	basemem:genericFullyAssociativeMemoryNoData_Operator
			generic map(tag_width => 30, 
					log_number_of_entries => SNOOP_CACHE_LOG_MEMORY_SIZE,
					ignore_collisions => true)
			port map(
					sample_req => sample_req,
					sample_ack => sample_ack_sig,
					update_req => update_req,
					update_ack => update_ack,
					clear_flag => zero_sig,
					erase_flag => erase,
					write_flag => update,
					write_tag => pa_of_line,
					lookup_flag => lookup,
					lookup_tag => pa_of_line,
					lookup_valid => tlb_hit,
					clk => clk, reset => reset);

	process(clk, reset)
	begin
		if(clk'event and (clk = '1')) then
			if(sample_ack_sig) then
				enable_reg <= enable;
				rwbar_reg  <= rwbar;
			end if;
		end if;
	end process;

	send_inval(0) <= enable_reg(0) and (not rwbar_reg(0)) and (not tlb_hit(0));
end Wrapper;

library std;
use std.standard.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library AjitCustom;
use AjitCustom.AjitCoreConfigurationPackage.all;
use AjitCustom.AjitCustomComponents.all;

entity snoopFilter_1_Operator is
  port ( -- 
    	sample_req: in boolean;
    	sample_ack: out boolean;
    	update_req: in boolean;
    	update_ack: out boolean;
	rwbar: in std_logic_vector(0 downto 0);
	enable: in std_logic_vector(0 downto 0);
        pa_of_line:  in std_logic_vector(29 downto 0);
	send_inval: out std_logic_vector(0 downto 0);
        clk, reset: in std_logic);
end entity;

architecture TrivArch of snoopFilter_1_Operator is
begin
	sf: snoopFilter_Operator 
		port map (
    			sample_req,
    			sample_ack,
    			update_req,
    			update_ack,
			rwbar,
			enable,
        		pa_of_line,
			send_inval,
        		clk, reset);
end TrivArch;

library std;
use std.standard.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library AjitCustom;
use AjitCustom.AjitCoreConfigurationPackage.all;
use AjitCustom.AjitCustomComponents.all;

entity snoopFilter_2_Operator is
  port ( -- 
    	sample_req: in boolean;
    	sample_ack: out boolean;
    	update_req: in boolean;
    	update_ack: out boolean;
	rwbar: in std_logic_vector(0 downto 0);
	enable: in std_logic_vector(0 downto 0);
        pa_of_line:  in std_logic_vector(29 downto 0);
	send_inval: out std_logic_vector(0 downto 0);
        clk, reset: in std_logic);
end entity;

architecture TrivArch of snoopFilter_2_Operator is
begin
	sf: snoopFilter_Operator 
		port map (
    			sample_req,
    			sample_ack,
    			update_req,
    			update_ack,
			rwbar,
			enable,
        		pa_of_line,
			send_inval,
        		clk, reset);
end TrivArch;

library std;
use std.standard.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library AjitCustom;
use AjitCustom.AjitCoreConfigurationPackage.all;
use AjitCustom.AjitCustomComponents.all;

entity snoopFilter_4_Operator is
  port ( -- 
    	sample_req: in boolean;
    	sample_ack: out boolean;
    	update_req: in boolean;
    	update_ack: out boolean;
	rwbar: in std_logic_vector(0 downto 0);
	enable: in std_logic_vector(0 downto 0);
        pa_of_line:  in std_logic_vector(29 downto 0);
	send_inval: out std_logic_vector(0 downto 0);
        clk, reset: in std_logic);
end entity;

architecture TrivArch of snoopFilter_4_Operator is
begin
	sf: snoopFilter_Operator 
		port map (
    			sample_req,
    			sample_ack,
    			update_req,
    			update_ack,
			rwbar,
			enable,
        		pa_of_line,
			send_inval,
        		clk, reset);
end TrivArch;
library std;
use std.standard.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.mem_component_pack.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

library AjitCustom;
use AjitCustom.AjitCustomComponents.all;

entity asr_daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    iunit_asr_access_command_pipe_read_req : out  std_logic_vector(0 downto 0);
    iunit_asr_access_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
    iunit_asr_access_command_pipe_read_data : in   std_logic_vector(43 downto 0);
    iunit_asr_access_response_pipe_write_req : out  std_logic_vector(0 downto 0);
    iunit_asr_access_response_pipe_write_ack : in   std_logic_vector(0 downto 0);
    iunit_asr_access_response_pipe_write_data : out  std_logic_vector(33 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity asr_daemon;
architecture asr_daemon_arch of asr_daemon is -- 
	signal write_reg_id, read_reg_id, read_reg_id_reg : std_logic_vector(4 downto 0);
	signal write_reg_value : std_logic_vector(31 downto 0);
	signal write_valid, read_valid: std_logic;


	type FsmState is (ResetState, IdleState, ReadState, ResponseState);
        signal fsm_state, next_fsm_state: FsmState;

	signal mem_addr: std_logic_vector(4 downto 0);
	signal mem_write_data, mem_read_data: std_logic_vector(31 downto 0);
	signal mem_enable, mem_read_writebar: std_logic;

	signal counter_reg: integer range  0 to 31;
	signal read_valid_reg, write_valid_reg: std_logic_vector(0 downto 0);

	signal read_data: std_logic_vector(31 downto 0);

	--
	-- 64-bit cycle count will be returned in ASR30 and ASR31
	--
	signal cycle_count_register: unsigned(63 downto 0);

-- see comment above..
--##decl_synopsys_sync_set_reset##
begin

	-- daemon can start any time, but never finishes.
	start_ack <= '1';
	fin_ack <= '0';
        tag_out <= tag_in;

	-- input side unpacking.
	read_valid <= iunit_asr_access_command_pipe_read_data(0);
	read_reg_id <= iunit_asr_access_command_pipe_read_data(5 downto 1);
	write_valid <= iunit_asr_access_command_pipe_read_data(6);
	write_reg_value <= iunit_asr_access_command_pipe_read_data(38 downto 7);
	write_reg_id <= iunit_asr_access_command_pipe_read_data(43 downto 39);

	-- output side packing.
	iunit_asr_access_response_pipe_write_data <= 
				write_valid_reg & read_data & read_valid_reg;	

	-- state machine.
	process(clk, reset, 
			fsm_state,
			counter_reg, cycle_count_register,
			read_valid, read_reg_id, read_reg_id_reg, write_valid, write_reg_value, write_reg_id,
			read_valid_reg, write_valid_reg,
			mem_read_data,
			iunit_asr_access_command_pipe_read_ack,
			iunit_asr_access_response_pipe_write_ack)

		variable next_fsm_state_var: FsmState;
		variable mem_addr_var: std_logic_vector(4 downto 0);
		variable mem_write_data_var: std_logic_vector(31 downto 0);
		variable mem_enable_var, mem_read_writebar_var: std_logic;
	
		variable next_counter_var : integer range 0 to 31;
		variable next_cycle_count_register_var: unsigned(63 downto 0);

		variable read_req_var, write_req_var : std_logic;
		variable next_read_valid_reg_var, next_write_valid_reg_var : std_logic_vector(0 downto 0);

		variable read_data_var : std_logic_vector(31 downto 0);
		variable next_read_reg_id_reg_var : std_logic_vector(4 downto 0);

		
	begin

		next_fsm_state_var := fsm_state;
		next_counter_var := counter_reg;
		next_read_reg_id_reg_var := read_reg_id_reg;

		read_req_var := '0';
		next_read_valid_reg_var := read_valid_reg;
		next_cycle_count_register_var := cycle_count_register + 1;

		write_req_var := '0';
		next_write_valid_reg_var := write_valid_reg;

		mem_write_data_var := (others => '0');
		mem_addr_var := (others => '0');
		mem_enable_var := '0';
		mem_read_writebar_var := '1';

		read_data_var := (others => '0');

		case fsm_state is
			when ResetState =>
				mem_enable_var := '1';
				mem_read_writebar_var 	 := '0';
				mem_write_data_var := (others => '0');
				mem_addr_var := std_logic_vector(to_unsigned(counter_reg, 5));
				if (counter_reg = 31) then
				    next_fsm_state_var := IdleState;
				    next_counter_var := 0;
				else
				    next_counter_var := counter_reg + 1;
				end if;
			when IdleState =>
				read_req_var := '1';
				if(iunit_asr_access_command_pipe_read_ack(0) = '1') then
					next_read_reg_id_reg_var := read_reg_id;
					if(write_valid = '1') then
						mem_enable_var := '1';
						mem_read_writebar_var := '0';
						mem_addr_var := write_reg_id;
						mem_write_data_var := write_reg_value;
						next_write_valid_reg_var(0) := '1';
						if (read_valid = '1') then 	
							next_fsm_state_var := ReadState;
							next_read_valid_reg_var(0) := '1';
						else
							next_fsm_state_var := ResponseState;
							next_read_valid_reg_var(0) := '0';
						end if;
					elsif (read_valid = '1') then
						next_read_valid_reg_var(0) := '1';
						next_write_valid_reg_var(0) := '0';
						mem_enable_var := '1';
						mem_read_writebar_var := '1';
						mem_addr_var := read_reg_id;
						mem_write_data_var := (others => '0');
						next_fsm_state_var := ResponseState;
					else
						next_read_valid_reg_var(0) := '0';
						next_write_valid_reg_var(0) := '0';
					end if;
				end if;
			when ReadState =>

				mem_enable_var := '1';
				mem_read_writebar_var := '1';
				mem_addr_var := read_reg_id_reg;
				mem_write_data_var := (others => '0');
				next_fsm_state_var := ResponseState;
				
			when ResponseState =>
				write_req_var := '1';
				if(read_valid_reg(0) = '1') then
					if(read_reg_id_reg = "11110") then
						read_data_var := std_logic_vector(cycle_count_register(63 downto 32));
					elsif(read_reg_id_reg = "11111") then
						read_data_var := std_logic_vector(cycle_count_register(31 downto 0));
					else
						read_data_var := mem_read_data;	
					end if;
				else
					read_data_var := (others => '0');
				end if;
				if(iunit_asr_access_response_pipe_write_ack(0) = '1') then
					next_fsm_state_var := IdleState;
				end if;
		end case;

		read_data <= read_data_var;
		iunit_asr_access_command_pipe_read_req(0) <= read_req_var;
		iunit_asr_access_response_pipe_write_req(0) <= write_req_var;

		mem_addr <= mem_addr_var;
		mem_write_data <= mem_write_data_var;
		mem_enable <= mem_enable_var;
		mem_read_writebar <= mem_read_writebar_var;


		if(clk'event and clk = '1') then
			if(reset = '1') then
				fsm_state <= ResetState;
				read_valid_reg <= "0";
				write_valid_reg <= "0";
				counter_reg <= 0;
				read_reg_id_reg <= (others => '0');
				cycle_count_register <= (others => '0');
			else 
				fsm_state <= next_fsm_state_var;
				read_valid_reg <= next_read_valid_reg_var;
				write_valid_reg <= next_write_valid_reg_var;
				counter_reg <= next_counter_var;
				read_reg_id_reg <= next_read_reg_id_reg_var;
				cycle_count_register <= next_cycle_count_register_var;
			end if;
		end if;
	end process;
	

	bb: base_bank 
		generic map (name => "asr_daemon:base_bank",
				g_addr_width => 5, g_data_width => 32)
		port map (datain => mem_write_data, dataout => mem_read_data,
				addrin => mem_addr, enable => mem_enable,
					writebar => mem_read_writebar, clk => clk, reset => reset);

end asr_daemon_arch;
library std;
use std.standard.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.mem_component_pack.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

library AjitCustom;
use AjitCustom.AjitCustomComponents.all;

library AjitCustom;
use AjitCustom.AjitCoreConfigurationPackage.all;

entity asr_update_core is -- 
  port ( -- 
    core_id: in std_logic_vector(7 downto 0);
    thread_id: in std_logic_vector(7 downto 0);
    access_cmd : in  std_logic_vector(43 downto 0);
    read_val : out  std_logic_vector(31 downto 0);
    clk, reset: in std_logic;
    trigger : in boolean
  );
  -- 
end entity asr_update_core;

architecture asr_update_core_arch of asr_update_core is -- 

	signal write_reg_id, read_reg_id, read_reg_id_reg : std_logic_vector(4 downto 0);
	signal write_reg_value : std_logic_vector(31 downto 0);
	signal write_valid, read_valid: std_logic;

	signal read_data, mem_read_data: std_logic_vector(31 downto 0);

	--
	-- 64-bit cycle count will be returned in ASR30 and ASR31
	--
	signal cycle_count_register: unsigned(63 downto 0);
	signal read_valid_reg, write_valid_reg: std_logic;

	signal   thread_description_value: std_logic_vector(31 downto 0);
	constant MY_MAGIC_STRING: std_logic_vector(15 downto 0) := X"5052";

	signal is_special_read, is_special_read_reg: boolean;
	signal special_read_data, special_read_data_reg: std_logic_vector(31 downto 0);

-- see comment above..
--##decl_synopsys_sync_set_reset##
begin

	-- input side unpacking.
	-- write-reg-id write-reg-value write-valid read-reg-id read-valid
	--     5             32             1           5          1
	read_valid <= access_cmd(0) when trigger else '0';
	read_reg_id <= access_cmd(5 downto 1);
	write_valid <= access_cmd(6) when trigger else '0';
	write_reg_value <= access_cmd(38 downto 7);
	write_reg_id <= access_cmd(43 downto 39);

	-- output side packing.
	read_val <= special_read_data_reg when is_special_read_reg else mem_read_data;

	-- state machine.
	process(clk, reset, trigger, cycle_count_register)
		variable next_cycle_count_register_var: unsigned(63 downto 0);
	begin
		next_cycle_count_register_var := cycle_count_register + 1;

		if(clk'event and clk = '1') then
			if(reset = '1') then
				cycle_count_register <= (others => '0');
			else 
				cycle_count_register <= next_cycle_count_register_var;
				if(trigger) then
					is_special_read_reg <= is_special_read;
					special_read_data_reg <= special_read_data;
				end if;
			end if;
		end if;
	end process;
	

	bb: register_file_1w_1r_port
		generic map ("asr_update_core:register_file_1w_1r_port", g_addr_width => 5, g_data_width => 32)
			port map (
				-- write port 0
	 			datain_0 => write_reg_value,
         			addrin_0 => write_reg_id,
         			enable_0 => write_valid,
	 			-- read port 1
         			dataout_1 => mem_read_data,
         			addrin_1  => read_reg_id,
         			enable_1  => read_valid,
         			clk => clk,
         			reset => reset);

	process(read_reg_id, cycle_count_register, thread_description_value)
	     variable read_data_var: std_logic_vector(31 downto 0);
	     variable is_special_read_var : boolean;
	begin
	     read_data_var := (others => '0');
	     is_special_read_var := false;
             if(read_reg_id= "11110") then
                   read_data_var := std_logic_vector(cycle_count_register(63 downto 32));
		   is_special_read_var := true;
             elsif(read_reg_id = "11111") then
                    read_data_var := std_logic_vector(cycle_count_register(31 downto 0));
		   is_special_read_var := true;
             -- core_id, cpu_id mapped to asr 29 
             elsif (read_reg_id  = "11101")  then
                   read_data_var := MY_MAGIC_STRING & core_id & thread_id;
		   is_special_read_var := true;
             -- thread description information register mapped to asr 28.
             elsif (read_reg_id = "11100")  then
                   read_data_var := thread_description_value;
		   is_special_read_var := true;
	     end if;
	     is_special_read   <= is_special_read_var;
	     special_read_data <= read_data_var;
	end process;
     
	
        -- Thread description value.....
	thread_description_value(31 downto 30) <=
			"11" when (LOG_DCACHE_SIZE_IN_BLOCKS = 9) 
			else "10" when (LOG_DCACHE_SIZE_IN_BLOCKS = 8)
			else "01" when (LOG_DCACHE_SIZE_IN_BLOCKS = 7)
			else "00";
	thread_description_value(29 downto 28) <=
			"11" when (LOG_ICACHE_SIZE_IN_BLOCKS = 9) 
			else "10" when (LOG_ICACHE_SIZE_IN_BLOCKS = 8)
			else "01" when (LOG_ICACHE_SIZE_IN_BLOCKS = 7)
			else "00";
	thread_description_value(27 downto 26) <=
			"00" when LOG_DCACHE_SET_ASSOCIATIVITY = 0 
				else "01" when LOG_DCACHE_SET_ASSOCIATIVITY = 1
				else "10" when LOG_DCACHE_SET_ASSOCIATIVITY = 2
				else "11";
	thread_description_value(25 downto 24) <=
			"00" when LOG_ICACHE_SET_ASSOCIATIVITY = 0 
				else "01" when LOG_ICACHE_SET_ASSOCIATIVITY = 1
				else "10" when LOG_ICACHE_SET_ASSOCIATIVITY = 2
				else "11";
	thread_description_value(23 downto 20) <=
			std_logic_vector(to_unsigned(DCACHE_HIT_LATENCY,4));
	thread_description_value(19 downto 16) <=
			std_logic_vector(to_unsigned(ICACHE_HIT_LATENCY,4));
	thread_description_value(15 downto 12) <=
			std_logic_vector(to_unsigned(TLB_NEW_3_LOG_MEM_SIZE,4));
	thread_description_value(11 downto 9) <=
			std_logic_vector(to_unsigned(TLB_NEW_2_LOG_MEM_SIZE,3));
	thread_description_value(8 downto 7) <=
			std_logic_vector(to_unsigned(TLB_NEW_1_LOG_MEM_SIZE,2));
	thread_description_value(6 downto 5) <=
			std_logic_vector(to_unsigned(TLB_NEW_0_LOG_MEM_SIZE,2));
	thread_description_value(4 downto 3) <= "00";
	thread_description_value(2) <= '1' when TREAT_NONCACHEABLE_AS_BYPASS = 1 else '0';
	thread_description_value(1) <= '1' when TWO_THREADS_IN_CORE = 1 else '0';
	thread_description_value(0) <= '1' when THREAD_IS_ISA_64 = 1 else '0';

end asr_update_core_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.BaseComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;

entity asr_update_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    core_id: in std_logic_vector(7 downto 0);
    thread_id: in std_logic_vector(7 downto 0);
    access_cmd : in  std_logic_vector(43 downto 0);
    read_val : out  std_logic_vector(31 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity asr_update_Operator;

architecture MpdIsAKlutz of asr_update_Operator is
	signal trigger, trigger_reg: boolean;

    	signal core_read_val : std_logic_vector(31 downto 0);
    	signal core_read_val_reg : std_logic_vector(31 downto 0);
    	signal access_cmd_reg, access_cmd_qualified : std_logic_vector(43 downto 0);
begin

   trig_join: join2 generic map (name => "bpbV2:trig-join", bypass => true)
			port map (pred0 => sample_req, pred1 => update_req,
					symbol_out => trigger, clk => clk, reset => reset);

    sample_ack <= trigger;
    
    process(clk, reset)
    begin
	if(clk'event and (clk = '1')) then
		if(reset = '1') then
			update_ack <= false;
			access_cmd_reg <= (others => '0');
		else
    			update_ack <= trigger;
			trigger_reg <= trigger;
			if(trigger_reg) then
				core_read_val_reg <= core_read_val;
			end if;

			if(sample_req) then
				access_cmd_reg <= access_cmd;
			end if;
		end if;
	end if;
    end process;

    access_cmd_qualified <= access_cmd when sample_req else access_cmd_reg;


  
   core: asr_update_core
  	port map ( -- 
			core_id => core_id,
			thread_id => thread_id,
			trigger => trigger,
			access_cmd => access_cmd_qualified,
			read_val => core_read_val,
    			clk => clk,
    			reset => reset
  		);

   read_val <= core_read_val when trigger_reg else core_read_val_reg;

end architecture MpdIsAKlutz;
-- Pipe multiplexor at input end of iu-register file
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.mem_component_pack.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;

entity iunit_writeback_in_mux_ajit_64_daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    iunit_64_exec_fast_alu_result_to_writeback_pipe_read_req : out  std_logic_vector(0 downto 0);
    iunit_64_exec_fast_alu_result_to_writeback_pipe_read_ack : in   std_logic_vector(0 downto 0);
    iunit_64_exec_fast_alu_result_to_writeback_pipe_read_data : in   std_logic_vector(140 downto 0);
    iunit_64_exec_to_writeback_pipe_read_req : out  std_logic_vector(0 downto 0);
    iunit_64_exec_to_writeback_pipe_read_ack : in   std_logic_vector(0 downto 0);
    iunit_64_exec_to_writeback_pipe_read_data : in   std_logic_vector(157 downto 0);
    noblock_teu_idispatch_to_iunit_writeback_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_teu_idispatch_to_iunit_writeback_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_teu_idispatch_to_iunit_writeback_pipe_read_data : in   std_logic_vector(83 downto 0);
    teu_fpunit_trap_to_iunit_pipe_read_req : out  std_logic_vector(0 downto 0);
    teu_fpunit_trap_to_iunit_pipe_read_ack : in   std_logic_vector(0 downto 0);
    teu_fpunit_trap_to_iunit_pipe_read_data : in   std_logic_vector(12 downto 0);
    teu_loadstore_to_iunit_pipe_read_req : out  std_logic_vector(0 downto 0);
    teu_loadstore_to_iunit_pipe_read_ack : in   std_logic_vector(0 downto 0);
    teu_loadstore_to_iunit_pipe_read_data : in   std_logic_vector(77 downto 0);
    teu_stream_corrector_to_iunit_pipe_read_req : out  std_logic_vector(0 downto 0);
    teu_stream_corrector_to_iunit_pipe_read_ack : in   std_logic_vector(0 downto 0);
    teu_stream_corrector_to_iunit_pipe_read_data : in   std_logic_vector(17 downto 0);
    noblock_iunit_64_writeback_in_args_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_iunit_64_writeback_in_args_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_iunit_64_writeback_in_args_pipe_pipe_write_data : out  std_logic_vector(436 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity iunit_writeback_in_mux_ajit_64_daemon;
architecture iunit_writeback_in_mux_ajit_64_daemon_arch of 
		iunit_writeback_in_mux_ajit_64_daemon is -- 
	signal dispatch_rdy, sc_rdy, ls_rdy, fp_rdy, exec_rdy, exec_fast_rdy : boolean;
	signal iuregs_rdy: boolean;

	signal get_from_sc, get_from_ls, get_from_fp, get_from_exec, get_from_exec_fast: boolean;

	signal do_transfer: boolean;

    	signal data_from_exec_fast : std_logic_vector(140 downto 0);
    	signal data_from_exec : std_logic_vector(157 downto 0);
    	signal from_dispatch, data_from_dispatch : std_logic_vector(83 downto 0);
    	signal data_from_fp : std_logic_vector(12 downto 0);
    	signal data_from_ls : std_logic_vector(77 downto 0);
    	signal data_from_sc : std_logic_vector(17 downto 0);
    	signal data_to_iuregs : std_logic_vector(436 downto 0);

	signal pop_req_to_dispatch,
		pop_req_to_exec_fast, pop_req_to_exec, pop_req_to_sc, pop_req_to_ls, pop_req_to_fp: std_logic;

	signal pop_ack_from_dispatch, pop_ack_from_exec_fast, 
			pop_ack_from_exec, pop_ack_from_sc, pop_ack_from_ls, pop_ack_from_fp: std_logic;

	signal get_flags: std_logic_vector(4 downto 0);

	signal data_from_sc_to_wb: std_logic_vector ( 5 downto 0);
	signal data_from_ls_to_wb : std_logic_vector (65 downto 0);
	signal data_from_fp_to_wb : std_logic_vector (0 downto 0);
	signal data_from_exec_slow_to_wb : std_logic_vector (145 downto 0);
	signal data_from_exec_fast_to_wb : std_logic_vector (128 downto 0);

	

begin --  
	tag_out <= tag_in;
	start_ack <= '1';
	fin_ack <= '0';

	-- dispatch side information.
	--    queue-depth = 0 since dispatch->iu-writeback is not a p2p pipe.
	qbDispatch: QueueBase
		generic map (name => "iu_wb_in_mux_qbDispatch", queue_depth => 0, data_width => 84)
		port map (
			clk => clk, reset => reset,
			data_in => noblock_teu_idispatch_to_iunit_writeback_pipe_read_data ,
			push_req => noblock_teu_idispatch_to_iunit_writeback_pipe_read_ack(0) ,
			push_ack => noblock_teu_idispatch_to_iunit_writeback_pipe_read_req(0) ,
			data_out => data_from_dispatch,
			pop_req  => pop_req_to_dispatch,
			pop_ack  => pop_ack_from_dispatch);
	-- dispatch_rdy <= (pop_ack_from_dispatch = '1') and (data_from_dispatch(83) = '1'); 
	--  no need to check bit 83.. we are not using the nonblocking nature of the access.
	dispatch_rdy <= (pop_ack_from_dispatch = '1');
	from_dispatch <= data_from_dispatch when dispatch_rdy else (others => '0');

	get_from_fp 	   <= dispatch_rdy and (from_dispatch(34) = '1');
	get_from_ls 	   <= dispatch_rdy and (from_dispatch(35) = '1');
	get_from_sc 	   <= dispatch_rdy and (from_dispatch(36) = '1');
	get_from_exec 	   <= dispatch_rdy and (from_dispatch(37) = '1');
	get_from_exec_fast <= dispatch_rdy and (from_dispatch(38) = '1');

	-- consistent with writeback-in-mux in Aa.
	get_flags(2) <= from_dispatch(34);   -- fp
	get_flags(3) <= from_dispatch(35);   -- ls
	get_flags(4) <= from_dispatch(36);   -- sc
	get_flags(1) <= from_dispatch(37);   -- iu
	get_flags(0) <= from_dispatch(38);-- iu-fast

	-- from exec-fast, bypassed..
	qbExecFast: QueueWithBypass
		generic map (name => "iu_wb_in_mux_qbExecFast", queue_depth => 2, data_width => 141)
		port map (
			clk => clk, reset => reset,
			data_in => iunit_64_exec_fast_alu_result_to_writeback_pipe_read_data,
			push_req => iunit_64_exec_fast_alu_result_to_writeback_pipe_read_ack(0),
			push_ack => iunit_64_exec_fast_alu_result_to_writeback_pipe_read_req(0),
			data_out => data_from_exec_fast,
			pop_req  => pop_req_to_exec_fast,
			pop_ack  => pop_ack_from_exec_fast);

	exec_fast_rdy <= pop_ack_from_exec_fast= '1';
	data_from_exec_fast_to_wb <= data_from_exec_fast(128 downto 0) when get_from_exec_fast else (others => '0');

	-- from exec, bypassed..
	qbExec: QueueWithBypass
		generic map (name => "iu_wb_in_mux_qbExec", queue_depth => 2, data_width => 158)
		port map (
			clk => clk, reset => reset,
			data_in => iunit_64_exec_to_writeback_pipe_read_data,
			push_req => iunit_64_exec_to_writeback_pipe_read_ack(0),
			push_ack => iunit_64_exec_to_writeback_pipe_read_req(0),
			data_out => data_from_exec,
			pop_req  => pop_req_to_exec,
			pop_ack  => pop_ack_from_exec);

	exec_rdy <= pop_ack_from_exec = '1';
	data_from_exec_slow_to_wb <= data_from_exec(145 downto 0)  when get_from_exec else (others => '0');


	-- from sc: bypassing gives boost? check.
	qbSC: QueueWithBypass
		generic map (name => "iu_wb_in_mux_qbSC", queue_depth => 2, data_width => 18)
		port map (
			clk => clk, reset => reset,
			data_in => teu_stream_corrector_to_iunit_pipe_read_data,
			push_req => teu_stream_corrector_to_iunit_pipe_read_ack(0),
			push_ack => teu_stream_corrector_to_iunit_pipe_read_req(0),
			data_out => data_from_sc,
			pop_req  => pop_req_to_sc,
			pop_ack  => pop_ack_from_sc);


	sc_rdy <= pop_ack_from_sc = '1';
	data_from_sc_to_wb <= data_from_sc(5 downto 0)  when get_from_sc else (others => '0');


	-- from ls: try bypass... if critical path is ok.
	qbLS: QueueWithBypass
		generic map (name => "iu_wb_in_mux_qbLS", queue_depth => 2, data_width => 78)
		port map (
			clk => clk, reset => reset,
			data_in => teu_loadstore_to_iunit_pipe_read_data,
			push_req => teu_loadstore_to_iunit_pipe_read_ack(0),
			push_ack => teu_loadstore_to_iunit_pipe_read_req(0),
			data_out => data_from_ls,
			pop_req  => pop_req_to_ls,
			pop_ack  => pop_ack_from_ls);

	ls_rdy <= pop_ack_from_ls = '1';
	data_from_ls_to_wb <= data_from_ls(65 downto 0)  when get_from_ls else (others => '0');

	-- from fpunit
	qbFP: QueueWithBypass
		generic map (name => "iu_wb_in_mux_qbFP", queue_depth => 3, data_width => 13)
		port map (
			clk => clk, reset => reset,
			data_in => teu_fpunit_trap_to_iunit_pipe_read_data,
			push_req => teu_fpunit_trap_to_iunit_pipe_read_ack(0),
			push_ack => teu_fpunit_trap_to_iunit_pipe_read_req(0),
			data_out => data_from_fp,
			pop_req  => pop_req_to_fp,
			pop_ack  => pop_ack_from_fp);

	fp_rdy <= pop_ack_from_fp = '1';
	data_from_fp_to_wb(0) <= data_from_fp(0)  when get_from_fp else '0';


	data_to_iuregs <= from_dispatch & get_flags & 
				data_from_sc_to_wb & data_from_ls_to_wb & data_from_fp_to_wb & data_from_exec_slow_to_wb & data_from_exec_fast_to_wb;
	iuregs_rdy <= noblock_iunit_64_writeback_in_args_pipe_pipe_write_ack (0) = '1';

	do_transfer <= (dispatch_rdy 
				and iuregs_rdy
				and ((not get_from_sc) or sc_rdy)
				and ((not get_from_ls) or ls_rdy)
				and ((not get_from_fp) or fp_rdy)
				and ((not get_from_exec) or exec_rdy)
				and ((not get_from_exec_fast) or exec_fast_rdy));
	

	-- requests to writers.
    	pop_req_to_dispatch  <= '1' when do_transfer else '0';

    	pop_req_to_exec_fast <= '1' when (do_transfer and get_from_exec_fast) else '0';
    	pop_req_to_exec <= '1' when (do_transfer and get_from_exec) else '0';
    	pop_req_to_fp <= '1' when (do_transfer and get_from_fp) else '0';
    	pop_req_to_ls <= '1' when (do_transfer and get_from_ls) else '0';
    	pop_req_to_sc <= '1' when (do_transfer and get_from_sc) else '0';

	-- requests to reader.
    	noblock_iunit_64_writeback_in_args_pipe_pipe_write_req(0) <= '1' when do_transfer else '0';

	-- data to reader.
    	noblock_iunit_64_writeback_in_args_pipe_pipe_write_data <= data_to_iuregs;

end iunit_writeback_in_mux_ajit_64_daemon_arch;
-- Pipe multiplexor at input end of iu-register file
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.mem_component_pack.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;

entity iunit_writeback_in_mux_daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    iunit_exec_fast_alu_result_to_writeback_pipe_read_req : out  std_logic_vector(0 downto 0);
    iunit_exec_fast_alu_result_to_writeback_pipe_read_ack : in   std_logic_vector(0 downto 0);
    iunit_exec_fast_alu_result_to_writeback_pipe_read_data : in   std_logic_vector(108 downto 0);
    iunit_exec_to_writeback_pipe_read_req : out  std_logic_vector(0 downto 0);
    iunit_exec_to_writeback_pipe_read_ack : in   std_logic_vector(0 downto 0);
    iunit_exec_to_writeback_pipe_read_data : in   std_logic_vector(125 downto 0);
    noblock_teu_idispatch_to_iunit_writeback_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_teu_idispatch_to_iunit_writeback_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_teu_idispatch_to_iunit_writeback_pipe_read_data : in   std_logic_vector(83 downto 0);
    teu_fpunit_trap_to_iunit_pipe_read_req : out  std_logic_vector(0 downto 0);
    teu_fpunit_trap_to_iunit_pipe_read_ack : in   std_logic_vector(0 downto 0);
    teu_fpunit_trap_to_iunit_pipe_read_data : in   std_logic_vector(12 downto 0);
    teu_loadstore_to_iunit_pipe_read_req : out  std_logic_vector(0 downto 0);
    teu_loadstore_to_iunit_pipe_read_ack : in   std_logic_vector(0 downto 0);
    teu_loadstore_to_iunit_pipe_read_data : in   std_logic_vector(77 downto 0);
    teu_stream_corrector_to_iunit_pipe_read_req : out  std_logic_vector(0 downto 0);
    teu_stream_corrector_to_iunit_pipe_read_ack : in   std_logic_vector(0 downto 0);
    teu_stream_corrector_to_iunit_pipe_read_data : in   std_logic_vector(17 downto 0);
    noblock_iunit_writeback_in_args_pipe_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_iunit_writeback_in_args_pipe_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_iunit_writeback_in_args_pipe_pipe_write_data : out  std_logic_vector(372 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity iunit_writeback_in_mux_daemon;
architecture iunit_writeback_in_mux_daemon_arch of iunit_writeback_in_mux_daemon is -- 
	signal dispatch_rdy, sc_rdy, ls_rdy, fp_rdy, exec_rdy, exec_fast_rdy : boolean;
	signal iuregs_rdy: boolean;

	signal get_from_sc, get_from_ls, get_from_fp, get_from_exec, get_from_exec_fast: boolean;

	signal do_transfer: boolean;

    	signal data_from_exec_fast : std_logic_vector(108 downto 0);
    	signal data_from_exec : std_logic_vector(125 downto 0);
    	signal from_dispatch, data_from_dispatch : std_logic_vector(83 downto 0);
    	signal data_from_fp : std_logic_vector(12 downto 0);
    	signal data_from_ls : std_logic_vector(77 downto 0);
    	signal data_from_sc : std_logic_vector(17 downto 0);
    	signal data_to_iuregs : std_logic_vector(372 downto 0);

	signal pop_req_to_dispatch,
		pop_req_to_exec_fast, pop_req_to_exec, pop_req_to_sc, pop_req_to_ls, pop_req_to_fp: std_logic;

	signal pop_ack_from_dispatch, pop_ack_from_exec_fast, 
			pop_ack_from_exec, pop_ack_from_sc, pop_ack_from_ls, pop_ack_from_fp: std_logic;

	signal get_flags: std_logic_vector(4 downto 0);

	signal data_from_sc_to_wb: std_logic_vector ( 5 downto 0);
	signal data_from_ls_to_wb : std_logic_vector (65 downto 0);
	signal data_from_fp_to_wb : std_logic_vector (0 downto 0);
	signal data_from_exec_slow_to_wb : std_logic_vector (113 downto 0);
	signal data_from_exec_fast_to_wb : std_logic_vector (96 downto 0);

	

begin --  
	tag_out <= tag_in;
	start_ack <= '1';
	fin_ack <= '0';

	-- dispatch side information.
	--    queue-depth = 0 since dispatch->iu-writeback is not a p2p pipe.
	qbDispatch: QueueBase
		generic map (name => "iu_wb_in_mux_qbDispatch", queue_depth => 0, data_width => 84)
		port map (
			clk => clk, reset => reset,
			data_in => noblock_teu_idispatch_to_iunit_writeback_pipe_read_data ,
			push_req => noblock_teu_idispatch_to_iunit_writeback_pipe_read_ack(0) ,
			push_ack => noblock_teu_idispatch_to_iunit_writeback_pipe_read_req(0) ,
			data_out => data_from_dispatch,
			pop_req  => pop_req_to_dispatch,
			pop_ack  => pop_ack_from_dispatch);
	-- dispatch_rdy <= (pop_ack_from_dispatch = '1') and (data_from_dispatch(83) = '1'); 
	--  no need to check bit 83.. we are not using the nonblocking nature of the access.
	dispatch_rdy <= (pop_ack_from_dispatch = '1');
	from_dispatch <= data_from_dispatch when dispatch_rdy else (others => '0');

	get_from_fp 	   <= dispatch_rdy and (from_dispatch(34) = '1');
	get_from_ls 	   <= dispatch_rdy and (from_dispatch(35) = '1');
	get_from_sc 	   <= dispatch_rdy and (from_dispatch(36) = '1');
	get_from_exec 	   <= dispatch_rdy and (from_dispatch(37) = '1');
	get_from_exec_fast <= dispatch_rdy and (from_dispatch(38) = '1');

	-- consistent with writeback-in-mux in Aa.
	get_flags(2) <= from_dispatch(34);   -- fp
	get_flags(3) <= from_dispatch(35);   -- ls
	get_flags(4) <= from_dispatch(36);   -- sc
	get_flags(1) <= from_dispatch(37);   -- iu
	get_flags(0) <= from_dispatch(38);-- iu-fast

	-- from exec-fast, bypassed..
	qbExecFast: QueueWithBypass
		generic map (name => "iu_wb_in_mux_qbExecFast", queue_depth => 2, data_width => 109)
		port map (
			clk => clk, reset => reset,
			data_in => iunit_exec_fast_alu_result_to_writeback_pipe_read_data,
			push_req => iunit_exec_fast_alu_result_to_writeback_pipe_read_ack(0),
			push_ack => iunit_exec_fast_alu_result_to_writeback_pipe_read_req(0),
			data_out => data_from_exec_fast,
			pop_req  => pop_req_to_exec_fast,
			pop_ack  => pop_ack_from_exec_fast);

	exec_fast_rdy <= pop_ack_from_exec_fast= '1';
	data_from_exec_fast_to_wb <= data_from_exec_fast(96 downto 0) when get_from_exec_fast else (others => '0');

	-- from exec, bypassed..
	qbExec: QueueWithBypass
		generic map (name => "iu_wb_in_mux_qbExec", queue_depth => 2, data_width => 126)
		port map (
			clk => clk, reset => reset,
			data_in => iunit_exec_to_writeback_pipe_read_data,
			push_req => iunit_exec_to_writeback_pipe_read_ack(0),
			push_ack => iunit_exec_to_writeback_pipe_read_req(0),
			data_out => data_from_exec,
			pop_req  => pop_req_to_exec,
			pop_ack  => pop_ack_from_exec);

	exec_rdy <= pop_ack_from_exec = '1';
	data_from_exec_slow_to_wb <= data_from_exec(113 downto 0)  when get_from_exec else (others => '0');


	-- from sc: bypassing gives boost? check.
	qbSC: QueueWithBypass
		generic map (name => "iu_wb_in_mux_qbSC", queue_depth => 2, data_width => 18)
		port map (
			clk => clk, reset => reset,
			data_in => teu_stream_corrector_to_iunit_pipe_read_data,
			push_req => teu_stream_corrector_to_iunit_pipe_read_ack(0),
			push_ack => teu_stream_corrector_to_iunit_pipe_read_req(0),
			data_out => data_from_sc,
			pop_req  => pop_req_to_sc,
			pop_ack  => pop_ack_from_sc);


	sc_rdy <= pop_ack_from_sc = '1';
	data_from_sc_to_wb <= data_from_sc(5 downto 0)  when get_from_sc else (others => '0');


	-- from ls: try bypass... if critical path is ok.
	qbLS: QueueWithBypass
		generic map (name => "iu_wb_in_mux_qbLS", queue_depth => 2, data_width => 78)
		port map (
			clk => clk, reset => reset,
			data_in => teu_loadstore_to_iunit_pipe_read_data,
			push_req => teu_loadstore_to_iunit_pipe_read_ack(0),
			push_ack => teu_loadstore_to_iunit_pipe_read_req(0),
			data_out => data_from_ls,
			pop_req  => pop_req_to_ls,
			pop_ack  => pop_ack_from_ls);

	ls_rdy <= pop_ack_from_ls = '1';
	data_from_ls_to_wb <= data_from_ls(65 downto 0)  when get_from_ls else (others => '0');

	-- from fpunit
	qbFP: QueueWithBypass
		generic map (name => "iu_wb_in_mux_qbFP", queue_depth => 3, data_width => 13)
		port map (
			clk => clk, reset => reset,
			data_in => teu_fpunit_trap_to_iunit_pipe_read_data,
			push_req => teu_fpunit_trap_to_iunit_pipe_read_ack(0),
			push_ack => teu_fpunit_trap_to_iunit_pipe_read_req(0),
			data_out => data_from_fp,
			pop_req  => pop_req_to_fp,
			pop_ack  => pop_ack_from_fp);

	fp_rdy <= pop_ack_from_fp = '1';
	data_from_fp_to_wb(0) <= data_from_fp(0)  when get_from_fp else '0';


	data_to_iuregs <= from_dispatch & get_flags & 
				data_from_sc_to_wb & data_from_ls_to_wb & data_from_fp_to_wb & data_from_exec_slow_to_wb & data_from_exec_fast_to_wb;
	iuregs_rdy <= noblock_iunit_writeback_in_args_pipe_pipe_write_ack (0) = '1';

	do_transfer <= (dispatch_rdy 
				and iuregs_rdy
				and ((not get_from_sc) or sc_rdy)
				and ((not get_from_ls) or ls_rdy)
				and ((not get_from_fp) or fp_rdy)
				and ((not get_from_exec) or exec_rdy)
				and ((not get_from_exec_fast) or exec_fast_rdy));
	

	-- requests to writers.
    	pop_req_to_dispatch  <= '1' when do_transfer else '0';

    	pop_req_to_exec_fast <= '1' when (do_transfer and get_from_exec_fast) else '0';
    	pop_req_to_exec <= '1' when (do_transfer and get_from_exec) else '0';
    	pop_req_to_fp <= '1' when (do_transfer and get_from_fp) else '0';
    	pop_req_to_ls <= '1' when (do_transfer and get_from_ls) else '0';
    	pop_req_to_sc <= '1' when (do_transfer and get_from_sc) else '0';

	-- requests to reader.
    	noblock_iunit_writeback_in_args_pipe_pipe_write_req(0) <= '1' when do_transfer else '0';

	-- data to reader.
    	noblock_iunit_writeback_in_args_pipe_pipe_write_data <= data_to_iuregs;

end iunit_writeback_in_mux_daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.mem_component_pack.all;

library AjitCustom;
use AjitCustom.AjitCustomComponents.all;

-- two ports 
--    port 1 for reads
--    port 0 for writes
--
-- Note: on write/read collision,
--     the written value is available as read_data_0
--     and maintained until the next enable.
-- 
entity window_registers_bank is
	generic (name : string := "anon");
	port (trigger: in boolean; 
		write_enable_0: in std_logic;
		address_0, address_1: in std_logic_vector(5 downto 0);
		read_data_1 : out std_logic_vector(31 downto 0);
		write_data_0: in std_logic_vector(31 downto 0);
		clk, reset: in std_logic);
end entity window_registers_bank;
architecture Simple of window_registers_bank is
	signal mem_data_out_1, mem_data_in_0, bypass_data_reg, mem_data_out_1_reg: std_logic_vector(31 downto 0);
	signal use_bypass_reg, trigger_reg, collision: boolean;
	signal mem_enable_0, mem_enable_1: std_logic;
begin
	collision <= (write_enable_0 = '1') and (address_0 = address_1);
	-- The whole bypass angle..
	process(clk, reset, trigger, trigger_reg, collision, write_enable_0, write_data_0)
	begin
		if(clk'event and (clk = '1')) then
			if(reset = '1') then
				use_bypass_reg <= false;
			else
				if(trigger) then 
					use_bypass_reg <= collision;
					bypass_data_reg    <= write_data_0;
				end if;

				trigger_reg <= trigger;

				if(trigger_reg) then
					mem_data_out_1_reg <= mem_data_out_1;
				end if;	
			end if;
		end if;
	end process;


	mem_data_in_0 <= write_data_0;
	mem_enable_0  <= write_enable_0 when trigger else '0';
	mem_enable_1  <= '1'  when (trigger and (not collision)) else '0';


	bb: register_file_1w_1r_port
		generic map (name & ":register_file_1w_1r_port", g_addr_width => 6, g_data_width => 32)
			port map (
				-- write port 0
	 			datain_0 => mem_data_in_0,
         			addrin_0 => address_0,
         			enable_0 => mem_enable_0,
	 			-- read port 1
         			dataout_1 => mem_data_out_1,
         			addrin_1  => address_1,
         			enable_1  => mem_enable_1,
         			clk => clk,
         			reset => reset);

	-- either from bypass data or from mem data (note use of mem_data_out_reg.
	read_data_1 <= bypass_data_reg when use_bypass_reg else mem_data_out_1 when trigger_reg else 
				mem_data_out_1_reg;
end Simple;


library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.basecomponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
entity iu_registers_3r_1w_port_register_file_inner is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    rs1 : in  std_logic_vector(4 downto 0);
    rs2 : in  std_logic_vector(4 downto 0);
    read_rd : in  std_logic_vector(4 downto 0);
    read_cwp : in  std_logic_vector(4 downto 0);
    write_gpr_even : in  std_logic_vector(0 downto 0);
    write_gpr_odd : in  std_logic_vector(0 downto 0);
    write_rd : in  std_logic_vector(4 downto 0);
    write_gpr_value_even : in  std_logic_vector(31 downto 0);
    write_gpr_value_odd : in  std_logic_vector(31 downto 0);
    write_cwp : in  std_logic_vector(4 downto 0);
    reg_pair_values : out  std_logic_vector(191 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity iu_registers_3r_1w_port_register_file_inner;
architecture iu_registers_3r_1w_port_register_file_inner_arch of iu_registers_3r_1w_port_register_file_inner is -- 

	signal trigger:boolean;

	signal mem_enable_rs1_even, mem_enable_rs1_odd,
			mem_enable_rs2_even, mem_enable_rs2_odd,
				mem_enable_rd_even, mem_enable_rd_odd: std_logic;
	signal mem_rs1_read_address, mem_rs2_read_address,
			mem_read_rd_read_address, mem_write_rd_write_address : std_logic_vector (5 downto 0);

	signal mem_rs1_read_data, mem_rs2_read_data,
			mem_read_rd_read_data, mem_write_rd_write_data : std_logic_vector (63 downto 0);
			
	signal mem_writebar_rs1_even, mem_writebar_rs1_odd,
			mem_writebar_rs2_even, mem_writebar_rs2_odd,
				mem_writebar_rd_even, mem_writebar_rd_odd: std_logic;

	type RegArray is array (natural range <>) of std_logic_vector(31 downto 0);

	-- global_registers are handled separately.
	signal global_registers : RegArray (0 to 7);


	signal rs1_data_reg_even, 
		rs1_data_reg_odd,
		rs2_data_reg_even, 
		rs2_data_reg_odd,
		rd_data_reg_even, 
		rd_data_reg_odd: std_logic_vector(31 downto 0);

	signal g_rs1_data_reg_even, 
		g_rs1_data_reg_odd,
		g_rs2_data_reg_even, 
		g_rs2_data_reg_odd,
		g_read_rd_data_reg_even, 
		g_read_rd_data_reg_odd: std_logic_vector(31 downto 0);


	signal rs1_index, rs2_index, read_rd_index, write_rd_index: integer range 0 to 31;
	signal rs1_even_index, rs2_even_index, read_rd_even_index, write_rd_even_index: integer range 0 to 31;
	signal rs1_odd_index, rs2_odd_index, read_rd_odd_index, write_rd_odd_index: integer range 0 to 31;
	signal rs1_pair_index, rs2_pair_index, read_rd_pair_index, write_rd_pair_index: integer range 0 to 15;

	signal use_rs1_global, use_rs2_global, use_read_rd_global, use_write_rd_global: boolean;
	signal use_rs1_global_reg, use_rs2_global_reg, use_read_rd_global_reg, use_write_rd_global_reg: boolean;
	
	signal write_enable_even, write_enable_odd: std_logic;

	signal bypass_global_to_rs1_even, bypass_global_to_rs2_even, bypass_global_to_read_rd_even: boolean;
	signal bypass_global_to_rs1_odd, bypass_global_to_rs2_odd, bypass_global_to_read_rd_odd: boolean;
	
	signal g_rs1_index_match, g_rs2_index_match, g_read_rd_index_match: boolean;

	signal rs1_pair_value, rs2_pair_value, rd_pair_value: std_logic_vector(63 downto 0);
begin --  

	-------------------------------------------------------------------------------
	-- trigger logic
	-------------------------------------------------------------------------------
        trig_join: join2 generic map (name => "iu_3r_1w:trig-join", bypass => true)
			port map (pred0 => sample_req, pred1 => update_req,
					symbol_out => trigger, clk => clk, reset => reset);
	sample_ack <= trigger;
	process(clk, reset)
	begin
		if(clk'event and (clk = '1')) then
			if(reset = '1') then
				update_ack <= false;
			else
				update_ack <= trigger;
			end if;
		end if;
	end process;

	-------------------------------------------------------------------------------
	-- Globals.
	-------------------------------------------------------------------------------
	rs1_index          <= to_integer(unsigned(rs1));
	rs1_even_index     <= to_integer(unsigned(rs1 and "11110"));
	rs1_odd_index      <= to_integer(unsigned(rs1 or  "00001"));
	rs1_pair_index     <= to_integer(unsigned(rs1(4 downto 1)));

	use_rs1_global <= (rs1_index < 8);

	rs2_index      <= to_integer(unsigned(rs2));
	rs2_even_index     <= to_integer(unsigned(rs2 and "11110"));
	rs2_odd_index      <= to_integer(unsigned(rs2 or  "00001"));
	rs2_pair_index     <= to_integer(unsigned(rs2(4 downto 1)));

	use_rs2_global <= (rs2_index < 8);

	read_rd_index  <= to_integer(unsigned(read_rd));
	read_rd_even_index     <= to_integer(unsigned(read_rd and "11110"));
	read_rd_odd_index      <= to_integer(unsigned(read_rd or  "00001"));
	read_rd_pair_index     <= to_integer(unsigned(read_rd(4 downto 1)));

	use_read_rd_global <= (read_rd_index < 8);

	write_rd_index <= to_integer(unsigned(write_rd));
	write_rd_even_index     <= to_integer(unsigned(write_rd and "11110"));
	write_rd_odd_index      <= to_integer(unsigned(write_rd or  "00001"));
	write_rd_pair_index     <= to_integer(unsigned(write_rd(4 downto 1)));

	use_write_rd_global <= (write_rd_index < 8);

	-- bypass the global write to global read..
	g_rs1_index_match <= (rs1_pair_index = write_rd_pair_index);
	g_rs2_index_match <= (rs2_pair_index = write_rd_pair_index);
	g_read_rd_index_match <= (read_rd_pair_index = write_rd_pair_index);

	-- do not bypass to register 0!!
	bypass_global_to_rs1_even     <= use_rs1_global     and  g_rs1_index_match     and (write_gpr_even(0) = '1') and (write_rd_pair_index /= 0);
	bypass_global_to_rs2_even     <= use_rs2_global     and  g_rs2_index_match     and (write_gpr_even(0) = '1') and (write_rd_pair_index /= 0);
	bypass_global_to_read_rd_even <= use_read_rd_global and  g_read_rd_index_match and (write_gpr_even(0) = '1') and (write_rd_pair_index /= 0);

	bypass_global_to_rs1_odd     <= use_rs1_global     and g_rs1_index_match     and (write_gpr_odd(0) = '1');
	bypass_global_to_rs2_odd     <= use_rs2_global     and g_rs2_index_match     and (write_gpr_odd(0) = '1');
	bypass_global_to_read_rd_odd <= use_read_rd_global and g_read_rd_index_match and (write_gpr_odd(0) = '1');

	-------------------------------------------------------------------------------
	-- Mux and Reg.
	-------------------------------------------------------------------------------
	process(clk, reset)
	begin
		if(clk'event and (clk = '1')) then
			if(reset = '1') then
				-- register 0 is always 0!
				global_registers(0) <= (others => '0');
			elsif(trigger) then
				use_rs1_global_reg  <= use_rs1_global;
				use_rs2_global_reg  <= use_rs2_global;
				use_read_rd_global_reg  <= use_read_rd_global;
				use_write_rd_global_reg  <= use_write_rd_global;

				if(use_rs1_global) then 
					if(bypass_global_to_rs1_even) then
						g_rs1_data_reg_even <= write_gpr_value_even;
					else
						g_rs1_data_reg_even <= global_registers(rs1_even_index);
					end if;

					if(bypass_global_to_rs1_odd) then
						g_rs1_data_reg_odd <= write_gpr_value_odd;
					else
						g_rs1_data_reg_odd <= global_registers(rs1_odd_index);
					end if;
				end if;

				if(use_rs2_global) then 
					if(bypass_global_to_rs2_even) then
						g_rs2_data_reg_even <= write_gpr_value_even;
					else
						g_rs2_data_reg_even <= global_registers(rs2_even_index);
					end if;

					if(bypass_global_to_rs2_odd) then
						g_rs2_data_reg_odd <= write_gpr_value_odd;
					else
						g_rs2_data_reg_odd <= global_registers(rs2_odd_index);
					end if;
				end if;

				if(use_read_rd_global) then 
					if(bypass_global_to_read_rd_even) then
						g_read_rd_data_reg_even <= write_gpr_value_even;
					else
						g_read_rd_data_reg_even <= global_registers(read_rd_even_index);
					end if;

					if(bypass_global_to_read_rd_odd) then
						g_read_rd_data_reg_odd <= write_gpr_value_odd;
					else
						g_read_rd_data_reg_odd <= global_registers(read_rd_odd_index);
					end if;
				end if;

				if(use_write_rd_global) then 
					if(write_gpr_even(0) = '1') then
						if(write_rd_even_index /= 0) then
						    global_registers(write_rd_even_index) <= write_gpr_value_even;
						end if;
					end if;
					if(write_gpr_odd(0) = '1') then
						global_registers(write_rd_odd_index)  <= write_gpr_value_odd;
					end if;
				end if;
			end if;
		end if;
	end process;
	
	-------------------------------------------------------------------------------
	-- window bank address calculation
	-------------------------------------------------------------------------------
	rs1_addr_calc:
		window_address_calculator_Volatile
			port map (cwp => read_cwp, reg_id => rs1, reg_address => mem_rs1_read_address);

	rs2_addr_calc:
		window_address_calculator_Volatile
			port map (cwp => read_cwp, reg_id => rs2, reg_address => mem_rs2_read_address);

	read_rd_addr_calc:
		window_address_calculator_Volatile
			port map (cwp => read_cwp, reg_id => read_rd, reg_address => mem_read_rd_read_address);

	write_rd_addr_calc:
		window_address_calculator_Volatile
			port map (cwp => write_cwp, reg_id => write_rd, reg_address => mem_write_rd_write_address);

	-------------------------------------------------------------------------------
	-- window banks: note that write->read bypass is already included in the bank.
	--       also, if global_registers are used, these will not be read from.
	-------------------------------------------------------------------------------
	write_enable_even <= '1' when ((not use_write_rd_global) and (write_gpr_even(0) = '1')) else '0';
	write_enable_odd  <= '1' when ((not use_write_rd_global) and (write_gpr_odd(0)  = '1')) else '0';

	rs1_even_bank: window_registers_bank
				port map (trigger => trigger,
						write_enable_0 => write_enable_even,
						address_0 => mem_write_rd_write_address,
						write_data_0 => write_gpr_value_even,
						address_1 => mem_rs1_read_address,
						read_data_1 => mem_rs1_read_data(63 downto 32),
						clk => clk, reset => reset);

	rs1_odd_bank: window_registers_bank
				port map (trigger => trigger,
						write_enable_0 => write_enable_odd,
						address_0 => mem_write_rd_write_address,
						write_data_0 => write_gpr_value_odd,
						address_1 => mem_rs1_read_address,
						read_data_1 => mem_rs1_read_data(31 downto 0),
						clk => clk, reset => reset);

	rs2_even_bank: window_registers_bank
				port map (trigger => trigger,
						write_enable_0 => write_enable_even,
						address_0 => mem_write_rd_write_address,
						write_data_0 => write_gpr_value_even,
						address_1 => mem_rs2_read_address,
						read_data_1 => mem_rs2_read_data(63 downto 32),
						clk => clk, reset => reset);

	rs2_odd_bank: window_registers_bank
				port map (trigger => trigger,
						write_enable_0 => write_enable_odd,
						address_0 => mem_write_rd_write_address,
						write_data_0 => write_gpr_value_odd,
						address_1 => mem_rs2_read_address,
						read_data_1 => mem_rs2_read_data(31 downto 0),
						clk => clk, reset => reset);
		
	read_rd_even_bank: window_registers_bank
				port map (trigger => trigger,
						write_enable_0 => write_enable_even,
						address_0 => mem_write_rd_write_address,
						write_data_0 => write_gpr_value_even,
						address_1 => mem_read_rd_read_address,
						read_data_1 => mem_read_rd_read_data(63 downto 32),
						clk => clk, reset => reset);

	read_rd_odd_bank: window_registers_bank
				port map (trigger => trigger,
						write_enable_0 => write_enable_odd,
						address_0 => mem_write_rd_write_address,
						write_data_0 => write_gpr_value_odd,
						address_1 => mem_read_rd_read_address,
						read_data_1 => mem_read_rd_read_data(31 downto 0),
						clk => clk, reset => reset);
		
	-------------------------------------------------------------------------------
	-- final muxing between global_registers and window banks.
	-------------------------------------------------------------------------------
    	rs1_pair_value(63 downto 32) <= g_rs1_data_reg_even when use_rs1_global_reg else mem_rs1_read_data (63 downto 32);
    	rs1_pair_value(31 downto 0)  <= g_rs1_data_reg_odd  when use_rs1_global_reg else mem_rs1_read_data (31 downto 0);

    	rs2_pair_value(63 downto 32) <= g_rs2_data_reg_even when use_rs2_global_reg else mem_rs2_read_data (63 downto 32);
    	rs2_pair_value(31 downto 0)  <= g_rs2_data_reg_odd  when use_rs2_global_reg else mem_rs2_read_data (31 downto 0);
			
    	rd_pair_value(63 downto 32)  <= g_read_rd_data_reg_even when use_read_rd_global_reg else mem_read_rd_read_data (63 downto 32);
    	rd_pair_value(31 downto 0)   <= g_read_rd_data_reg_odd  when use_read_rd_global_reg else mem_read_rd_read_data (31 downto 0);

	reg_pair_values <= rs1_pair_value & rs2_pair_value & rd_pair_value;
end iu_registers_3r_1w_port_register_file_inner_arch;

library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.basecomponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
entity iu_registers_3r_1w_port_register_file_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    rs1 : in  std_logic_vector(4 downto 0);
    rs2 : in  std_logic_vector(4 downto 0);
    read_rd : in  std_logic_vector(4 downto 0);
    read_cwp : in  std_logic_vector(4 downto 0);
    write_gpr_even : in  std_logic_vector(0 downto 0);
    write_gpr_odd : in  std_logic_vector(0 downto 0);
    write_rd : in  std_logic_vector(4 downto 0);
    write_gpr_value_even : in  std_logic_vector(31 downto 0);
    write_gpr_value_odd : in  std_logic_vector(31 downto 0);
    write_cwp : in  std_logic_vector(4 downto 0);
    reg_pair_values : out  std_logic_vector(191 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity iu_registers_3r_1w_port_register_file_Operator;
architecture iu_registers_3r_1w_port_register_file_Operator_arch of iu_registers_3r_1w_port_register_file_Operator is -- 
    signal rs1_reg : std_logic_vector(4 downto 0);
    signal rs2_reg : std_logic_vector(4 downto 0);
    signal read_rd_reg : std_logic_vector(4 downto 0);
    signal read_cwp_reg : std_logic_vector(4 downto 0);
    signal write_gpr_even_reg : std_logic_vector(0 downto 0);
    signal write_gpr_odd_reg : std_logic_vector(0 downto 0);
    signal write_rd_reg : std_logic_vector(4 downto 0);
    signal write_gpr_value_even_reg : std_logic_vector(31 downto 0);
    signal write_gpr_value_odd_reg : std_logic_vector(31 downto 0);
    signal write_cwp_reg : std_logic_vector(4 downto 0);

    signal rs1_qual : std_logic_vector(4 downto 0);
    signal rs2_qual : std_logic_vector(4 downto 0);
    signal read_rd_qual : std_logic_vector(4 downto 0);
    signal read_cwp_qual : std_logic_vector(4 downto 0);
    signal write_gpr_even_qual : std_logic_vector(0 downto 0);
    signal write_gpr_odd_qual : std_logic_vector(0 downto 0);
    signal write_rd_qual : std_logic_vector(4 downto 0);
    signal write_gpr_value_even_qual : std_logic_vector(31 downto 0);
    signal write_gpr_value_odd_qual : std_logic_vector(31 downto 0);
    signal write_cwp_qual : std_logic_vector(4 downto 0);

begin --  
	baseInst: iu_registers_3r_1w_port_register_file_inner
		port map (clk => clk, reset => reset,
				sample_req => sample_req, sample_ack => sample_ack,
				update_req => update_req, update_ack => update_ack,
    				rs1 => rs1_qual,
    				rs2 => rs2_qual,
    				read_rd  => read_rd_qual,
    				read_cwp => read_cwp_qual,
    				write_gpr_even => write_gpr_even_qual,
    				write_gpr_odd => write_gpr_odd_qual,
    				write_rd => write_rd_qual,
    				write_gpr_value_even => write_gpr_value_even_qual,
    				write_gpr_value_odd => write_gpr_value_odd_qual,
    				write_cwp => write_cwp_qual,
    				reg_pair_values => reg_pair_values
			);

	process(clk,reset)
	begin
		if(clk'event and (clk = '1')) then
		  if(sample_req) then
			rs1_reg <= rs1;
			rs2_reg <= rs2;
			read_rd_reg <= read_rd;
			read_cwp_reg <= read_cwp;
			write_gpr_even_reg <= write_gpr_even;
			write_gpr_odd_reg <= write_gpr_odd;
    			write_rd_reg <= write_rd;
    			write_gpr_value_even_reg <= write_gpr_value_even;
    			write_gpr_value_odd_reg <= write_gpr_value_odd;
    			write_cwp_reg <= write_cwp;
		  end if;
		end if;
	end process;

	rs1_qual <= rs1 when sample_req else rs1_reg;
	rs2_qual <= rs2 when sample_req else rs2_reg;
	read_rd_qual <= read_rd when sample_req else read_rd_reg;
	read_cwp_qual <= read_cwp when sample_req else read_cwp_reg;
	write_gpr_even_qual <= write_gpr_even when sample_req else write_gpr_even_reg;
	write_gpr_odd_qual <= write_gpr_odd when sample_req else write_gpr_odd_reg;
	write_rd_qual <= write_rd when sample_req else write_rd_reg;
	write_gpr_value_even_qual <= write_gpr_value_even when sample_req else write_gpr_value_even_reg;
	write_gpr_value_odd_qual <= write_gpr_value_odd when sample_req else write_gpr_value_odd_reg;
	write_cwp_qual <= write_cwp when sample_req else write_cwp_reg;
				
end iu_registers_3r_1w_port_register_file_Operator_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
use AjitCustom.UsefulFunctions.all;

entity update_registers_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    next_registers : in  std_logic_vector(1023 downto 0);
    window_update_command : in  std_logic_vector(50 downto 0);
    new_cwp_and_updated_registers : out  std_logic_vector(1028 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity update_registers_Operator;
architecture MpdIsSometimesAKlutz of update_registers_Operator is
	signal start_req, start_ack, fin_req, fin_ack: std_logic;
	
	type FsmState is (IDLE, WINWAIT);
	signal fsm_state : FsmState;

	signal wu_flag : boolean;

	signal wu_save, wu_restore, wu_write_psr: std_logic;
	signal wu_rd, wu_old_cwp, wu_new_cwp: std_logic_vector(4 downto 0);
	signal wu_rd_val: std_logic_vector(31 downto 0);
	
	signal trigger, done_wu, trigger_to_wu, joined_sig: boolean;

	constant ZERO_5: std_logic_vector(4 downto 0) := (others=> '0');

	
   	signal incoming_globals, incoming_outs, incoming_locals, incoming_ins: std_logic_vector(255 downto 0);

   	signal outgoing_globals_reg, outgoing_outs_reg, outgoing_locals_reg, outgoing_ins_reg: std_logic_vector(255 downto 0);
   	signal outgoing_outs_wu, outgoing_locals_wu, outgoing_ins_wu: std_logic_vector(255 downto 0);

   	signal updated_globals: std_logic_vector(255 downto 0);
	signal outgoing_cwp_reg, outgoing_cwp_wu : std_logic_vector(4 downto 0); 

	signal latch_outs_wu, latch_locals_wu, latch_ins_wu, latch_outgoing_cwp_wu: boolean;

	constant z32: std_logic_vector(31 downto 0) := (others => '0');
begin

   
   trig_join: join2 generic map (name => "bpbV2:trig-join", bypass => true)
			port map (pred0 => sample_req, pred1 => update_req,
					symbol_out => trigger, clk => clk, reset => reset);

   wu_flag    <= (window_update_command(50) = '1');
   wu_save    <= window_update_command(49);
   wu_restore <= window_update_command(48);
   wu_write_psr    <= window_update_command(47); 
   wu_rd 	    <= window_update_command(46 downto 42);
   wu_rd_val  <= window_update_command(41 downto 10);
   wu_old_cwp    <= window_update_command(9 downto 5);
   wu_new_cwp    <= window_update_command(4 downto 0);

   incoming_ins <= next_registers(255 downto 0);
   incoming_locals <= next_registers(255+256 downto 256);
   incoming_outs <= next_registers(255+256+256 downto 256+256);
   incoming_globals <= next_registers(255+256+256+256 downto 256+256+256);

   updated_globals <= InsertRdVal(0, wu_save, wu_restore, wu_rd, wu_rd_val, incoming_globals);
	
   core: window_update_core
		port map (
				incoming_outs => incoming_outs,
				incoming_locals => incoming_locals,
				incoming_ins => incoming_ins,
				save      => wu_save, 
				restore   => wu_restore, 
				write_psr => wu_write_psr,
				rd        => wu_rd, 
				rd_val    => wu_rd_val, 
				old_cwp   => wu_old_cwp, 
				new_cwp   => wu_new_cwp,
				outgoing_outs => outgoing_outs_wu, 
				outgoing_locals => outgoing_locals_wu, 
				outgoing_ins => outgoing_ins_wu, 
				outgoing_cwp => outgoing_cwp_wu,
				trigger => trigger_to_wu,
				done => done_wu,
				latch_outs => latch_outs_wu,
				latch_ins => latch_ins_wu,
				latch_locals => latch_locals_wu,
				latch_outgoing_cwp => latch_outgoing_cwp_wu,
				clk => clk,
				reset => reset
			);


   process(clk, reset, fsm_state, 
		wu_flag,
		trigger, 
		done_wu,
		updated_globals, 
		outgoing_outs_wu,
		outgoing_locals_wu, 
		outgoing_ins_wu,
		outgoing_cwp_wu,
		next_registers, 
		latch_outs_wu,
		latch_locals_wu,
		latch_ins_wu,
		latch_outgoing_cwp_wu,
		window_update_command)
	variable next_fsm_state_var: FsmState;
	variable tr_wu_var, sa_var, next_ua_var: boolean;

	variable latch_non_wu_outputs_var:  boolean;
	variable latch_globals_var: boolean;
   begin
	next_fsm_state_var := fsm_state;
	latch_non_wu_outputs_var:= false;
	latch_globals_var := false;

	tr_wu_var := false;
	sa_var := false;
	next_ua_var := false;

	case fsm_state is 
		when IDLE  =>
			if trigger then
				if(wu_flag) then
					next_fsm_state_var := WINWAIT;
					tr_wu_var := true;
					latch_globals_var := true;
				else
					next_fsm_state_var := IDLE;
					next_ua_var   := true;
					sa_var := true;
					latch_non_wu_outputs_var := true;
				end if;
			end if;
		when WINWAIT =>
			if done_wu then
				sa_var := true;
				next_ua_var   := true;
				next_fsm_state_var := IDLE;
			end if;
	end case;

	sample_ack <= sa_var;
	trigger_to_wu <= tr_wu_var;

	if(clk'event and clk = '1') then
		if(reset = '1') then
			update_ack <= false;
			fsm_state <= IDLE;
		else
			update_ack <= next_ua_var;
			fsm_state <= next_fsm_state_var;
		end if;

		if(wu_flag and latch_outs_wu) then
			outgoing_outs_reg <= outgoing_outs_wu;
		end if;

		if(wu_flag and latch_locals_wu) then
			outgoing_locals_reg <= outgoing_locals_wu;
		end if;

		if(wu_flag and latch_ins_wu) then
			outgoing_ins_reg <= outgoing_ins_wu;
		end if;

		if(wu_flag and latch_outgoing_cwp_wu) then
			outgoing_cwp_reg <= outgoing_cwp_wu;
		end if;

		if(wu_flag and latch_globals_var) then
			outgoing_globals_reg <= updated_globals;
		end if;

		if(latch_non_wu_outputs_var) then

			outgoing_globals_reg <= incoming_globals;
			outgoing_outs_reg   <= incoming_outs;
			outgoing_locals_reg <= incoming_locals;
			outgoing_ins_reg    <= incoming_ins;
			outgoing_cwp_reg    <= ZERO_5;

		end if;
	end if;
   end process;

   
   new_cwp_and_updated_registers <= (outgoing_cwp_reg & z32 & outgoing_globals_reg((255-32) downto 0)  & outgoing_outs_reg & outgoing_locals_reg & outgoing_ins_reg);
    
end MpdIsSometimesAKlutz;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;

entity window_address_calculator_Volatile is -- 
  port ( -- 
    cwp : in  std_logic_vector(4 downto 0);
    reg_id : in  std_logic_vector(4 downto 0);
    reg_address : out  std_logic_vector(5 downto 0)-- 
  );
  -- 
end entity window_address_calculator_Volatile;
architecture window_address_calculator_Volatile_arch of window_address_calculator_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(10-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal cwp_buffer :  std_logic_vector(4 downto 0);
  signal reg_id_buffer :  std_logic_vector(4 downto 0);
  -- output port buffer signals
  signal reg_address_buffer :  std_logic_vector(5 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  cwp_buffer <= cwp;
  reg_id_buffer <= reg_id;
  -- output handling  -------------------------------------------------------
  reg_address <= reg_address_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal ADD_u5_u5_25_wire : std_logic_vector(4 downto 0);
    signal SUB_u5_u5_38_wire : std_logic_vector(4 downto 0);
    signal ULT_u5_u1_75_wire : std_logic_vector(0 downto 0);
    signal cwp_6_19 : std_logic_vector(5 downto 0);
    signal incr_cwp_6_28 : std_logic_vector(5 downto 0);
    signal ireg_addr_71 : std_logic_vector(5 downto 0);
    signal ireg_base_61 : std_logic_vector(5 downto 0);
    signal ireg_offset_66 : std_logic_vector(5 downto 0);
    signal konst_24_wire_constant : std_logic_vector(4 downto 0);
    signal konst_37_wire_constant : std_logic_vector(4 downto 0);
    signal konst_44_wire_constant : std_logic_vector(5 downto 0);
    signal konst_49_wire_constant : std_logic_vector(5 downto 0);
    signal konst_59_wire_constant : std_logic_vector(5 downto 0);
    signal konst_64_wire_constant : std_logic_vector(5 downto 0);
    signal konst_74_wire_constant : std_logic_vector(4 downto 0);
    signal oreg_local_addr_56 : std_logic_vector(5 downto 0);
    signal oreg_local_base_46 : std_logic_vector(5 downto 0);
    signal oreg_local_offset_51 : std_logic_vector(5 downto 0);
    signal reg_pair_id_6_34 : std_logic_vector(5 downto 0);
    signal reg_pair_id_minus_16_6_41 : std_logic_vector(5 downto 0);
    signal slice_17_wire : std_logic_vector(2 downto 0);
    signal slice_26_wire : std_logic_vector(2 downto 0);
    signal slice_32_wire : std_logic_vector(3 downto 0);
    signal slice_39_wire : std_logic_vector(3 downto 0);
    signal type_cast_15_wire_constant : std_logic_vector(2 downto 0);
    signal type_cast_22_wire_constant : std_logic_vector(2 downto 0);
    -- 
  begin -- 
    konst_24_wire_constant <= "00001";
    konst_37_wire_constant <= "10000";
    konst_44_wire_constant <= "000011";
    konst_49_wire_constant <= "000100";
    konst_59_wire_constant <= "000011";
    konst_64_wire_constant <= "000100";
    konst_74_wire_constant <= "11000";
    type_cast_15_wire_constant <= "000";
    type_cast_22_wire_constant <= "000";
    -- flow-through select operator MUX_79_inst
    reg_address_buffer <= oreg_local_addr_56 when (ULT_u5_u1_75_wire(0) /=  '0') else ireg_addr_71;
    -- flow-through slice operator slice_17_inst
    slice_17_wire <= cwp_buffer(2 downto 0);
    -- flow-through slice operator slice_26_inst
    slice_26_wire <= ADD_u5_u5_25_wire(2 downto 0);
    -- flow-through slice operator slice_32_inst
    slice_32_wire <= reg_id_buffer(4 downto 1);
    -- flow-through slice operator slice_39_inst
    slice_39_wire <= SUB_u5_u5_38_wire(4 downto 1);
    -- interlock type_cast_33_inst
    process(slice_32_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 3 downto 0) := slice_32_wire(3 downto 0);
      reg_pair_id_6_34 <= tmp_var; -- 
    end process;
    -- interlock type_cast_40_inst
    process(slice_39_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 3 downto 0) := slice_39_wire(3 downto 0);
      reg_pair_id_minus_16_6_41 <= tmp_var; -- 
    end process;
    -- binary operator ADD_u5_u5_25_inst
    process(cwp_buffer) -- 
      variable tmp_var : std_logic_vector(4 downto 0); -- 
    begin -- 
      ApIntAdd_proc(cwp_buffer, konst_24_wire_constant, tmp_var);
      ADD_u5_u5_25_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u6_u6_55_inst
    process(oreg_local_base_46, oreg_local_offset_51) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(oreg_local_base_46, oreg_local_offset_51, tmp_var);
      oreg_local_addr_56 <= tmp_var; --
    end process;
    -- binary operator ADD_u6_u6_70_inst
    process(ireg_base_61, ireg_offset_66) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(ireg_base_61, ireg_offset_66, tmp_var);
      ireg_addr_71 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u3_u6_18_inst
    process(type_cast_15_wire_constant, slice_17_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_15_wire_constant, slice_17_wire, tmp_var);
      cwp_6_19 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u3_u6_27_inst
    process(type_cast_22_wire_constant, slice_26_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_22_wire_constant, slice_26_wire, tmp_var);
      incr_cwp_6_28 <= tmp_var; --
    end process;
    -- binary operator SHL_u6_u6_45_inst
    process(cwp_6_19) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntSHL_proc(cwp_6_19, konst_44_wire_constant, tmp_var);
      oreg_local_base_46 <= tmp_var; --
    end process;
    -- binary operator SHL_u6_u6_60_inst
    process(incr_cwp_6_28) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntSHL_proc(incr_cwp_6_28, konst_59_wire_constant, tmp_var);
      ireg_base_61 <= tmp_var; --
    end process;
    -- binary operator SUB_u5_u5_38_inst
    process(reg_id_buffer) -- 
      variable tmp_var : std_logic_vector(4 downto 0); -- 
    begin -- 
      ApIntSub_proc(reg_id_buffer, konst_37_wire_constant, tmp_var);
      SUB_u5_u5_38_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u6_u6_50_inst
    process(reg_pair_id_6_34) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntSub_proc(reg_pair_id_6_34, konst_49_wire_constant, tmp_var);
      oreg_local_offset_51 <= tmp_var; --
    end process;
    -- binary operator SUB_u6_u6_65_inst
    process(reg_pair_id_minus_16_6_41) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntSub_proc(reg_pair_id_minus_16_6_41, konst_64_wire_constant, tmp_var);
      ireg_offset_66 <= tmp_var; --
    end process;
    -- binary operator ULT_u5_u1_75_inst
    process(reg_id_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(reg_id_buffer, konst_74_wire_constant, tmp_var);
      ULT_u5_u1_75_wire <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end window_address_calculator_Volatile_arch;

library std;
use std.standard.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.mem_component_pack.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;

library AjitCustom;
use AjitCustom.UsefulFunctions.all;

entity window_update_core is -- 
  port ( -- 
    incoming_outs, incoming_locals, incoming_ins : in  std_logic_vector(255 downto 0);
    save, restore, write_psr: in std_logic;
    rd: in std_logic_vector(4 downto 0);
    rd_val: in std_logic_vector(31 downto 0);
    old_cwp, new_cwp : in std_logic_vector(4 downto 0);
    outgoing_outs, outgoing_locals, outgoing_ins : out  std_logic_vector(255 downto 0);
    outgoing_cwp : out std_logic_vector(4 downto 0);
    clk : in std_logic;
    reset : in std_logic;
    trigger : in boolean;
    done    : out boolean;
    latch_locals, latch_outs, latch_ins, latch_outgoing_cwp: out boolean
  );
  -- 
end entity window_update_core;

architecture MpdIsWhatCanISay of window_update_core is -- 
	type FsmState is (IdleState, FirstAccessState, SecondAccessState, ResponseDoneState);
	signal fsm_state: FsmState;
		

	signal rd_wp_reg, old_cwp_reg: std_logic_vector (4 downto 0);

	constant NWINDOWS_MOD_MASK_5  : std_logic_vector(4 downto 0) := "00111";
	constant uNWINDOWSx16_MOD_MASK_16: unsigned(15 downto 0) := "0000000001111111";
					
	constant const_one_1: std_logic_vector(0 downto 0) := "1";
						

	function DecrementStdLogicVector (X: std_logic_vector)
			return std_logic_vector is
		alias lx : std_logic_vector(1 to X'length) is X;
		variable ret_val : std_logic_vector(1 to X'length);
		variable lx_u, ret_val_u : unsigned (1 to X'length);
	begin
		lx_u := unsigned(lx);
		ret_val_u := lx_u - 1;
		ret_val := std_logic_vector(ret_val_u);
		return(ret_val);
	end function DecrementStdLogicVector;
	function IncrementStdLogicVector (X: std_logic_vector)
			return std_logic_vector is
		alias lx : std_logic_vector(1 to X'length) is X;
		variable ret_val : std_logic_vector(1 to X'length);
		variable lx_u, ret_val_u : unsigned (1 to X'length);
	begin
		lx_u := unsigned(lx);
		ret_val_u := lx_u + 1;
		ret_val := std_logic_vector(ret_val_u);
		return(ret_val);
	end function IncrementStdLogicVector;
	
	function RegBlockAddress(offset: integer; cwp: std_logic_vector(4 downto 0))
		return std_logic_vector is
		variable ret_val : std_logic_vector(3 downto 0);
		variable cwp_u : unsigned(4 downto 0);
		variable cwp_16 : unsigned (15 downto 0);
	begin
		cwp_u := unsigned (cwp);

		cwp_16 := resize(cwp_u, 16);
		cwp_16 := shift_right(((shift_left(cwp_16, 4) + offset) and uNWINDOWSx16_MOD_MASK_16), 3);
		ret_val := std_logic_vector(cwp_16(3 downto 0));

		return(ret_val);
	end function RegBlockAddress;


	signal dpmem_address_0 : std_logic_vector( 3 downto 0);
	signal dpmem_write_data_0, dpmem_read_data_0 : std_logic_vector (255 downto 0);
	signal dpmem_enable_0 : std_logic;
	signal dpmem_read_writebar_0 : std_logic;

	signal dpmem_address_1: std_logic_vector(3 downto 0);
	signal dpmem_write_data_1, dpmem_read_data_1: std_logic_vector(255 downto 0);
	signal dpmem_enable_1: std_logic;
	signal dpmem_read_writebar_1 : std_logic;
		
	signal address_0_reg, address_1_reg : std_logic_vector(3 downto 0);
    
	-- tried hard to eliminate these registers, but too complicated..
	signal incoming_outs_reg, incoming_locals_reg, incoming_ins_reg : std_logic_vector(255 downto 0);
    	signal save_reg, restore_reg, write_psr_reg: std_logic;
    	signal rd_reg: std_logic_vector(4 downto 0);
    	signal rd_val_reg: std_logic_vector(31 downto 0);

	constant OUTS_OFFSET:    integer := 8;
	constant LOCALS_OFFSET:  integer := 16;
	constant INS_OFFSET:     integer := 24;


-- see comment above..
--##decl_synopsys_sync_set_reset##
begin --  
	process(clk,reset,
		fsm_state, 
		trigger,
		rd_wp_reg, 
		save, restore,
		old_cwp, new_cwp,
		dpmem_read_data_0, dpmem_read_data_1,
		incoming_locals, rd, rd_val,
		incoming_outs, incoming_ins,
		address_0_reg, address_1_reg)
		
		variable next_fsm_state: FsmState;	
		variable done_var: boolean;

		variable cycle_count_var: std_logic_vector (15 downto 0);
		variable outgoing_outs_var, outgoing_locals_var, outgoing_ins_var: 
								std_logic_vector(255 downto 0);

		variable latch_rd_wp_var: boolean;

		-- windows memory is 32x256 dpram
		variable address_0_var, address_1_var : std_logic_vector(3 downto 0);
		variable enable_0_var, enable_1_var: std_logic;
		variable read_writebar_0_var, read_writebar_1_var: std_logic;

		variable write_data_0_var : std_logic_vector(255 downto 0);
		variable write_data_1_var : std_logic_vector(255 downto 0);

		variable rd_wp_var, outgoing_cwp_var  : std_logic_vector(4 downto 0);
		variable latch_ins_var, latch_outs_var, latch_locals_var, latch_outgoing_cwp_var : boolean;

		variable latch_incomings_var: boolean;
		
	begin
		outgoing_cwp_var := (others => '0');

		latch_outs_var := false;
		latch_locals_var := false;
		latch_ins_var := false;
		latch_outgoing_cwp_var := false;

		latch_incomings_var := false;

		latch_rd_wp_var := false;
		done_var := false;

		enable_0_var := '0';
		enable_1_var := '0';

		read_writebar_0_var := '0';
		read_writebar_1_var := '0';

		address_0_var := (others => '0');
		address_1_var := (others => '0');

		write_data_0_var := (others => '0');
		write_data_1_var := (others => '0');
	
		rd_wp_var := (others => '0');


								
		next_fsm_state := fsm_state;
		
		outgoing_outs_var   :=  (others => '0');
		outgoing_locals_var    :=  (others => '0');
		outgoing_ins_var    :=  (others => '0');
		
		-- Cycle 1:  
		--    If save
		--        new_ins <- old_outs, read-locals, read-outs... 
		--    If restore
		--        new_outs <- old_ins, read-locals, read-ins... 
		--    If write-psr
		--        write-outs, write-ins, 
				-- register incoming outs, locals, ins.

		-- Cycle 2: 
		--    If save/restore
		--        write-locals, write-ins.
		--    If write-psr
		--        write-locals, read-locals.
		-- 
		-- Cycle 3:  
		--     If save/restore
		--        write-outs.
		--     If write-psr
		--        latch-locals,  read-outs, read-ins.
		case fsm_state is
			when IdleState =>
				if trigger then
					next_fsm_state := FirstAccessState;
					latch_incomings_var := true;

					if(save = '1') then
						rd_wp_var := DecrementStdLogicVector(old_cwp) and
								NWINDOWS_MOD_MASK_5;
					elsif (restore = '1') then
						rd_wp_var := IncrementStdLogicVector(old_cwp) and
								NWINDOWS_MOD_MASK_5;
					else
						rd_wp_var := new_cwp and NWINDOWS_MOD_MASK_5;
					end if;

					latch_outgoing_cwp_var := true;
					outgoing_cwp_var := rd_wp_var;

					if ((save = '1') or (restore = '1')) then
						-- read new locals on port 0
						address_0_var  := RegBlockAddress(8, rd_wp_var);
						enable_0_var   := '1';
						read_writebar_0_var  := '1';
						next_fsm_state := SecondAccessState;


						if (save = '1') then
							-- read new outs on port 1
							address_1_var := RegBlockAddress(0, rd_wp_var);
							enable_1_var  := '1';
							read_writebar_1_var  := '1';
	
							outgoing_ins_var := InsertRdVal(INS_OFFSET, save, restore, rd, rd_val, incoming_outs);
							latch_ins_var := true;
						end if;

						if (restore = '1') then
							-- read new ins on port 1
							address_1_var := RegBlockAddress(16, rd_wp_var);
							enable_1_var  := '1';
							read_writebar_1_var  := '1';
	
							outgoing_outs_var := InsertRdVal(OUTS_OFFSET, save, restore, rd, rd_val, incoming_ins);
							latch_outs_var := true;
						end if;
					else -- (write_psr = '1')

						-- write outs on port 0
						address_0_var := RegBlockAddress(0, old_cwp);
						write_data_0_var    := incoming_outs;
						enable_0_var  := '1';
						read_writebar_0_var  := '0';

						-- write ins on port 1
						address_1_var := RegBlockAddress(16, old_cwp);
						write_data_1_var    := incoming_ins;
						enable_1_var  := '1';
						read_writebar_1_var  := '0';
					end if;

					latch_rd_wp_var  := true;
					next_fsm_state :=  FirstAccessState;

				   end if;
			when FirstAccessState =>

				outgoing_cwp_var := rd_wp_reg;
				if((save_reg = '1') or (restore_reg = '1')) then

					-- initiated in previous cycle, available
					-- now on port 0.
					outgoing_locals_var := InsertRdVal(LOCALS_OFFSET, save_reg, restore_reg, rd_reg, rd_val_reg, dpmem_read_data_0);
					-- indicate that locals should be latched.
					latch_locals_var := true;


					-- write old locals on port 0.
					address_0_var := RegBlockAddress(8, old_cwp_reg);
					write_data_0_var    := incoming_locals_reg;
					enable_0_var  := '1';
					read_writebar_0_var  := '0';

					

					-- write old ins on port 1.
					address_1_var := RegBlockAddress(16, old_cwp_reg);
					write_data_1_var    := incoming_ins_reg;
					enable_1_var  := '1';
					read_writebar_1_var  := '0';

					if(save_reg = '1') then
						-- outs available on port 1.
						outgoing_outs_var := InsertRdVal(OUTS_OFFSET, save_reg, restore_reg, rd_reg, rd_val_reg, dpmem_read_data_1);
						latch_outs_var := true;
					end if;

					if(restore_reg = '1') then
						-- ins available on port 1
						outgoing_ins_var := InsertRdVal(INS_OFFSET, save_reg, restore_reg, rd_reg, rd_val_reg, dpmem_read_data_1);
						latch_ins_var := true;
					end if;

					-- done... move on.
					done_var := true;

				else -- (write_psr_reg = '1')

					-- read new locals on port 0
					address_0_var  := RegBlockAddress(8, rd_wp_reg);
					enable_0_var   := '1';
					read_writebar_0_var  := '1';
						
					-- write old locals on port 1
					address_1_var := RegBlockAddress(8, old_cwp_reg);
					write_data_1_var    := incoming_locals_reg;
					enable_1_var  := '1';
					read_writebar_1_var  := '0';
				
					next_fsm_state :=  SecondAccessState;
				end if;
					
				next_fsm_state :=  SecondAccessState;


			when SecondAccessState =>

				outgoing_cwp_var := rd_wp_reg;
				if((save_reg = '1') or (restore_reg = '1')) then
					-- write old outs on port 1
					address_1_var := RegBlockAddress(0, old_cwp_reg);
					write_data_1_var    := incoming_outs_reg;
					enable_1_var  := '1';
					read_writebar_1_var  := '0';


					next_fsm_state := IdleState;

				else -- (write_psr_reg = '1') 
					-- read new outs on port 0
					address_0_var := RegBlockAddress(0, rd_wp_reg);
					enable_0_var  := '1';
					read_writebar_0_var  := '1';

					-- read new ins on port 1
					address_1_var := RegBlockAddress(16, rd_wp_reg);
					enable_1_var  := '1';
					read_writebar_1_var  := '1';
	
					-- locals are available on port 0.
					latch_locals_var  := true;
					outgoing_locals_var := InsertRdVal(LOCALS_OFFSET, save_reg, restore_reg, rd_reg, rd_val_reg, dpmem_read_data_0);

					next_fsm_state :=  ResponseDoneState;

				end if;
			when ResponseDoneState =>

				outgoing_cwp_var := rd_wp_reg;
				done_var := true;

				-- outs available on port 0.
				outgoing_outs_var := InsertRdVal(OUTS_OFFSET, save_reg, restore_reg, rd_reg, rd_val_reg, dpmem_read_data_0);
				latch_outs_var := true;

				-- ins available on port 1.	
				outgoing_ins_var := InsertRdVal(INS_OFFSET, save_reg, restore_reg, rd_reg, rd_val_reg, dpmem_read_data_1);
				latch_ins_var := true;

				next_fsm_state := IdleState;
		end case;

		done <= done_var;

		latch_locals <= latch_locals_var;
		latch_outs   <= latch_outs_var;
		latch_ins   <= latch_ins_var;
		latch_outgoing_cwp <= latch_outgoing_cwp_var;
		outgoing_cwp <= outgoing_cwp_var;
		
		dpmem_address_0 <= address_0_var;
		dpmem_write_data_0 <= write_data_0_var;
		dpmem_enable_0 <= enable_0_var;
		dpmem_read_writebar_0 <= read_writebar_0_var;

		dpmem_address_1 <= address_1_var;
		dpmem_write_data_1 <= write_data_1_var;
		dpmem_enable_1 <= enable_1_var;
		dpmem_read_writebar_1 <= read_writebar_1_var;

		outgoing_outs   <= outgoing_outs_var;
		outgoing_locals <= outgoing_locals_var;
		outgoing_ins    <= outgoing_ins_var;

		if(clk'event and clk = '1') then
			if(reset = '1') then
				fsm_state <= IdleState;
			else
				fsm_state <= next_fsm_state;
				if(latch_rd_wp_var) then
					rd_wp_reg <= rd_wp_var;
				end if;
				if(latch_incomings_var) then

					incoming_outs_reg <= incoming_outs;
					incoming_locals_reg <= incoming_locals;
					incoming_ins_reg <= incoming_ins;
					old_cwp_reg <= old_cwp;

					save_reg <= save;
					restore_reg <= restore;
					write_psr_reg <= write_psr;
					rd_reg <= rd;
					rd_val_reg <= rd_val;

				end if;
			end if;
		end if;
	end process;

	dpmem: base_bank_dual_port
			generic map (name => "window_update_daemon:dpmem",
					g_addr_width => 4,
					g_data_width => 256)
			port map ( datain_0 => dpmem_write_data_0,
					dataout_0 => dpmem_read_data_0,
					enable_0 => dpmem_enable_0,
					writebar_0 => dpmem_read_writebar_0,
					addrin_0 => dpmem_address_0, 
					datain_1 => dpmem_write_data_1,
					dataout_1 => dpmem_read_data_1,
					enable_1 => dpmem_enable_1,
					writebar_1 => dpmem_read_writebar_1,
					addrin_1 => dpmem_address_1, 
					clk => clk, reset => reset);

end MpdIsWhatCanISay;

library std;
use std.standard.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.mem_component_pack.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;

entity window_update_daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    iunit_register_file_window_update_command_pipe_read_req : out  std_logic_vector(0 downto 0);
    iunit_register_file_window_update_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
    iunit_register_file_window_update_command_pipe_read_data : in   std_logic_vector(1090 downto 0);
    iunit_register_file_window_update_response_pipe_write_req : out  std_logic_vector(0 downto 0);
    iunit_register_file_window_update_response_pipe_write_ack : in   std_logic_vector(0 downto 0);
    iunit_register_file_window_update_response_pipe_write_data : out  std_logic_vector(1045 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity window_update_daemon;
architecture window_update_daemon_arch of window_update_daemon is -- 
	type FsmState is (IdleState, FirstAccessState, SecondAccessState, WaitResponsePipeState);
	signal fsm_state: FsmState;
		
	signal cycle_count_reg: std_logic_vector (15 downto 0);
	signal wr_wp_reg: std_logic_vector (4 downto 0);
	signal globals_reg, outs_reg, locals_reg, ins_reg: std_logic_vector(255 downto 0);
	signal fetched_locals_reg: std_logic_vector(255 downto 0);
	signal new_globals, new_outs, new_locals, new_ins: std_logic_vector(255 downto 0);
	signal write_psr_reg, save_reg, restore_reg: std_logic;
	signal rd_reg: std_logic_vector (4 downto 0);
	signal rd_val_reg: std_logic_vector (31 downto 0);
	signal valid_reg: std_logic;
									
	signal rd_wp_reg: std_logic_vector (4 downto 0);

	constant NWINDOWS_MOD_MASK_5  : std_logic_vector(4 downto 0) := "00111";
	constant uNWINDOWSx16_MOD_MASK_16: unsigned(15 downto 0) := "0000000001111111";
					
	constant const_one_1: std_logic_vector(0 downto 0) := "1";
						

	function DecrementStdLogicVector (X: std_logic_vector)
			return std_logic_vector is
		alias lx : std_logic_vector(1 to X'length) is X;
		variable ret_val : std_logic_vector(1 to X'length);
		variable lx_u, ret_val_u : unsigned (1 to X'length);
	begin
		lx_u := unsigned(lx);
		ret_val_u := lx_u - 1;
		ret_val := std_logic_vector(ret_val_u);
		return(ret_val);
	end function DecrementStdLogicVector;
	function IncrementStdLogicVector (X: std_logic_vector)
			return std_logic_vector is
		alias lx : std_logic_vector(1 to X'length) is X;
		variable ret_val : std_logic_vector(1 to X'length);
		variable lx_u, ret_val_u : unsigned (1 to X'length);
	begin
		lx_u := unsigned(lx);
		ret_val_u := lx_u + 1;
		ret_val := std_logic_vector(ret_val_u);
		return(ret_val);
	end function IncrementStdLogicVector;
	
	function RegBlockAddress(offset: integer; cwp: std_logic_vector(4 downto 0))
		return std_logic_vector is
		variable ret_val : std_logic_vector(4 downto 0);
		variable cwp_u : unsigned(4 downto 0);
		variable cwp_16 : unsigned (15 downto 0);
	begin
		cwp_u := unsigned (cwp);

		cwp_16 := resize(cwp_u, 16);
		cwp_16 := shift_right(((shift_left(cwp_16, 4) + offset) and uNWINDOWSx16_MOD_MASK_16), 3);
		ret_val := std_logic_vector(cwp_16(4 downto 0));

		return(ret_val);
	end function RegBlockAddress;

	function InsertRdVal(offset: integer; save, restore : std_logic;
						rd: std_logic_vector(4 downto 0);
						rd_val: std_logic_vector(31 downto 0);
						reg_256: std_logic_vector(255 downto 0))
		return std_logic_vector is
		variable ret_val : std_logic_vector(255 downto 0);
		variable wr_val : std_logic_vector(31 downto 0);
		variable w0,w1,w2,w3,w4,w5,w6,w7: std_logic_vector(31 downto 0);

		variable reg_index : integer range 0 to 31;
	begin
		w7 := reg_256 (31 downto 0);
		w6 := reg_256 (63 downto 32);
		w5 := reg_256 (95 downto 64);
		w4 := reg_256 (127 downto 96);
		w3 := reg_256 (159 downto 128);
		w2 := reg_256 (191 downto 160);
		w1 := reg_256 (223 downto 192);
		w0 := reg_256 (255 downto 224);

		reg_index := to_integer(unsigned(rd));

		-- register 0 always contains 0.
		if(reg_index = 0) then
			wr_val := (others => '0');
		else
			wr_val := rd_val;
		end if;

		if(((save = '1')  or (restore = '1')) and (reg_index >= offset)) then
			
			reg_index := reg_index - offset;

			if(reg_index < 8) then

				
				if (reg_index = 0) then
					w0 := wr_val;
				elsif reg_index = 1 then
					w1 := wr_val;
				elsif reg_index = 2 then
					w2 := wr_val;
				elsif reg_index = 3 then
					w3 := wr_val;
				elsif reg_index = 4 then
					w4 := wr_val;
				elsif reg_index = 5 then
					w5 := wr_val;
				elsif reg_index = 6 then
					w6 := wr_val;
				elsif reg_index = 7 then
					w7 := wr_val;
				end if;
			end if;
		end if;

		ret_val := w0 & w1 & w2 & w3 & w4 & w5 & w6 & w7;
		return(ret_val);
	end function InsertRdVal;

	signal dpmem_address_0 : std_logic_vector( 4 downto 0);
	signal dpmem_write_data_0, dpmem_read_data_0 : std_logic_vector (255 downto 0);
	signal dpmem_enable_0 : std_logic;
	signal dpmem_read_writebar_0 : std_logic;

	signal dpmem_address_1: std_logic_vector(4 downto 0);
	signal dpmem_write_data_1, dpmem_read_data_1: std_logic_vector(255 downto 0);
	signal dpmem_enable_1: std_logic;
	signal dpmem_read_writebar_1 : std_logic;
		
	signal cycle_count: std_logic_vector (15 downto 0);
	signal oldcwp: std_logic_vector (4 downto 0);
	signal oldcwp_reg: std_logic_vector (4 downto 0);
	signal newcwp: std_logic_vector (4 downto 0);
	signal newcwp_reg: std_logic_vector (4 downto 0);
		
	signal address_0_reg, address_1_reg : std_logic_vector(4 downto 0);
-- see comment above..
--##decl_synopsys_sync_set_reset##
begin --  

	start_ack <= '1';
	fin_ack <= '0';

	process(clk,reset,
		fsm_state, 
		iunit_register_file_window_update_command_pipe_read_ack,
		iunit_register_file_window_update_response_pipe_write_ack,
		iunit_register_file_window_update_command_pipe_read_data,
		rd_wp_reg, wr_wp_reg, save_reg, restore_reg,
		oldcwp_reg, newcwp_reg,
		globals_reg, dpmem_read_data_0, dpmem_read_data_1, fetched_locals_reg,
		locals_reg, rd_reg, rd_val_reg,
		outs_reg, ins_reg,
		address_0_reg, address_1_reg)
		
		variable next_fsm_state: FsmState;	
		variable read_req_var, write_req_var: std_logic;

		variable cycle_count_var: std_logic_vector (15 downto 0);
		variable oldcwp_var: std_logic_vector (4 downto 0);
		variable newcwp_var: std_logic_vector (4 downto 0);
		variable globals_var, outs_var, locals_var, ins_var: std_logic_vector(255 downto 0);
		variable new_globals_var, new_outs_var, new_locals_var, new_ins_var: 
								std_logic_vector(255 downto 0);
		variable write_psr_var, save_var, restore_var: std_logic;
		variable rd_var: std_logic_vector (4 downto 0);
		variable rd_val_var: std_logic_vector (31 downto 0);
		variable valid_var: std_logic;

		variable latch_inputs_var: boolean;
		variable latch_rd_wp_var: boolean;

		variable latch_fetched_locals_var: boolean;
		variable latch_new_window_regs_var: boolean;

		-- windows memory is 32x256 dpram
		variable address_0_var, address_1_var : std_logic_vector(4 downto 0);
		variable enable_0_var, enable_1_var: std_logic;
		variable read_writebar_0_var, read_writebar_1_var: std_logic;

		variable write_data_0_var : std_logic_vector(255 downto 0);
		variable write_data_1_var : std_logic_vector(255 downto 0);

		variable rd_wp_var  : std_logic_vector(4 downto 0);
		variable latch_addresses_var : boolean;
	begin

		latch_addresses_var := false;

		latch_inputs_var := false;
		latch_rd_wp_var := false;
		latch_fetched_locals_var := false;
		latch_new_window_regs_var := false;

		enable_0_var := '0';
		enable_1_var := '0';

		read_writebar_0_var := '0';
		read_writebar_1_var := '0';

		address_0_var := (others => '0');
		address_1_var := (others => '0');

		write_data_0_var := (others => '0');
		write_data_1_var := (others => '0');
	
		rd_wp_var := (others => '0');

		valid_var   := iunit_register_file_window_update_command_pipe_read_data(0);
		rd_val_var  := iunit_register_file_window_update_command_pipe_read_data(32 downto 1);
		rd_var 	    := iunit_register_file_window_update_command_pipe_read_data(37 downto 33);
		restore_var := iunit_register_file_window_update_command_pipe_read_data(38);
		save_var    := iunit_register_file_window_update_command_pipe_read_data(39);
		write_psr_var    := iunit_register_file_window_update_command_pipe_read_data(40);
		--variable globals_var, outs_var, locals_vr, ins_var: std_logic_vector(255 downto 0);
		ins_var    := iunit_register_file_window_update_command_pipe_read_data(296 downto 41);
		locals_var    := iunit_register_file_window_update_command_pipe_read_data(552 downto 297);
		outs_var    := iunit_register_file_window_update_command_pipe_read_data(808 downto 553);
		globals_var    := iunit_register_file_window_update_command_pipe_read_data(1064 downto 809);
		newcwp_var    := iunit_register_file_window_update_command_pipe_read_data(1069 downto 1065);
		oldcwp_var    := iunit_register_file_window_update_command_pipe_read_data(1074 downto 1070);
		cycle_count_var  := iunit_register_file_window_update_command_pipe_read_data(1090 downto 1075);

		cycle_count <= cycle_count_var;
		oldcwp <= oldcwp_var;
		newcwp <= newcwp_var;

		
								
		next_fsm_state := fsm_state;
		read_req_var := '0';
		write_req_var := '0';
		
		new_globals_var := InsertRdVal(0, save_reg, restore_reg,
								rd_reg, rd_val_reg, 
									globals_reg);
		new_outs_var := InsertRdVal(8, save_reg, restore_reg,
								rd_reg, rd_val_reg, 
									dpmem_read_data_0);
		new_locals_var := InsertRdVal(16,save_reg,restore_reg,
								rd_reg, rd_val_reg, 
									fetched_locals_reg);
		new_ins_var := InsertRdVal(24, save_reg, restore_reg,
								rd_reg, rd_val_reg, 
											dpmem_read_data_1);
		case fsm_state is
			when IdleState =>
				read_req_var := '1';
				if(iunit_register_file_window_update_command_pipe_read_ack(0) = '1') then
				   if(valid_var = '1') then
					latch_inputs_var := true;
					next_fsm_state := FirstAccessState;
					
					if(save_var = '1') then
						rd_wp_var := DecrementStdLogicVector(oldcwp_var) and
								NWINDOWS_MOD_MASK_5;
					elsif (restore_var = '1') then
						rd_wp_var := IncrementStdLogicVector(oldcwp_var) and
								NWINDOWS_MOD_MASK_5;
					else
						rd_wp_var := newcwp_var and NWINDOWS_MOD_MASK_5;
					end if;

					-- write outs
					address_0_var := RegBlockAddress(0, oldcwp_var);
					write_data_0_var    := outs_var;
					enable_0_var  := '1';
					read_writebar_0_var  := '0';
	
					-- write ins.
					address_1_var := RegBlockAddress(16, oldcwp_var);
					write_data_1_var    := ins_var;
					enable_1_var  := '1';
					read_writebar_1_var  := '0';
	
					latch_rd_wp_var  := true;
					next_fsm_state :=  FirstAccessState;
				  end if;
				end if;
			when FirstAccessState =>
				-- write old locals
				address_0_var := RegBlockAddress(8, wr_wp_reg);
				write_data_0_var    := locals_reg;
				enable_0_var  := '1';
				read_writebar_0_var  := '0';

				-- read new locals
				address_1_var  := RegBlockAddress(8, rd_wp_reg);
				enable_1_var   := '1';
				read_writebar_1_var  := '1';

				next_fsm_state :=  SecondAccessState;

			when SecondAccessState =>

				-- read new outs
				address_0_var := RegBlockAddress(0, rd_wp_reg);
				enable_0_var  := '1';
				read_writebar_0_var  := '1';

				-- read new ins
				address_1_var := RegBlockAddress(16, rd_wp_reg);
				enable_1_var  := '1';
				read_writebar_1_var  := '1';


				next_fsm_state :=  WaitResponsePipeState;

				latch_fetched_locals_var  := true;
				latch_addresses_var := true;

			when WaitResponsePipeState =>
	
				-- continue presenting latched addresses so that
				-- dpmem outputs are held stable
				address_0_var := address_0_reg;
				address_1_var := address_1_reg;

	
				next_fsm_state := WaitResponsePipeState;
				latch_new_window_regs_var := true;
				
				write_req_var := '1';
				if(iunit_register_file_window_update_response_pipe_write_ack(0) = '1') then
					next_fsm_state := IdleState;
				end if;
		end case;

		iunit_register_file_window_update_response_pipe_write_req(0) <= write_req_var;
		iunit_register_file_window_update_command_pipe_read_req(0)  <= read_req_var;

		
		dpmem_address_0 <= address_0_var;
		dpmem_write_data_0 <= write_data_0_var;
		dpmem_enable_0 <= enable_0_var;
		dpmem_read_writebar_0 <= read_writebar_0_var;

		dpmem_address_1 <= address_1_var;
		dpmem_write_data_1 <= write_data_1_var;
		dpmem_enable_1 <= enable_1_var;
		dpmem_read_writebar_1 <= read_writebar_1_var;

		new_globals<= new_globals_var;
		new_outs<= new_outs_var;
		new_locals<= new_locals_var;
		new_ins<= new_ins_var;

		if(clk'event and clk = '1') then
			if(reset = '1') then
				fsm_state <= IdleState;
			else
				fsm_state <= next_fsm_state;
				if(latch_inputs_var) then
					valid_reg  <= valid_var;
					rd_val_reg <= rd_val_var;
					rd_reg <= rd_var;
					restore_reg <= restore_var;
					save_reg <= save_var;
					write_psr_reg <= write_psr_var;
					ins_reg  <= ins_var;
					locals_reg <= locals_var;
					outs_reg <= outs_var;
					globals_reg <= globals_var;
					wr_wp_reg <= oldcwp_var;
					cycle_count_reg <= cycle_count_var;
					tag_out <= tag_in;
					oldcwp_reg <= oldcwp_var;
					newcwp_reg <= newcwp_var;
				end if;

				if(latch_rd_wp_var) then
					rd_wp_reg <= rd_wp_var;
				end if;

				if(latch_fetched_locals_var) then
					fetched_locals_reg <= dpmem_read_data_1;
				end if;

				if(latch_addresses_var) then
					address_0_reg <= address_0_var;
					address_1_reg <= address_1_var;
				end if;

			end if;
		end if;
	end process;

	
				
    	iunit_register_file_window_update_response_pipe_write_data <=
			cycle_count_reg & new_globals & new_outs & new_locals & new_ins & rd_wp_reg & const_one_1;

				
	dpmem: base_bank_dual_port
			generic map (name => "window_update_daemon:dpmem",
					g_addr_width => 5,
					g_data_width => 256)
			port map ( datain_0 => dpmem_write_data_0,
					dataout_0 => dpmem_read_data_0,
					enable_0 => dpmem_enable_0,
					writebar_0 => dpmem_read_writebar_0,
					addrin_0 => dpmem_address_0, 
					datain_1 => dpmem_write_data_1,
					dataout_1 => dpmem_read_data_1,
					enable_1 => dpmem_enable_1,
					writebar_1 => dpmem_read_writebar_1,
					addrin_1 => dpmem_address_1, 
					clk => clk, reset => reset);

end window_update_daemon_arch;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library AjitCustom;
use AjitCustom.AjitCustomComponents.all;

-- singl port memory to model dcache.
entity cpu_test_setup_memory_dcache  is
	generic (tag_length: integer := 2);
	port ( 
		read_write_bar : in std_logic_vector (0 downto 0);
		enable : in std_logic_vector (0 downto 0);
		byte_mask  : in std_logic_vector (7 downto 0);
		address    : in  std_logic_vector (12 downto 0); -- 16kwords.
		datain : in std_logic_vector (63 downto 0);
		dataout  : out  std_logic_vector (63 downto 0);
 	   	tag_in: in std_logic_vector(tag_length-1 downto 0);
      	   	tag_out: out std_logic_vector(tag_length-1 downto 0);
		clk, reset: in std_logic;
		start_req: in std_logic;
		start_ack: out std_logic;
		fin_req: in std_logic;
		fin_ack: out std_logic
	     );
end entity cpu_test_setup_memory_dcache;


architecture Mixed of cpu_test_setup_memory_dcache is
	signal fin_ack_sig: std_logic;
	signal enable_sig, enable_mem : std_logic;
begin
	enable_mem <= enable_sig and enable(0);
	

	memInst: generic_single_port_memory_with_byte_mask_and_init
			generic map (init_file_name => "cpu_test_setup_memmap_dcache.txt",
					g_addr_width => 13,
					g_data_width => 64)
			port map (
					datain => datain,
					dataout => dataout,
					addrin => address(12 downto 0),
					bytemask => byte_mask,
					enable => enable_mem,
					writebar => read_write_bar(0),
					clk => clk, 
					reset => reset);


	-- state machine! Assuming that the memory is one-cycle.
	process(clk, reset, fin_req, start_req, fin_ack_sig, tag_in, enable_sig)
		variable next_fin_ack_sig: std_logic;
	begin 
		next_fin_ack_sig :=
			((not fin_ack_sig) and start_req)
				or
			(fin_ack_sig and (not fin_req))
				or
			(fin_ack_sig and fin_req and start_req);

		enable_sig <= 
			((not fin_ack_sig) and start_req) 
				or
			(fin_ack_sig and fin_req and start_req);

		if(clk'event and (clk = '1')) then
			if(reset = '1') then
				fin_ack_sig <= '0';
				tag_out <= (others => '0');
			else
				if (enable_sig = '1') then
					tag_out <= tag_in;
				end if;

				fin_ack_sig <= next_fin_ack_sig;
			end if;

		end if;
	end process;

	fin_ack <= fin_ack_sig;
	start_ack <= enable_sig;
end Mixed;
		
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library AjitCustom;
use AjitCustom.AjitCustomComponents.all;

-- single port memory to model icache.
entity cpu_test_setup_memory_icache  is
	generic (tag_length: integer := 2);
	port ( 
		read_write_bar : in std_logic_vector (0 downto 0);
		enable : in std_logic_vector (0 downto 0);
		byte_mask  : in std_logic_vector (7 downto 0);
		address    : in  std_logic_vector (12 downto 0); -- 16kwords.
		datain : in std_logic_vector (63 downto 0);
		dataout  : out  std_logic_vector (63 downto 0);
 	   	tag_in: in std_logic_vector(tag_length-1 downto 0);
      	   	tag_out: out std_logic_vector(tag_length-1 downto 0);
		clk, reset: in std_logic;
		start_req: in std_logic;
		start_ack: out std_logic;
		fin_req: in std_logic;
		fin_ack: out std_logic
	     );
end entity cpu_test_setup_memory_icache;


architecture Mixed of cpu_test_setup_memory_icache is
	signal fin_ack_sig: std_logic;
	signal enable_sig, enable_mem : std_logic;
begin
	
	enable_mem <= enable_sig and enable(0);

	memInst: generic_single_port_memory_with_byte_mask_and_init
			generic map (init_file_name => "cpu_test_setup_memmap_icache.txt",
					g_addr_width => 13,
					g_data_width => 64)
			port map (
					datain => datain,
					dataout => dataout,
					addrin => address(12 downto 0),
					bytemask => byte_mask,
					enable => enable_mem,
					writebar => read_write_bar(0),
					clk => clk, 
					reset => reset);

	-- state machine! Assuming that the memory is one-cycle.
	process(clk, reset, fin_req, start_req, fin_ack_sig, tag_in)
		variable next_fin_ack_sig: std_logic;
	begin 
		next_fin_ack_sig :=
			((not fin_ack_sig) and start_req)
				or
			(fin_ack_sig and (not fin_req))
				or
			(fin_ack_sig and fin_req and start_req);

		enable_sig <= 
			((not fin_ack_sig) and start_req) 
				or
			(fin_ack_sig and fin_req and start_req);

		if(clk'event and (clk = '1')) then
			if(reset = '1') then
				fin_ack_sig <= '0';
				tag_out <= (others => '0');
			else
				if (enable_sig = '1') then
					tag_out <= tag_in;
				end if;

				fin_ack_sig <= next_fin_ack_sig;
			end if;
		end if;
	end process;

	fin_ack <= fin_ack_sig;
	start_ack <= enable_sig;
end Mixed;
		
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.BaseComponents.all;

library AjitCustom;
use AjitCustom.AjitCustomComponents.all;

-- dual port memory to model icache/dcache.
entity cpu_test_setup_memory_Operator  is
	port ( 
		read_write_bar_0 : in std_logic_vector (0 downto 0);
		enable_0 : in std_logic_vector (0 downto 0);
		byte_mask_0  : in std_logic_vector (7 downto 0);
		address_0    : in  std_logic_vector (11 downto 0); -- 8kwords.
		datain_0 : in std_logic_vector (63 downto 0);
		dataout_0  : out  std_logic_vector (63 downto 0);
		read_write_bar_1 : in std_logic_vector (0 downto 0);
		enable_1 : in std_logic_vector (0 downto 0);
		byte_mask_1  : in std_logic_vector (7 downto 0);
		address_1    : in  std_logic_vector (11 downto 0); -- 8kwords.
		datain_1 : in std_logic_vector (63 downto 0);
		dataout_1  : out  std_logic_vector (63 downto 0);
		clk, reset: in std_logic;
		sample_req: in boolean;
		sample_ack: out boolean;
		update_req: in boolean;
		update_ack: out boolean
	     );
end entity cpu_test_setup_memory_Operator;


architecture Mixed of cpu_test_setup_memory_Operator is
	signal start_req, start_ack, fin_req, fin_ack: std_logic;
	signal tag_in, tag_out : std_logic_vector(0 downto 0);
begin
   tag_in(0) <= '0';

   p2l: Sample_Pulse_To_Level_Translate_Entity
		generic map(name => "cpu_test_setup_memory-Operator-p2l")
		port map (rL => sample_req, rR => start_req,
				aL => sample_ack, aR => start_ack,
					clk => clk, reset => reset);
   l2p: Level_To_Pulse_Translate_Entity
		generic map(name => "cpu_test_setup_memory-Operator-l2p")
		port map (rL => fin_req, rR => update_req,
				aL => fin_ack, aR => update_ack, clk => clk, reset => reset);
				

    dpmem: cpu_test_setup_memory
		generic map (tag_length => 1)
		port map 
		(
			read_write_bar_0  => read_write_bar_0 ,
			enable_0  => enable_0 ,
			byte_mask_0  => byte_mask_0 ,
			address_0     => address_0    ,
			datain_0  => datain_0 ,
			dataout_0   => dataout_0  ,
			read_write_bar_1  => read_write_bar_1 ,
			enable_1  => enable_1 ,
			byte_mask_1   => byte_mask_1  ,
			address_1     => address_1    ,
			datain_1  => datain_1 ,
			dataout_1   => dataout_1  ,
 	   		tag_in => tag_in,
      	   		tag_out => tag_out,
			clk => clk, reset => reset,
			start_req => start_req,
			start_ack => start_ack,
			fin_req => fin_req,
			fin_ack => fin_ack
		);
end Mixed;
		
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library AjitCustom;
use AjitCustom.AjitCustomComponents.all;

-- dual port memory to model icache/dcache.
entity cpu_test_setup_memory  is
	generic (tag_length: integer := 2);
	port ( 
		read_write_bar_0 : in std_logic_vector (0 downto 0);
		enable_0 : in std_logic_vector (0 downto 0);
		byte_mask_0  : in std_logic_vector (7 downto 0);
		address_0    : in  std_logic_vector (11 downto 0); -- 8kwords.
		datain_0 : in std_logic_vector (63 downto 0);
		dataout_0  : out  std_logic_vector (63 downto 0);
		read_write_bar_1 : in std_logic_vector (0 downto 0);
		enable_1 : in std_logic_vector (0 downto 0);
		byte_mask_1  : in std_logic_vector (7 downto 0);
		address_1    : in  std_logic_vector (11 downto 0); -- 8kwords.
		datain_1 : in std_logic_vector (63 downto 0);
		dataout_1  : out  std_logic_vector (63 downto 0);
 	   	tag_in: in std_logic_vector(tag_length-1 downto 0);
      	   	tag_out: out std_logic_vector(tag_length-1 downto 0);
		clk, reset: in std_logic;
		start_req: in std_logic;
		start_ack: out std_logic;
		fin_req: in std_logic;
		fin_ack: out std_logic
	     );
end entity cpu_test_setup_memory;

-------------- BROKEN  DO NOT USE
architecture Mixed of cpu_test_setup_memory is
	signal stall_signal: std_logic;
	signal fin_ack_sig: std_logic;
	signal enable_sig : std_logic;
begin
	
	stall_signal <= (fin_ack_sig and (not fin_req));
	enable_sig <= (not stall_signal) and start_req;
	start_ack <= enable_sig;

	memInst: generic_dual_port_memory_with_byte_mask
			generic map (name => "GenericMem64KB",
					g_addr_width => 12,
					g_data_width => 64)
			port map (
					datain_0 => datain_0,
					dataout_0 => dataout_0,
					addrin_0 => address_0(11 downto 0),
					bytemask_0 => byte_mask_0,
					enable_0 => enable_0(0),
					writebar_0 => read_write_bar_0(0),
					datain_1 => datain_1,
					dataout_1 => dataout_1,
					addrin_1 => address_1(11 downto 0),
					bytemask_1 => byte_mask_1,
					enable_1 => enable_1(0),
					writebar_1 => read_write_bar_1(0),
					clk => clk, 
					reset => reset);

	process(clk)
	begin 
		if(clk'event and (clk = '1')) then
			if(reset = '1') then
				fin_ack_sig <= '0';
				tag_out <= (others => '0');
			elsif (enable_sig = '1') then
				tag_out <= tag_in;
				fin_ack_sig <= '1';
			elsif (fin_req = '1') then
				fin_ack_sig <= '0';
			end if;
		end if;
	end process;

	fin_ack <= fin_ack_sig;
end Mixed;
		
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
entity dcache_stub_daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    NOBLOCK_CPU_to_DCACHE_command_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_command_pipe_read_data : in   std_logic_vector(120 downto 0);
    NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_data : in   std_logic_vector(120 downto 0);
    DCACHE_to_CPU_response_pipe_write_req : out  std_logic_vector(0 downto 0);
    DCACHE_to_CPU_response_pipe_write_ack : in   std_logic_vector(0 downto 0);
    DCACHE_to_CPU_response_pipe_write_data : out  std_logic_vector(71 downto 0);
    DCACHE_to_CPU_slow_response_pipe_write_req : out  std_logic_vector(0 downto 0);
    DCACHE_to_CPU_slow_response_pipe_write_ack : in   std_logic_vector(0 downto 0);
    DCACHE_to_CPU_slow_response_pipe_write_data : out  std_logic_vector(71 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity dcache_stub_daemon;
architecture dcache_stub_daemon_arch of dcache_stub_daemon is -- 

	signal dcache_cmd : std_logic_vector(120 downto 0);
	signal dcache_cmd_valid: std_logic;
	signal dcache_cmd_req_type : std_logic_vector(7 downto 0);
	signal dcache_cmd_asi: std_logic_vector(7 downto 0);
	signal dcache_cmd_byte_mask: std_logic_vector(7 downto 0);
	signal dcache_cmd_addr: std_logic_vector(31 downto 0);
	signal dcache_cmd_data: std_logic_vector(63 downto 0);

	signal mem_enable, mem_read_writebar : std_logic;
	signal mem_addr: std_logic_vector(12 downto 0);
	signal mem_datain, mem_dataout: std_logic_vector(63 downto 0);
	signal mem_byte_mask : std_logic_vector (7 downto 0);

	signal dcache_response : std_logic_vector(71 downto 0);
	constant ccc_zero_8: std_logic_vector(7 downto 0) := "00000000";
	signal m_tag_in, m_tag_out: std_logic_vector(0 downto 0);

	signal m_start_req, m_start_ack, m_fin_req, m_fin_ack: std_logic;

	signal do_fast, do_slow: std_logic;

begin --  


	start_ack <= '1';
	fin_ack <= '0';

	do_fast <= NOBLOCK_CPU_to_DCACHE_command_pipe_read_ack(0);
	do_slow <= (NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_ack(0) and (not do_fast));
	m_tag_in(0) <= do_fast;
	
	m_start_req <= do_fast or do_slow;
	NOBLOCK_CPU_to_DCACHE_command_pipe_read_req(0)      <= m_start_ack when do_fast = '1' else '0';
	NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_req(0) <= m_start_ack when do_slow = '1' else '0';


	dcache_cmd <= NOBLOCK_CPU_to_DCACHE_command_pipe_read_data when do_fast = '1' else
						NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_data;
	dcache_cmd_data <= dcache_cmd (63 downto 0);
	dcache_cmd_addr <= dcache_cmd (95 downto 64);
	dcache_cmd_byte_mask <= dcache_cmd (103 downto 96);
	dcache_cmd_asi <= dcache_cmd (111 downto 104);
	dcache_cmd_req_type <= dcache_cmd (119 downto 112);
	dcache_cmd_valid <= dcache_cmd(120);

	mem_enable <= dcache_cmd_valid when 
				((dcache_cmd_asi(6 downto 0) = "0001010") 
					or (dcache_cmd_asi(6 downto 0) = "0100000")
					or (dcache_cmd_asi(6 downto 0) = "0001011")) else '0';
	mem_read_writebar <= '0' when (dcache_cmd_req_type(3 downto 0) = "0110") or
					(dcache_cmd_req_type(3 downto 0) = "0010") else '1';
	mem_addr <=  dcache_cmd_addr (15 downto 3);
	mem_datain <= dcache_cmd_data;
	mem_byte_mask <= dcache_cmd_byte_mask;
	
	dcacheMem: cpu_test_setup_memory_dcache
			generic map (tag_length => 1)
			port map (
				read_write_bar(0) => mem_read_writebar,
				enable(0) => mem_enable,
				byte_mask => mem_byte_mask,
				address => mem_addr,
				datain => mem_datain,
				dataout => mem_dataout,
				tag_in => m_tag_in,
				tag_out => m_tag_out,
				clk => clk, reset => reset,
				start_req => m_start_req,
				start_ack => m_start_ack,
				fin_req => m_fin_req,
				fin_ack => m_fin_ack);

	-- whose turn is it?
	m_fin_req <= DCACHE_to_CPU_response_pipe_write_ack(0) when ((m_fin_ack = '1') and (m_tag_out(0) = '1'))
				else DCACHE_to_CPU_slow_response_pipe_write_ack(0) when (m_fin_ack ='1')  else '0';
	DCACHE_to_CPU_response_pipe_write_req(0) <= (m_fin_ack and m_tag_out(0));
	DCACHE_to_CPU_slow_response_pipe_write_req(0) <= (m_fin_ack and (not m_tag_out(0)));

	DCACHE_to_CPU_response_pipe_write_data <= ccc_zero_8 & mem_dataout;
	DCACHE_to_CPU_slow_response_pipe_write_data <= ccc_zero_8 & mem_dataout;

end dcache_stub_daemon_arch;
-- A tightly coupled memory for use in the stupid dhrystone and coremark benchmarks..
library std;
use std.textio.all;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.BaseComponents.all;
use ahir.mem_component_pack.all;
use ahir.Utilities.all;

entity dual_port_u64_mem_64KB_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    read_0 : in  std_logic_vector(0 downto 0);
    addr_0 : in  std_logic_vector(12 downto 0);
    read_1 : in  std_logic_vector(0 downto 0);
    write_1 : in  std_logic_vector(0 downto 0);
    byte_mask : in  std_logic_vector(7 downto 0);
    addr_1 : in  std_logic_vector(12 downto 0);
    write_data_1 : in  std_logic_vector(63 downto 0);
    read_data_0 : out  std_logic_vector(63 downto 0);
    read_data_1 : out  std_logic_vector(63 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity dual_port_u64_mem_64KB_Operator;

architecture dual_port_u64_mem_64KB_Operator_arch of dual_port_u64_mem_64KB_Operator is -- 
	signal joined_sig: boolean;	
        signal memory_enable: std_logic;
	signal z8: std_logic_vector(7 downto 0);
        signal osig: std_logic;
begin --  

    trig_join: join2 generic map (name => "dual_port_u64_mem_Operator:trig-join", bypass => true)
			port map (pred0 => sample_req, pred1 => update_req,
					symbol_out => joined_sig, clk => clk, reset => reset);
   
    sample_ack <= joined_sig;

    process(clk, reset)
    begin
	if(clk'event and clk='1') then
		if(reset = '1') then
			update_ack <= false;
		else
			update_ack <= joined_sig;
		end if;
	end if;
    end process;

    memory_enable <= '1' when joined_sig else '0';
    z8 <= (others => '0');
    osig <= '1';

    -- instantiate base bank dual port....... (generate 8 banks).
    bankgen: for B in 0 to 7 generate
     bank: block
         signal local_enable_0, local_enable_1: std_logic;
	 signal writebar_1: std_logic;
     begin
	  writebar_1 <= not write_1(0);

          local_enable_0 <= memory_enable and read_0(0);
	  local_enable_1 <= memory_enable and (read_1(0) or (write_1(0) and byte_mask(B)));
	
	  bb: base_bank_dual_port
		generic map (name => "dual_port_u64_bb", g_addr_width => 13, g_data_width => 8)
		port map (
	 		datain_0 => z8,
         		dataout_0 => read_data_0((8*(B+1))-1 downto 8*B),
         		addrin_0 => addr_0,
         		enable_0 => local_enable_0,
         		writebar_0 => osig,
	 		datain_1  => write_data_1((8*(B+1))-1 downto 8*B),
         		dataout_1 => read_data_1((8*(B+1))-1 downto 8*B),
         		addrin_1 => addr_1,
         		enable_1 => local_enable_1,
         		writebar_1 => writebar_1,
         		clk => clk, reset => reset);
    end block;
  end generate bankgen;

end dual_port_u64_mem_64KB_Operator_arch;
-- THIS IS TO BE USED ONLY FOR SIMULATIONS!
library std;
use std.textio.all;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.BaseComponents.all;
use ahir.mem_component_pack.all;
use ahir.Utilities.all;

library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
use AjitCustom.MemmapPackage.all;

-- NOTE: only for simulations.
entity dual_port_u64_mem_with_init_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    first_time : in  std_logic_vector(0 downto 0);
    read_0 : in  std_logic_vector(0 downto 0);
    addr_0 : in  std_logic_vector(28 downto 0);
    read_1 : in  std_logic_vector(0 downto 0);
    write_1 : in  std_logic_vector(0 downto 0);
    byte_mask : in  std_logic_vector(7 downto 0);
    addr_1 : in  std_logic_vector(28 downto 0);
    write_data_1 : in  std_logic_vector(63 downto 0);
    read_data_0 : out  std_logic_vector(63 downto 0);
    read_data_1 : out  std_logic_vector(63 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity dual_port_u64_mem_with_init_Operator;

architecture dual_port_u64_mem_with_init_Operator_arch of dual_port_u64_mem_with_init_Operator is -- 
	type MemArray is array (natural range <>) of std_logic_vector(63 downto 0);
	
	signal joined_sig: boolean;	
begin --  

    trig_join: join2 generic map (name => "dual_port_u64_mem_with_init_Operator:trig-join", bypass => true)
			port map (pred0 => sample_req, pred1 => update_req,
					symbol_out => joined_sig, clk => clk, reset => reset);
   
    sample_ack <= joined_sig;

    process(clk, reset)
    begin
	if(clk'event and clk='1') then
		if(reset = '1') then
			update_ack <= false;
		else
			update_ack <= joined_sig;
		end if;
	end if;
    end process;

    -- ports
    process(clk, reset, joined_sig, first_time, read_0, addr_0, read_1, write_1, addr_1, byte_mask, write_data_1)
	-- 8k X 64B.  double word address is 13 bits (truncated).
	variable mem_array: MemArray (0 to 8191);
	variable tval: std_logic_vector(63 downto 0);
	variable address_var, u64_address_var, offset_var: integer;
    	variable data_var : bit_vector(7 downto 0);
    	variable slv_data_var : std_logic_vector(7 downto 0);
    	File INFILE: text open read_mode is "cpu_test_setup_memmap.txt";
        variable INPUT_LINE: Line;
    begin
	if(clk'event and clk = '1') then
		if(reset = '1') then
			read_data_0 <= (others => '0');
			read_data_1 <= (others => '0');
		else
			if(first_time(0) = '1') then
				-- read file and populate array.
    				while not endfile(INFILE) loop
          				readLine (INFILE, INPUT_LINE);
          				read (INPUT_LINE, address_var);
          				read (INPUT_LINE, data_var);
          				slv_data_var := to_std_logic_vector(data_var);
					u64_address_var := (address_var/8);
					offset_var      := (address_var - (u64_address_var * 8));
					tval := mem_array(u64_address_var);
					mem_array(u64_address_var) := 
						insertByteIntoU64(tval, offset_var, slv_data_var);
					assert false report "Info: byte mem_array[" &
								Convert_To_String(address_var) & "] = "
								& Convert_SLV_to_string(slv_data_var)
							severity note;
    				end loop;
          		end if; -- first_time
			
			if(joined_sig) then
				if(read_0(0) = '1') then
					read_data_0 <= mem_array(to_integer(unsigned(addr_0(12 downto 0))));
				end if; -- read_0
				if(read_1(0) = '1') then
					read_data_1 <=  mem_array(to_integer(unsigned(addr_1(12 downto 0))));
				end if; -- read_1
				if(write_1(0) = '1') then
					tval :=  mem_array(to_integer(unsigned(addr_1(12 downto 0))));
					mem_array(to_integer(unsigned(addr_1(12 downto 0)))) :=
							updateU64UsingByteMask(tval, byte_mask, write_data_1);
				end if; -- write_1
			end if; -- joined_sig
		end if;
	end if;
    end process;

end dual_port_u64_mem_with_init_Operator_arch;
-- Generic memory for use in proto-board.
--  Uses base_bank.vhd in AHIR.
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.BaseComponents.all;
use ahir.mem_component_pack.all;
use ahir.Utilities.all;

library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
use AjitCustom.MemmapPackage.all;


entity generic_dual_port_memory_with_byte_mask is
   generic ( name: string; 
		g_addr_width: natural := 10; 
		g_data_width : natural := 16);
   port (
	   datain_0 : in std_logic_vector(g_data_width-1 downto 0);
           dataout_0: out std_logic_vector(g_data_width-1 downto 0);
           addrin_0: in std_logic_vector(g_addr_width-1 downto 0);
	   bytemask_0: in std_logic_vector((g_data_width/8)-1 downto 0);
           enable_0: in std_logic;
           writebar_0 : in std_logic;
	   datain_1 : in std_logic_vector(g_data_width-1 downto 0);
           dataout_1: out std_logic_vector(g_data_width-1 downto 0);
           addrin_1: in std_logic_vector(g_addr_width-1 downto 0);
	   bytemask_1: in std_logic_vector((g_data_width/8)-1 downto 0);
           enable_1: in std_logic;
           writebar_1 : in std_logic;
           clk: in std_logic;
           reset : in std_logic);
end entity generic_dual_port_memory_with_byte_mask;


architecture Mixed of generic_dual_port_memory_with_byte_mask is
	constant init_byte_array : ByteArray(0 to (2**(g_addr_width+3))-1) :=
			construct_init_byte_array("cpu_test_setup_memmap.txt", (2**(g_addr_width+3)));
begin  -- XilinxBramInfer


  genByteMem: for I in 0 to (g_data_width/8)-1 generate

	memBlock: block
		signal local_enable_sig_0 : std_logic;
		signal local_enable_sig_1 : std_logic;
		constant local_init_byte_array : ByteArray(0 to (2**g_addr_width)-1) :=
			Select_Byte_Init_Value_By_Position_In_Double_Word (I, init_byte_array);
		constant J: integer := ((g_data_width/8)-1)-I;
	begin
		local_enable_sig_0 <= enable_0 and (writebar_0 or bytemask_0(J));
		local_enable_sig_1 <= enable_1 and (writebar_1 or bytemask_1(J));
		
		bb: dual_port_byte_ram_with_init
			generic map (byte_position => I,
					g_addr_width => g_addr_width,
					init_byte_array => local_init_byte_array)
			port map(
					datain_0 => datain_0((8*(J+1))-1 downto (8*J)),
					dataout_0 => dataout_0((8*(J+1))-1 downto (8*J)),
					addrin_0 => addrin_0,
					enable_0 => local_enable_sig_0,
					writebar_0 => writebar_0,
					datain_1 => datain_1((8*(J+1))-1 downto (8*J)),
					dataout_1 => dataout_1((8*(J+1))-1 downto (8*J)),
					addrin_1 => addrin_1,
					enable_1 => local_enable_sig_1,
					writebar_1 => writebar_1,
					clk => clk,
					reset => reset);

	end block memBlock;
  end generate genByteMem;

end Mixed;
-- Generic memory for use in proto-board.
--  Uses base_bank.vhd in AHIR.
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.BaseComponents.all;
use ahir.mem_component_pack.all;
use ahir.Utilities.all;

library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
use AjitCustom.MemmapPackage.all;

entity generic_single_port_memory_with_byte_mask_and_init is
   generic ( init_file_name: string; 
		g_addr_width: natural := 10; 
		g_data_width : natural := 16);
   port (
	   datain : in std_logic_vector(g_data_width-1 downto 0);
           dataout: out std_logic_vector(g_data_width-1 downto 0);
           addrin: in std_logic_vector(g_addr_width-1 downto 0);
	   bytemask: in std_logic_vector((g_data_width/8)-1 downto 0);
           enable: in std_logic;
           writebar : in std_logic;
           clk: in std_logic;
           reset : in std_logic);
end entity generic_single_port_memory_with_byte_mask_and_init;


architecture Mixed of generic_single_port_memory_with_byte_mask_and_init is
	constant init_byte_array : ByteArray(0 to (2**(g_addr_width+3))-1) :=
			construct_init_byte_array(init_file_name, (2**(g_addr_width+3)));
begin  -- XilinxBramInfer

  genByteMem: for I in 0 to (g_data_width/8)-1 generate

	memBlock: block
		signal local_enable_sig : std_logic;
		constant local_init_byte_array : ByteArray(0 to (2**g_addr_width)-1) :=
			Select_Byte_Init_Value_By_Position_In_Double_Word (I, init_byte_array);
		constant J: integer := ((g_data_width/8)-1)-I;
	begin
		local_enable_sig <= enable and (writebar or bytemask(J));
		
		bb: single_port_byte_ram_with_init
			generic map (byte_position => I,
					g_addr_width => g_addr_width,
					init_byte_array => local_init_byte_array)
			port map(
					datain => datain((8*(J+1))-1 downto (8*J)),
					dataout => dataout((8*(J+1))-1 downto (8*J)),
					addrin => addrin,
					enable => local_enable_sig,
					writebar => writebar,
					clk => clk,
					reset => reset);

	end block memBlock;
  end generate genByteMem;
end Mixed;
-- Generic memory for use in proto-board.
--  Uses base_bank.vhd in AHIR.
--
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.BaseComponents.all;
use ahir.mem_component_pack.all;
use ahir.Utilities.all;


entity generic_single_port_memory_with_byte_mask is
   generic ( name: string; 
		g_addr_width: natural := 10; 
		g_data_width : natural := 16);
   port (
	   datain : in std_logic_vector(g_data_width-1 downto 0);
           dataout: out std_logic_vector(g_data_width-1 downto 0);
           addrin: in std_logic_vector(g_addr_width-1 downto 0);
	   bytemask: in std_logic_vector((g_data_width/8)-1 downto 0);
           enable: in std_logic;
           writebar : in std_logic;
           clk: in std_logic;
           reset : in std_logic);
end entity generic_single_port_memory_with_byte_mask;


architecture Mixed of generic_single_port_memory_with_byte_mask is
begin  -- XilinxBramInfer

  genByteMem: for I in 0 to (g_data_width/8)-1 generate

	memBlock: block
		signal local_enable_sig : std_logic;
	begin
		local_enable_sig <= enable and (writebar or bytemask(I));
		
		bb: base_bank
			generic map (name => "BB_" & Convert_To_String(I),
					g_addr_width => g_addr_width,
					g_data_width => 8)
			port map(
					datain => datain((8*(I+1))-1 downto (8*I)),
					dataout => dataout((8*(I+1))-1 downto (8*I)),
					addrin => addrin,
					enable => local_enable_sig,
					writebar => writebar,
					clk => clk,
					reset => reset);

	end block memBlock;
  end generate genByteMem;

end Mixed;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
entity icache_stub_daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    NOBLOCK_CPU_to_ICACHE_command_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_ICACHE_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_ICACHE_command_pipe_read_data : in   std_logic_vector(40 downto 0);
    ICACHE_to_CPU_response_pipe_write_req : out  std_logic_vector(0 downto 0);
    ICACHE_to_CPU_response_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ICACHE_to_CPU_response_pipe_write_data : out  std_logic_vector(89 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity icache_stub_daemon;
architecture icache_stub_daemon_arch of icache_stub_daemon is -- 

	signal icache_cmd : std_logic_vector(40 downto 0);
	signal icache_cmd_valid: std_logic;
	signal icache_cmd_asi: std_logic_vector(7 downto 0);
	signal icache_cmd_addr: std_logic_vector(31 downto 0);

	signal mem_enable, mem_read_writebar : std_logic;
	signal mem_addr: std_logic_vector(12 downto 0);
	signal mem_datain, mem_dataout: std_logic_vector(63 downto 0);
	signal mem_byte_mask: std_logic_vector(7 downto 0);

	constant ccc_zero_26: std_logic_vector(25 downto 0) := (others => '0');
	signal m_tag_in, m_tag_out: std_logic_vector(0 downto 0);

	signal m_start_req, m_start_ack, m_fin_req, m_fin_ack: std_logic;

        function my_to_01 (x: std_logic_vector) return std_logic_vector is
          alias lx: std_logic_vector(1 to x'length) is x;
          variable ret_var : std_logic_vector(1 to x'length);
        begin
          for I in 1 to lx'length loop
            if(lx(I) = '0') then
               ret_var (I) := '0';
            elsif (lx(I) = '1') then
               ret_var (I) := '1';
            else
               ret_var (I) := '0';
            end if;
          end loop;
          return ret_var;
        end function;

begin --  
	mem_byte_mask <= "11111111";
	m_tag_in(0) <= '0';
	start_ack <= '1';
	fin_ack <= '0';
	
	m_start_req <= NOBLOCK_CPU_to_ICACHE_command_pipe_read_ack(0);
	NOBLOCK_CPU_to_ICACHE_command_pipe_read_req(0) <= m_start_ack;

	m_fin_req <= ICACHE_to_CPU_response_pipe_write_ack(0);
	ICACHE_to_CPU_response_pipe_write_req(0) <= m_fin_ack;

	icache_cmd <= NOBLOCK_CPU_to_ICACHE_command_pipe_read_data;
	icache_cmd_addr <= icache_cmd (31 downto 0);
	icache_cmd_asi <= icache_cmd (39 downto 32);
	icache_cmd_valid <= icache_cmd(40);

	mem_enable <= icache_cmd_valid;
	mem_read_writebar <= '1';
	mem_addr <=  icache_cmd_addr(15 downto 3);
	mem_datain <= (others => '0');
	
	icacheMem: cpu_test_setup_memory_icache
			generic map (tag_length => 1)
			port map (
				read_write_bar(0) => mem_read_writebar,
				enable(0) => mem_enable,
				byte_mask => mem_byte_mask,
				address => mem_addr,
				datain => mem_datain,
				dataout => mem_dataout,
				tag_in => m_tag_in,
				tag_out => m_tag_out,
				clk => clk, reset => reset,
				start_req => m_start_req,
				start_ack => m_start_ack,
				fin_req => m_fin_req,
				fin_ack => m_fin_ack);

	ICACHE_to_CPU_response_pipe_write_data <= ccc_zero_26 & my_to_01(mem_dataout);

end icache_stub_daemon_arch;
--
-- has all the interfaces necessary for initialization and access.
-- 
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity mem_test_setup_memory  is
	generic (tag_length: integer := 2);
	port ( 

		read_write_bar : in std_logic_vector (0 downto 0);
		byte_mask  : in std_logic_vector (7 downto 0);
		-- 2048 x 64
		address    : in  std_logic_vector (10 downto 0);
		write_data : in std_logic_vector (63 downto 0);
		read_data  : out  std_logic_vector (63 downto 0);
 	   	tag_in: in std_logic_vector(tag_length-1 downto 0);
      	   	tag_out: out std_logic_vector(tag_length-1 downto 0);
		clk, reset: in std_logic;
		start_req: in std_logic;
		start_ack: out std_logic;
		fin_req: in std_logic;
		fin_ack: out std_logic
	     );
end entity mem_test_setup_memory;


architecture Mixed of mem_test_setup_memory is
	signal stall_signal: std_logic;
	signal fin_ack_sig: std_logic;
	signal enable_sig : std_logic;
   
	component generic_single_port_memory_with_byte_mask is
   	generic ( name: string; 
		g_addr_width: natural := 10; 
		g_data_width : natural := 16);
   	port (
	   datain : in std_logic_vector(g_data_width-1 downto 0);
           dataout: out std_logic_vector(g_data_width-1 downto 0);
           addrin: in std_logic_vector(g_addr_width-1 downto 0);
	   bytemask: in std_logic_vector((g_data_width/8)-1 downto 0);
           enable: in std_logic;
           writebar : in std_logic;
           clk: in std_logic;
           reset : in std_logic);
	end component;
begin
	
	stall_signal <= (fin_ack_sig and (not fin_req));
	enable_sig <= (not stall_signal) and start_req;
	start_ack  <= enable_sig;

	memInst: generic_single_port_memory_with_byte_mask
			generic map (name => "GenericMem2MB",
					g_addr_width => 11,
					g_data_width => 64)
			port map (
					datain => write_data,
					dataout => read_data,
					addrin => address,
					bytemask => byte_mask,
					enable => enable_sig,
					writebar => read_write_bar(0),
					clk => clk, 
					reset => reset);

	process(clk)
	begin 
		if(clk'event and (clk = '1')) then
			if(reset = '1') then
				fin_ack_sig <= '0';
				tag_out <= (others => '0');
			elsif (enable_sig = '1') then
				tag_out <= tag_in;
				fin_ack_sig <= '1';
			else
				fin_ack_sig <= '0';
			end if;
		end if;
	end process;

	fin_ack <= fin_ack_sig;
end Mixed;
		
--
-- has all the interfaces necessary for initialization and access.
-- 
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity protoBoardMemX2MB  is
	generic (tag_length: integer := 2);
	port ( 

		read_write_bar : in std_logic_vector (0 downto 0);
		byte_mask  : in std_logic_vector (7 downto 0);
		address    : in  std_logic_vector (18 downto 0);
		write_data : in std_logic_vector (63 downto 0);
		read_data  : out  std_logic_vector (63 downto 0);
 	   	tag_in: in std_logic_vector(tag_length-1 downto 0);
      	   	tag_out: out std_logic_vector(tag_length-1 downto 0);
		clk, reset: in std_logic;
		start_req: in std_logic;
		start_ack: out std_logic;
		fin_req: in std_logic;
		fin_ack: out std_logic
	     );
end entity protoBoardMemX2MB;


architecture Mixed of protoBoardMemX2MB is
	signal stall_signal: std_logic;
	signal fin_ack_sig: std_logic;
	signal enable_sig : std_logic;
   
	component generic_single_port_memory_with_byte_mask is
   	generic ( name: string; 
		g_addr_width: natural := 10; 
		g_data_width : natural := 16);
   	port (
	   datain : in std_logic_vector(g_data_width-1 downto 0);
           dataout: out std_logic_vector(g_data_width-1 downto 0);
           addrin: in std_logic_vector(g_addr_width-1 downto 0);
	   bytemask: in std_logic_vector((g_data_width/8)-1 downto 0);
           enable: in std_logic;
           writebar : in std_logic;
           clk: in std_logic;
           reset : in std_logic);
	end component;
begin
	
	stall_signal <= (fin_ack_sig and (not fin_req));
	enable_sig <= (not stall_signal) and start_req;
	start_ack  <= enable_sig;

	memInst: generic_single_port_memory_with_byte_mask
			generic map (name => "GenericMem2MB",
					g_addr_width => 19,
					g_data_width => 64)
			port map (
					datain => write_data,
					dataout => read_data,
					addrin => address(18 downto 0),
					bytemask => byte_mask,
					enable => enable_sig,
					writebar => read_write_bar(0),
					clk => clk, 
					reset => reset);

	process(clk)
	begin 
		if(clk'event and (clk = '1')) then
			if(reset = '1') then
				fin_ack_sig <= '0';
				tag_out <= (others => '0');
			elsif (enable_sig = '1') then
				tag_out <= tag_in;
				fin_ack_sig <= '1';
			else
				fin_ack_sig <= '0';
			end if;
		end if;
	end process;

	fin_ack <= fin_ack_sig;
end Mixed;
		
-- THIS IS TO BE USED ONLY FOR SIMULATIONS!
library std;
use std.textio.all;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.BaseComponents.all;
use ahir.mem_component_pack.all;
use ahir.Utilities.all;

library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
use AjitCustom.MemmapPackage.all;

entity single_port_16kX64_memory_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    read : in  std_logic_vector(0 downto 0);
    -- 16K dwords..= 128KB
    addr : in  std_logic_vector(16 downto 0);
    byte_mask : in  std_logic_vector(7 downto 0);
    write_data : in  std_logic_vector(63 downto 0);
    read_data : out  std_logic_vector(63 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity single_port_16kX64_memory_Operator;

architecture single_port_16kX64_memory_Operator_arch of single_port_16kX64_memory_Operator is -- 
	signal joined_sig: boolean;	
 	signal enable: std_logic;
begin --  

    trig_join: join2 generic map (name => "single_port_16xK64_memory_Operator:trig-join", bypass => true)
			port map (pred0 => sample_req, pred1 => update_req,
					symbol_out => joined_sig, clk => clk, reset => reset);
   
    sample_ack <= joined_sig;

    process(clk, reset)
    begin
	if(clk'event and clk='1') then
		if(reset = '1') then
			update_ack <= false;
		else
			update_ack <= joined_sig;
		end if;
	end if;
    end process;

    enable <= '1' when joined_sig else '0';

    -- the base-bank
    bb:  generic_single_port_memory_with_byte_mask
		generic map (name => "single_port_16kX64_memory_Operator:bb",
				g_addr_width => 14, g_data_width => 64)
		port map (
	   		datain => write_data,
           		dataout => read_data,
			-- dword address!
           		addrin => addr(16 downto 3),
	   		bytemask => byte_mask,
           		enable => enable,
           		writebar => read(0),
           		clk => clk, 
           		reset => reset);
			

end single_port_16kX64_memory_Operator_arch;
-- THIS IS TO BE USED ONLY FOR SIMULATIONS!
library std;
use std.textio.all;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.BaseComponents.all;
use ahir.mem_component_pack.all;
use ahir.Utilities.all;

library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
use AjitCustom.MemmapPackage.all;

-- NOTE: only for simulations.
entity single_port_u64_mem_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    read : in  std_logic_vector(0 downto 0);
    -- 8K dwords..= 64KB
    addr : in  std_logic_vector(12 downto 0);
    byte_mask : in  std_logic_vector(7 downto 0);
    write_data : in  std_logic_vector(63 downto 0);
    read_data : out  std_logic_vector(63 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity single_port_u64_mem_Operator;

architecture single_port_u64_mem_Operator_arch of single_port_u64_mem_Operator is -- 
	type MemArray is array (natural range <>) of std_logic_vector(63 downto 0);
	signal joined_sig: boolean;	
begin --  

    trig_join: join2 generic map (name => "single_port_u64_mem_Operator:trig-join", bypass => true)
			port map (pred0 => sample_req, pred1 => update_req,
					symbol_out => joined_sig, clk => clk, reset => reset);
   
    sample_ack <= joined_sig;

    process(clk, reset)
    begin
	if(clk'event and clk='1') then
		if(reset = '1') then
			update_ack <= false;
		else
			update_ack <= joined_sig;
		end if;
	end if;
    end process;

    -- ports
    process(clk, reset, joined_sig, read, addr, byte_mask, write_data)
	-- 8k X 64B.  double word address is 13 bits (truncated).
	variable mem_array: MemArray (0 to 8191);
	variable tval: std_logic_vector(63 downto 0);
    begin
	if(clk'event and clk = '1') then
		if(reset = '1') then
			read_data <= (others => '0');
		else
			if(joined_sig) then
				if(read(0) = '1') then
					read_data <= mem_array(to_integer(unsigned(addr(12 downto 0))));
				else
					tval :=  mem_array(to_integer(unsigned(addr(12 downto 0))));
					mem_array(to_integer(unsigned(addr(12 downto 0)))) :=
							updateU64UsingByteMask(tval, byte_mask, write_data);
				end if;  
			end if; -- joined_sig
		end if;
	end if;
    end process;

end single_port_u64_mem_Operator_arch;
--
-- ROMs Using Block RAM Resources.
-- VHDL code for a ROM with registered output (template 1)
--   Adapted from Xilinx xst user guide by Madhav Desai.
--
library ieee;                                                         
use ieee.std_logic_1164.all;                                          
use ieee.numeric_std.all; 

library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
use AjitCustom.RomPackage.all;

-- 64 KB ROM.
entity ajit_64kB_rom is                                                     
    port (clk  : in std_logic;                                                   
          en   : in std_logic;                                                    
          addr : in std_logic_vector(15 downto 0);                               
          data : out std_logic_vector(7 downto 0));                             
end ajit_64kB_rom;                                                          

architecture xilinx_rom_infer of ajit_64kB_rom is                                        
    signal ROM :  AJIT_ROM_TYPE := ROM_INITIAL_VALUE; -- from RomPackage
begin                                                                 
    process (clk)                                                         
    begin                                                                 
        if (clk'event and clk = '1') then                                     
            if (en = '1') then                                                    
                data <= ROM(to_integer(unsigned(addr)));                                       
            end if;                                                               
        end if;                                                               
    end process;
end xilinx_rom_infer;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library AjitCustom;
use AjitCustom.MemmapPackage.all;

entity dual_port_byte_ram_with_init is
   generic (byte_position: integer; g_addr_width: natural := 10; init_byte_array: ByteArray);
   port (
    	 datain_0 : in std_logic_vector(8-1 downto 0);
         dataout_0: out std_logic_vector(8-1 downto 0);
         addrin_0: in std_logic_vector(g_addr_width-1 downto 0);
         enable_0: in std_logic;
         writebar_0 : in std_logic;
    	 datain_1 : in std_logic_vector(8-1 downto 0);
         dataout_1: out std_logic_vector(8-1 downto 0);
         addrin_1: in std_logic_vector(g_addr_width-1 downto 0);
         enable_1: in std_logic;
         writebar_1 : in std_logic;
         clk: in std_logic;
         reset : in std_logic);
end entity dual_port_byte_ram_with_init;


architecture XilinxBramInfer of dual_port_byte_ram_with_init is

  signal mem_array : ByteArray(0 to (2**g_addr_width)-1) :=  init_byte_array;
  signal addr_reg_0, addr_reg_1 : std_logic_vector(g_addr_width-1 downto 0);
  signal rd_enable_reg_0, rd_enable_reg_1 : std_logic;
  signal read_data_0, read_data_reg_0: std_logic_vector(8-1 downto 0);
  signal read_data_1, read_data_reg_1: std_logic_vector(8-1 downto 0);
begin  -- XilinxBramInfer

  -- read/write process
  process(clk,addrin_0,enable_0,writebar_0, datain_0, addrin_1, enable_1, writebar_1, datain_1)
  begin

    -- synch read-write memory
    if(clk'event and clk ='1') then

     	-- register the address
	-- and use it in a separate assignment
	-- for the delayed read.
      addr_reg_0 <= addrin_0;
      addr_reg_1 <= addrin_1;

	-- generate a registered read enable
      if(reset = '1') then
	rd_enable_reg_0 <= '0';
	rd_enable_reg_1 <= '0';
      else
	rd_enable_reg_0 <= enable_0 and writebar_0;
	rd_enable_reg_1 <= enable_1 and writebar_1;
      end if;

      if(enable_0 = '1' and writebar_0 = '0') then
        mem_array(To_Integer(unsigned(addrin_0))) <= datain_0;
      end if;
      if(enable_1 = '1' and writebar_1 = '0') then
        mem_array(To_Integer(unsigned(addrin_1))) <= datain_1;
      end if;
    end if;
  end process;

  -- read data.
  read_data_0 <= mem_array(To_Integer(unsigned(addr_reg_0)));
  read_data_1 <= mem_array(To_Integer(unsigned(addr_reg_1)));
  process(clk) 
  begin
	if(clk'event and clk = '1') then
		if(rd_enable_reg_0 = '1') then
			read_data_reg_0 <= read_data_0;
		end if;
		if(rd_enable_reg_1 = '1') then
			read_data_reg_1 <= read_data_1;
		end if;
	end if;
  end process;

  -- to maintain dataout to the last value that was read!
  dataout_0 <= read_data_0 when (rd_enable_reg_0 = '1') else read_data_reg_0;
  dataout_1 <= read_data_1 when (rd_enable_reg_1 = '1') else read_data_reg_1;

end XilinxBramInfer;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library AjitCustom;
use AjitCustom.MemmapPackage.all;

entity single_port_byte_ram_with_init is
   generic (byte_position: integer; g_addr_width: natural := 10; init_byte_array: ByteArray);
   port (
    	 datain : in std_logic_vector(8-1 downto 0);
         dataout: out std_logic_vector(8-1 downto 0);
         addrin: in std_logic_vector(g_addr_width-1 downto 0);
         enable: in std_logic;
         writebar : in std_logic;
         clk: in std_logic;
         reset : in std_logic);
end entity single_port_byte_ram_with_init;


architecture XilinxBramInfer of single_port_byte_ram_with_init is

  signal mem_array : ByteArray(0 to (2**g_addr_width)-1) :=  init_byte_array;
  signal addr_reg: std_logic_vector(g_addr_width-1 downto 0);
  signal rd_enable_reg: std_logic;
  signal read_data, read_data_reg: std_logic_vector(8-1 downto 0);
begin  -- XilinxBramInfer

  -- read/write process
  process(clk,addrin,enable,writebar, datain, addrin)
  begin

    -- synch read-write memory
    if(clk'event and clk ='1') then

     	-- register the address
	-- and use it in a separate assignment
	-- for the delayed read.
      addr_reg <= addrin;

	-- generate a registered read enable
      if(reset = '1') then
	rd_enable_reg <= '0';
      else
	rd_enable_reg <= enable and writebar;
      end if;

      if(enable = '1' and writebar = '0') then
        mem_array(To_Integer(unsigned(addrin))) <= datain;
      end if;
    end if;
  end process;

  -- read data.
  read_data <= mem_array(To_Integer(unsigned(addr_reg)));
  process(clk) 
  begin
	if(clk'event and clk = '1') then
		if(rd_enable_reg = '1') then
			read_data_reg <= read_data;
		end if;
	end if;
  end process;

  -- to maintain dataout to the last value that was read!
  dataout <= read_data when (rd_enable_reg = '1') else read_data_reg;

end XilinxBramInfer;
library std;
use std.textio.all;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.utilities.all;

library AjitCustom;
use AjitCustom.MemmapPackage.all;


entity byte_ram_with_mmap_init is
   generic (mmap_file_name: string; g_addr_width: natural := 10);
   port (datain : in std_logic_vector(8-1 downto 0);
         dataout: out std_logic_vector(8-1 downto 0);
         addrin: in std_logic_vector(g_addr_width-1 downto 0);
         enable: in std_logic;
         writebar : in std_logic;
         clk: in std_logic;
         reset : in std_logic);
end entity byte_ram_with_mmap_init;


architecture XilinxBramInfer of byte_ram_with_mmap_init is

  signal addr_reg : std_logic_vector(g_addr_width-1 downto 0);
  signal rd_enable_reg : std_logic;
  signal read_data, read_data_reg: std_logic_vector(8-1 downto 0);
  

begin  -- XilinxBramInfer

  -- read/write process
  process(clk,addrin,enable,writebar,addr_reg)
    
  	-- will be initialized below... 
  	variable mem_array : ByteArray(0 to (2**g_addr_width)-1);
    	variable bit_data_var : bit_vector(7 downto 0);
    	variable slv_data_var : std_logic_vector(7 downto 0);
	variable address_var: integer;

    	File INFILE: text open read_mode is mmap_file_name;
    	variable INPUT_LINE: Line;
    	variable r_line_count: integer;
  	variable init_done: std_logic := '0';
  begin

    -- initialization, one time.
    if(init_done = '0') then
		init_done := '1';

		assert false report "Reading MMAP file " & mmap_file_name severity note;
    		r_line_count := 0;
		while not endfile (INFILE) loop
	  		readLine (INFILE, INPUT_LINE);
         		read (INPUT_LINE, address_var);
          		read (INPUT_LINE, bit_data_var);
			
			slv_data_var := to_std_logic_vector(bit_data_var);
	 
  	  		if((address_var >= 0) and (address_var < mem_array'length)) then
				mem_array(address_var) := slv_data_var;
			end if;
			-- assert false report "mem[" & Convert_To_String(address_var) & "] = " & 
		 	--	Convert_SLV_To_String (slv_data_var) severity note;

 	  		r_line_count := r_line_count + 1;
		end loop;
		assert false report "Finished Reading MMAP file " & mmap_file_name  & ": read  " &
					Convert_To_String(r_line_count)  & " lines"
										severity note;
    end if;

    -- read-data..
    read_data <= mem_array(To_Integer(unsigned(addr_reg)));

    if(clk'event and clk ='1') then
     	-- register the address
	-- and use it in a separate assignment
	-- for the delayed read.
      addr_reg <= addrin;

	-- generate a registered read enable
      if(reset = '1') then
	rd_enable_reg <= '0';
      else
	rd_enable_reg <= enable and writebar;
      end if;

      if(enable = '1' and writebar = '0') then
        mem_array(To_Integer(unsigned(addrin))) := datain;
      end if;
    end if;
  end process;

  -- read data.
  process(clk) 
  begin
	if(clk'event and clk = '1') then
		if(rd_enable_reg = '1') then
			read_data_reg <= read_data;
		end if;
	end if;
  end process;

  -- to maintain dataout to the last value that was read!
  dataout <= read_data when (rd_enable_reg = '1') else read_data_reg;

end XilinxBramInfer;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.OperatorPackage.all;
entity isIcacheFlushAsi_VVV is -- 
  port ( -- 
    asi : in  std_logic_vector(7 downto 0);
    ret_val : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity isIcacheFlushAsi_VVV;
architecture isIcacheFlushAsi_VVV_arch of isIcacheFlushAsi_VVV is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(8-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal asi_buffer :  std_logic_vector(7 downto 0);
  -- output port buffer signals
  signal ret_val_buffer :  std_logic_vector(0 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  asi_buffer <= asi;
  -- output handling  -------------------------------------------------------
  ret_val <= ret_val_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal UGE_u8_u1_623_wire : std_logic_vector(0 downto 0);
    signal ULE_u8_u1_626_wire : std_logic_vector(0 downto 0);
    signal konst_622_wire_constant : std_logic_vector(7 downto 0);
    signal konst_625_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    konst_622_wire_constant <= "00011000";
    konst_625_wire_constant <= "00011100";
    -- binary operator AND_u1_u1_627_inst
    process(UGE_u8_u1_623_wire, ULE_u8_u1_626_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(UGE_u8_u1_623_wire, ULE_u8_u1_626_wire, tmp_var);
      ret_val_buffer <= tmp_var; -- 
    end process;
    -- binary operator UGE_u8_u1_623_inst
    process(asi_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUge_proc(asi_buffer, konst_622_wire_constant, tmp_var);
      UGE_u8_u1_623_wire <= tmp_var; -- 
    end process;
    -- binary operator ULE_u8_u1_626_inst
    process(asi_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUle_proc(asi_buffer, konst_625_wire_constant, tmp_var);
      ULE_u8_u1_626_wire <= tmp_var; -- 
    end process;
    -- 
  end Block; -- data_path
  -- 
end isIcacheFlushAsi_VVV_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.operatorpackage.all;
entity isIcacheFlushLineOnly_VVV is -- 
  port ( -- 
    asi : in  std_logic_vector(7 downto 0);
    flush_line_only : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity isIcacheFlushLineOnly_VVV;
architecture isIcacheFlushLineOnly_VVV_arch of isIcacheFlushLineOnly_VVV is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(8-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal asi_buffer :  std_logic_vector(7 downto 0);
  -- output port buffer signals
  signal flush_line_only_buffer :  std_logic_vector(0 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  asi_buffer <= asi;
  -- output handling  -------------------------------------------------------
  flush_line_only <= flush_line_only_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal EQ_u8_u1_850_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_853_wire : std_logic_vector(0 downto 0);
    signal R_ASI_FLUSH_I_D_USER_852_wire_constant : std_logic_vector(7 downto 0);
    signal R_ASI_FLUSH_I_USER_849_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    R_ASI_FLUSH_I_D_USER_852_wire_constant <= "00010100";
    R_ASI_FLUSH_I_USER_849_wire_constant <= "00011100";
    -- binary operator EQ_u8_u1_850_inst
    process(asi_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(asi_buffer, R_ASI_FLUSH_I_USER_849_wire_constant, tmp_var);
      EQ_u8_u1_850_wire <= tmp_var; -- 
    end process;
    -- binary operator EQ_u8_u1_853_inst
    process(asi_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(asi_buffer, R_ASI_FLUSH_I_D_USER_852_wire_constant, tmp_var);
      EQ_u8_u1_853_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_854_inst
    process(EQ_u8_u1_850_wire, EQ_u8_u1_853_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u8_u1_850_wire, EQ_u8_u1_853_wire, tmp_var);
      flush_line_only_buffer <= tmp_var; -- 
    end process;
    -- 
  end Block; -- data_path
  -- 
end isIcacheFlushLineOnly_VVV_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library ahir;
use ahir.OperatorPackage.all;

entity isIcacheInstructionFetch_VVV is -- 
  port ( -- 
    asi : in  std_logic_vector(7 downto 0);
    ret_val : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity isIcacheInstructionFetch_VVV;
architecture isIcacheInstructionFetch_VVV_arch of isIcacheInstructionFetch_VVV is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(8-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal asi_buffer :  std_logic_vector(7 downto 0);
  -- output port buffer signals
  signal ret_val_buffer :  std_logic_vector(0 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  asi_buffer <= asi;
  -- output handling  -------------------------------------------------------
  ret_val <= ret_val_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal EQ_u8_u1_610_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_613_wire : std_logic_vector(0 downto 0);
    signal R_ASI_SUPERVISOR_INSTRUCTION_612_wire_constant : std_logic_vector(7 downto 0);
    signal R_ASI_USER_INSTRUCTION_609_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    R_ASI_SUPERVISOR_INSTRUCTION_612_wire_constant <= "00001001";
    R_ASI_USER_INSTRUCTION_609_wire_constant <= "00001000";
    -- binary operator EQ_u8_u1_610_inst
    process(asi_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(asi_buffer, R_ASI_USER_INSTRUCTION_609_wire_constant, tmp_var);
      EQ_u8_u1_610_wire <= tmp_var; -- 
    end process;
    -- binary operator EQ_u8_u1_613_inst
    process(asi_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(asi_buffer, R_ASI_SUPERVISOR_INSTRUCTION_612_wire_constant, tmp_var);
      EQ_u8_u1_613_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_614_inst
    process(EQ_u8_u1_610_wire, EQ_u8_u1_613_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u8_u1_610_wire, EQ_u8_u1_613_wire, tmp_var);
      ret_val_buffer <= tmp_var; -- 
    end process;
    -- 
  end Block; -- data_path
  -- 
end isIcacheInstructionFetch_VVV_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.operatorpackage.all;
entity isIcacheSupervisorAsi_VVV is -- 
  port ( -- 
    asi : in  std_logic_vector(7 downto 0);
    ret_val : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity isIcacheSupervisorAsi_VVV;
architecture isIcacheSupervisorAsi_VVV_arch of isIcacheSupervisorAsi_VVV is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(8-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal asi_buffer :  std_logic_vector(7 downto 0);
  -- output port buffer signals
  signal ret_val_buffer :  std_logic_vector(0 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  asi_buffer <= asi;
  -- output handling  -------------------------------------------------------
  ret_val <= ret_val_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal R_ASI_SUPERVISOR_INSTRUCTION_635_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    R_ASI_SUPERVISOR_INSTRUCTION_635_wire_constant <= "00001001";
    -- binary operator EQ_u8_u1_636_inst
    process(asi_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(asi_buffer, R_ASI_SUPERVISOR_INSTRUCTION_635_wire_constant, tmp_var);
      ret_val_buffer <= tmp_var; -- 
    end process;
    -- 
  end Block; -- data_path
  -- 
end isIcacheSupervisorAsi_VVV_arch;

library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.operatorpackage.all;

entity analyzeBeResponse is -- 
  port ( -- 
    from_backend : in  std_logic_vector(101 downto 0);
    be_valid : out  std_logic_vector(0 downto 0);
    be_counter : out  std_logic_vector(2 downto 0);
    be_dword_id : out  std_logic_vector(2 downto 0);
    be_last_dword : out  std_logic_vector(0 downto 0);
    be_mae : out  std_logic_vector(0 downto 0);
    be_access_error : out  std_logic_vector(0 downto 0);
    be_acc : out  std_logic_vector(2 downto 0);
    be_tag_cmd : out  std_logic_vector(2 downto 0);
    be_array_cmd : out  std_logic_vector(2 downto 0);
    be_mmu_fsr : out  std_logic_vector(17 downto 0);
    be_dword : out  std_logic_vector(63 downto 0)-- 
  );
  -- 
end entity analyzeBeResponse;

architecture analyze_backend_response_Volatile_arch of analyzeBeResponse is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(102-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal from_backend_buffer :  std_logic_vector(101 downto 0);
  -- output port buffer signals
  signal be_valid_buffer :  std_logic_vector(0 downto 0);
  signal be_counter_buffer :  std_logic_vector(2 downto 0);
  signal be_dword_id_buffer :  std_logic_vector(2 downto 0);
  signal be_last_dword_buffer :  std_logic_vector(0 downto 0);
  signal be_mae_buffer :  std_logic_vector(0 downto 0);
  signal be_access_error_buffer :  std_logic_vector(0 downto 0);
  signal be_acc_buffer :  std_logic_vector(2 downto 0);
  signal be_tag_cmd_buffer :  std_logic_vector(2 downto 0);
  signal be_array_cmd_buffer :  std_logic_vector(2 downto 0);
  signal be_mmu_fsr_buffer :  std_logic_vector(17 downto 0);
  signal be_dword_buffer :  std_logic_vector(63 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  from_backend_buffer <= from_backend;
  -- output handling  -------------------------------------------------------
  be_valid <= be_valid_buffer;
  be_counter <= be_counter_buffer;
  be_dword_id <= be_dword_id_buffer;
  be_last_dword <= be_last_dword_buffer;
  be_mae <= be_mae_buffer;
  be_access_error <= be_access_error_buffer;
  be_acc <= be_acc_buffer;
  be_tag_cmd <= be_tag_cmd_buffer;
  be_array_cmd <= be_array_cmd_buffer;
  be_mmu_fsr <= be_mmu_fsr_buffer;
  be_dword <= be_dword_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal be_cacheable_1013 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    -- flow-through slice operator slice_1000_inst
    be_dword_id_buffer <= from_backend_buffer(91 downto 89);
    -- flow-through slice operator slice_1004_inst
    be_last_dword_buffer <= from_backend_buffer(88 downto 88);
    -- flow-through slice operator slice_1008_inst
    be_acc_buffer <= from_backend_buffer(87 downto 85);
    -- flow-through slice operator slice_1012_inst
    be_cacheable_1013 <= from_backend_buffer(84 downto 84);
    -- flow-through slice operator slice_1016_inst
    be_mae_buffer <= from_backend_buffer(83 downto 83);
    -- flow-through slice operator slice_1020_inst
    be_access_error_buffer <= from_backend_buffer(82 downto 82);
    -- flow-through slice operator slice_1024_inst
    be_mmu_fsr_buffer <= from_backend_buffer(81 downto 64);
    -- flow-through slice operator slice_1028_inst
    be_dword_buffer <= from_backend_buffer(63 downto 0);
    -- flow-through slice operator slice_984_inst
    be_valid_buffer <= from_backend_buffer(101 downto 101);
    -- flow-through slice operator slice_988_inst
    be_counter_buffer <= from_backend_buffer(100 downto 98);
    -- flow-through slice operator slice_992_inst
    be_tag_cmd_buffer <= from_backend_buffer(97 downto 95);
    -- flow-through slice operator slice_996_inst
    be_array_cmd_buffer <= from_backend_buffer(94 downto 92);
    -- 
  end Block; -- data_path
  -- 
end analyze_backend_response_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.operatorpackage.all;
entity classifyCpuSideRequests is -- 
  port ( -- 
    from_cpu_ifetch : in  std_logic_vector(40 downto 0);
    cpu_valid : out  std_logic_vector(0 downto 0);
    cpu_ifetch_valid : out  std_logic_vector(0 downto 0);
    exec_cpu_ifetch : out  std_logic_vector(0 downto 0);
    exec_cpu_new_stream_flush : out  std_logic_vector(0 downto 0);
    exec_cpu_flush : out  std_logic_vector(0 downto 0);
    exec_cpu_S : out  std_logic_vector(0 downto 0);
    exec_cpu_tag_command : out  std_logic_vector(2 downto 0);
    exec_cpu_array_command : out  std_logic_vector(2 downto 0);
    exec_cpu_asi : out  std_logic_vector(7 downto 0);
    exec_cpu_addr : out  std_logic_vector(31 downto 0)-- 
  );
  -- 
end entity classifyCpuSideRequests;
architecture classify_cpu_side_requests_VVV_arch of classifyCpuSideRequests is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(41-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal from_cpu_ifetch_buffer :  std_logic_vector(40 downto 0);
  -- output port buffer signals
  signal cpu_valid_buffer :  std_logic_vector(0 downto 0);
  signal cpu_ifetch_valid_buffer :  std_logic_vector(0 downto 0);
  signal exec_cpu_ifetch_buffer :  std_logic_vector(0 downto 0);
  signal exec_cpu_new_stream_flush_buffer :  std_logic_vector(0 downto 0);
  signal exec_cpu_flush_buffer :  std_logic_vector(0 downto 0);
  signal exec_cpu_S_buffer :  std_logic_vector(0 downto 0);
  signal exec_cpu_tag_command_buffer :  std_logic_vector(2 downto 0);
  signal exec_cpu_array_command_buffer :  std_logic_vector(2 downto 0);
  signal exec_cpu_asi_buffer :  std_logic_vector(7 downto 0);
  signal exec_cpu_addr_buffer :  std_logic_vector(31 downto 0);
  -- volatile/operator module components. 
  component isIcacheFlushLineOnly_VVV is -- 
    port ( -- 
      asi : in  std_logic_vector(7 downto 0);
      flush_line_only : out  std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component; 
  component isIcacheInstructionFetch_VVV is -- 
    port ( -- 
      asi : in  std_logic_vector(7 downto 0);
      ret_val : out  std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component; 
  component isIcacheFlushAsi_VVV is -- 
    port ( -- 
      asi : in  std_logic_vector(7 downto 0);
      ret_val : out  std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component; 
  component isIcacheSupervisorAsi_VVV is -- 
    port ( -- 
      asi : in  std_logic_vector(7 downto 0);
      ret_val : out  std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component; 
  -- 
begin --  
  -- input handling ------------------------------------------------
  from_cpu_ifetch_buffer <= from_cpu_ifetch;
  -- output handling  -------------------------------------------------------
  cpu_valid <= cpu_valid_buffer;
  cpu_ifetch_valid <= cpu_ifetch_valid_buffer;
  exec_cpu_ifetch <= exec_cpu_ifetch_buffer;
  exec_cpu_new_stream_flush <= exec_cpu_new_stream_flush_buffer;
  exec_cpu_flush <= exec_cpu_flush_buffer;
  exec_cpu_S <= exec_cpu_S_buffer;
  exec_cpu_tag_command <= exec_cpu_tag_command_buffer;
  exec_cpu_array_command <= exec_cpu_array_command_buffer;
  exec_cpu_asi <= exec_cpu_asi_buffer;
  exec_cpu_addr <= exec_cpu_addr_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal MUX_941_wire : std_logic_vector(2 downto 0);
    signal MUX_945_wire : std_logic_vector(2 downto 0);
    signal MUX_956_wire : std_logic_vector(2 downto 0);
    signal OR_u1_u1_937_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_951_wire : std_logic_vector(0 downto 0);
    signal R_CACHE_ARRAY_NOP_952_wire_constant : std_logic_vector(2 downto 0);
    signal R_CACHE_ARRAY_NOP_955_wire_constant : std_logic_vector(2 downto 0);
    signal R_CACHE_ARRAY_READ_DWORD_954_wire_constant : std_logic_vector(2 downto 0);
    signal R_CACHE_TAG_CLEAR_ALL_940_wire_constant : std_logic_vector(2 downto 0);
    signal R_CACHE_TAG_CLEAR_LINE_939_wire_constant : std_logic_vector(2 downto 0);
    signal R_CACHE_TAG_LOOKUP_943_wire_constant : std_logic_vector(2 downto 0);
    signal R_CACHE_TAG_NOP_944_wire_constant : std_logic_vector(2 downto 0);
    signal cpu_S_904 : std_logic_vector(0 downto 0);
    signal cpu_ifetch_addr_880 : std_logic_vector(31 downto 0);
    signal flush_line_933 : std_logic_vector(0 downto 0);
    signal flush_line_only_910 : std_logic_vector(0 downto 0);
    signal is_flush_asi_907 : std_logic_vector(0 downto 0);
    signal is_ifetch_asi_913 : std_logic_vector(0 downto 0);
    signal konst_891_wire_constant : std_logic_vector(7 downto 0);
    signal konst_896_wire_constant : std_logic_vector(7 downto 0);
    signal r_cpu_ifetch_asi_876 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    R_CACHE_ARRAY_NOP_952_wire_constant <= "100";
    R_CACHE_ARRAY_NOP_955_wire_constant <= "100";
    R_CACHE_ARRAY_READ_DWORD_954_wire_constant <= "001";
    R_CACHE_TAG_CLEAR_ALL_940_wire_constant <= "100";
    R_CACHE_TAG_CLEAR_LINE_939_wire_constant <= "011";
    R_CACHE_TAG_LOOKUP_943_wire_constant <= "001";
    R_CACHE_TAG_NOP_944_wire_constant <= "101";
    konst_891_wire_constant <= "01111111";
    konst_896_wire_constant <= "00000111";
    -- flow-through select operator MUX_941_inst
    MUX_941_wire <= R_CACHE_TAG_CLEAR_LINE_939_wire_constant when (flush_line_933(0) /=  '0') else R_CACHE_TAG_CLEAR_ALL_940_wire_constant;
    -- flow-through select operator MUX_945_inst
    MUX_945_wire <= R_CACHE_TAG_LOOKUP_943_wire_constant when (exec_cpu_ifetch_buffer(0) /=  '0') else R_CACHE_TAG_NOP_944_wire_constant;
    -- flow-through select operator MUX_946_inst
    exec_cpu_tag_command_buffer <= MUX_941_wire when (OR_u1_u1_937_wire(0) /=  '0') else MUX_945_wire;
    -- flow-through select operator MUX_956_inst
    MUX_956_wire <= R_CACHE_ARRAY_READ_DWORD_954_wire_constant when (exec_cpu_ifetch_buffer(0) /=  '0') else R_CACHE_ARRAY_NOP_955_wire_constant;
    -- flow-through select operator MUX_957_inst
    exec_cpu_array_command_buffer <= R_CACHE_ARRAY_NOP_952_wire_constant when (OR_u1_u1_951_wire(0) /=  '0') else MUX_956_wire;
    -- flow-through slice operator slice_871_inst
    cpu_ifetch_valid_buffer <= from_cpu_ifetch_buffer(40 downto 40);
    -- flow-through slice operator slice_875_inst
    r_cpu_ifetch_asi_876 <= from_cpu_ifetch_buffer(39 downto 32);
    -- flow-through slice operator slice_879_inst
    cpu_ifetch_addr_880 <= from_cpu_ifetch_buffer(31 downto 0);
    -- interlock W_cpu_valid_886_inst
    process(cpu_ifetch_valid_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := cpu_ifetch_valid_buffer(0 downto 0);
      cpu_valid_buffer <= tmp_var; -- 
    end process;
    -- interlock W_exec_cpu_addr_899_inst
    process(cpu_ifetch_addr_880) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := cpu_ifetch_addr_880(31 downto 0);
      exec_cpu_addr_buffer <= tmp_var; -- 
    end process;
    -- binary operator AND_u1_u1_917_inst
    process(cpu_valid_buffer, is_flush_asi_907) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cpu_valid_buffer, is_flush_asi_907, tmp_var);
      exec_cpu_flush_buffer <= tmp_var; -- 
    end process;
    -- binary operator AND_u1_u1_922_inst
    process(cpu_valid_buffer, is_ifetch_asi_913) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cpu_valid_buffer, is_ifetch_asi_913, tmp_var);
      exec_cpu_ifetch_buffer <= tmp_var; -- 
    end process;
    -- binary operator AND_u1_u1_927_inst
    process(cpu_valid_buffer, cpu_S_904) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(cpu_valid_buffer, cpu_S_904, tmp_var);
      exec_cpu_S_buffer <= tmp_var; -- 
    end process;
    -- binary operator AND_u1_u1_932_inst
    process(exec_cpu_flush_buffer, flush_line_only_910) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(exec_cpu_flush_buffer, flush_line_only_910, tmp_var);
      flush_line_933 <= tmp_var; -- 
    end process;
    -- binary operator AND_u8_u8_892_inst
    process(r_cpu_ifetch_asi_876) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAnd_proc(r_cpu_ifetch_asi_876, konst_891_wire_constant, tmp_var);
      exec_cpu_asi_buffer <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_897_inst
    process(r_cpu_ifetch_asi_876) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(r_cpu_ifetch_asi_876, konst_896_wire_constant, tmp_var);
      exec_cpu_new_stream_flush_buffer <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_937_inst
    process(exec_cpu_new_stream_flush_buffer, exec_cpu_flush_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(exec_cpu_new_stream_flush_buffer, exec_cpu_flush_buffer, tmp_var);
      OR_u1_u1_937_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_951_inst
    process(exec_cpu_flush_buffer, exec_cpu_new_stream_flush_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(exec_cpu_flush_buffer, exec_cpu_new_stream_flush_buffer, tmp_var);
      OR_u1_u1_951_wire <= tmp_var; -- 
    end process;
    volatile_operator_isIcacheSupervisorAsi_1021: isIcacheSupervisorAsi_VVV port map(asi => exec_cpu_asi_buffer, ret_val => cpu_S_904); 
    volatile_operator_isIcacheFlushAsi_1022: isIcacheFlushAsi_VVV port map(asi => exec_cpu_asi_buffer, ret_val => is_flush_asi_907); 
    volatile_operator_isIcacheFlushLineOnly_1023: isIcacheFlushLineOnly_VVV port map(asi => exec_cpu_asi_buffer, flush_line_only => flush_line_only_910); 
    volatile_operator_isIcacheInstructionFetch_1024: isIcacheInstructionFetch_VVV port map(asi => exec_cpu_asi_buffer, ret_val => is_ifetch_asi_913); 
    -- 
  end Block; -- data_path
  -- 
end classify_cpu_side_requests_VVV_arch;
-- A front-end for the icache.  Can provide response in 1 clock cycle
-- if there is a hit!

library ieee;
use ieee.std_logic_1164.all;
package icache_global_package is -- 
  constant ASI_AJIT_BRIDGE_CONFIG : std_logic_vector(7 downto 0) := "00110000";
  constant ASI_BLOCK_COPY : std_logic_vector(7 downto 0) := "00010111";
  constant ASI_BLOCK_FILL : std_logic_vector(7 downto 0) := "00011111";
  constant ASI_CACHE_DATA_I : std_logic_vector(7 downto 0) := "00001101";
  constant ASI_CACHE_DATA_I_D : std_logic_vector(7 downto 0) := "00001111";
  constant ASI_CACHE_TAG_I : std_logic_vector(7 downto 0) := "00001100";
  constant ASI_CACHE_TAG_I_D : std_logic_vector(7 downto 0) := "00001110";
  constant ASI_FLUSH_I_CONTEXT : std_logic_vector(7 downto 0) := "00011011";
  constant ASI_FLUSH_I_D_CONTEXT : std_logic_vector(7 downto 0) := "00010011";
  constant ASI_FLUSH_I_D_PAGE : std_logic_vector(7 downto 0) := "00010000";
  constant ASI_FLUSH_I_D_REGION : std_logic_vector(7 downto 0) := "00010010";
  constant ASI_FLUSH_I_D_SEGMENT : std_logic_vector(7 downto 0) := "00010001";
  constant ASI_FLUSH_I_D_USER : std_logic_vector(7 downto 0) := "00010100";
  constant ASI_FLUSH_I_PAGE : std_logic_vector(7 downto 0) := "00011000";
  constant ASI_FLUSH_I_REGION : std_logic_vector(7 downto 0) := "00011010";
  constant ASI_FLUSH_I_SEGMENT : std_logic_vector(7 downto 0) := "00011001";
  constant ASI_FLUSH_I_USER : std_logic_vector(7 downto 0) := "00011100";
  constant ASI_MMU_DIAGNOSTIC_I : std_logic_vector(7 downto 0) := "00000101";
  constant ASI_MMU_DIAGNOSTIC_IO : std_logic_vector(7 downto 0) := "00000111";
  constant ASI_MMU_DIAGNOSTIC_I_D : std_logic_vector(7 downto 0) := "00000110";
  constant ASI_MMU_FLUSH_PROBE : std_logic_vector(7 downto 0) := "00000011";
  constant ASI_MMU_REGISTER : std_logic_vector(7 downto 0) := "00000100";
  constant ASI_SUPERVISOR_DATA : std_logic_vector(7 downto 0) := "00001011";
  constant ASI_SUPERVISOR_INSTRUCTION : std_logic_vector(7 downto 0) := "00001001";
  constant ASI_USER_DATA : std_logic_vector(7 downto 0) := "00001010";
  constant ASI_USER_INSTRUCTION : std_logic_vector(7 downto 0) := "00001000";
  constant CACHE_ARRAY_READ_DWORD : std_logic_vector(2 downto 0) := "001";
  constant CACHE_ARRAY_WRITE_DWORD : std_logic_vector(2 downto 0) := "010";
  constant CACHE_ARRAY_NOP : std_logic_vector(2 downto 0) := "011";
  constant CACHE_TAG_CLEAR_ALL : std_logic_vector(2 downto 0) := "100";
  constant CACHE_TAG_CLEAR_LINE : std_logic_vector(2 downto 0) := "011";
  constant CACHE_TAG_INSERT : std_logic_vector(2 downto 0) := "010";
  constant CACHE_TAG_LOOKUP : std_logic_vector(2 downto 0) := "001";
  constant CACHE_TAG_NOP : std_logic_vector(2 downto 0) := "101";
  constant MMU_PASS_THROUGH_HLIMIT : std_logic_vector(7 downto 0) := "00101111";
  constant MMU_PASS_THROUGH_LLIMIT : std_logic_vector(7 downto 0) := "00100000";
  constant MMU_READ_DWORD : std_logic_vector(7 downto 0) := "00000010";
  constant MMU_READ_LINE : std_logic_vector(7 downto 0) := "00000011";
  constant MMU_WRITE_DWORD : std_logic_vector(7 downto 0) := "00000001";
  constant MMU_WRITE_DWORD_NO_RESPONSE : std_logic_vector(7 downto 0) := "00000101";
  constant MMU_WRITE_FSR : std_logic_vector(7 downto 0) := "00000100";
  constant REQUEST_TYPE_BRIDGE_CONFIG_READ : std_logic_vector(3 downto 0) := "1001";
  constant REQUEST_TYPE_BRIDGE_CONFIG_WRITE : std_logic_vector(3 downto 0) := "1000";
  constant REQUEST_TYPE_CCU_CACHE_READ : std_logic_vector(3 downto 0) := "0101";
  constant REQUEST_TYPE_CCU_CACHE_WRITE : std_logic_vector(3 downto 0) := "0110";
  constant REQUEST_TYPE_IFETCH : std_logic_vector(3 downto 0) := "0000";
  constant REQUEST_TYPE_NOP : std_logic_vector(3 downto 0) := "0111";
  constant REQUEST_TYPE_READ : std_logic_vector(3 downto 0) := "0001";
  constant REQUEST_TYPE_STBAR : std_logic_vector(3 downto 0) := "0011";
  constant REQUEST_TYPE_WRFSRFAR : std_logic_vector(3 downto 0) := "0100";
  constant REQUEST_TYPE_WRITE : std_logic_vector(3 downto 0) := "0010";
  constant FE_BE_COMMAND_SIZE :integer := 42; -- will be changed.
  constant BE_FE_RESPONSE_SIZE :integer := 102; -- will be changed.

  component classifyCpuSideRequests is -- 
    port ( -- 
      from_cpu_ifetch : in  std_logic_vector(40 downto 0);
      cpu_valid : out  std_logic_vector(0 downto 0);
      cpu_ifetch_valid : out  std_logic_vector(0 downto 0);
      exec_cpu_ifetch : out  std_logic_vector(0 downto 0);
      exec_cpu_new_stream_flush : out  std_logic_vector(0 downto 0);
      exec_cpu_flush : out  std_logic_vector(0 downto 0);
      exec_cpu_S : out  std_logic_vector(0 downto 0);
      exec_cpu_tag_command : out  std_logic_vector(2 downto 0);
      exec_cpu_array_command : out  std_logic_vector(2 downto 0);
      exec_cpu_asi : out  std_logic_vector(7 downto 0);
      exec_cpu_addr : out  std_logic_vector(31 downto 0)-- 
    );
    -- 
  end component; 

  component analyzeBeResponse  is -- 
   port ( -- 
    from_backend : in  std_logic_vector(101 downto 0);
    be_valid : out  std_logic_vector(0 downto 0);
    be_counter : out  std_logic_vector(2 downto 0);
    be_dword_id : out  std_logic_vector(2 downto 0);
    be_last_dword : out  std_logic_vector(0 downto 0);
    be_mae : out  std_logic_vector(0 downto 0);
    be_access_error : out  std_logic_vector(0 downto 0);
    be_acc : out  std_logic_vector(2 downto 0);
    be_tag_cmd : out  std_logic_vector(2 downto 0);
    be_array_cmd : out  std_logic_vector(2 downto 0);
    be_mmu_fsr : out  std_logic_vector(17 downto 0);
    be_dword : out  std_logic_vector(63 downto 0)-- 
   );
  end component; 

end package icache_global_package;

library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

library AjitCustom;

use AjitCustom.AjitGlobalConfigurationPackage.all;
use AjitCustom.AjitCoreConfigurationPackage.all;
use AjitCustom.icache_global_package.all;
use AjitCustom.AjitCustomComponents.all;

entity IcacheFrontendCoreDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    NOBLOCK_CPU_to_ICACHE_command_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_ICACHE_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_ICACHE_command_pipe_read_data : in   std_logic_vector(40 downto 0);
    NOBLOCK_CPU_to_ICACHE_reset_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_ICACHE_reset_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_ICACHE_reset_pipe_read_data : in   std_logic_vector(0 downto 0);
    noblock_icache_backend_to_frontend_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_icache_backend_to_frontend_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_icache_backend_to_frontend_pipe_read_data : in   std_logic_vector(101 downto 0);
    ICACHE_to_CPU_reset_ack_pipe_write_req : out  std_logic_vector(0 downto 0);
    ICACHE_to_CPU_reset_ack_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ICACHE_to_CPU_reset_ack_pipe_write_data : out  std_logic_vector(0 downto 0);
    ICACHE_to_CPU_response_pipe_write_req : out  std_logic_vector(0 downto 0);
    ICACHE_to_CPU_response_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ICACHE_to_CPU_response_pipe_write_data : out  std_logic_vector(89 downto 0);
    icache_frontend_to_backend_pipe_write_req : out  std_logic_vector(0 downto 0);
    icache_frontend_to_backend_pipe_write_ack : in   std_logic_vector(0 downto 0);
    icache_frontend_to_backend_pipe_write_data : out  std_logic_vector(41 downto 0);
    MMU_TO_ICACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_req: out std_logic_vector(0 downto 0);
    MMU_TO_ICACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_ack: in std_logic_vector(0 downto 0);
    MMU_TO_ICACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_data: in std_logic_vector(26 downto 0);
    NOBLOCK_MMU_TO_ICACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_req: out std_logic_vector(0 downto 0);
    NOBLOCK_MMU_TO_ICACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_ack: in std_logic_vector(0 downto 0);
    NOBLOCK_MMU_TO_ICACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_data: in std_logic_vector(26 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity IcacheFrontendCoreDaemon;
architecture IcacheFrontendCoreArch  of IcacheFrontEndCoreDaemon is -- system-architecture 

	constant ZERO_64 : std_logic_vector(63 downto 0) := (others => '0');
	constant ZERO_18 : std_logic_vector(17 downto 0) := (others => '0');
	constant ZERO_5 : std_logic_vector(4 downto 0) := (others => '0');
	constant mZERO_1 : std_logic_vector(0 downto 0) := (others => '0');

	Type IcacheState is (IDLE, CHECK_HIT_OR_MISS, SYN_INVALIDATE, SEND_WAIT_ON_CPU, SEND_WAIT_ON_BE, 
							RECV_WAIT_ON_BE_FIRST_DWORD, 
							RECV_WAIT_ON_BE_REMAINING_DWORDS);
	signal icache_state : IcacheState;

	-------------------------------------------------------------------------------------------
	-- predicates/inputs
	-------------------------------------------------------------------------------------------
	signal  cpu_command_available  : boolean;
	signal  cpu_reset	       : boolean;

	signal  be_is_needed	       : boolean;
	signal  expect_be_response     : boolean;
	signal  be_has_completed       : boolean;

	signal  be_ready_for_command   : boolean;
	signal  be_response_available  : boolean;
	signal  be_response_can_be_applied : boolean;
	signal  first_be_response_can_be_applied : boolean;

	signal  cpu_ready_for_response : boolean;
	signal  init_or_reset, init_or_reset_reg: boolean;

	-------------------------------------------------------------------------------------------
	-- actions/outputs
	-------------------------------------------------------------------------------------------
	signal accept_cpu_commands  : boolean;
	signal latch_cpu_commands  : boolean;
	signal clear_cpu_commands  : boolean;
	signal latch_tag_results   : boolean;
	signal latch_to_cpu	   : boolean;
	signal latch_to_be	   : boolean;
	signal accept_be_response  : boolean;
	signal write_to_be	   : boolean;
	signal write_to_cpu	   : boolean;
	signal be_latch_last_dword : boolean;
	

	signal latch_to_cpu_registered	   : boolean;
	signal latch_to_be_registered	   : boolean;

	signal send_cpu_reset_ack: boolean;
	signal accept_cpu_reset  :   boolean;

	-------------------------------------------------------------------------------------------
	-- signals, registers
	-------------------------------------------------------------------------------------------
	signal cpu_command : std_logic_vector(40 downto 0);
	signal cpu_reset_registered : boolean;
      
      	signal cpu_valid : std_logic_vector(0 downto 0);
      	signal cpu_ifetch_valid : std_logic_vector(0 downto 0);
      	signal exec_cpu_ifetch : std_logic_vector(0 downto 0);
      	signal exec_cpu_new_stream_flush : std_logic_vector(0 downto 0);
      	signal exec_cpu_flush : std_logic_vector(0 downto 0);
      	signal exec_cpu_S : std_logic_vector(0 downto 0);
      	signal exec_cpu_tag_command : std_logic_vector(2 downto 0);
      	signal exec_cpu_array_command : std_logic_vector(2 downto 0);
      	signal exec_cpu_asi : std_logic_vector(7 downto 0);
      	signal exec_cpu_addr : std_logic_vector(31 downto 0);

        -- need to remember some things about the incoming cpu command!
      	signal exec_cpu_ifetch_reg : std_logic_vector(0 downto 0);
      	signal exec_cpu_asi_reg : std_logic_vector(7 downto 0);
      	signal exec_cpu_addr_reg : std_logic_vector(31 downto 0);
      	signal exec_cpu_S_reg : std_logic_vector(0 downto 0);
      	signal cpu_ifetch_valid_reg : std_logic_vector(0 downto 0);
      	signal cpu_valid_reg: std_logic_vector(0 downto 0);
      
	signal from_backend : std_logic_vector(101 downto 0);
      	signal be_S : std_logic_vector(0 downto 0);
      	signal be_acc, access_tags_acc : std_logic_vector(2 downto 0);
      	signal be_tag_cmd : std_logic_vector(2 downto 0);
      	signal be_array_cmd : std_logic_vector(2 downto 0);
      	signal be_addr : std_logic_vector(31 downto 0);
    	signal be_counter : std_logic_vector(2 downto 0);
    	signal be_dword_id : std_logic_vector(2 downto 0);
    	signal be_last_dword : std_logic_vector(0 downto 0);
    	signal be_dword : std_logic_vector(63 downto 0);

	signal tags_arrays_trigger,  tags_arrays_done: std_logic;
	signal wait_on_tags_arrays: boolean;
	signal waiting_on_tags_arrays: boolean;

	signal access_is_read, access_is_ifetch : std_logic;

    	signal is_hit: std_logic_vector(0 downto 0);
    	signal cpu_permissions_ok: std_logic_vector(0 downto 0);
    	signal dword_out, 
			dword_out_registered, 
			instr_pair_to_cpu : std_logic_vector(63 downto 0);

	signal is_a_hit, is_a_hit_registered, is_a_hit_to_cpu, mae_to_cpu, access_error_to_cpu : std_logic_vector(0 downto 0);
	signal cacheable_to_cpu: std_logic_vector(0 downto 0);
	signal acc_to_cpu : std_logic_vector(2 downto 0);

	signal cpu_tag_lookup, cpu_tag_lookup_reg: boolean;

      	signal be_valid, be_valid_registered : std_logic_vector(0 downto 0);
      	signal be_mmu_fsr, be_mmu_fsr_registered : std_logic_vector(17 downto 0);
      	signal mmu_fsr_to_cpu: std_logic_vector(17 downto 0);
      	signal be_mae, be_mae_registered : std_logic_vector(0 downto 0);
	signal mae_8_to_cpu: std_logic_vector (7 downto 0);
      	signal be_access_error, be_access_error_registered : std_logic_vector(0 downto 0);
	
    	signal to_cpu, to_cpu_registered: std_logic_vector(89 downto 0);
    	signal to_be, to_be_registered :  std_logic_vector(FE_BE_COMMAND_SIZE-1 downto 0);

	signal access_byte_mask: std_logic_vector((2**LOG_BYTES_PER_DWORD)-1 downto 0); 

	constant LOG2_NUMBER_OF_BLOCKS: integer := LOG_ICACHE_SIZE_IN_BLOCKS;
        constant LOG2_BLOCK_SIZE_IN_BYTES: integer := 6;

    	signal access_mae : std_logic;
    	signal access_S : std_logic;
	signal tags_start_req, arrays_start_req, 
					tags_start_ack, 
					arrays_fin_req, 
					tags_fin_ack: std_logic;
	signal array_fin_ack, array_start_ack: std_logic;
	signal init_flag: std_logic;

	signal syn_inval_ready, coherence_inval_ready: boolean;
	signal syn_inval_accept, coherence_inval_accept: boolean;
	signal syn_inval_applicable, coherence_inval_applicable: boolean;

	signal tag_invalidate_apply: std_logic_vector(0 downto 0);
	signal tag_invalidate_line_address : std_logic_vector(25 downto 0);

	signal cpu_command_is_not_a_clear_or_flush: boolean;
	signal lookup_acc: std_logic_vector(2 downto 0);

-- see comment above..
--##decl_synopsys_sync_set_reset##
begin -- 
	-- once started, never finish!
	start_ack <= '1';
	fin_ack <= '0'; 
	tag_out <= tag_in;

	--------------------------------------------------------------------------------------------
	-- invalidate logic.
	--------------------------------------------------------------------------------------------
    	MMU_TO_ICACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_req(0) <= '1' when syn_inval_accept else '0';
	syn_inval_ready <= (MMU_TO_ICACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_ack(0) = '1');
	syn_inval_applicable <= syn_inval_ready and
					(MMU_TO_ICACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_data(26) = '1');
	syn_inval_accept <= (icache_state = SYN_INVALIDATE);


    	NOBLOCK_MMU_TO_ICACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_req(0) <= 
			'1' when coherence_inval_accept else '0';
    	coherence_inval_ready <= (NOBLOCK_MMU_TO_ICACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_ack(0) = '1');
    	coherence_inval_applicable <= 
			coherence_inval_ready and 
			     (NOBLOCK_MMU_TO_ICACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_data(26) = '1');
	coherence_inval_accept <=  cpu_command_is_not_a_clear_or_flush; 

	tag_invalidate_apply(0) <= 
		'1' when ((syn_inval_accept and syn_inval_applicable) or 
				(coherence_inval_accept and coherence_inval_applicable))
											else '0'; 
	tag_invalidate_line_address
		<= MMU_TO_ICACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_data(25 downto 0)
				when (syn_inval_accept and syn_inval_applicable) else
					NOBLOCK_MMU_TO_ICACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_data(25 downto 0);
	
	cpu_command_is_not_a_clear_or_flush <=
			latch_cpu_commands and (cpu_valid(0) = '1') and 
					(exec_cpu_flush(0) = '0') and (exec_cpu_new_stream_flush(0) = '0');
	--------------------------------------------------------------------------------------------

	-- for GenericCacheTags.
	access_is_read <= '1';
	access_is_ifetch <= '1';

	

	-- byte mask is always  0xff
 	access_byte_mask  <= (others => '1');
	-------------------------------------------------------------------------------------------
	-- registers, muxes.
	-------------------------------------------------------------------------------------------
	process(clk,reset)
	begin
		if(clk'event and clk = '1') then
	   	   if reset = '1' then
			cpu_reset_registered <= false;
			is_a_hit_registered <= (others => '0');
			dword_out_registered <= (others => '0');
			be_valid_registered(0)  <= '0';
			to_cpu_registered <= (others => '0');
			to_be_registered  <= (others => '0');
			latch_to_cpu_registered <= false;
			latch_to_be_registered <= false;
			init_or_reset_reg <= false;
      			exec_cpu_ifetch_reg <= (others => '0');
      			exec_cpu_asi_reg <= (others => '0');
			exec_cpu_S_reg <= (others => '0');
      			exec_cpu_addr_reg <= (others => '0');
			cpu_tag_lookup_reg <= false;
      			cpu_ifetch_valid_reg (0) <= '0';
			cpu_valid_reg(0) <= '0';
		   else
			
			latch_to_cpu_registered <= latch_to_cpu;
			latch_to_be_registered <= latch_to_be;

			if(latch_cpu_commands) then
				cpu_reset_registered <= cpu_reset;
				init_or_reset_reg <= init_or_reset;
      				exec_cpu_ifetch_reg <= exec_cpu_ifetch;
      				exec_cpu_asi_reg <= exec_cpu_asi;
				exec_cpu_S_reg <= exec_cpu_S;
      				exec_cpu_addr_reg <= exec_cpu_addr;
				cpu_tag_lookup_reg <= cpu_tag_lookup;
      				cpu_ifetch_valid_reg  <= cpu_ifetch_valid;
				cpu_valid_reg <= cpu_valid;
			elsif clear_cpu_commands then
				init_or_reset_reg <= false;
      				exec_cpu_ifetch_reg <= (others => '0');
      				exec_cpu_asi_reg <= (others => '0');
      				exec_cpu_addr_reg <= (others => '0');
				cpu_tag_lookup_reg <= false;
      				cpu_ifetch_valid_reg (0) <= '0';
				cpu_reset_registered <= false;
				cpu_valid_reg(0) <= '0';
			end if;
			if(latch_tag_results) then
				is_a_hit_registered <= is_a_hit;
				dword_out_registered <= dword_out;
			end if;
			if latch_cpu_commands then
				-- accept a new cpu command? Then clean up the
				-- be information.  
				be_valid_registered(0)  <= '0';
			end if;
			if(latch_to_cpu) then
				to_cpu_registered <= to_cpu;
			end if;
			if(latch_to_be) then
				to_be_registered <= to_be;
			end if;
                  end if;
		end if;
	end process;


	instr_pair_to_cpu  <= dword_out when  (icache_state = CHECK_HIT_OR_MISS) and (exec_cpu_ifetch_reg(0) = '1') 
				else be_dword when (first_be_response_can_be_applied and (exec_cpu_ifetch_reg(0) = '1')) 
					else ZERO_64;
	is_a_hit_to_cpu(0) <= is_a_hit(0) when (icache_state = CHECK_HIT_OR_MISS) else '0';
	mae_to_cpu(0)   <= be_mae(0) when first_be_response_can_be_applied else '0';
	access_error_to_cpu(0)  <= be_access_error(0) when first_be_response_can_be_applied else '0';
	
	-- insert into instruction buffer if relevant ....
	cacheable_to_cpu(0) <= 
		'1' when ((is_a_hit_to_cpu(0) = '1') or 
				(first_be_response_can_be_applied and (be_tag_cmd = CACHE_TAG_INSERT)))
				 								else '0';
	acc_to_cpu <= be_acc when first_be_response_can_be_applied else 
				lookup_acc when (is_a_hit_to_cpu(0) = '1') else (others => '0');


	mae_8_to_cpu <= (cacheable_to_cpu & acc_to_cpu & mZERO_1 & 
					is_a_hit_to_cpu & access_error_to_cpu & mae_to_cpu);
	mmu_fsr_to_cpu <= be_mmu_fsr  when first_be_response_can_be_applied else ZERO_18;

	to_cpu <= (mmu_fsr_to_cpu & mae_8_to_cpu & instr_pair_to_cpu);

	-------------------------------------------------------------------------------------------
	-- the command to the be will be generated after tag look up
	--   (note the use of registered values from the cpu).
	-------------------------------------------------------------------------------------------
	to_be  <= is_hit & cpu_permissions_ok & exec_cpu_asi_reg & exec_cpu_addr_reg;

	-------------------------------------------------------------------------------------------
	-- decoders.
	-------------------------------------------------------------------------------------------

  	classifyCmd : classifyCpuSideRequests 
    		port map ( -- 
      			from_cpu_ifetch => cpu_command,
      			cpu_valid => cpu_valid,
      			cpu_ifetch_valid => cpu_ifetch_valid,
      			exec_cpu_ifetch => exec_cpu_ifetch,
      			exec_cpu_new_stream_flush => exec_cpu_new_stream_flush,
      			exec_cpu_flush => exec_cpu_flush,
      			exec_cpu_S => exec_cpu_S,
      			exec_cpu_tag_command => exec_cpu_tag_command,
      			exec_cpu_array_command => exec_cpu_array_command,
      			exec_cpu_asi => exec_cpu_asi,
      			exec_cpu_addr => exec_cpu_addr);
	cpu_tag_lookup <= ((not init_or_reset) and (cpu_valid(0) = '1') and (exec_cpu_ifetch(0) = '1'));

    	beAnalyz: analyzeBeResponse  
    		port map ( -- 
      				from_backend => from_backend,
      				be_valid => be_valid,
				be_counter => be_counter,
				be_dword_id => be_dword_id,
				be_last_dword => be_last_dword,
      				be_mae  => be_mae,
      				be_access_error => be_access_error,
				be_acc => be_acc,
      				be_tag_cmd => be_tag_cmd,
      				be_array_cmd => be_array_cmd,
      				be_mmu_fsr => be_mmu_fsr,
     				be_dword => be_dword);

	-------------------------------------------------------------------------------------------
	-- construct predicates/inputs
	-------------------------------------------------------------------------------------------
	is_a_hit <= is_hit  and cpu_permissions_ok;

	cpu_reset <= ((NOBLOCK_CPU_to_ICACHE_reset_pipe_read_ack(0) = '1') and 
				  (NOBLOCK_CPU_to_ICACHE_reset_pipe_read_data(0) = '1'));
	cpu_command_available <= 
			((NOBLOCK_CPU_to_ICACHE_command_pipe_read_ack(0) = '1') and 
				  (NOBLOCK_CPU_to_ICACHE_command_pipe_read_data(40) = '1'));
	be_response_available <= 
			((noblock_icache_backend_to_frontend_pipe_read_ack(0) = '1') and 
				  (noblock_icache_backend_to_frontend_pipe_read_data(BE_FE_RESPONSE_SIZE-1) = '1'));
	be_ready_for_command  <= (icache_frontend_to_backend_pipe_write_ack(0) = '1');

	cpu_ready_for_response  <= 
			((cpu_ifetch_valid_reg(0) = '1') and (ICACHE_to_CPU_response_pipe_write_ack(0) = '1'))
				or
			(cpu_reset_registered and (ICACHE_to_CPU_reset_ack_pipe_write_ack(0) = '1'));


	-- be is needed is computed one cycle  after command is seen.
	be_is_needed <= (cpu_tag_lookup_reg and (is_a_hit(0) = '0'));
	expect_be_response <= true;

	init_or_reset <=  cpu_reset;
	---------------------------------------------------------------------------------------------
	-- control state machine
	---------------------------------------------------------------------------------------------
	process(clk, reset, icache_state, 
			cpu_command_available,
			cpu_reset,
			be_ready_for_command,
			be_is_needed,
			be_has_completed,
			expect_be_response,
			be_last_dword,
			be_response_available,
			cpu_ready_for_response)
		variable next_icache_state : IcacheState;
		variable accept_cpu_commands_var  : boolean;
		variable latch_cpu_commands_var  : boolean;
		variable clear_cpu_commands_var  : boolean;
		variable latch_tag_results_var  : boolean;
		variable latch_to_be_var	: boolean;
		variable latch_to_cpu_var	: boolean;
		variable accept_be_response_var  : boolean;
		variable write_to_be_var	 : boolean;
		variable write_to_cpu_var	 : boolean;
		variable next_be_has_completed_var	 : boolean;

		variable accept_cpu_reset_var: boolean;
		variable send_cpu_reset_ack_var: boolean;

	begin
		next_icache_state := icache_state;
		accept_cpu_commands_var  := false;
		latch_cpu_commands_var  := false;
		accept_be_response_var  := false;
		latch_to_be_var := false;
		latch_to_cpu_var := false;
		write_to_be_var	 := false;
		write_to_cpu_var	 := false;
		next_be_has_completed_var := false;
		clear_cpu_commands_var := false;

		send_cpu_reset_ack_var := false;
		accept_cpu_reset_var   := false;
	

		case icache_state is 
			when IDLE => 
			    if (not waiting_on_tags_arrays) then 
			      accept_cpu_reset_var := true;
			      -- important: it is assumed that there is always room
			      -- for the reset ack to the cpu..
			      if (cpu_reset) then
				  send_cpu_reset_ack_var := true;
			      else
				  accept_cpu_commands_var := true;
				  if(cpu_command_available) then
					  latch_cpu_commands_var := true;
					  next_icache_state := CHECK_HIT_OR_MISS;
				  end if;
			      end if;
			    end if;
			when CHECK_HIT_OR_MISS =>
				if(waiting_on_tags_arrays) then
					next_icache_state := CHECK_HIT_OR_MISS;
				elsif (be_is_needed) then
					write_to_be_var := true;
					if be_ready_for_command then
						if expect_be_response then
							next_icache_state := SYN_INVALIDATE;	
						else
							-- can send response to CPU!
							write_to_cpu_var := true;
							if(cpu_ready_for_response) then
							-- CPU has accepted.. see if it has a command..

			    					accept_cpu_reset_var := true;
			    					-- important: it is assumed that there is always room
			    					-- for the reset ack to the cpu..
			    					if (cpu_reset) then
									send_cpu_reset_ack_var := true;
									next_icache_state := IDLE;
			    					else
									accept_cpu_commands_var := true;
									if(cpu_command_available) then
										latch_cpu_commands_var := true;
									else
										clear_cpu_commands_var := true;
										next_icache_state := IDLE;
									end if;
								end if;
							else
								-- latch to_cpu!
								latch_to_cpu_var := true;
								next_icache_state := SEND_WAIT_ON_CPU;
							end if;
							-- no be response expected..
							-- be has completed.
							next_be_has_completed_var := true;
						end if;
					else
						-- be not ready to be receiver, latch to_be!
						latch_to_be_var := true;
						-- cpu will be responded to later..
						-- need to register the return values to cpu
						-- as well!
						latch_to_cpu_var := true;
						next_icache_state := SEND_WAIT_ON_BE;	
					end if;
				elsif cpu_ready_for_response then 
					write_to_cpu_var := true;
			    		accept_cpu_reset_var := true;
			    		-- important: it is assumed that there is always room
			    		-- for the reset ack to the cpu..
			    		if (cpu_reset) then
						send_cpu_reset_ack_var := true;
						next_icache_state := IDLE;
					else
						accept_cpu_commands_var := true;
						if cpu_command_available then
							latch_cpu_commands_var := true;
						else
							clear_cpu_commands_var := true;
							next_icache_state := IDLE;
						end if;
					end if;
				else
					-- not sending cpu response in CHECK-HIT?
					-- latch to_cpu!
					latch_to_cpu_var := true;
					next_icache_state := SEND_WAIT_ON_CPU;	
					-- no be needed, ergo it has completed..
					next_be_has_completed_var := true;
				end if;
			when SEND_WAIT_ON_BE =>
				-- to_be_registered will be used to send to be.
				write_to_be_var := true;
				if be_ready_for_command then
					if(expect_be_response) then
						next_icache_state := SYN_INVALIDATE;	
					else
						-- can send response to CPU!
						write_to_cpu_var := true;
						if(cpu_ready_for_response) then
						-- CPU has accepted.. see if it has a command..

			    				accept_cpu_reset_var := true;
			    				-- important: it is assumed that there is always room
			    				-- for the reset ack to the cpu..
			    				if (cpu_reset) then
								send_cpu_reset_ack_var := true;
								next_icache_state := IDLE;
							else
								accept_cpu_commands_var := true;
								if(cpu_command_available) then
									latch_cpu_commands_var := true;
								else
									clear_cpu_commands_var := true;
									next_icache_state := IDLE;
								end if;
							end if;
						else
							-- no response expected from be..
						        -- to_cpu_reg has already been updated.	
							next_icache_state := SEND_WAIT_ON_CPU;	
						end if;
						next_be_has_completed_var := true;
					end if;
				end if;
			when SYN_INVALIDATE =>
				if(syn_inval_ready) then
					next_icache_state := RECV_WAIT_ON_BE_FIRST_DWORD;
				end if;
			when RECV_WAIT_ON_BE_FIRST_DWORD =>
			   if (not waiting_on_tags_arrays) then
				-- Wait for the first dword from the BE.
				-- (Note that this could be the last also!)
				accept_be_response_var := true;
				if (be_response_available) then
					-- we will be doing tag access.
					-- and also writing dword to memory.
					latch_to_cpu_var := true;
					next_icache_state := SEND_WAIT_ON_CPU;

					if (be_last_dword(0) = '1') then
						next_be_has_completed_var := true;
					end if;
				end if;
                            end if;
			when SEND_WAIT_ON_CPU =>
				if(waiting_on_tags_arrays) then
					-- if be has completed, it stays completed.
					next_be_has_completed_var := be_has_completed;
				else
				   write_to_cpu_var := true;
				   if cpu_ready_for_response then
					if(be_has_completed) then 
			    			accept_cpu_reset_var := true;
			    			-- important: it is assumed that there is always room
			    			-- for the reset ack to the cpu..
			    			if (cpu_reset) then
							send_cpu_reset_ack_var := true;
							next_icache_state := IDLE;
						else
							accept_cpu_commands_var := true;
							if cpu_command_available then
								latch_cpu_commands_var := true;
								next_icache_state := CHECK_HIT_OR_MISS;
							else
								clear_cpu_commands_var := true;
								next_icache_state := IDLE;
							end if;
						end if;
					else
						next_icache_state := RECV_WAIT_ON_BE_REMAINING_DWORDS;
					end if;
				   else
					-- if be has completed, it stays completed.
					next_be_has_completed_var := be_has_completed;
				   end if;
				end if;
			when RECV_WAIT_ON_BE_REMAINING_DWORDS =>
			        if (waiting_on_tags_arrays) then
				 	next_be_has_completed_var := be_has_completed; 
				else
				  -- wait for the remaining dwords from the backend.
				  accept_be_response_var := true;
				  if (be_response_available) then
				     if (be_last_dword(0) = '1') then
					  next_be_has_completed_var := true; 
					  clear_cpu_commands_var := true;
					  next_icache_state := IDLE;
				      end if;
                                  end if;
				end if;
		end case;

		accept_cpu_commands <= accept_cpu_commands_var;
		latch_cpu_commands <= latch_cpu_commands_var;
		clear_cpu_commands <= clear_cpu_commands_var;
		latch_to_be  <= latch_to_be_var;
		latch_to_cpu  <= latch_to_cpu_var;
		accept_be_response <= accept_be_response_var;
		write_to_be	   <= write_to_be_var;
		write_to_cpu	   <= write_to_cpu_var;

		accept_cpu_reset <= accept_cpu_reset_var;
		send_cpu_reset_ack <= send_cpu_reset_ack_var;
		

		if clk'event and clk = '1' then
			if reset = '1' then	
				icache_state <= IDLE;
				be_has_completed <= false;
			else
				icache_state <= next_icache_state;
				be_has_completed <= next_be_has_completed_var;
			end if;
		end if;	
	end process;


	------------------------------------------------------------------------------------------------------
	-- BE response will be digested using the registered cpu address.
	------------------------------------------------------------------------------------------------------
        be_addr <= exec_cpu_addr_reg (31 downto 6) & be_dword_id & "000";
        be_S    <= exec_cpu_S_reg;
	be_response_can_be_applied <= 
		(not waiting_on_tags_arrays) and (be_valid(0) = '1') and 
			((icache_state = RECV_WAIT_ON_BE_FIRST_DWORD)
					or
			  (icache_state = RECV_WAIT_ON_BE_REMAINING_DWORDS));

	first_be_response_can_be_applied <= 
			(not waiting_on_tags_arrays) and
				((icache_state = RECV_WAIT_ON_BE_FIRST_DWORD) and (be_valid(0) = '1')); 

	------------------------------------------------------------------------------------------------------
	-- accessIcache
	------------------------------------------------------------------------------------------------------
	arrays_start_req  <= '1' when (send_cpu_reset_ack or latch_cpu_commands  or  
							be_response_can_be_applied) else '0';
	tags_start_req <= arrays_start_req or tag_invalidate_apply(0);
	tags_arrays_trigger <= tags_start_req or arrays_start_req;

	init_flag  <= '1' when send_cpu_reset_ack else '0';
	access_mae <= be_mae(0) when be_response_can_be_applied else '0';
	access_S <= be_S(0) when be_response_can_be_applied else exec_cpu_S(0);
	access_tags_acc <= be_acc when be_response_can_be_applied else (others => '0');

	TagsArraysBlock: block
    		signal access_tag_command : std_logic_vector(2 downto 0);
    		signal access_tag_lookup, access_tag_insert, 
				access_tag_clear_line,
				access_tag_clear_all : std_logic;
    		signal access_array_command : std_logic_vector(2 downto 0);
    		signal access_addr : std_logic_vector(31 downto 0);
    		signal access_dword : std_logic_vector((2**log2_block_size_in_bytes)-1 downto 0);

	begin
	   access_tag_command <=  CACHE_TAG_CLEAR_LINE
					when (((be_mae(0) = '1') or (be_access_error(0) = '1')) and be_response_can_be_applied)
					else be_tag_cmd when first_be_response_can_be_applied
					else exec_cpu_tag_command when (latch_cpu_commands and (cpu_valid(0) = '1'))
					else CACHE_TAG_CLEAR_ALL when send_cpu_reset_ack
					else CACHE_TAG_NOP;
	   access_tag_lookup <= '1' when ((exec_cpu_tag_command = CACHE_TAG_LOOKUP) and
						latch_cpu_commands and (cpu_valid(0) = '1')) else '0';
	   access_tag_insert <= '1' when ((be_tag_cmd = CACHE_TAG_INSERT) and first_be_response_can_be_applied)
						else '0';
	   access_tag_clear_line <= '1' when (access_tag_command = CACHE_TAG_CLEAR_LINE) else '0';
	   access_tag_clear_all <= '1' when (access_tag_command = CACHE_TAG_CLEAR_ALL) else '0';
 
	   access_addr <= be_addr when be_response_can_be_applied else exec_cpu_addr;

	   access_array_command <=  CACHE_ARRAY_NOP when (((be_mae(0) = '1') or (be_access_error(0) = '1')) and be_response_can_be_applied)
					else be_array_cmd when be_response_can_be_applied
					else exec_cpu_array_command when latch_cpu_commands and (cpu_valid(0) = '1')
					else CACHE_ARRAY_NOP;
	   access_dword      <= be_dword when be_response_can_be_applied else (others => '0');

           directMappedGen: if (LOG_ICACHE_SET_ASSOCIATIVITY = 0) generate 
	      tagsArraysInst: 
		GenericIcacheTagsArraysWithInvalidate
                        generic map (name => "icache-tags-arrays",
                                        log2_number_of_blocks => LOG2_NUMBER_OF_BLOCKS, -- 9  
                                        log2_block_size_in_bytes => LOG2_BLOCK_SIZE_IN_BYTES, -- 6
                                        address_width => 32,
                                        log2_data_width_in_bytes => 3)
			port map (
					trigger => tags_arrays_trigger,	
					done => tags_arrays_done,	
					init_flag => init_flag,
					access_mae => access_mae,
					access_S => access_S,
					access_is_read => access_is_read,
					access_is_ifetch => access_is_ifetch,
					access_acc => access_tags_acc,
					access_tag_command => access_tag_command,
					invalidate => tag_invalidate_apply,
					invalidate_line_address => tag_invalidate_line_address,
					is_hit => is_hit,
					permissions_ok => cpu_permissions_ok,
					lookup_acc => lookup_acc,
    					access_array_command  => access_array_command ,
    					access_addr  => access_addr ,
    					access_dword  => access_dword ,
    					dword_out  => dword_out ,
    					clk => clk,
					reset => reset
				);
			waiting_on_tags_arrays <= false;
		end generate directMappedGen;


    		setAssociativeGen: if (LOG_ICACHE_SET_ASSOCIATIVITY > 0) generate 
	   	   tagsArraysInst: 
			GenericSetAssociativeCacheTagsArraysWithInvalidate
                             generic map (name => "dcache-tags-arrays",
                                        log2_number_of_blocks => LOG2_NUMBER_OF_BLOCKS, 	-- 9  
                                        log2_block_size_in_bytes => LOG2_BLOCK_SIZE_IN_BYTES, 	-- 6
					log2_associativity => LOG_ICACHE_SET_ASSOCIATIVITY, 	-- as specified.
                                        address_width => 32,
                                        log2_data_width_in_bytes => 3,
					icache_flag => true)
		 	     port map (
					trigger => tags_arrays_trigger,	
					done => tags_arrays_done,	
					init_flag => init_flag,
					access_mae => access_mae,
					access_S => access_S,
					access_is_read => access_is_read,
					access_is_ifetch => access_is_ifetch,
					access_acc => access_tags_acc,
					access_tag_lookup => access_tag_lookup,
					access_tag_insert => access_tag_insert,
					access_tag_clear_line => access_tag_clear_line,
					access_tag_clear_all => access_tag_clear_all,
    					access_array_command  => access_array_command ,
					access_addr => access_addr,
    					access_byte_mask  => access_byte_mask ,
    					access_dword  => access_dword ,
					-- invalidation...
					invalidate => tag_invalidate_apply,
					invalidate_line_address => tag_invalidate_line_address,
					-- outputs.
					is_hit => is_hit,
					permissions_ok => cpu_permissions_ok,
					lookup_acc => lookup_acc,
    					dword_out  => dword_out ,
    					clk => clk,
					-- clock, reset.
					reset => reset
				);
	
			process(clk, reset, tags_arrays_trigger, tags_arrays_done)
			begin
				if(clk'event and (clk = '1')) then
					if(reset = '1') then
						wait_on_tags_arrays <= false;
					else
						if(tags_arrays_trigger = '1')  then
							wait_on_tags_arrays <= true;
						elsif (wait_on_tags_arrays and (tags_arrays_done = '1')) then
							wait_on_tags_arrays <= false;
						end if;
					end if;
				end if;
		
			end process;
			waiting_on_tags_arrays <= wait_on_tags_arrays and (tags_arrays_done = '0');
		end generate setAssociativeGen;
	end block TagsArraysBlock;

	-------------------------------------------------------------------------------------------
	-- pipe access logic.
	-------------------------------------------------------------------------------------------
	NOBLOCK_CPU_to_ICACHE_command_pipe_read_req (0) <= '1' when accept_cpu_commands else '0';
	cpu_command <= NOBLOCK_CPU_to_ICACHE_command_pipe_read_data when NOBLOCK_CPU_to_ICACHE_command_pipe_read_ack(0) = '1' 
					else (others => '0');

	NOBLOCK_CPU_to_ICACHE_reset_pipe_read_req (0) <= '1' when accept_cpu_reset else '0';

	noblock_icache_backend_to_frontend_pipe_read_req (0) <= '1' when accept_be_response else '0';
	from_backend <= noblock_icache_backend_to_frontend_pipe_read_data when
				noblock_icache_backend_to_frontend_pipe_read_ack(0) = '1' else
					(others => '0');

	icache_frontend_to_backend_pipe_write_req (0) <= '1' when write_to_be else '0';
	icache_frontend_to_backend_pipe_write_data  <= to_be_registered when (icache_state = SEND_WAIT_ON_BE) else to_be;

	ICACHE_to_CPU_response_pipe_write_req(0) <= '1' when (cpu_valid_reg(0) = '1') and write_to_cpu else '0';
	ICACHE_to_CPU_response_pipe_write_data <= to_cpu when (icache_state = CHECK_HIT_OR_MISS) else to_cpu_registered;

	ICACHE_to_CPU_reset_ack_pipe_write_req(0) <= '1' when send_cpu_reset_ack else '0';
	ICACHE_to_CPU_reset_ack_pipe_write_data(0) <= '1';
end IcacheFrontendCoreArch;

library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.basecomponents.all;

library AjitCustom;

use AjitCustom.AjitGlobalConfigurationPackage.all;
use AjitCustom.AjitCoreConfigurationPackage.all;
use AjitCustom.AjitCustomComponents.all;
use AjitCustom.CachePackage.all;

entity IcacheFrontendDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    NOBLOCK_CPU_to_ICACHE_command_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_ICACHE_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_ICACHE_command_pipe_read_data : in   std_logic_vector(40 downto 0);
    NOBLOCK_CPU_to_ICACHE_reset_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_ICACHE_reset_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_ICACHE_reset_pipe_read_data : in   std_logic_vector(0 downto 0);
    noblock_icache_backend_to_frontend_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_icache_backend_to_frontend_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_icache_backend_to_frontend_pipe_read_data : in   std_logic_vector(101 downto 0);
    ICACHE_to_CPU_reset_ack_pipe_write_req : out  std_logic_vector(0 downto 0);
    ICACHE_to_CPU_reset_ack_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ICACHE_to_CPU_reset_ack_pipe_write_data : out  std_logic_vector(0 downto 0);
    ICACHE_to_CPU_response_pipe_write_req : out  std_logic_vector(0 downto 0);
    ICACHE_to_CPU_response_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ICACHE_to_CPU_response_pipe_write_data : out  std_logic_vector(89 downto 0);
    icache_frontend_to_backend_pipe_write_req : out  std_logic_vector(0 downto 0);
    icache_frontend_to_backend_pipe_write_ack : in   std_logic_vector(0 downto 0);
    icache_frontend_to_backend_pipe_write_data : out  std_logic_vector(41 downto 0);
    MMU_TO_ICACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_req: out std_logic_vector(0 downto 0);
    MMU_TO_ICACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_ack: in std_logic_vector(0 downto 0);
    MMU_TO_ICACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_data: in std_logic_vector(26 downto 0);
    NOBLOCK_MMU_TO_ICACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_req: out std_logic_vector(0 downto 0);
    NOBLOCK_MMU_TO_ICACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_ack: in std_logic_vector(0 downto 0);
    NOBLOCK_MMU_TO_ICACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_data: in std_logic_vector(26 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity IcacheFrontendDaemon;

architecture IcacheFrontendArch  of IcacheFrontEndDaemon is -- system-architecture 

    signal NOBLOCK_BUFFERED_CPU_to_ICACHE_command_pipe_read_req : std_logic_vector(0 downto 0);
    signal NOBLOCK_BUFFERED_CPU_to_ICACHE_command_pipe_read_ack : std_logic_vector(0 downto 0);
    signal NOBLOCK_BUFFERED_CPU_to_ICACHE_command_pipe_read_data : std_logic_vector(40 downto 0);

begin -- 
	ifBuffer: if (ICACHE_BUFFER_REQUEST > 0) generate
		qBuf: QueueBase
			generic map (name => "IcacheRequestQueue", queue_depth => 2,
						data_width => 41, save_one_slot => false)
			port map (
				clk => clk,
				reset => reset,
				data_in => NOBLOCK_CPU_to_ICACHE_command_pipe_read_data,
				push_req => NOBLOCK_CPU_to_ICACHE_command_pipe_read_ack(0),
				push_ack => NOBLOCK_CPU_to_ICACHE_command_pipe_read_req(0),
				data_out => NOBLOCK_BUFFERED_CPU_to_ICACHE_command_pipe_read_data,
				pop_req =>  NOBLOCK_BUFFERED_CPU_to_ICACHE_command_pipe_read_req(0),
				pop_ack =>  NOBLOCK_BUFFERED_CPU_to_ICACHE_command_pipe_read_ack(0)
			);
	end generate ifBuffer;

	ifNoBuffer: if (ICACHE_BUFFER_REQUEST = 0) generate

		NOBLOCK_CPU_to_ICACHE_command_pipe_read_req <= NOBLOCK_BUFFERED_CPU_to_ICACHE_command_pipe_read_req;
    		NOBLOCK_BUFFERED_CPU_to_ICACHE_command_pipe_read_ack <= NOBLOCK_CPU_to_ICACHE_command_pipe_read_ack;
    		NOBLOCK_BUFFERED_CPU_to_ICACHE_command_pipe_read_data <= NOBLOCK_CPU_to_ICACHE_command_pipe_read_data;
	end generate ifNoBuffer;


	coreInst: IcacheFrontendCoreDaemon 
  		generic map (tag_length => tag_length)
  		port map ( -- 
    			NOBLOCK_BUFFERED_CPU_to_ICACHE_command_pipe_read_req ,
    			NOBLOCK_BUFFERED_CPU_to_ICACHE_command_pipe_read_ack ,
    			NOBLOCK_BUFFERED_CPU_to_ICACHE_command_pipe_read_data ,
    			NOBLOCK_CPU_to_ICACHE_reset_pipe_read_req ,
    			NOBLOCK_CPU_to_ICACHE_reset_pipe_read_ack ,
    			NOBLOCK_CPU_to_ICACHE_reset_pipe_read_data ,
    			noblock_icache_backend_to_frontend_pipe_read_req ,
    			noblock_icache_backend_to_frontend_pipe_read_ack ,
    			noblock_icache_backend_to_frontend_pipe_read_data ,
    			ICACHE_to_CPU_reset_ack_pipe_write_req ,
    			ICACHE_to_CPU_reset_ack_pipe_write_ack ,
    			ICACHE_to_CPU_reset_ack_pipe_write_data ,
    			ICACHE_to_CPU_response_pipe_write_req ,
    			ICACHE_to_CPU_response_pipe_write_ack ,
    			ICACHE_to_CPU_response_pipe_write_data ,
    			icache_frontend_to_backend_pipe_write_req ,
    			icache_frontend_to_backend_pipe_write_ack ,
    			icache_frontend_to_backend_pipe_write_data ,
    			MMU_TO_ICACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_req,
    			MMU_TO_ICACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_ack,
    			MMU_TO_ICACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_data,
    			NOBLOCK_MMU_TO_ICACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_req,
    			NOBLOCK_MMU_TO_ICACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_ack,
    			NOBLOCK_MMU_TO_ICACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_data,
    			tag_in,
    			tag_out,
    			clk ,
    			reset ,
    			start_req ,
    			start_ack ,
    			fin_req ,
    			fin_ack   
  			);

end IcacheFrontendArch;

library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
entity createCacheLineFromDword_VVD is -- 
  port ( -- 
    be_write_data : in  std_logic_vector(63 downto 0);
    be_offset_in_line : in  std_logic_vector(3 downto 0);
    be_cache_line : out  std_logic_vector(511 downto 0)-- 
  );
  -- 
end entity createCacheLineFromDword_VVD;
architecture createCacheLineFromDword_VVD_arch of createCacheLineFromDword_VVD is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(68-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal be_write_data_buffer :  std_logic_vector(63 downto 0);
  signal be_offset_in_line_buffer :  std_logic_vector(3 downto 0);
  -- output port buffer signals
  signal be_cache_line_buffer :  std_logic_vector(511 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  be_write_data_buffer <= be_write_data;
  be_offset_in_line_buffer <= be_offset_in_line;
  -- output handling  -------------------------------------------------------
  be_cache_line <= be_cache_line_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u128_u256_860_wire : std_logic_vector(255 downto 0);
    signal CONCAT_u128_u256_867_wire : std_logic_vector(255 downto 0);
    signal CONCAT_u64_u128_856_wire : std_logic_vector(127 downto 0);
    signal CONCAT_u64_u128_859_wire : std_logic_vector(127 downto 0);
    signal CONCAT_u64_u128_863_wire : std_logic_vector(127 downto 0);
    signal CONCAT_u64_u128_866_wire : std_logic_vector(127 downto 0);
    signal EQ_u3_u1_792_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_800_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_808_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_816_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_824_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_832_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_840_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_848_wire : std_logic_vector(0 downto 0);
    signal konst_791_wire_constant : std_logic_vector(2 downto 0);
    signal konst_794_wire_constant : std_logic_vector(63 downto 0);
    signal konst_799_wire_constant : std_logic_vector(2 downto 0);
    signal konst_802_wire_constant : std_logic_vector(63 downto 0);
    signal konst_807_wire_constant : std_logic_vector(2 downto 0);
    signal konst_810_wire_constant : std_logic_vector(63 downto 0);
    signal konst_815_wire_constant : std_logic_vector(2 downto 0);
    signal konst_818_wire_constant : std_logic_vector(63 downto 0);
    signal konst_823_wire_constant : std_logic_vector(2 downto 0);
    signal konst_826_wire_constant : std_logic_vector(63 downto 0);
    signal konst_831_wire_constant : std_logic_vector(2 downto 0);
    signal konst_834_wire_constant : std_logic_vector(63 downto 0);
    signal konst_839_wire_constant : std_logic_vector(2 downto 0);
    signal konst_842_wire_constant : std_logic_vector(63 downto 0);
    signal konst_847_wire_constant : std_logic_vector(2 downto 0);
    signal konst_850_wire_constant : std_logic_vector(63 downto 0);
    signal o7_788 : std_logic_vector(2 downto 0);
    signal w0_796 : std_logic_vector(63 downto 0);
    signal w1_804 : std_logic_vector(63 downto 0);
    signal w2_812 : std_logic_vector(63 downto 0);
    signal w3_820 : std_logic_vector(63 downto 0);
    signal w4_828 : std_logic_vector(63 downto 0);
    signal w5_836 : std_logic_vector(63 downto 0);
    signal w6_844 : std_logic_vector(63 downto 0);
    signal w7_852 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    konst_791_wire_constant <= "000";
    konst_794_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_799_wire_constant <= "001";
    konst_802_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_807_wire_constant <= "010";
    konst_810_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_815_wire_constant <= "011";
    konst_818_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_823_wire_constant <= "100";
    konst_826_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_831_wire_constant <= "101";
    konst_834_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_839_wire_constant <= "110";
    konst_842_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_847_wire_constant <= "111";
    konst_850_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    -- flow-through select operator MUX_795_inst
    w0_796 <= be_write_data_buffer when (EQ_u3_u1_792_wire(0) /=  '0') else konst_794_wire_constant;
    -- flow-through select operator MUX_803_inst
    w1_804 <= be_write_data_buffer when (EQ_u3_u1_800_wire(0) /=  '0') else konst_802_wire_constant;
    -- flow-through select operator MUX_811_inst
    w2_812 <= be_write_data_buffer when (EQ_u3_u1_808_wire(0) /=  '0') else konst_810_wire_constant;
    -- flow-through select operator MUX_819_inst
    w3_820 <= be_write_data_buffer when (EQ_u3_u1_816_wire(0) /=  '0') else konst_818_wire_constant;
    -- flow-through select operator MUX_827_inst
    w4_828 <= be_write_data_buffer when (EQ_u3_u1_824_wire(0) /=  '0') else konst_826_wire_constant;
    -- flow-through select operator MUX_835_inst
    w5_836 <= be_write_data_buffer when (EQ_u3_u1_832_wire(0) /=  '0') else konst_834_wire_constant;
    -- flow-through select operator MUX_843_inst
    w6_844 <= be_write_data_buffer when (EQ_u3_u1_840_wire(0) /=  '0') else konst_842_wire_constant;
    -- flow-through select operator MUX_851_inst
    w7_852 <= be_write_data_buffer when (EQ_u3_u1_848_wire(0) /=  '0') else konst_850_wire_constant;
    -- flow-through slice operator slice_787_inst
    o7_788 <= be_offset_in_line_buffer(2 downto 0);
    -- binary operator CONCAT_u128_u256_860_inst
    process(CONCAT_u64_u128_856_wire, CONCAT_u64_u128_859_wire) -- 
      variable tmp_var : std_logic_vector(255 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u64_u128_856_wire, CONCAT_u64_u128_859_wire, tmp_var);
      CONCAT_u128_u256_860_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u128_u256_867_inst
    process(CONCAT_u64_u128_863_wire, CONCAT_u64_u128_866_wire) -- 
      variable tmp_var : std_logic_vector(255 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u64_u128_863_wire, CONCAT_u64_u128_866_wire, tmp_var);
      CONCAT_u128_u256_867_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u256_u512_868_inst
    process(CONCAT_u128_u256_860_wire, CONCAT_u128_u256_867_wire) -- 
      variable tmp_var : std_logic_vector(511 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u128_u256_860_wire, CONCAT_u128_u256_867_wire, tmp_var);
      be_cache_line_buffer <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u64_u128_856_inst
    process(w0_796, w1_804) -- 
      variable tmp_var : std_logic_vector(127 downto 0); -- 
    begin -- 
      ApConcat_proc(w0_796, w1_804, tmp_var);
      CONCAT_u64_u128_856_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u64_u128_859_inst
    process(w2_812, w3_820) -- 
      variable tmp_var : std_logic_vector(127 downto 0); -- 
    begin -- 
      ApConcat_proc(w2_812, w3_820, tmp_var);
      CONCAT_u64_u128_859_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u64_u128_863_inst
    process(w4_828, w5_836) -- 
      variable tmp_var : std_logic_vector(127 downto 0); -- 
    begin -- 
      ApConcat_proc(w4_828, w5_836, tmp_var);
      CONCAT_u64_u128_863_wire <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u64_u128_866_inst
    process(w6_844, w7_852) -- 
      variable tmp_var : std_logic_vector(127 downto 0); -- 
    begin -- 
      ApConcat_proc(w6_844, w7_852, tmp_var);
      CONCAT_u64_u128_866_wire <= tmp_var; -- 
    end process;
    -- binary operator EQ_u3_u1_792_inst
    process(o7_788) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(o7_788, konst_791_wire_constant, tmp_var);
      EQ_u3_u1_792_wire <= tmp_var; -- 
    end process;
    -- binary operator EQ_u3_u1_800_inst
    process(o7_788) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(o7_788, konst_799_wire_constant, tmp_var);
      EQ_u3_u1_800_wire <= tmp_var; -- 
    end process;
    -- binary operator EQ_u3_u1_808_inst
    process(o7_788) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(o7_788, konst_807_wire_constant, tmp_var);
      EQ_u3_u1_808_wire <= tmp_var; -- 
    end process;
    -- binary operator EQ_u3_u1_816_inst
    process(o7_788) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(o7_788, konst_815_wire_constant, tmp_var);
      EQ_u3_u1_816_wire <= tmp_var; -- 
    end process;
    -- binary operator EQ_u3_u1_824_inst
    process(o7_788) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(o7_788, konst_823_wire_constant, tmp_var);
      EQ_u3_u1_824_wire <= tmp_var; -- 
    end process;
    -- binary operator EQ_u3_u1_832_inst
    process(o7_788) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(o7_788, konst_831_wire_constant, tmp_var);
      EQ_u3_u1_832_wire <= tmp_var; -- 
    end process;
    -- binary operator EQ_u3_u1_840_inst
    process(o7_788) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(o7_788, konst_839_wire_constant, tmp_var);
      EQ_u3_u1_840_wire <= tmp_var; -- 
    end process;
    -- binary operator EQ_u3_u1_848_inst
    process(o7_788) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(o7_788, konst_847_wire_constant, tmp_var);
      EQ_u3_u1_848_wire <= tmp_var; -- 
    end process;
    -- 
  end Block; -- data_path
  -- 
end createCacheLineFromDword_VVD_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
entity create_cpu_cache_line_VVD is -- 
  port ( -- 
    cpu_addr : in  std_logic_vector(31 downto 0);
    cpu_write_data : in  std_logic_vector(63 downto 0);
    cpu_cache_line : out  std_logic_vector(511 downto 0)-- 
  );
  -- 
end entity create_cpu_cache_line_VVD;
architecture create_cpu_cache_line_VVD_arch of create_cpu_cache_line_VVD is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(96-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal cpu_addr_buffer :  std_logic_vector(31 downto 0);
  signal cpu_write_data_buffer :  std_logic_vector(63 downto 0);
  -- output port buffer signals
  signal cpu_cache_line_buffer :  std_logic_vector(511 downto 0);
  -- volatile/operator module components. 
  component createCacheLineFromDword_VVD is -- 
    port ( -- 
      be_write_data : in  std_logic_vector(63 downto 0);
      be_offset_in_line : in  std_logic_vector(3 downto 0);
      be_cache_line : out  std_logic_vector(511 downto 0)-- 
    );
    -- 
  end component; 
  component offsetInLine_VVD is -- 
    port ( -- 
      addr : in  std_logic_vector(31 downto 0);
      ret_val : out  std_logic_vector(3 downto 0)-- 
    );
    -- 
  end component; 
  -- 
begin --  
  -- input handling ------------------------------------------------
  cpu_addr_buffer <= cpu_addr;
  cpu_write_data_buffer <= cpu_write_data;
  -- output handling  -------------------------------------------------------
  cpu_cache_line <= cpu_cache_line_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal cpu_offset_in_line_1496 : std_logic_vector(3 downto 0);
    -- 
  begin -- 
    volatile_operator_offsetInLine_1873: offsetInLine_VVD port map(addr => cpu_addr_buffer, ret_val => cpu_offset_in_line_1496); 
    volatile_operator_createCacheLineFromDword_1874: createCacheLineFromDword_VVD port map(be_write_data => cpu_write_data_buffer, be_offset_in_line => cpu_offset_in_line_1496, be_cache_line => cpu_cache_line_buffer); 
    -- 
  end Block; -- data_path
  -- 
end create_cpu_cache_line_VVD_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
entity dcacheNeedsToBeFlushed_VVD is -- 
  port ( -- 
    asi : in  std_logic_vector(7 downto 0);
    req_type : in  std_logic_vector(3 downto 0);
    is_flush_asi : out  std_logic_vector(0 downto 0);
    is_mmu_ctrl_reg_write : out  std_logic_vector(0 downto 0);
    flush_line_only : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity dcacheNeedsToBeFlushed_VVD;
architecture dcacheNeedsToBeFlushed_VVD_arch of dcacheNeedsToBeFlushed_VVD is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(12-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal asi_buffer :  std_logic_vector(7 downto 0);
  signal req_type_buffer :  std_logic_vector(3 downto 0);
  -- output port buffer signals
  signal is_flush_asi_buffer :  std_logic_vector(0 downto 0);
  signal is_mmu_ctrl_reg_write_buffer :  std_logic_vector(0 downto 0);
  signal flush_line_only_buffer :  std_logic_vector(0 downto 0);
  -- volatile/operator module components. 
  component isDcacheFlushAsi_VVD is -- 
    port ( -- 
      asi : in  std_logic_vector(7 downto 0);
      ret_val : out  std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component; 
  -- 
begin --  
  -- input handling ------------------------------------------------
  asi_buffer <= asi;
  req_type_buffer <= req_type;
  -- output handling  -------------------------------------------------------
  is_flush_asi <= is_flush_asi_buffer;
  is_mmu_ctrl_reg_write <= is_mmu_ctrl_reg_write_buffer;
  flush_line_only <= flush_line_only_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal EQ_u4_u1_1236_wire : std_logic_vector(0 downto 0);
    signal EQ_u4_u1_1239_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_1249_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_1255_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_1258_wire : std_logic_vector(0 downto 0);
    signal R_ASI_FLUSH_I_D_USER_1254_wire_constant : std_logic_vector(7 downto 0);
    signal R_ASI_FLUSH_I_USER_1257_wire_constant : std_logic_vector(7 downto 0);
    signal R_ASI_MMU_REGISTER_1248_wire_constant : std_logic_vector(7 downto 0);
    signal R_REQUEST_TYPE_CCU_CACHE_WRITE_1238_wire_constant : std_logic_vector(3 downto 0);
    signal R_REQUEST_TYPE_WRITE_1235_wire_constant : std_logic_vector(3 downto 0);
    signal asi_without_head_bit_1232 : std_logic_vector(7 downto 0);
    signal is_write_1241 : std_logic_vector(0 downto 0);
    signal konst_1230_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    R_ASI_FLUSH_I_D_USER_1254_wire_constant <= "00010100";
    R_ASI_FLUSH_I_USER_1257_wire_constant <= "00011100";
    R_ASI_MMU_REGISTER_1248_wire_constant <= "00000100";
    R_REQUEST_TYPE_CCU_CACHE_WRITE_1238_wire_constant <= "0110";
    R_REQUEST_TYPE_WRITE_1235_wire_constant <= "0010";
    konst_1230_wire_constant <= "01111111";
    -- binary operator AND_u1_u1_1250_inst
    process(is_write_1241, EQ_u8_u1_1249_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(is_write_1241, EQ_u8_u1_1249_wire, tmp_var);
      is_mmu_ctrl_reg_write_buffer <= tmp_var; -- 
    end process;
    -- binary operator AND_u8_u8_1231_inst
    process(asi_buffer) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAnd_proc(asi_buffer, konst_1230_wire_constant, tmp_var);
      asi_without_head_bit_1232 <= tmp_var; -- 
    end process;
    -- binary operator EQ_u4_u1_1236_inst
    process(req_type_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(req_type_buffer, R_REQUEST_TYPE_WRITE_1235_wire_constant, tmp_var);
      EQ_u4_u1_1236_wire <= tmp_var; -- 
    end process;
    -- binary operator EQ_u4_u1_1239_inst
    process(req_type_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(req_type_buffer, R_REQUEST_TYPE_CCU_CACHE_WRITE_1238_wire_constant, tmp_var);
      EQ_u4_u1_1239_wire <= tmp_var; -- 
    end process;
    -- binary operator EQ_u8_u1_1249_inst
    process(asi_without_head_bit_1232) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(asi_without_head_bit_1232, R_ASI_MMU_REGISTER_1248_wire_constant, tmp_var);
      EQ_u8_u1_1249_wire <= tmp_var; -- 
    end process;
    -- binary operator EQ_u8_u1_1255_inst
    process(asi_without_head_bit_1232) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(asi_without_head_bit_1232, R_ASI_FLUSH_I_D_USER_1254_wire_constant, tmp_var);
      EQ_u8_u1_1255_wire <= tmp_var; -- 
    end process;
    -- binary operator EQ_u8_u1_1258_inst
    process(asi_without_head_bit_1232) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(asi_without_head_bit_1232, R_ASI_FLUSH_I_USER_1257_wire_constant, tmp_var);
      EQ_u8_u1_1258_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_1240_inst
    process(EQ_u4_u1_1236_wire, EQ_u4_u1_1239_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u4_u1_1236_wire, EQ_u4_u1_1239_wire, tmp_var);
      is_write_1241 <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_1259_inst
    process(EQ_u8_u1_1255_wire, EQ_u8_u1_1258_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u8_u1_1255_wire, EQ_u8_u1_1258_wire, tmp_var);
      flush_line_only_buffer <= tmp_var; -- 
    end process;
    volatile_operator_isDcacheFlushAsi_1702: isDcacheFlushAsi_VVD port map(asi => asi_without_head_bit_1232, ret_val => is_flush_asi_buffer); 
    -- 
  end Block; -- data_path
  -- 
end dcacheNeedsToBeFlushed_VVD_arch;

library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
entity isDcacheFlushAsi_VVD is -- 
  port ( -- 
    asi : in  std_logic_vector(7 downto 0);
    ret_val : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity isDcacheFlushAsi_VVD;
architecture isDcacheFlushAsi_VVD_arch of isDcacheFlushAsi_VVD is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(8-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal asi_buffer :  std_logic_vector(7 downto 0);
  -- output port buffer signals
  signal ret_val_buffer :  std_logic_vector(0 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  asi_buffer <= asi;
  -- output handling  -------------------------------------------------------
  ret_val <= ret_val_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal UGE_u8_u1_1215_wire : std_logic_vector(0 downto 0);
    signal ULE_u8_u1_1218_wire : std_logic_vector(0 downto 0);
    signal konst_1214_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1217_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    konst_1214_wire_constant <= "00010000";
    konst_1217_wire_constant <= "00010100";
    -- binary operator AND_u1_u1_1219_inst
    process(UGE_u8_u1_1215_wire, ULE_u8_u1_1218_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(UGE_u8_u1_1215_wire, ULE_u8_u1_1218_wire, tmp_var);
      ret_val_buffer <= tmp_var; -- 
    end process;
    -- binary operator UGE_u8_u1_1215_inst
    process(asi_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUge_proc(asi_buffer, konst_1214_wire_constant, tmp_var);
      UGE_u8_u1_1215_wire <= tmp_var; -- 
    end process;
    -- binary operator ULE_u8_u1_1218_inst
    process(asi_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUle_proc(asi_buffer, konst_1217_wire_constant, tmp_var);
      ULE_u8_u1_1218_wire <= tmp_var; -- 
    end process;
    -- 
  end Block; -- data_path
  -- 
end isDcacheFlushAsi_VVD_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
entity isMmuAccessAsi_VVD is -- 
  port ( -- 
    asi : in  std_logic_vector(7 downto 0);
    ret_val : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity isMmuAccessAsi_VVD;
architecture isMmuAccessAsi_VVD_arch of isMmuAccessAsi_VVD is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(8-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal asi_buffer :  std_logic_vector(7 downto 0);
  -- output port buffer signals
  signal ret_val_buffer :  std_logic_vector(0 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  asi_buffer <= asi;
  -- output handling  -------------------------------------------------------
  ret_val <= ret_val_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_1296_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_1274_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_1277_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_1281_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_1284_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_1289_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_1300_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1278_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1285_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1286_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1297_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1301_wire : std_logic_vector(0 downto 0);
    signal R_ASI_AJIT_BRIDGE_CONFIG_1299_wire_constant : std_logic_vector(7 downto 0);
    signal R_ASI_MMU_DIAGNOSTIC_IO_1288_wire_constant : std_logic_vector(7 downto 0);
    signal R_ASI_MMU_DIAGNOSTIC_I_1280_wire_constant : std_logic_vector(7 downto 0);
    signal R_ASI_MMU_DIAGNOSTIC_I_D_1283_wire_constant : std_logic_vector(7 downto 0);
    signal R_ASI_MMU_FLUSH_PROBE_1273_wire_constant : std_logic_vector(7 downto 0);
    signal R_ASI_MMU_REGISTER_1276_wire_constant : std_logic_vector(7 downto 0);
    signal UGE_u8_u1_1292_wire : std_logic_vector(0 downto 0);
    signal ULE_u8_u1_1295_wire : std_logic_vector(0 downto 0);
    signal konst_1291_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1294_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    R_ASI_AJIT_BRIDGE_CONFIG_1299_wire_constant <= "00110000";
    R_ASI_MMU_DIAGNOSTIC_IO_1288_wire_constant <= "00000111";
    R_ASI_MMU_DIAGNOSTIC_I_1280_wire_constant <= "00000101";
    R_ASI_MMU_DIAGNOSTIC_I_D_1283_wire_constant <= "00000110";
    R_ASI_MMU_FLUSH_PROBE_1273_wire_constant <= "00000011";
    R_ASI_MMU_REGISTER_1276_wire_constant <= "00000100";
    konst_1291_wire_constant <= "00100000";
    konst_1294_wire_constant <= "00101111";
    -- binary operator AND_u1_u1_1296_inst
    process(UGE_u8_u1_1292_wire, ULE_u8_u1_1295_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(UGE_u8_u1_1292_wire, ULE_u8_u1_1295_wire, tmp_var);
      AND_u1_u1_1296_wire <= tmp_var; -- 
    end process;
    -- binary operator EQ_u8_u1_1274_inst
    process(asi_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(asi_buffer, R_ASI_MMU_FLUSH_PROBE_1273_wire_constant, tmp_var);
      EQ_u8_u1_1274_wire <= tmp_var; -- 
    end process;
    -- binary operator EQ_u8_u1_1277_inst
    process(asi_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(asi_buffer, R_ASI_MMU_REGISTER_1276_wire_constant, tmp_var);
      EQ_u8_u1_1277_wire <= tmp_var; -- 
    end process;
    -- binary operator EQ_u8_u1_1281_inst
    process(asi_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(asi_buffer, R_ASI_MMU_DIAGNOSTIC_I_1280_wire_constant, tmp_var);
      EQ_u8_u1_1281_wire <= tmp_var; -- 
    end process;
    -- binary operator EQ_u8_u1_1284_inst
    process(asi_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(asi_buffer, R_ASI_MMU_DIAGNOSTIC_I_D_1283_wire_constant, tmp_var);
      EQ_u8_u1_1284_wire <= tmp_var; -- 
    end process;
    -- binary operator EQ_u8_u1_1289_inst
    process(asi_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(asi_buffer, R_ASI_MMU_DIAGNOSTIC_IO_1288_wire_constant, tmp_var);
      EQ_u8_u1_1289_wire <= tmp_var; -- 
    end process;
    -- binary operator EQ_u8_u1_1300_inst
    process(asi_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(asi_buffer, R_ASI_AJIT_BRIDGE_CONFIG_1299_wire_constant, tmp_var);
      EQ_u8_u1_1300_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_1278_inst
    process(EQ_u8_u1_1274_wire, EQ_u8_u1_1277_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u8_u1_1274_wire, EQ_u8_u1_1277_wire, tmp_var);
      OR_u1_u1_1278_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_1285_inst
    process(EQ_u8_u1_1281_wire, EQ_u8_u1_1284_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u8_u1_1281_wire, EQ_u8_u1_1284_wire, tmp_var);
      OR_u1_u1_1285_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_1286_inst
    process(OR_u1_u1_1278_wire, OR_u1_u1_1285_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_1278_wire, OR_u1_u1_1285_wire, tmp_var);
      OR_u1_u1_1286_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_1297_inst
    process(EQ_u8_u1_1289_wire, AND_u1_u1_1296_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u8_u1_1289_wire, AND_u1_u1_1296_wire, tmp_var);
      OR_u1_u1_1297_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_1301_inst
    process(OR_u1_u1_1297_wire, EQ_u8_u1_1300_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_1297_wire, EQ_u8_u1_1300_wire, tmp_var);
      OR_u1_u1_1301_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_1302_inst
    process(OR_u1_u1_1286_wire, OR_u1_u1_1301_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_1286_wire, OR_u1_u1_1301_wire, tmp_var);
      ret_val_buffer <= tmp_var; -- 
    end process;
    -- binary operator UGE_u8_u1_1292_inst
    process(asi_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUge_proc(asi_buffer, konst_1291_wire_constant, tmp_var);
      UGE_u8_u1_1292_wire <= tmp_var; -- 
    end process;
    -- binary operator ULE_u8_u1_1295_inst
    process(asi_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUle_proc(asi_buffer, konst_1294_wire_constant, tmp_var);
      ULE_u8_u1_1295_wire <= tmp_var; -- 
    end process;
    -- 
  end Block; -- data_path
  -- 
end isMmuAccessAsi_VVD_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
entity isSupervisorAsi_VVD is -- 
  port ( -- 
    asi : in  std_logic_vector(7 downto 0);
    ret_val : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity isSupervisorAsi_VVD;
architecture isSupervisorAsi_VVD_arch of isSupervisorAsi_VVD is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(8-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal asi_buffer :  std_logic_vector(7 downto 0);
  -- output port buffer signals
  signal ret_val_buffer :  std_logic_vector(0 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  asi_buffer <= asi;
  -- output handling  -------------------------------------------------------
  ret_val <= ret_val_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal EQ_u8_u1_657_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_660_wire : std_logic_vector(0 downto 0);
    signal R_ASI_SUPERVISOR_DATA_659_wire_constant : std_logic_vector(7 downto 0);
    signal R_ASI_SUPERVISOR_INSTRUCTION_656_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    R_ASI_SUPERVISOR_DATA_659_wire_constant <= "00001011";
    R_ASI_SUPERVISOR_INSTRUCTION_656_wire_constant <= "00001001";
    -- binary operator EQ_u8_u1_657_inst
    process(asi_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(asi_buffer, R_ASI_SUPERVISOR_INSTRUCTION_656_wire_constant, tmp_var);
      EQ_u8_u1_657_wire <= tmp_var; -- 
    end process;
    -- binary operator EQ_u8_u1_660_inst
    process(asi_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(asi_buffer, R_ASI_SUPERVISOR_DATA_659_wire_constant, tmp_var);
      EQ_u8_u1_660_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_661_inst
    process(EQ_u8_u1_657_wire, EQ_u8_u1_660_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u8_u1_657_wire, EQ_u8_u1_660_wire, tmp_var);
      ret_val_buffer <= tmp_var; -- 
    end process;
    -- 
  end Block; -- data_path
  -- 
end isSupervisorAsi_VVD_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
entity merge_and_decode_from_cpu_VVD is -- 
  port ( -- 
    from_cpu_fast : in  std_logic_vector(120 downto 0);
    from_cpu_slow : in  std_logic_vector(120 downto 0);
    is_thread_head : out  std_logic_vector(0 downto 0);
    lock_bus : out  std_logic_vector(0 downto 0);
    cpu_valid : out  std_logic_vector(0 downto 0);
    cpu_valid_fast : out  std_logic_vector(0 downto 0);
    cpu_valid_slow : out  std_logic_vector(0 downto 0);
    cpu_req_type : out  std_logic_vector(7 downto 0);
    cpu_asi : out  std_logic_vector(7 downto 0);
    cpu_byte_mask : out  std_logic_vector(7 downto 0);
    cpu_addr : out  std_logic_vector(31 downto 0);
    cpu_write_data : out  std_logic_vector(63 downto 0);
    is_flush_asi : out  std_logic_vector(0 downto 0);
    is_mmu_ctrl_reg_write : out  std_logic_vector(0 downto 0);
    flush_line_only : out  std_logic_vector(0 downto 0);
    is_supervisor_asi : out  std_logic_vector(0 downto 0);
    is_mmu_access_asi : out  std_logic_vector(0 downto 0);
    dcache_needs_to_be_flushed : out  std_logic_vector(0 downto 0);
    is_memory_read : out  std_logic_vector(0 downto 0);
    is_memory_write : out  std_logic_vector(0 downto 0);
    is_mmu_fsr_write : out  std_logic_vector(0 downto 0);
    is_stbar : out  std_logic_vector(0 downto 0);
    is_ccu_request : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity merge_and_decode_from_cpu_VVD;
architecture merge_and_decode_from_cpu_VVD_arch of merge_and_decode_from_cpu_VVD is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(242-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal from_cpu_fast_buffer :  std_logic_vector(120 downto 0);
  signal from_cpu_slow_buffer :  std_logic_vector(120 downto 0);
  -- output port buffer signals
  signal is_thread_head_buffer :  std_logic_vector(0 downto 0);
  signal lock_bus_buffer :  std_logic_vector(0 downto 0);
  signal cpu_valid_buffer :  std_logic_vector(0 downto 0);
  signal cpu_valid_fast_buffer :  std_logic_vector(0 downto 0);
  signal cpu_valid_slow_buffer :  std_logic_vector(0 downto 0);
  signal cpu_req_type_buffer :  std_logic_vector(7 downto 0);
  signal cpu_asi_buffer :  std_logic_vector(7 downto 0);
  signal cpu_byte_mask_buffer :  std_logic_vector(7 downto 0);
  signal cpu_addr_buffer :  std_logic_vector(31 downto 0);
  signal cpu_write_data_buffer :  std_logic_vector(63 downto 0);
  signal is_flush_asi_buffer :  std_logic_vector(0 downto 0);
  signal is_mmu_ctrl_reg_write_buffer :  std_logic_vector(0 downto 0);
  signal flush_line_only_buffer :  std_logic_vector(0 downto 0);
  signal is_supervisor_asi_buffer :  std_logic_vector(0 downto 0);
  signal is_mmu_access_asi_buffer :  std_logic_vector(0 downto 0);
  signal dcache_needs_to_be_flushed_buffer :  std_logic_vector(0 downto 0);
  signal is_memory_read_buffer :  std_logic_vector(0 downto 0);
  signal is_memory_write_buffer :  std_logic_vector(0 downto 0);
  signal is_mmu_fsr_write_buffer :  std_logic_vector(0 downto 0);
  signal is_stbar_buffer :  std_logic_vector(0 downto 0);
  signal is_ccu_request_buffer :  std_logic_vector(0 downto 0);
  -- volatile/operator module components. 
  component isMmuAccessAsi_VVD is -- 
    port ( -- 
      asi : in  std_logic_vector(7 downto 0);
      ret_val : out  std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component; 
  component isSupervisorAsi_VVD is -- 
    port ( -- 
      asi : in  std_logic_vector(7 downto 0);
      ret_val : out  std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component; 
  component dcacheNeedsToBeFlushed_VVD is -- 
    port ( -- 
      asi : in  std_logic_vector(7 downto 0);
      req_type : in  std_logic_vector(3 downto 0);
      is_flush_asi : out  std_logic_vector(0 downto 0);
      is_mmu_ctrl_reg_write : out  std_logic_vector(0 downto 0);
      flush_line_only : out  std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component; 
  -- 
begin --  
  -- input handling ------------------------------------------------
  from_cpu_fast_buffer <= from_cpu_fast;
  from_cpu_slow_buffer <= from_cpu_slow;
  -- output handling  -------------------------------------------------------
  is_thread_head <= is_thread_head_buffer;
  lock_bus <= lock_bus_buffer;
  cpu_valid <= cpu_valid_buffer;
  cpu_valid_fast <= cpu_valid_fast_buffer;
  cpu_valid_slow <= cpu_valid_slow_buffer;
  cpu_req_type <= cpu_req_type_buffer;
  cpu_asi <= cpu_asi_buffer;
  cpu_byte_mask <= cpu_byte_mask_buffer;
  cpu_addr <= cpu_addr_buffer;
  cpu_write_data <= cpu_write_data_buffer;
  is_flush_asi <= is_flush_asi_buffer;
  is_mmu_ctrl_reg_write <= is_mmu_ctrl_reg_write_buffer;
  flush_line_only <= flush_line_only_buffer;
  is_supervisor_asi <= is_supervisor_asi_buffer;
  is_mmu_access_asi <= is_mmu_access_asi_buffer;
  dcache_needs_to_be_flushed <= dcache_needs_to_be_flushed_buffer;
  is_memory_read <= is_memory_read_buffer;
  is_memory_write <= is_memory_write_buffer;
  is_mmu_fsr_write <= is_mmu_fsr_write_buffer;
  is_stbar <= is_stbar_buffer;
  is_ccu_request <= is_ccu_request_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal EQ_u4_u1_1455_wire : std_logic_vector(0 downto 0);
    signal EQ_u4_u1_1458_wire : std_logic_vector(0 downto 0);
    signal EQ_u4_u1_1464_wire : std_logic_vector(0 downto 0);
    signal EQ_u4_u1_1467_wire : std_logic_vector(0 downto 0);
    signal EQ_u4_u1_1483_wire : std_logic_vector(0 downto 0);
    signal EQ_u4_u1_1486_wire : std_logic_vector(0 downto 0);
    signal R_REQUEST_TYPE_CCU_CACHE_READ_1457_wire_constant : std_logic_vector(3 downto 0);
    signal R_REQUEST_TYPE_CCU_CACHE_READ_1482_wire_constant : std_logic_vector(3 downto 0);
    signal R_REQUEST_TYPE_CCU_CACHE_WRITE_1466_wire_constant : std_logic_vector(3 downto 0);
    signal R_REQUEST_TYPE_CCU_CACHE_WRITE_1485_wire_constant : std_logic_vector(3 downto 0);
    signal R_REQUEST_TYPE_READ_1454_wire_constant : std_logic_vector(3 downto 0);
    signal R_REQUEST_TYPE_STBAR_1477_wire_constant : std_logic_vector(3 downto 0);
    signal R_REQUEST_TYPE_WRFSRFAR_1472_wire_constant : std_logic_vector(3 downto 0);
    signal R_REQUEST_TYPE_WRITE_1463_wire_constant : std_logic_vector(3 downto 0);
    signal cpu_addr_fast_1348 : std_logic_vector(31 downto 0);
    signal cpu_addr_slow_1379 : std_logic_vector(31 downto 0);
    signal cpu_asi_fast_1340 : std_logic_vector(7 downto 0);
    signal cpu_asi_slow_1371 : std_logic_vector(7 downto 0);
    signal cpu_byte_mask_fast_1344 : std_logic_vector(7 downto 0);
    signal cpu_byte_mask_slow_1375 : std_logic_vector(7 downto 0);
    signal cpu_req_type_fast_1336 : std_logic_vector(7 downto 0);
    signal cpu_req_type_slow_1367 : std_logic_vector(7 downto 0);
    signal cpu_write_data_fast_1352 : std_logic_vector(63 downto 0);
    signal cpu_write_data_slow_1383 : std_logic_vector(63 downto 0);
    signal eff_crq_4_1434 : std_logic_vector(3 downto 0);
    signal from_cpu_1396 : std_logic_vector(120 downto 0);
    signal konst_1423_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1428_wire_constant : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    R_REQUEST_TYPE_CCU_CACHE_READ_1457_wire_constant <= "0101";
    R_REQUEST_TYPE_CCU_CACHE_READ_1482_wire_constant <= "0101";
    R_REQUEST_TYPE_CCU_CACHE_WRITE_1466_wire_constant <= "0110";
    R_REQUEST_TYPE_CCU_CACHE_WRITE_1485_wire_constant <= "0110";
    R_REQUEST_TYPE_READ_1454_wire_constant <= "0001";
    R_REQUEST_TYPE_STBAR_1477_wire_constant <= "0011";
    R_REQUEST_TYPE_WRFSRFAR_1472_wire_constant <= "0100";
    R_REQUEST_TYPE_WRITE_1463_wire_constant <= "0010";
    konst_1423_wire_constant <= "00000111";
    konst_1428_wire_constant <= "00000110";
    -- flow-through select operator MUX_1395_inst
    from_cpu_1396 <= from_cpu_fast_buffer when (cpu_valid_fast_buffer(0) /=  '0') else from_cpu_slow_buffer;
    -- flow-through slice operator slice_1331_inst
    cpu_valid_fast_buffer <= from_cpu_fast_buffer(120 downto 120);
    -- flow-through slice operator slice_1335_inst
    cpu_req_type_fast_1336 <= from_cpu_fast_buffer(119 downto 112);
    -- flow-through slice operator slice_1339_inst
    cpu_asi_fast_1340 <= from_cpu_fast_buffer(111 downto 104);
    -- flow-through slice operator slice_1343_inst
    cpu_byte_mask_fast_1344 <= from_cpu_fast_buffer(103 downto 96);
    -- flow-through slice operator slice_1347_inst
    cpu_addr_fast_1348 <= from_cpu_fast_buffer(95 downto 64);
    -- flow-through slice operator slice_1351_inst
    cpu_write_data_fast_1352 <= from_cpu_fast_buffer(63 downto 0);
    -- flow-through slice operator slice_1362_inst
    cpu_valid_slow_buffer <= from_cpu_slow_buffer(120 downto 120);
    -- flow-through slice operator slice_1366_inst
    cpu_req_type_slow_1367 <= from_cpu_slow_buffer(119 downto 112);
    -- flow-through slice operator slice_1370_inst
    cpu_asi_slow_1371 <= from_cpu_slow_buffer(111 downto 104);
    -- flow-through slice operator slice_1374_inst
    cpu_byte_mask_slow_1375 <= from_cpu_slow_buffer(103 downto 96);
    -- flow-through slice operator slice_1378_inst
    cpu_addr_slow_1379 <= from_cpu_slow_buffer(95 downto 64);
    -- flow-through slice operator slice_1382_inst
    cpu_write_data_slow_1383 <= from_cpu_slow_buffer(63 downto 0);
    -- flow-through slice operator slice_1399_inst
    cpu_valid_buffer <= from_cpu_1396(120 downto 120);
    -- flow-through slice operator slice_1403_inst
    cpu_req_type_buffer <= from_cpu_1396(119 downto 112);
    -- flow-through slice operator slice_1407_inst
    cpu_asi_buffer <= from_cpu_1396(111 downto 104);
    -- flow-through slice operator slice_1411_inst
    cpu_byte_mask_buffer <= from_cpu_1396(103 downto 96);
    -- flow-through slice operator slice_1415_inst
    cpu_addr_buffer <= from_cpu_1396(95 downto 64);
    -- flow-through slice operator slice_1419_inst
    cpu_write_data_buffer <= from_cpu_1396(63 downto 0);
    -- flow-through slice operator slice_1433_inst
    eff_crq_4_1434 <= cpu_req_type_buffer(3 downto 0);
    -- binary operator BITSEL_u8_u1_1424_inst
    process(cpu_req_type_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(cpu_req_type_buffer, konst_1423_wire_constant, tmp_var);
      is_thread_head_buffer <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u8_u1_1429_inst
    process(cpu_req_type_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(cpu_req_type_buffer, konst_1428_wire_constant, tmp_var);
      lock_bus_buffer <= tmp_var; -- 
    end process;
    -- binary operator EQ_u4_u1_1455_inst
    process(eff_crq_4_1434) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(eff_crq_4_1434, R_REQUEST_TYPE_READ_1454_wire_constant, tmp_var);
      EQ_u4_u1_1455_wire <= tmp_var; -- 
    end process;
    -- binary operator EQ_u4_u1_1458_inst
    process(eff_crq_4_1434) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(eff_crq_4_1434, R_REQUEST_TYPE_CCU_CACHE_READ_1457_wire_constant, tmp_var);
      EQ_u4_u1_1458_wire <= tmp_var; -- 
    end process;
    -- binary operator EQ_u4_u1_1464_inst
    process(eff_crq_4_1434) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(eff_crq_4_1434, R_REQUEST_TYPE_WRITE_1463_wire_constant, tmp_var);
      EQ_u4_u1_1464_wire <= tmp_var; -- 
    end process;
    -- binary operator EQ_u4_u1_1467_inst
    process(eff_crq_4_1434) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(eff_crq_4_1434, R_REQUEST_TYPE_CCU_CACHE_WRITE_1466_wire_constant, tmp_var);
      EQ_u4_u1_1467_wire <= tmp_var; -- 
    end process;
    -- binary operator EQ_u4_u1_1473_inst
    process(eff_crq_4_1434) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(eff_crq_4_1434, R_REQUEST_TYPE_WRFSRFAR_1472_wire_constant, tmp_var);
      is_mmu_fsr_write_buffer <= tmp_var; -- 
    end process;
    -- binary operator EQ_u4_u1_1478_inst
    process(eff_crq_4_1434) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(eff_crq_4_1434, R_REQUEST_TYPE_STBAR_1477_wire_constant, tmp_var);
      is_stbar_buffer <= tmp_var; -- 
    end process;
    -- binary operator EQ_u4_u1_1483_inst
    process(eff_crq_4_1434) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(eff_crq_4_1434, R_REQUEST_TYPE_CCU_CACHE_READ_1482_wire_constant, tmp_var);
      EQ_u4_u1_1483_wire <= tmp_var; -- 
    end process;
    -- binary operator EQ_u4_u1_1486_inst
    process(eff_crq_4_1434) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(eff_crq_4_1434, R_REQUEST_TYPE_CCU_CACHE_WRITE_1485_wire_constant, tmp_var);
      EQ_u4_u1_1486_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_1450_inst
    process(is_flush_asi_buffer, is_mmu_ctrl_reg_write_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(is_flush_asi_buffer, is_mmu_ctrl_reg_write_buffer, tmp_var);
      dcache_needs_to_be_flushed_buffer <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_1459_inst
    process(EQ_u4_u1_1455_wire, EQ_u4_u1_1458_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u4_u1_1455_wire, EQ_u4_u1_1458_wire, tmp_var);
      is_memory_read_buffer <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_1468_inst
    process(EQ_u4_u1_1464_wire, EQ_u4_u1_1467_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u4_u1_1464_wire, EQ_u4_u1_1467_wire, tmp_var);
      is_memory_write_buffer <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_1487_inst
    process(EQ_u4_u1_1483_wire, EQ_u4_u1_1486_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u4_u1_1483_wire, EQ_u4_u1_1486_wire, tmp_var);
      is_ccu_request_buffer <= tmp_var; -- 
    end process;
    volatile_operator_dcacheNeedsToBeFlushed_1849: dcacheNeedsToBeFlushed_VVD port map(asi => cpu_asi_buffer, req_type => eff_crq_4_1434, is_flush_asi => is_flush_asi_buffer, is_mmu_ctrl_reg_write => is_mmu_ctrl_reg_write_buffer, flush_line_only => flush_line_only_buffer); 
    volatile_operator_isSupervisorAsi_1850: isSupervisorAsi_VVD port map(asi => cpu_asi_buffer, ret_val => is_supervisor_asi_buffer); 
    volatile_operator_isMmuAccessAsi_1851: isMmuAccessAsi_VVD port map(asi => cpu_asi_buffer, ret_val => is_mmu_access_asi_buffer); 
    -- 
  end Block; -- data_path
  -- 
end merge_and_decode_from_cpu_VVD_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
entity offsetInLine_VVD is -- 
  port ( -- 
    addr : in  std_logic_vector(31 downto 0);
    ret_val : out  std_logic_vector(3 downto 0)-- 
  );
  -- 
end entity offsetInLine_VVD;
architecture offsetInLine_VVD_arch of offsetInLine_VVD is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(32-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal addr_buffer :  std_logic_vector(31 downto 0);
  -- output port buffer signals
  signal ret_val_buffer :  std_logic_vector(3 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  addr_buffer <= addr;
  -- output handling  -------------------------------------------------------
  ret_val <= ret_val_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal konst_777_wire_constant : std_logic_vector(3 downto 0);
    signal slice_776_wire : std_logic_vector(3 downto 0);
    -- 
  begin -- 
    konst_777_wire_constant <= "0111";
    -- flow-through slice operator slice_776_inst
    slice_776_wire <= addr_buffer(6 downto 3);
    -- binary operator AND_u4_u4_778_inst
    process(slice_776_wire) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApIntAnd_proc(slice_776_wire, konst_777_wire_constant, tmp_var);
      ret_val_buffer <= tmp_var; -- 
    end process;
    -- 
  end Block; -- data_path
  -- 
end offsetInLine_VVD_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
entity identify_cpu_actions_VVD is -- 
  port ( -- 
    exec_cpu : in  std_logic_vector(0 downto 0);
    next_dcache_trapped : in  std_logic_vector(0 downto 0);
    is_ccu_request : in  std_logic_vector(0 downto 0);
    is_a_hit : in  std_logic_vector(0 downto 0);
    skip_tag_lookup : in  std_logic_vector(0 downto 0);
    is_memory_write : in  std_logic_vector(0 downto 0);
    is_memory_read : in  std_logic_vector(0 downto 0);
    is_flush_asi : in  std_logic_vector(0 downto 0);
    is_stbar : in  std_logic_vector(0 downto 0);
    is_mmu_access_asi : in  std_logic_vector(0 downto 0);
    is_mmu_fsr_write : in  std_logic_vector(0 downto 0);
    write_dword_hit : out  std_logic_vector(0 downto 0);
    write_dword_miss : out  std_logic_vector(0 downto 0);
    read_dword_hit : out  std_logic_vector(0 downto 0);
    read_dword_miss : out  std_logic_vector(0 downto 0);
    finished_flush_or_nop : out  std_logic_vector(0 downto 0);
    write_to_mmu_or_bypass : out  std_logic_vector(0 downto 0);
    read_from_mmu_or_bypass : out  std_logic_vector(0 downto 0);
    write_to_mmu_fsr : out  std_logic_vector(0 downto 0);
    send_to_be : out  std_logic_vector(0 downto 0);
    no_response_from_be : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity identify_cpu_actions_VVD;
architecture identify_cpu_actions_VVD_arch of identify_cpu_actions_VVD is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(11-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal exec_cpu_buffer :  std_logic_vector(0 downto 0);
  signal next_dcache_trapped_buffer :  std_logic_vector(0 downto 0);
  signal is_ccu_request_buffer :  std_logic_vector(0 downto 0);
  signal is_a_hit_buffer :  std_logic_vector(0 downto 0);
  signal skip_tag_lookup_buffer :  std_logic_vector(0 downto 0);
  signal is_memory_write_buffer :  std_logic_vector(0 downto 0);
  signal is_memory_read_buffer :  std_logic_vector(0 downto 0);
  signal is_flush_asi_buffer :  std_logic_vector(0 downto 0);
  signal is_stbar_buffer :  std_logic_vector(0 downto 0);
  signal is_mmu_access_asi_buffer :  std_logic_vector(0 downto 0);
  signal is_mmu_fsr_write_buffer :  std_logic_vector(0 downto 0);
  -- output port buffer signals
  signal write_dword_hit_buffer :  std_logic_vector(0 downto 0);
  signal write_dword_miss_buffer :  std_logic_vector(0 downto 0);
  signal read_dword_hit_buffer :  std_logic_vector(0 downto 0);
  signal read_dword_miss_buffer :  std_logic_vector(0 downto 0);
  signal finished_flush_or_nop_buffer :  std_logic_vector(0 downto 0);
  signal write_to_mmu_or_bypass_buffer :  std_logic_vector(0 downto 0);
  signal read_from_mmu_or_bypass_buffer :  std_logic_vector(0 downto 0);
  signal write_to_mmu_fsr_buffer :  std_logic_vector(0 downto 0);
  signal send_to_be_buffer :  std_logic_vector(0 downto 0);
  signal no_response_from_be_buffer :  std_logic_vector(0 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  exec_cpu_buffer <= exec_cpu;
  next_dcache_trapped_buffer <= next_dcache_trapped;
  is_ccu_request_buffer <= is_ccu_request;
  is_a_hit_buffer <= is_a_hit;
  skip_tag_lookup_buffer <= skip_tag_lookup;
  is_memory_write_buffer <= is_memory_write;
  is_memory_read_buffer <= is_memory_read;
  is_flush_asi_buffer <= is_flush_asi;
  is_stbar_buffer <= is_stbar;
  is_mmu_access_asi_buffer <= is_mmu_access_asi;
  is_mmu_fsr_write_buffer <= is_mmu_fsr_write;
  -- output handling  -------------------------------------------------------
  write_dword_hit <= write_dword_hit_buffer;
  write_dword_miss <= write_dword_miss_buffer;
  read_dword_hit <= read_dword_hit_buffer;
  read_dword_miss <= read_dword_miss_buffer;
  finished_flush_or_nop <= finished_flush_or_nop_buffer;
  write_to_mmu_or_bypass <= write_to_mmu_or_bypass_buffer;
  read_from_mmu_or_bypass <= read_from_mmu_or_bypass_buffer;
  write_to_mmu_fsr <= write_to_mmu_fsr_buffer;
  send_to_be <= send_to_be_buffer;
  no_response_from_be <= no_response_from_be_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_2199_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_2202_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_2211_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_2215_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_2224_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_2227_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_2236_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_2240_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_2248_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_2251_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_2257_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_2264_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_2190_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_2198_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_2210_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_2213_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_2223_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_2235_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_2238_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_2192_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_2276_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_2278_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_2281_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_2283_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_2289_wire : std_logic_vector(0 downto 0);
    signal run_this_transaction_2194 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    -- binary operator AND_u1_u1_2193_inst
    process(exec_cpu_buffer, OR_u1_u1_2192_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(exec_cpu_buffer, OR_u1_u1_2192_wire, tmp_var);
      run_this_transaction_2194 <= tmp_var; -- 
    end process;
    -- binary operator AND_u1_u1_2199_inst
    process(run_this_transaction_2194, NOT_u1_u1_2198_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(run_this_transaction_2194, NOT_u1_u1_2198_wire, tmp_var);
      AND_u1_u1_2199_wire <= tmp_var; -- 
    end process;
    -- binary operator AND_u1_u1_2202_inst
    process(is_a_hit_buffer, is_memory_write_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(is_a_hit_buffer, is_memory_write_buffer, tmp_var);
      AND_u1_u1_2202_wire <= tmp_var; -- 
    end process;
    -- binary operator AND_u1_u1_2203_inst
    process(AND_u1_u1_2199_wire, AND_u1_u1_2202_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_2199_wire, AND_u1_u1_2202_wire, tmp_var);
      write_dword_hit_buffer <= tmp_var; -- 
    end process;
    -- binary operator AND_u1_u1_2211_inst
    process(run_this_transaction_2194, NOT_u1_u1_2210_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(run_this_transaction_2194, NOT_u1_u1_2210_wire, tmp_var);
      AND_u1_u1_2211_wire <= tmp_var; -- 
    end process;
    -- binary operator AND_u1_u1_2215_inst
    process(NOT_u1_u1_2213_wire, is_memory_write_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_2213_wire, is_memory_write_buffer, tmp_var);
      AND_u1_u1_2215_wire <= tmp_var; -- 
    end process;
    -- binary operator AND_u1_u1_2216_inst
    process(AND_u1_u1_2211_wire, AND_u1_u1_2215_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_2211_wire, AND_u1_u1_2215_wire, tmp_var);
      write_dword_miss_buffer <= tmp_var; -- 
    end process;
    -- binary operator AND_u1_u1_2224_inst
    process(run_this_transaction_2194, NOT_u1_u1_2223_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(run_this_transaction_2194, NOT_u1_u1_2223_wire, tmp_var);
      AND_u1_u1_2224_wire <= tmp_var; -- 
    end process;
    -- binary operator AND_u1_u1_2227_inst
    process(is_a_hit_buffer, is_memory_read_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(is_a_hit_buffer, is_memory_read_buffer, tmp_var);
      AND_u1_u1_2227_wire <= tmp_var; -- 
    end process;
    -- binary operator AND_u1_u1_2228_inst
    process(AND_u1_u1_2224_wire, AND_u1_u1_2227_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_2224_wire, AND_u1_u1_2227_wire, tmp_var);
      read_dword_hit_buffer <= tmp_var; -- 
    end process;
    -- binary operator AND_u1_u1_2236_inst
    process(run_this_transaction_2194, NOT_u1_u1_2235_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(run_this_transaction_2194, NOT_u1_u1_2235_wire, tmp_var);
      AND_u1_u1_2236_wire <= tmp_var; -- 
    end process;
    -- binary operator AND_u1_u1_2240_inst
    process(NOT_u1_u1_2238_wire, is_memory_read_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_2238_wire, is_memory_read_buffer, tmp_var);
      AND_u1_u1_2240_wire <= tmp_var; -- 
    end process;
    -- binary operator AND_u1_u1_2241_inst
    process(AND_u1_u1_2236_wire, AND_u1_u1_2240_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_2236_wire, AND_u1_u1_2240_wire, tmp_var);
      read_dword_miss_buffer <= tmp_var; -- 
    end process;
    -- binary operator AND_u1_u1_2248_inst
    process(run_this_transaction_2194, exec_cpu_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(run_this_transaction_2194, exec_cpu_buffer, tmp_var);
      AND_u1_u1_2248_wire <= tmp_var; -- 
    end process;
    -- binary operator AND_u1_u1_2251_inst
    process(is_flush_asi_buffer, is_stbar_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(is_flush_asi_buffer, is_stbar_buffer, tmp_var);
      AND_u1_u1_2251_wire <= tmp_var; -- 
    end process;
    -- binary operator AND_u1_u1_2252_inst
    process(AND_u1_u1_2248_wire, AND_u1_u1_2251_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_2248_wire, AND_u1_u1_2251_wire, tmp_var);
      finished_flush_or_nop_buffer <= tmp_var; -- 
    end process;
    -- binary operator AND_u1_u1_2257_inst
    process(run_this_transaction_2194, is_mmu_access_asi_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(run_this_transaction_2194, is_mmu_access_asi_buffer, tmp_var);
      AND_u1_u1_2257_wire <= tmp_var; -- 
    end process;
    -- binary operator AND_u1_u1_2259_inst
    process(AND_u1_u1_2257_wire, is_memory_write_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_2257_wire, is_memory_write_buffer, tmp_var);
      write_to_mmu_or_bypass_buffer <= tmp_var; -- 
    end process;
    -- binary operator AND_u1_u1_2264_inst
    process(run_this_transaction_2194, is_mmu_access_asi_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(run_this_transaction_2194, is_mmu_access_asi_buffer, tmp_var);
      AND_u1_u1_2264_wire <= tmp_var; -- 
    end process;
    -- binary operator AND_u1_u1_2266_inst
    process(AND_u1_u1_2264_wire, is_memory_read_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_2264_wire, is_memory_read_buffer, tmp_var);
      read_from_mmu_or_bypass_buffer <= tmp_var; -- 
    end process;
    -- binary operator AND_u1_u1_2271_inst
    process(exec_cpu_buffer, is_mmu_fsr_write_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(exec_cpu_buffer, is_mmu_fsr_write_buffer, tmp_var);
      write_to_mmu_fsr_buffer <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_2190_inst
    process(next_dcache_trapped_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", next_dcache_trapped_buffer, tmp_var);
      NOT_u1_u1_2190_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_2198_inst
    process(skip_tag_lookup_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_tag_lookup_buffer, tmp_var);
      NOT_u1_u1_2198_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_2210_inst
    process(skip_tag_lookup_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_tag_lookup_buffer, tmp_var);
      NOT_u1_u1_2210_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_2213_inst
    process(is_a_hit_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", is_a_hit_buffer, tmp_var);
      NOT_u1_u1_2213_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_2223_inst
    process(skip_tag_lookup_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_tag_lookup_buffer, tmp_var);
      NOT_u1_u1_2223_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_2235_inst
    process(skip_tag_lookup_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", skip_tag_lookup_buffer, tmp_var);
      NOT_u1_u1_2235_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_2238_inst
    process(is_a_hit_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", is_a_hit_buffer, tmp_var);
      NOT_u1_u1_2238_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_2192_inst
    process(NOT_u1_u1_2190_wire, is_ccu_request_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_2190_wire, is_ccu_request_buffer, tmp_var);
      OR_u1_u1_2192_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_2276_inst
    process(read_dword_miss_buffer, write_dword_miss_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(read_dword_miss_buffer, write_dword_miss_buffer, tmp_var);
      OR_u1_u1_2276_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_2278_inst
    process(OR_u1_u1_2276_wire, write_dword_hit_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_2276_wire, write_dword_hit_buffer, tmp_var);
      OR_u1_u1_2278_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_2281_inst
    process(write_to_mmu_or_bypass_buffer, read_from_mmu_or_bypass_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(write_to_mmu_or_bypass_buffer, read_from_mmu_or_bypass_buffer, tmp_var);
      OR_u1_u1_2281_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_2283_inst
    process(OR_u1_u1_2281_wire, write_to_mmu_fsr_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_2281_wire, write_to_mmu_fsr_buffer, tmp_var);
      OR_u1_u1_2283_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_2284_inst
    process(OR_u1_u1_2278_wire, OR_u1_u1_2283_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_2278_wire, OR_u1_u1_2283_wire, tmp_var);
      send_to_be_buffer <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_2289_inst
    process(write_dword_hit_buffer, write_to_mmu_or_bypass_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(write_dword_hit_buffer, write_to_mmu_or_bypass_buffer, tmp_var);
      OR_u1_u1_2289_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_2291_inst
    process(OR_u1_u1_2289_wire, write_to_mmu_fsr_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_2289_wire, write_to_mmu_fsr_buffer, tmp_var);
      no_response_from_be_buffer <= tmp_var; -- 
    end process;
    -- 
  end Block; -- data_path
  -- 
end identify_cpu_actions_VVD_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
entity parse_from_backend_Volatile is -- 
  port ( -- 
    from_be : in  std_logic_vector(83 downto 0);
    be_valid : out  std_logic_vector(0 downto 0);
    be_counter : out  std_logic_vector(2 downto 0);
    be_tag_command : out  std_logic_vector(2 downto 0);
    be_array_command : out  std_logic_vector(2 downto 0);
    be_dword_id : out  std_logic_vector(2 downto 0);
    be_last_dword : out  std_logic_vector(0 downto 0);
    be_acc : out  std_logic_vector(2 downto 0);
    be_cacheable : out  std_logic_vector(0 downto 0);
    be_mae : out  std_logic_vector(0 downto 0);
    be_access_error : out  std_logic_vector(0 downto 0);
    be_dword : out  std_logic_vector(63 downto 0)-- 
  );
  -- 
end entity parse_from_backend_Volatile;
architecture parse_from_backend_Volatile_arch of parse_from_backend_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(84-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal from_be_buffer :  std_logic_vector(83 downto 0);
  -- output port buffer signals
  signal be_valid_buffer :  std_logic_vector(0 downto 0);
  signal be_counter_buffer :  std_logic_vector(2 downto 0);
  signal be_tag_command_buffer :  std_logic_vector(2 downto 0);
  signal be_array_command_buffer :  std_logic_vector(2 downto 0);
  signal be_dword_id_buffer :  std_logic_vector(2 downto 0);
  signal be_last_dword_buffer :  std_logic_vector(0 downto 0);
  signal be_acc_buffer :  std_logic_vector(2 downto 0);
  signal be_cacheable_buffer :  std_logic_vector(0 downto 0);
  signal be_mae_buffer :  std_logic_vector(0 downto 0);
  signal be_access_error_buffer :  std_logic_vector(0 downto 0);
  signal be_dword_buffer :  std_logic_vector(63 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  from_be_buffer <= from_be;
  -- output handling  -------------------------------------------------------
  be_valid <= be_valid_buffer;
  be_counter <= be_counter_buffer;
  be_tag_command <= be_tag_command_buffer;
  be_array_command <= be_array_command_buffer;
  be_dword_id <= be_dword_id_buffer;
  be_last_dword <= be_last_dword_buffer;
  be_acc <= be_acc_buffer;
  be_cacheable <= be_cacheable_buffer;
  be_mae <= be_mae_buffer;
  be_access_error <= be_access_error_buffer;
  be_dword <= be_dword_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    -- 
  begin -- 
    -- flow-through slice operator slice_1550_inst
    be_valid_buffer <= from_be_buffer(83 downto 83);
    -- flow-through slice operator slice_1554_inst
    be_counter_buffer <= from_be_buffer(82 downto 80);
    -- flow-through slice operator slice_1558_inst
    be_tag_command_buffer <= from_be_buffer(79 downto 77);
    -- flow-through slice operator slice_1562_inst
    be_array_command_buffer <= from_be_buffer(76 downto 74);
    -- flow-through slice operator slice_1566_inst
    be_dword_id_buffer <= from_be_buffer(73 downto 71);
    -- flow-through slice operator slice_1570_inst
    be_last_dword_buffer <= from_be_buffer(70 downto 70);
    -- flow-through slice operator slice_1574_inst
    be_acc_buffer <= from_be_buffer(69 downto 67);
    -- flow-through slice operator slice_1578_inst
    be_cacheable_buffer <= from_be_buffer(66 downto 66);
    -- flow-through slice operator slice_1582_inst
    be_mae_buffer <= from_be_buffer(65 downto 65);
    -- flow-through slice operator slice_1586_inst
    be_access_error_buffer <= from_be_buffer(64 downto 64);
    -- flow-through slice operator slice_1590_inst
    be_dword_buffer <= from_be_buffer(63 downto 0);
    -- 
  end Block; -- data_path
  -- 
end parse_from_backend_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
entity parse_from_frontend_Volatile is -- 
  port ( -- 
    from_frontend : in  std_logic_vector(119 downto 0);
    no_response_to_fe : out  std_logic_vector(0 downto 0);
    lock_bus : out  std_logic_vector(0 downto 0);
    read_miss : out  std_logic_vector(0 downto 0);
    write_miss : out  std_logic_vector(0 downto 0);
    write_hit : out  std_logic_vector(0 downto 0);
    read_bypass : out  std_logic_vector(0 downto 0);
    write_bypass : out  std_logic_vector(0 downto 0);
    write_fsr : out  std_logic_vector(0 downto 0);
    asi : out  std_logic_vector(7 downto 0);
    byte_mask : out  std_logic_vector(7 downto 0);
    addr : out  std_logic_vector(31 downto 0);
    write_data : out  std_logic_vector(63 downto 0)-- 
  );
  -- 
end entity parse_from_frontend_Volatile;
architecture parse_from_frontend_Volatile_arch of parse_from_frontend_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(120-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal from_frontend_buffer :  std_logic_vector(119 downto 0);
  -- output port buffer signals
  signal no_response_to_fe_buffer :  std_logic_vector(0 downto 0);
  signal lock_bus_buffer :  std_logic_vector(0 downto 0);
  signal read_miss_buffer :  std_logic_vector(0 downto 0);
  signal write_miss_buffer :  std_logic_vector(0 downto 0);
  signal write_hit_buffer :  std_logic_vector(0 downto 0);
  signal read_bypass_buffer :  std_logic_vector(0 downto 0);
  signal write_bypass_buffer :  std_logic_vector(0 downto 0);
  signal write_fsr_buffer :  std_logic_vector(0 downto 0);
  signal asi_buffer :  std_logic_vector(7 downto 0);
  signal byte_mask_buffer :  std_logic_vector(7 downto 0);
  signal addr_buffer :  std_logic_vector(31 downto 0);
  signal write_data_buffer :  std_logic_vector(63 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  from_frontend_buffer <= from_frontend;
  -- output handling  -------------------------------------------------------
  no_response_to_fe <= no_response_to_fe_buffer;
  lock_bus <= lock_bus_buffer;
  read_miss <= read_miss_buffer;
  write_miss <= write_miss_buffer;
  write_hit <= write_hit_buffer;
  read_bypass <= read_bypass_buffer;
  write_bypass <= write_bypass_buffer;
  write_fsr <= write_fsr_buffer;
  asi <= asi_buffer;
  byte_mask <= byte_mask_buffer;
  addr <= addr_buffer;
  write_data <= write_data_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    -- 
  begin -- 
    -- flow-through slice operator slice_676_inst
    no_response_to_fe_buffer <= from_frontend_buffer(119 downto 119);
    -- flow-through slice operator slice_680_inst
    lock_bus_buffer <= from_frontend_buffer(118 downto 118);
    -- flow-through slice operator slice_684_inst
    read_miss_buffer <= from_frontend_buffer(117 downto 117);
    -- flow-through slice operator slice_688_inst
    write_miss_buffer <= from_frontend_buffer(116 downto 116);
    -- flow-through slice operator slice_692_inst
    write_hit_buffer <= from_frontend_buffer(115 downto 115);
    -- flow-through slice operator slice_696_inst
    read_bypass_buffer <= from_frontend_buffer(114 downto 114);
    -- flow-through slice operator slice_700_inst
    write_bypass_buffer <= from_frontend_buffer(113 downto 113);
    -- flow-through slice operator slice_704_inst
    write_fsr_buffer <= from_frontend_buffer(112 downto 112);
    -- flow-through slice operator slice_708_inst
    asi_buffer <= from_frontend_buffer(111 downto 104);
    -- flow-through slice operator slice_712_inst
    byte_mask_buffer <= from_frontend_buffer(103 downto 96);
    -- flow-through slice operator slice_716_inst
    addr_buffer <= from_frontend_buffer(95 downto 64);
    -- flow-through slice operator slice_720_inst
    write_data_buffer <= from_frontend_buffer(63 downto 0);
    -- 
  end Block; -- data_path
  -- 
end parse_from_frontend_Volatile_arch;
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.basecomponents.all;


-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

entity DcacheBypassController is -- 
  port ( -- 

    cpu_bypass_command_available: in  boolean; 
    cpu_bypass_command_accept   : out boolean;

    cpu_fast_valid		: in std_logic;
    cpu_slow_valid		: in std_logic;

    is_memory_write		: in std_logic;
    locked_access		: in std_logic;

    cpu_asi		        : in std_logic_vector(7 downto 0);
    cpu_byte_mask	        : in std_logic_vector(7 downto 0);
    cpu_address			: in std_logic_vector(31 downto 0);
    cpu_write_data		: in std_logic_vector(63 downto 0);

    cpu_slow_ready_for_bypass_response      : in boolean;
    write_to_cpu_slow		            : out boolean;

    cpu_fast_ready_for_bypass_response      : in boolean;
    write_to_cpu_fast		            : out boolean;

    response_to_cpu		: out std_logic_vector(71 downto 0);

    be_ready_for_request	: in boolean;
    be_write		       	: out boolean;
    to_be_from_bypass 		: out  std_logic_vector(119 downto 0);

    be_response_ready		: in boolean;
    be_read			: out boolean;
    be_dword			: in std_logic_vector(63 downto 0);

    bypass_response_pending : out boolean;

    clk : in std_logic;
    reset : in std_logic
  );
  -- 
end entity DcacheBypassController;

architecture DcacheBypassController_arch of DcacheBypassController is -- 
    
	-------------------------------------------------------------------------
	-- initial registering
	-------------------------------------------------------------------------
	signal cpu_fast_valid_reg		: std_logic;
    	signal cpu_slow_valid_reg		: std_logic;

    	signal is_memory_write_reg		: std_logic;
    	signal locked_access_reg		: std_logic;

    	signal cpu_asi_reg		        : std_logic_vector(7 downto 0);
    	signal cpu_byte_mask_reg	        : std_logic_vector(7 downto 0);
    	signal cpu_address_reg			: std_logic_vector(31 downto 0);
    	signal cpu_write_data_reg		: std_logic_vector(63 downto 0);

	-------------------------------------------------------------------------
	-- forwarding the response...
	-------------------------------------------------------------------------
	signal forward_bypass_response, forward_bypass_to_fast, forward_bypass_to_slow: boolean;
	signal forward_zero_bypass_response: boolean;

	-------------------------------------------------------------------------
	-- bypass assist logic
	-------------------------------------------------------------------------
	signal bypass_queue_push_req, bypass_queue_push_ack: std_logic;
	signal bypass_queue_pop_req, bypass_queue_pop_ack: std_logic;

	-- fields
	-- [2] = cpu_fast_valid
	-- [1] = cpu_slow_valid
	-- [0] = send_zero_response
	signal bypass_queue_push_data, bypass_queue_pop_data: std_logic_vector(2 downto 0);

	signal data_to_cpu: std_logic_vector(63 downto 0);
	constant MAE8: std_logic_vector(7 downto 0) := (others => '0');
	constant ZERO_1: std_logic_vector(0 downto 0) := (others => '0');
	constant ZERO_64: std_logic_vector(63 downto 0) := (others => '0');
	

	type FsmState is (IDLE, READY_TO_SEND);
	signal fsm_state : FsmState;

	signal cpu_command_available_to_be: boolean;
    		

-- see comment above..
--##decl_synopsys_sync_set_reset##

begin
	--------------------------------------------------------------------------------------
	-- control FSM and registering: need to delay by one cycle to ensure that
	-- the bypass timing is aligned with the normal timing (fixing a bug!).
	--------------------------------------------------------------------------------------
	process(clk, reset, cpu_bypass_command_available, be_ready_for_request, 
			bypass_queue_push_ack, fsm_state)
		variable next_fsm_state_var: FsmState;
		variable command_ready_var, command_accept_var: boolean;
		variable latch_cpu_info_var: boolean;
	begin
		next_fsm_state_var := fsm_state;
		command_ready_var  := false;
		command_accept_var := false;
		latch_cpu_info_var := false;

		case fsm_state is 
			when IDLE =>
				command_accept_var := true;
				if(cpu_bypass_command_available) then
					next_fsm_state_var := READY_TO_SEND;
					latch_cpu_info_var := true;
				end if;
			when READY_TO_SEND =>
				command_ready_var := true;
				if(be_ready_for_request and (bypass_queue_push_ack = '1')) then
					command_accept_var := true;
					if(cpu_bypass_command_available) then
						latch_cpu_info_var := true;
					else
						next_fsm_state_var := IDLE;
					end if;
				end if;
		end case;
		
		cpu_bypass_command_accept <= command_accept_var;
		cpu_command_available_to_be   <= command_ready_var;


		if (clk'event and (clk = '1')) then
			if(reset = '1') then
				fsm_state <= IDLE;
			else
				fsm_state <= next_fsm_state_var;
				if(latch_cpu_info_var) then
					cpu_fast_valid_reg <= cpu_fast_valid;
					cpu_slow_valid_reg <= cpu_slow_valid;
					is_memory_write_reg <= is_memory_write;
					locked_access_reg <= locked_access;
					cpu_asi_reg <= cpu_asi;
					cpu_byte_mask_reg <= cpu_byte_mask;
					cpu_address_reg <= cpu_address;
					cpu_write_data_reg <= cpu_write_data;
				end if;
			end if;
		end if;
	end process;
	
	--------------------------------------------------------------------------------------
	-- bypass..
	--------------------------------------------------------------------------------------
	bypass_response_pending <= (fsm_state = READY_TO_SEND) or (bypass_queue_pop_ack = '1');

	-- BE, COMMAND, QUEUE interaction.
	
	-- push into the queue when BE, CMD are ready.
	bypass_queue_push_req <= '1' when cpu_command_available_to_be and be_ready_for_request else '0';
	-- Write to BE when CMD, Queue are ready. 
	be_write <= cpu_command_available_to_be and (bypass_queue_push_ack = '1');


	-- fields
	-- [2] = cpu_fast_valid
	-- [1] = cpu_slow_valid
	-- [0] = send_zero_response
	bypass_queue_push_data(2) <=  cpu_fast_valid_reg;
	bypass_queue_push_data(1) <=  cpu_slow_valid_reg;
	bypass_queue_push_data(0) <=  is_memory_write_reg;
	
	to_be_from_bypass <= 
			( is_memory_write_reg &
				locked_access_reg & 
				ZERO_1 & -- read miss
				ZERO_1 & -- write miss
				ZERO_1 & -- write hit
				(not is_memory_write_reg)	&
				is_memory_write_reg &
				ZERO_1 & -- write fsr
				cpu_asi_reg & 
				cpu_byte_mask_reg &
				cpu_address_reg &
				cpu_write_data_reg);

	bypQueue: QueueBase generic map
				(name => "DcacheBypassResponseQueue",
					queue_depth => 8,
					data_width  => 3, save_one_slot => false)
			port map (
				clk => clk, reset => reset,
				push_req => bypass_queue_push_req,
				push_ack => bypass_queue_push_ack,
				pop_req =>  bypass_queue_pop_req,
				pop_ack =>  bypass_queue_pop_ack,
				data_in =>  bypass_queue_push_data,
				data_out => bypass_queue_pop_data
			);

	forward_bypass_response <= 
			((bypass_queue_pop_ack = '1')  and (bypass_queue_pop_data(0) = '0'));
	forward_zero_bypass_response <=
			((bypass_queue_pop_ack = '1')  and (bypass_queue_pop_data(0) = '1'));

	forward_bypass_to_fast <= 
			(forward_bypass_response or forward_zero_bypass_response) and 
								(bypass_queue_pop_data(2) = '1');
	forward_bypass_to_slow <= 
			(forward_bypass_response or forward_zero_bypass_response)  and 
					(bypass_queue_pop_data(2) = '0') and
								(bypass_queue_pop_data(1) = '1');

	-- pop when cpu, be are both ready.
	bypass_queue_pop_req <= '1' when 
		((forward_bypass_to_fast and cpu_fast_ready_for_bypass_response) or
			(forward_bypass_to_slow and cpu_slow_ready_for_bypass_response)) and 
						(forward_zero_bypass_response or be_response_ready)   
								else '0';

	be_read <= (bypass_queue_pop_req = '1')  and (bypass_queue_pop_ack = '1')  and forward_bypass_response;
        write_to_cpu_fast <= (bypass_queue_pop_req = '1') and (bypass_queue_pop_ack = '1') and 
										forward_bypass_to_fast;
        write_to_cpu_slow <= (bypass_queue_pop_req = '1') and (bypass_queue_pop_ack = '1') and 
										forward_bypass_to_slow;

	data_to_cpu <= be_dword when forward_bypass_response  else ZERO_64;
        response_to_cpu <= MAE8 & data_to_cpu;

end DcacheBypassController_arch;
library ieee;
use ieee.std_logic_1164.all;

library std;
use std.standard.all;

library AjitCustom;
use AjitCustom.AjitCustomComponents.all;

entity DcacheFrontendDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    NOBLOCK_CPU_to_DCACHE_command_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_command_pipe_read_data : in   std_logic_vector(142 downto 0);
    NOBLOCK_CPU_to_DCACHE_reset_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_reset_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_reset_pipe_read_data : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_data : in   std_logic_vector(120 downto 0);
    noblock_dcache_backend_to_frontend_command_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_dcache_backend_to_frontend_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_dcache_backend_to_frontend_command_pipe_read_data : in   std_logic_vector(83 downto 0);
    -----------------------------------------------------------------------------------------------
    NOBLOCK_DCACHE_TO_CPU_IU_BYPASS_pipe_write_req: out std_logic_vector(0 downto 0);
    NOBLOCK_DCACHE_TO_CPU_IU_BYPASS_pipe_write_ack: in std_logic_vector(0 downto 0);
    NOBLOCK_DCACHE_TO_CPU_IU_BYPASS_pipe_write_data: out std_logic_vector(92 downto 0);
    -----------------------------------------------------------------------------------------------
    NOBLOCK_DCACHE_TO_CPU_FU_BYPASS_pipe_write_req:  out std_logic_vector(0 downto 0);
    NOBLOCK_DCACHE_TO_CPU_FU_BYPASS_pipe_write_ack:  in std_logic_vector(0 downto 0);
    NOBLOCK_DCACHE_TO_CPU_FU_BYPASS_pipe_write_data: out std_logic_vector(92 downto 0);
    -----------------------------------------------------------------------------------------------
    DCACHE_to_CPU_reset_ack_pipe_write_req : out  std_logic_vector(0 downto 0);
    DCACHE_to_CPU_reset_ack_pipe_write_ack : in   std_logic_vector(0 downto 0);
    DCACHE_to_CPU_reset_ack_pipe_write_data : out  std_logic_vector(0 downto 0);
    DCACHE_to_CPU_response_pipe_write_req : out  std_logic_vector(0 downto 0);
    DCACHE_to_CPU_response_pipe_write_ack : in   std_logic_vector(0 downto 0);
    DCACHE_to_CPU_response_pipe_write_data : out  std_logic_vector(71 downto 0);
    DCACHE_to_CPU_slow_response_pipe_write_req : out  std_logic_vector(0 downto 0);
    DCACHE_to_CPU_slow_response_pipe_write_ack : in   std_logic_vector(0 downto 0);
    DCACHE_to_CPU_slow_response_pipe_write_data : out  std_logic_vector(71 downto 0);
    MMU_TO_DCACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_req: out std_logic_vector(0 downto 0);
    MMU_TO_DCACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_ack: in std_logic_vector(0 downto 0);
    MMU_TO_DCACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_data: in std_logic_vector(26 downto 0);
    NOBLOCK_MMU_TO_DCACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_req: out std_logic_vector(0 downto 0);
    NOBLOCK_MMU_TO_DCACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_ack: in std_logic_vector(0 downto 0);
    NOBLOCK_MMU_TO_DCACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_data: in std_logic_vector(26 downto 0);
    dcache_frontend_to_backend_pipe_write_req : out  std_logic_vector(0 downto 0);
    dcache_frontend_to_backend_pipe_write_ack : in   std_logic_vector(0 downto 0);
    dcache_frontend_to_backend_pipe_write_data : out  std_logic_vector(119 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity DcacheFrontendDaemon;
architecture UseStall of DcacheFrontendDaemon is -- 
	signal CACHE_STALL_ENABLE: std_logic_vector(0 downto 0);
    	signal NOBLOCK_INVALIDATE_SLOT_RETURN_pipe_read_req : std_logic_vector(0 downto 0);
    	signal NOBLOCK_INVALIDATE_SLOT_RETURN_pipe_read_ack : std_logic_vector(0 downto 0);
    	signal NOBLOCK_INVALIDATE_SLOT_RETURN_pipe_read_data: std_logic_vector(0 downto 0);
begin
    NOBLOCK_INVALIDATE_SLOT_RETURN_pipe_read_ack(0) <= '0';
    NOBLOCK_INVALIDATE_SLOT_RETURN_pipe_read_data   <= (others => '0');
    CACHE_STALL_ENABLE(0)  <= '0';

    dcache_frontend_with_stall:
		DcacheFrontendWithStallDaemon
			generic map (tag_length => tag_length)
			port map (
    				NOBLOCK_CPU_to_DCACHE_command_pipe_read_req,
    				NOBLOCK_CPU_to_DCACHE_command_pipe_read_ack,
    				NOBLOCK_CPU_to_DCACHE_command_pipe_read_data,
    				NOBLOCK_CPU_to_DCACHE_reset_pipe_read_req,
    				NOBLOCK_CPU_to_DCACHE_reset_pipe_read_ack,
    				NOBLOCK_CPU_to_DCACHE_reset_pipe_read_data,
    				NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_req,
    				NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_ack,
    				NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_data,
    				noblock_dcache_backend_to_frontend_command_pipe_read_req,
    				noblock_dcache_backend_to_frontend_command_pipe_read_ack,
    				noblock_dcache_backend_to_frontend_command_pipe_read_data,
    				-----------------------------------------------------------------------------------------------
    				NOBLOCK_DCACHE_TO_CPU_IU_BYPASS_pipe_write_req,
    				NOBLOCK_DCACHE_TO_CPU_IU_BYPASS_pipe_write_ack,
    				NOBLOCK_DCACHE_TO_CPU_IU_BYPASS_pipe_write_data,
    				-----------------------------------------------------------------------------------------------
    				NOBLOCK_DCACHE_TO_CPU_FU_BYPASS_pipe_write_req,
    				NOBLOCK_DCACHE_TO_CPU_FU_BYPASS_pipe_write_ack,
    				NOBLOCK_DCACHE_TO_CPU_FU_BYPASS_pipe_write_data,
    				-----------------------------------------------------------------------------------------------
    				DCACHE_to_CPU_reset_ack_pipe_write_req,
    				DCACHE_to_CPU_reset_ack_pipe_write_ack,
    				DCACHE_to_CPU_reset_ack_pipe_write_data,
    				DCACHE_to_CPU_response_pipe_write_req,
    				DCACHE_to_CPU_response_pipe_write_ack,
    				DCACHE_to_CPU_response_pipe_write_data,
    				DCACHE_to_CPU_slow_response_pipe_write_req,
    				DCACHE_to_CPU_slow_response_pipe_write_ack,
    				DCACHE_to_CPU_slow_response_pipe_write_data,
    				MMU_TO_DCACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_req,
    				MMU_TO_DCACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_ack,
    				MMU_TO_DCACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_data,
    				NOBLOCK_MMU_TO_DCACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_req,
    				NOBLOCK_MMU_TO_DCACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_ack,
    				NOBLOCK_MMU_TO_DCACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_data,
    				CACHE_STALL_ENABLE,
    				NOBLOCK_INVALIDATE_SLOT_RETURN_pipe_read_req,
    				NOBLOCK_INVALIDATE_SLOT_RETURN_pipe_read_ack,
    				NOBLOCK_INVALIDATE_SLOT_RETURN_pipe_read_data,
    				dcache_frontend_to_backend_pipe_write_req,
    				dcache_frontend_to_backend_pipe_write_ack,
    				dcache_frontend_to_backend_pipe_write_data,
    				tag_in,
    				tag_out,
    				clk,
    				reset,
    				start_req,
    				start_ack,
    				fin_req,
    				fin_ack);

end UseStall;
-- VHDL global package produced by vc2vhdl from virtual circuit (vc) description 
--  Copyright: Madhav Desai
library ieee;
use ieee.std_logic_1164.all;
package dcache_global_package is -- 
  constant ASI_AJIT_BRIDGE_CONFIG : std_logic_vector(7 downto 0) := "00110000";
  constant ASI_BLOCK_COPY : std_logic_vector(7 downto 0) := "00010111";
  constant ASI_BLOCK_FILL : std_logic_vector(7 downto 0) := "00011111";
  constant ASI_CACHE_DATA_I : std_logic_vector(7 downto 0) := "00001101";
  constant ASI_CACHE_DATA_I_D : std_logic_vector(7 downto 0) := "00001111";
  constant ASI_CACHE_TAG_I : std_logic_vector(7 downto 0) := "00001100";
  constant ASI_CACHE_TAG_I_D : std_logic_vector(7 downto 0) := "00001110";
  constant ASI_FLUSH_I_CONTEXT : std_logic_vector(7 downto 0) := "00011011";
  constant ASI_FLUSH_I_D_CONTEXT : std_logic_vector(7 downto 0) := "00010011";
  constant ASI_FLUSH_I_D_PAGE : std_logic_vector(7 downto 0) := "00010000";
  constant ASI_FLUSH_I_D_REGION : std_logic_vector(7 downto 0) := "00010010";
  constant ASI_FLUSH_I_D_SEGMENT : std_logic_vector(7 downto 0) := "00010001";
  constant ASI_FLUSH_I_D_USER : std_logic_vector(7 downto 0) := "00010100";
  constant ASI_FLUSH_I_PAGE : std_logic_vector(7 downto 0) := "00011000";
  constant ASI_FLUSH_I_REGION : std_logic_vector(7 downto 0) := "00011010";
  constant ASI_FLUSH_I_SEGMENT : std_logic_vector(7 downto 0) := "00011001";
  constant ASI_FLUSH_I_USER : std_logic_vector(7 downto 0) := "00011100";
  constant ASI_MMU_DIAGNOSTIC_I : std_logic_vector(7 downto 0) := "00000101";
  constant ASI_MMU_DIAGNOSTIC_IO : std_logic_vector(7 downto 0) := "00000111";
  constant ASI_MMU_DIAGNOSTIC_I_D : std_logic_vector(7 downto 0) := "00000110";
  constant ASI_MMU_FLUSH_PROBE : std_logic_vector(7 downto 0) := "00000011";
  constant ASI_MMU_REGISTER : std_logic_vector(7 downto 0) := "00000100";
  constant ASI_SUPERVISOR_DATA : std_logic_vector(7 downto 0) := "00001011";
  constant ASI_SUPERVISOR_INSTRUCTION : std_logic_vector(7 downto 0) := "00001001";
  constant ASI_USER_DATA : std_logic_vector(7 downto 0) := "00001010";
  constant ASI_USER_INSTRUCTION : std_logic_vector(7 downto 0) := "00001000";
  
  -- corrected!
  constant CACHE_ARRAY_READ_DWORD : std_logic_vector(2 downto 0) := "001";
  constant CACHE_ARRAY_WRITE_DWORD : std_logic_vector(2 downto 0) := "010";
  constant CACHE_ARRAY_NOP : std_logic_vector(2 downto 0) := "011";

  -- corrected
  constant CACHE_TAG_CLEAR_ALL : std_logic_vector(2 downto 0) := "100";
  constant CACHE_TAG_CLEAR_LINE : std_logic_vector(2 downto 0) := "011";
  constant CACHE_TAG_INSERT : std_logic_vector(2 downto 0) := "010";
  constant CACHE_TAG_LOOKUP : std_logic_vector(2 downto 0) := "001";
  constant CACHE_TAG_NOP : std_logic_vector(2 downto 0) := "101";

  constant DCACHE_BE_FLUSH_ALL : std_logic_vector(7 downto 0) := "00001100";
  constant DCACHE_BE_FLUSH_LINE : std_logic_vector(7 downto 0) := "00001011";
  constant DCACHE_BE_MMU_READ_LINE : std_logic_vector(7 downto 0) := "00000011";
  constant DCACHE_BE_NOCACHE_READ_MMU_DWORD : std_logic_vector(7 downto 0) := "00010000";
  constant DCACHE_BE_NOCACHE_WRITE_MMU_DWORD : std_logic_vector(7 downto 0) := "00001111";
  constant DCACHE_BE_NOP : std_logic_vector(7 downto 0) := "00001110";
  constant DCACHE_BE_READ_DWORD : std_logic_vector(7 downto 0) := "00000001";
  constant DCACHE_BE_READ_MMU_BYPASS_DWORD : std_logic_vector(7 downto 0) := "00000110";
  constant DCACHE_BE_READ_MMU_CTRL_REGISTER : std_logic_vector(7 downto 0) := "00001000";
  constant DCACHE_BE_SEND_ERROR_RESPONSE : std_logic_vector(7 downto 0) := "00010010";
  constant DCACHE_BE_SEND_MAE_RESPONSE : std_logic_vector(7 downto 0) := "00001010";
  constant DCACHE_BE_SEND_ZERO_RESPONSE : std_logic_vector(7 downto 0) := "00001001";
  constant DCACHE_BE_UNLOCK_TAGS : std_logic_vector(7 downto 0) := "00001101";
  constant DCACHE_BE_UPDATE_LAST_LINE : std_logic_vector(7 downto 0) := "00010001";
  constant DCACHE_BE_WRITE_DWORD : std_logic_vector(7 downto 0) := "00000010";
  constant DCACHE_BE_WRITE_MISS : std_logic_vector(7 downto 0) := "00000100";
  constant DCACHE_BE_WRITE_MMU_BYPASS_DWORD : std_logic_vector(7 downto 0) := "00000101";
  constant DCACHE_BE_WRITE_MMU_CTRL_REGISTER : std_logic_vector(7 downto 0) := "00000111";
  constant DEBUG_MODE_MASK : std_logic_vector(7 downto 0) := "00000010";
  constant FOUR_3 : std_logic_vector(2 downto 0) := "100";
  constant GDB_DBG_CONNECT : std_logic_vector(7 downto 0) := "00001110";
  constant GDB_DBG_CONTINUE : std_logic_vector(7 downto 0) := "00010000";
  constant GDB_DBG_DETACH : std_logic_vector(7 downto 0) := "00001111";
  constant GDB_DBG_KILL : std_logic_vector(7 downto 0) := "00010011";
  constant GDB_DBG_READ_CONTROL_REG : std_logic_vector(7 downto 0) := "00001101";
  constant GDB_DBG_READ_CPUNIT_REG : std_logic_vector(7 downto 0) := "00010001";
  constant GDB_DBG_READ_FPUNIT_REG : std_logic_vector(7 downto 0) := "00000011";
  constant GDB_DBG_READ_IUNIT_REG : std_logic_vector(7 downto 0) := "00000001";
  constant GDB_DBG_READ_MEM : std_logic_vector(7 downto 0) := "00000110";
  constant GDB_DBG_REMOVE_BREAK_POINT : std_logic_vector(7 downto 0) := "00001001";
  constant GDB_DBG_REMOVE_WATCH_POINT : std_logic_vector(7 downto 0) := "00001011";
  constant GDB_DBG_SET_BREAK_POINT : std_logic_vector(7 downto 0) := "00001000";
  constant GDB_DBG_SET_WATCH_POINT : std_logic_vector(7 downto 0) := "00001010";
  constant GDB_DBG_WRITE_CONTROL_REG : std_logic_vector(7 downto 0) := "00010100";
  constant GDB_DBG_WRITE_CPUNIT_REG : std_logic_vector(7 downto 0) := "00010010";
  constant GDB_DBG_WRITE_FPUNIT_REG : std_logic_vector(7 downto 0) := "00000100";
  constant GDB_DBG_WRITE_IUNIT_REG : std_logic_vector(7 downto 0) := "00000010";
  constant GDB_DBG_WRITE_MEM : std_logic_vector(7 downto 0) := "00000111";
  constant HARD_RESET_MASK : std_logic_vector(7 downto 0) := "00000001";
  constant KILL_STREAM_MASK : std_logic_vector(7 downto 0) := "10000000";
  constant KILL_THREAD_MASK : std_logic_vector(7 downto 0) := "10000000";
  constant LOGGER_ACTIVE_MASK : std_logic_vector(7 downto 0) := "00001000";
  constant MMU_PASS_THROUGH_HLIMIT : std_logic_vector(7 downto 0) := "00101111";
  constant MMU_PASS_THROUGH_LLIMIT : std_logic_vector(7 downto 0) := "00100000";
  constant MMU_READ_DWORD : std_logic_vector(7 downto 0) := "00000010";
  constant MMU_READ_LINE : std_logic_vector(7 downto 0) := "00000011";
  constant MMU_WRITE_DWORD : std_logic_vector(7 downto 0) := "00000001";
  constant MMU_WRITE_DWORD_NO_RESPONSE : std_logic_vector(7 downto 0) := "00000101";
  constant MMU_WRITE_FSR : std_logic_vector(7 downto 0) := "00000100";
  constant NEW_STREAM_MASK : std_logic_vector(7 downto 0) := "10000000";
  constant NEW_THREAD_MASK : std_logic_vector(7 downto 0) := "10000000";
  constant NPC_RESET_VALUE : std_logic_vector(31 downto 0) := "00000000000000000000000000000100";
  constant NWINDOWS : std_logic_vector(31 downto 0) := "00000000000000000000000000001000";
  constant NWINDOWS_MOD_MASK_32 : std_logic_vector(31 downto 0) := "00000000000000000000000000000111";
  constant NWINDOWS_MOD_MASK_5 : std_logic_vector(4 downto 0) := "00111";
  constant NWINDOWSx16 : std_logic_vector(31 downto 0) := "00000000000000000000000010000000";
  constant NWINDOWSx16_MOD_MASK_32 : std_logic_vector(31 downto 0) := "00000000000000000000000001111111";
  constant NWINDOWSx2 : std_logic_vector(31 downto 0) := "00000000000000000000000000010000";
  constant ONE_1 : std_logic_vector(0 downto 0) := "1";
  constant ONE_10 : std_logic_vector(9 downto 0) := "0000000001";
  constant ONE_11 : std_logic_vector(10 downto 0) := "00000000001";
  constant ONE_12 : std_logic_vector(11 downto 0) := "000000000001";
  constant ONE_128 : std_logic_vector(127 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001";
  constant ONE_13 : std_logic_vector(12 downto 0) := "0000000000001";
  constant ONE_14 : std_logic_vector(13 downto 0) := "00000000000001";
  constant ONE_16 : std_logic_vector(15 downto 0) := "0000000000000001";
  constant ONE_17 : std_logic_vector(16 downto 0) := "00000000000000001";
  constant ONE_18 : std_logic_vector(17 downto 0) := "000000000000000001";
  constant ONE_19 : std_logic_vector(18 downto 0) := "0000000000000000001";
  constant ONE_2 : std_logic_vector(1 downto 0) := "01";
  constant ONE_23 : std_logic_vector(22 downto 0) := "00000000000000000000001";
  constant ONE_24 : std_logic_vector(23 downto 0) := "000000000000000000000001";
  constant ONE_25 : std_logic_vector(24 downto 0) := "0000000000000000000000001";
  constant ONE_256 : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000001";
  constant ONE_29 : std_logic_vector(28 downto 0) := "00000000000000000000000000001";
  constant ONE_3 : std_logic_vector(2 downto 0) := "001";
  constant ONE_31 : std_logic_vector(30 downto 0) := "0000000000000000000000000000001";
  constant ONE_32 : std_logic_vector(31 downto 0) := "00000000000000000000000000000001";
  constant ONE_36 : std_logic_vector(35 downto 0) := "000000000000000000000000000000000001";
  constant ONE_4 : std_logic_vector(3 downto 0) := "0001";
  constant ONE_48 : std_logic_vector(47 downto 0) := "000000000000000000000000000000000000000000000001";
  constant ONE_5 : std_logic_vector(4 downto 0) := "00001";
  constant ONE_6 : std_logic_vector(5 downto 0) := "000001";
  constant ONE_64 : std_logic_vector(63 downto 0) := "0000000000000000000000000000000000000000000000000000000000000001";
  constant ONE_7 : std_logic_vector(6 downto 0) := "0000001";
  constant ONE_8 : std_logic_vector(7 downto 0) := "00000001";
  constant ONE_9 : std_logic_vector(8 downto 0) := "000000001";
  constant PC_RESET_VALUE : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
  constant PROCESSOR_ERROR_MODE : std_logic_vector(1 downto 0) := "11";
  constant PROCESSOR_EXECUTE_MODE : std_logic_vector(1 downto 0) := "10";
  constant PROCESSOR_RESET_MODE : std_logic_vector(1 downto 0) := "01";
  constant PROCESSOR_UNDEFINED_MODE : std_logic_vector(1 downto 0) := "00";
  constant PSR_RESET_VALUE : std_logic_vector(31 downto 0) := "00000000000000000001000011000000";
  constant REQUEST_TYPE_BRIDGE_CONFIG_READ : std_logic_vector(3 downto 0) := "1001";
  constant REQUEST_TYPE_BRIDGE_CONFIG_WRITE : std_logic_vector(3 downto 0) := "1000";
  constant REQUEST_TYPE_CCU_CACHE_READ : std_logic_vector(3 downto 0) := "0101";
  constant REQUEST_TYPE_CCU_CACHE_WRITE : std_logic_vector(3 downto 0) := "0110";
  constant REQUEST_TYPE_IFETCH : std_logic_vector(3 downto 0) := "0000";
  constant REQUEST_TYPE_NOP : std_logic_vector(3 downto 0) := "0111";
  constant REQUEST_TYPE_READ : std_logic_vector(3 downto 0) := "0001";
  constant REQUEST_TYPE_STBAR : std_logic_vector(3 downto 0) := "0011";
  constant REQUEST_TYPE_WRFSRFAR : std_logic_vector(3 downto 0) := "0100";
  constant REQUEST_TYPE_WRITE : std_logic_vector(3 downto 0) := "0010";
  constant SINGLE_STEP_MASK : std_logic_vector(7 downto 0) := "00000100";
  constant THREE_2 : std_logic_vector(1 downto 0) := "11";
  constant THREE_3 : std_logic_vector(2 downto 0) := "011";
  constant TRACE_ON : std_logic_vector(0 downto 0) := "1";
  constant TWO_2 : std_logic_vector(1 downto 0) := "10";
  constant TWO_3 : std_logic_vector(2 downto 0) := "010";
  constant WIM_MASK : std_logic_vector(31 downto 0) := "00000000000000000000000011111111";
  constant ZADDR : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
  constant ZERO_1 : std_logic_vector(0 downto 0) := "0";
  constant ZERO_10 : std_logic_vector(9 downto 0) := "0000000000";
  constant ZERO_11 : std_logic_vector(10 downto 0) := "00000000000";
  constant ZERO_12 : std_logic_vector(11 downto 0) := "000000000000";
  constant ZERO_128 : std_logic_vector(127 downto 0) := "00000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant ZERO_13 : std_logic_vector(12 downto 0) := "0000000000000";
  constant ZERO_14 : std_logic_vector(13 downto 0) := "00000000000000";
  constant ZERO_16 : std_logic_vector(15 downto 0) := "0000000000000000";
  constant ZERO_17 : std_logic_vector(16 downto 0) := "00000000000000000";
  constant ZERO_18 : std_logic_vector(17 downto 0) := "000000000000000000";
  constant ZERO_19 : std_logic_vector(18 downto 0) := "0000000000000000000";
  constant ZERO_2 : std_logic_vector(1 downto 0) := "00";
  constant ZERO_23 : std_logic_vector(22 downto 0) := "00000000000000000000000";
  constant ZERO_24 : std_logic_vector(23 downto 0) := "000000000000000000000000";
  constant ZERO_25 : std_logic_vector(24 downto 0) := "0000000000000000000000000";
  constant ZERO_256 : std_logic_vector(255 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
  constant ZERO_29 : std_logic_vector(28 downto 0) := "00000000000000000000000000000";
  constant ZERO_3 : std_logic_vector(2 downto 0) := "000";
  constant ZERO_31 : std_logic_vector(30 downto 0) := "0000000000000000000000000000000";
  constant ZERO_32 : std_logic_vector(31 downto 0) := "00000000000000000000000000000000";
  constant ZERO_36 : std_logic_vector(35 downto 0) := "000000000000000000000000000000000000";
  constant ZERO_4 : std_logic_vector(3 downto 0) := "0000";
  constant ZERO_48 : std_logic_vector(47 downto 0) := "000000000000000000000000000000000000000000000000";
  constant ZERO_5 : std_logic_vector(4 downto 0) := "00000";
  constant ZERO_6 : std_logic_vector(5 downto 0) := "000000";
  constant ZERO_64 : std_logic_vector(63 downto 0) := "0000000000000000000000000000000000000000000000000000000000000000";
  constant ZERO_7 : std_logic_vector(6 downto 0) := "0000000";
  constant ZERO_8 : std_logic_vector(7 downto 0) := "00000000";
  constant ZERO_9 : std_logic_vector(8 downto 0) := "000000000";

  component parse_from_backend_Volatile is -- 
   port ( -- 
    from_be : in  std_logic_vector(83 downto 0);
    be_valid : out  std_logic_vector(0 downto 0);
    be_counter : out  std_logic_vector(2 downto 0);
    be_tag_command : out  std_logic_vector(2 downto 0);
    be_array_command : out  std_logic_vector(2 downto 0);
    be_dword_id : out  std_logic_vector(2 downto 0);
    be_last_dword : out  std_logic_vector(0 downto 0);
    be_acc : out  std_logic_vector(2 downto 0);
    be_cacheable : out  std_logic_vector(0 downto 0);
    be_mae : out  std_logic_vector(0 downto 0);
    be_access_error : out  std_logic_vector(0 downto 0);
    be_dword : out  std_logic_vector(63 downto 0)-- 
  );
  -- 
  end component parse_from_backend_Volatile;

  component merge_and_decode_from_cpu_VVD is -- 
  port ( -- 
    from_cpu_fast : in  std_logic_vector(120 downto 0);
    from_cpu_slow : in  std_logic_vector(120 downto 0);
    is_thread_head : out  std_logic_vector(0 downto 0);
    lock_bus : out  std_logic_vector(0 downto 0);
    cpu_valid : out  std_logic_vector(0 downto 0);
    cpu_valid_fast : out  std_logic_vector(0 downto 0);
    cpu_valid_slow : out  std_logic_vector(0 downto 0);
    cpu_req_type : out  std_logic_vector(7 downto 0);
    cpu_asi : out  std_logic_vector(7 downto 0);
    cpu_byte_mask : out  std_logic_vector(7 downto 0);
    cpu_addr : out  std_logic_vector(31 downto 0);
    cpu_write_data : out  std_logic_vector(63 downto 0);
    is_flush_asi : out  std_logic_vector(0 downto 0);
    is_mmu_ctrl_reg_write : out  std_logic_vector(0 downto 0);
    flush_line_only : out  std_logic_vector(0 downto 0);
    is_supervisor_asi : out  std_logic_vector(0 downto 0);
    is_mmu_access_asi : out  std_logic_vector(0 downto 0);
    dcache_needs_to_be_flushed : out  std_logic_vector(0 downto 0);
    is_memory_read : out  std_logic_vector(0 downto 0);
    is_memory_write : out  std_logic_vector(0 downto 0);
    is_mmu_fsr_write : out  std_logic_vector(0 downto 0);
    is_stbar : out  std_logic_vector(0 downto 0);
    is_ccu_request : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
  end component merge_and_decode_from_cpu_VVD;
  component offsetInLine_VVD is -- 
  port ( -- 
    addr : in  std_logic_vector(31 downto 0);
    ret_val : out  std_logic_vector(3 downto 0)-- 
  );
  -- 
  end component offsetInLine_VVD;
  component identify_cpu_actions_VVD is -- 
  port ( -- 
    exec_cpu : in  std_logic_vector(0 downto 0);
    next_dcache_trapped : in  std_logic_vector(0 downto 0);
    is_ccu_request : in  std_logic_vector(0 downto 0);
    is_a_hit : in  std_logic_vector(0 downto 0);
    skip_tag_lookup : in  std_logic_vector(0 downto 0);
    is_memory_write : in  std_logic_vector(0 downto 0);
    is_memory_read : in  std_logic_vector(0 downto 0);
    is_flush_asi : in  std_logic_vector(0 downto 0);
    is_stbar : in  std_logic_vector(0 downto 0);
    is_mmu_access_asi : in  std_logic_vector(0 downto 0);
    is_mmu_fsr_write : in  std_logic_vector(0 downto 0);
    write_dword_hit : out  std_logic_vector(0 downto 0);
    write_dword_miss : out  std_logic_vector(0 downto 0);
    read_dword_hit : out  std_logic_vector(0 downto 0);
    read_dword_miss : out  std_logic_vector(0 downto 0);
    finished_flush_or_nop : out  std_logic_vector(0 downto 0);
    write_to_mmu_or_bypass : out  std_logic_vector(0 downto 0);
    read_from_mmu_or_bypass : out  std_logic_vector(0 downto 0);
    write_to_mmu_fsr : out  std_logic_vector(0 downto 0);
    send_to_be : out  std_logic_vector(0 downto 0);
    no_response_from_be : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
  end component identify_cpu_actions_VVD;
  component dcacheNeedsToBeFlushed_VVD is -- 
  port ( -- 
    asi : in  std_logic_vector(7 downto 0);
    req_type : in  std_logic_vector(3 downto 0);
    is_flush_asi : out  std_logic_vector(0 downto 0);
    is_mmu_ctrl_reg_write : out  std_logic_vector(0 downto 0);
    flush_line_only : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
  end component dcacheNeedsToBeFlushed_VVD;
  component isDcacheFlushAsi_VVD is -- 
  port ( -- 
    asi : in  std_logic_vector(7 downto 0);
    ret_val : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
  end component isDcacheFlushAsi_VVD;
  component isMmuAccessAsi_VVD is -- 
  port ( -- 
    asi : in  std_logic_vector(7 downto 0);
    ret_val : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
  end component isMmuAccessAsi_VVD;

  component isSupervisorAsi_VVD is -- 
  port ( -- 
    asi : in  std_logic_vector(7 downto 0);
    ret_val : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
  end component isSupervisorAsi_VVD;

end package dcache_global_package;

library std;
use std.standard.all;

library ieee;
use ieee.std_logic_1164.all;

library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;

library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;

library AjitCustom;
use AjitCustom.AjitGlobalConfigurationPackage.all;
use AjitCustom.AjitCoreConfigurationPackage.all;
use AjitCustom.AjitCustomComponents.all;
use AjitCustom.dcache_global_package.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

entity DcacheFrontendWithStallCoreDaemon is -- 
  generic (tag_length : integer := 1); 
  port ( -- 
    NOBLOCK_CPU_to_DCACHE_command_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_command_pipe_read_data : in   std_logic_vector(142 downto 0);
    NOBLOCK_CPU_to_DCACHE_reset_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_reset_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_reset_pipe_read_data : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_data : in   std_logic_vector(120 downto 0);
    noblock_dcache_backend_to_frontend_command_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_dcache_backend_to_frontend_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_dcache_backend_to_frontend_command_pipe_read_data : in   std_logic_vector(83 downto 0);
    -----------------------------------------------------------------------------------------------
    NOBLOCK_DCACHE_TO_CPU_IU_BYPASS_pipe_write_req: out std_logic_vector(0 downto 0);
    NOBLOCK_DCACHE_TO_CPU_IU_BYPASS_pipe_write_ack: in std_logic_vector(0 downto 0);
    NOBLOCK_DCACHE_TO_CPU_IU_BYPASS_pipe_write_data: out std_logic_vector(92 downto 0);
    -----------------------------------------------------------------------------------------------
    NOBLOCK_DCACHE_TO_CPU_FU_BYPASS_pipe_write_req:  out std_logic_vector(0 downto 0);
    NOBLOCK_DCACHE_TO_CPU_FU_BYPASS_pipe_write_ack:  in std_logic_vector(0 downto 0);
    NOBLOCK_DCACHE_TO_CPU_FU_BYPASS_pipe_write_data: out std_logic_vector(92 downto 0);
    -----------------------------------------------------------------------------------------------
    DCACHE_to_CPU_reset_ack_pipe_write_req : out  std_logic_vector(0 downto 0);
    DCACHE_to_CPU_reset_ack_pipe_write_ack : in   std_logic_vector(0 downto 0);
    DCACHE_to_CPU_reset_ack_pipe_write_data : out  std_logic_vector(0 downto 0);
    DCACHE_to_CPU_response_pipe_write_req : out  std_logic_vector(0 downto 0);
    DCACHE_to_CPU_response_pipe_write_ack : in   std_logic_vector(0 downto 0);
    DCACHE_to_CPU_response_pipe_write_data : out  std_logic_vector(71 downto 0);
    DCACHE_to_CPU_slow_response_pipe_write_req : out  std_logic_vector(0 downto 0);
    DCACHE_to_CPU_slow_response_pipe_write_ack : in   std_logic_vector(0 downto 0);
    DCACHE_to_CPU_slow_response_pipe_write_data : out  std_logic_vector(71 downto 0);
    MMU_TO_DCACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_req: out std_logic_vector(0 downto 0);
    MMU_TO_DCACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_ack: in std_logic_vector(0 downto 0);
    MMU_TO_DCACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_data: in std_logic_vector(26 downto 0);
    NOBLOCK_MMU_TO_DCACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_req: out std_logic_vector(0 downto 0);
    NOBLOCK_MMU_TO_DCACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_ack: in std_logic_vector(0 downto 0);
    NOBLOCK_MMU_TO_DCACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_data: in std_logic_vector(26 downto 0);
    CACHE_STALL_ENABLE: in std_logic_vector(0 downto 0);
    NOBLOCK_INVALIDATE_SLOT_RETURN_pipe_read_req : out std_logic_vector(0 downto 0);
    NOBLOCK_INVALIDATE_SLOT_RETURN_pipe_read_ack : in std_logic_vector(0 downto 0);
    NOBLOCK_INVALIDATE_SLOT_RETURN_pipe_read_data: in std_logic_vector(0 downto 0);
    dcache_frontend_to_backend_pipe_write_req : out  std_logic_vector(0 downto 0);
    dcache_frontend_to_backend_pipe_write_ack : in   std_logic_vector(0 downto 0);
    dcache_frontend_to_backend_pipe_write_data : out  std_logic_vector(119 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity DcacheFrontendWithStallCoreDaemon;
architecture DcacheFrontendCoreDaemon_arch of DcacheFrontendWithStallCoreDaemon is -- 
	Type DcacheState is (IDLE,
					CHECK_HIT_OR_MISS, SYN_INVALIDATE, SEND_WAIT_ON_CPU, 
						SEND_WAIT_ON_BE, RECV_WAIT_ON_BE_FIRST_DWORD,
								RECV_WAIT_ON_BE_REMAINING_DWORDS);
	function StateToString(x:DcacheState) return string is
             variable ret_var: string (1 to 9);
        begin
            ret_var := "IdleState";
            if(x = CHECK_HIT_OR_MISS) then
               ret_var := "ChekHitSt";
            elsif(x = SEND_WAIT_ON_CPU) then
               ret_var := "SndWaitCp";
            elsif(x = SEND_WAIT_ON_BE) then
               ret_var := "SndWaitBe";
            elsif(x = RECV_WAIT_ON_BE_FIRST_DWORD) then
               ret_var := "RxFirstBe";
            elsif(x = RECV_WAIT_ON_BE_REMAINING_DWORDS) then
               ret_var := "RxRest_Be";
            elsif(x = SYN_INVALIDATE) then
               ret_var := "SynInvald";
	    end if;
	    return(ret_var);
        end StateToString;

	signal dcache_state : DcacheState;
	signal cpu_fast_command_valid : boolean;
	signal cpu_slow_command_valid : boolean;
	-------------------------------------------------------------------------------------------
	-- predicates/inputs
	-------------------------------------------------------------------------------------------
	signal  is_bypass_asi, bypass_case, normal_case: boolean;

	signal  cpu_command_available  : boolean;
	signal  cpu_bypass_command_available  : boolean;
	signal  cpu_bypass_command_accept  : boolean;

	signal  cpu_reset	       : boolean;

	signal  be_is_needed	       : boolean;
	signal  expect_be_response     : boolean;
	signal  expect_be_response_reg : boolean;
	signal  be_has_completed       : boolean;
	signal  be_has_exception       : boolean;

	signal  be_ready_for_command   	    : boolean;
	signal  be_response_available  	    : boolean;
	signal  be_response_can_be_applied  : boolean;
	signal  first_be_response_can_be_applied  : boolean;

	signal  cpu_ready_for_response : boolean;

	signal  cpu_slow_ready_for_bypass_response : boolean;
	signal  cpu_fast_ready_for_bypass_response : boolean;

	signal  write_bypass_to_cpu_slow: boolean;
	signal  write_bypass_to_cpu_fast: boolean;

	signal skip_tag_lookup, do_tag_lookup: boolean;
	signal skip_tag_lookup_slv, skip_tag_lookup_slv_reg: std_logic_vector(0 downto 0);

	signal exec_be: boolean;
	signal exec_tag_access_cpu: boolean;
	-------------------------------------------------------------------------------------------
	-- actions/outputs
	-------------------------------------------------------------------------------------------
	signal latch_cpu_commands  : boolean;
	signal accept_cpu_commands  : boolean;
	signal clear_cpu_commands  : boolean;
	signal latch_tag_results   : boolean;
	signal latch_be_info	   : boolean;
	signal latch_to_cpu	   : boolean;
	signal latch_to_be	   : boolean;
	signal latch_expect_be_response	   : boolean;
	signal accept_be_response  : boolean;
	signal accept_be_bypass_response: boolean;
	signal bypass_response_pending: boolean;	
	signal write_to_be	   : boolean;
	signal write_to_be_from_bypass : boolean;
	signal write_to_cpu	   : boolean;
	signal untrap_dcache	   : boolean;
	signal trap_dcache	   : boolean;
	signal do_write_to_arrays_if_applicable : boolean;
	

	signal latch_to_cpu_registered	   : boolean;
	signal latch_to_be_registered	   : boolean;
	-------------------------------------------------------------------------------------------
	-- signals, registers
	-------------------------------------------------------------------------------------------
	signal DCACHE_TRAPPED: boolean;

	-- is the cpu thread trapped.. for the two threads..
	signal dcache_trapped_vector: std_logic_vector(0 to 1);

	signal from_cpu_fast, from_cpu_slow, cpu_slow_command, 
					cpu_fast_command : std_logic_vector(120 downto 0);

	signal fast_command_bypass_control_info: std_logic_vector(21 downto 0);
	signal fast_command_bypass_control_info_reg: std_logic_vector(21 downto 0);

	signal cpu_thread_id: std_logic_vector(1 downto 0);
	signal cpu_thread_id_registered: std_logic_vector(1 downto 0);
	signal active_cpu_thread_id: std_logic_vector(1 downto 0);
	signal ACPU: integer range 0 to 1;

      
      	signal cpu_valid, cpu_valid_fast, cpu_valid_slow : std_logic_vector(0 downto 0);
	signal cpu_req_type, cpu_asi, cpu_byte_mask: std_logic_vector(7 downto 0);
	signal cpu_addr: std_logic_vector(31 downto 0);
	signal cpu_write_data: std_logic_vector(63 downto 0);
      	signal cpu_cache_line : std_logic_vector(511 downto 0);
	signal cpu_tag_command: std_logic_vector(2 downto 0);

      	signal cpu_valid_reg, cpu_valid_fast_reg, cpu_valid_slow_reg : std_logic_vector(0 downto 0);
	signal cpu_req_type_reg, cpu_asi_reg, cpu_byte_mask_reg: std_logic_vector(7 downto 0);
	signal cpu_addr_reg: std_logic_vector(31 downto 0);
	signal cpu_write_data_reg: std_logic_vector(63 downto 0);

	signal is_thread_head, lock_bus: std_logic_vector(0 downto 0);
	signal is_flush_asi, is_mmu_ctrl_reg_write, flush_line_only,
			is_supervisor_asi,
			is_mmu_access_asi,
			dcache_needs_to_be_flushed,
			is_memory_read,
			is_memory_write,
			is_mmu_fsr_write,
			is_stbar,
			is_ccu_request : std_logic_vector(0 downto 0);

	signal access_is_read, access_is_ifetch: std_logic;

	signal lock_bus_reg: std_logic_vector(0 downto 0);
	signal is_flush_asi_reg, is_mmu_ctrl_reg_write_reg, flush_line_only_reg,
			is_supervisor_asi_reg,
			is_mmu_access_asi_reg,
			is_memory_read_reg,
			is_memory_write_reg,
			is_mmu_fsr_write_reg,
			is_stbar_reg,
			is_ccu_request_reg : std_logic_vector(0 downto 0);


	signal from_backend : std_logic_vector(83 downto 0);
	signal be_valid : std_logic_vector(0 downto 0);
      	signal be_acc, access_tags_acc : std_logic_vector(2 downto 0);
      	signal be_mae : std_logic_vector(0 downto 0);
      	signal be_access_error: std_logic_vector(0 downto 0);
      	signal be_tag_command : std_logic_vector(2 downto 0);
      	signal be_array_command : std_logic_vector(2 downto 0);
      	signal be_counter : std_logic_vector(2 downto 0);
      	signal be_dword_id : std_logic_vector(2 downto 0);
      	signal be_last_dword : std_logic_vector(0 downto 0);
      	signal be_cacheable : std_logic_vector(0 downto 0);
	
      	signal be_dword : std_logic_vector(63 downto 0);

	

    	signal is_hit: std_logic_vector(0 downto 0);
    	signal cpu_permissions_ok: std_logic_vector(0 downto 0);
    	signal dword_out : std_logic_vector(63 downto 0);

	signal mae_8_to_cpu: std_logic_vector (7 downto 0);
	signal data_to_cpu: std_logic_vector (63 downto 0);
	signal is_a_hit, is_a_hit_to_cpu, mae_to_cpu, access_error_to_cpu : std_logic_vector(0 downto 0);
	signal cpu_tag_lookup: boolean;

	
    	signal to_cpu, to_cpu_registered: std_logic_vector(71 downto 0);
    	signal bypass_response_to_cpu:  std_logic_vector(71 downto 0);
    	signal to_be, to_be_registered, to_be_from_bypass :  std_logic_vector(119 downto 0);

	signal access_byte_mask: std_logic_vector(7 downto 0); 

	constant LOG2_NUMBER_OF_BLOCKS: integer := LOG_DCACHE_SIZE_IN_BLOCKS;
        constant LOG2_BLOCK_SIZE_IN_BYTES: integer := 6;
        constant LOG2_DATA_WIDTH_IN_BYTES: integer := 3;

    	signal access_mae : std_logic;
    	signal access_S : std_logic;

	signal tags_arrays_trigger,  tags_arrays_done: std_logic;
	signal wait_on_tags_arrays: boolean;
	signal waiting_on_tags_arrays: boolean;

	signal arrays_fin_ack, arrays_start_ack: std_logic;
	signal tags_start_req, arrays_start_req, tags_start_ack, 
				tags_fin_req, arrays_fin_req, tags_fin_ack: std_logic;
	signal init_flag: std_logic;


	signal write_dword_hit, write_dword_miss,
			read_dword_hit, read_dword_miss,
			finished_flush_or_nop, write_to_mmu_or_bypass,
			read_from_mmu_or_bypass, 
			write_to_mmu_fsr: std_logic_vector(0 downto 0);	
	signal send_to_be, no_response_from_be, exec_cpu, 
			dcache_in_trapped_state, dcache_in_trapped_state_reg: std_logic_vector(0 downto 0);

	signal exec_cpu_reg: std_logic_vector(0 downto 0);
	signal send_cpu_reset_ack : boolean;
	signal accept_cpu_reset: boolean;

	constant byte_mask_ff : std_logic_vector(7 downto 0) := (others => '1');

	signal syn_inval_ready, coherence_inval_ready: boolean;
	signal syn_inval_accept, coherence_inval_accept: boolean;
	signal syn_inval_applicable, coherence_inval_applicable: boolean;

	signal tag_invalidate_apply: std_logic_vector(0 downto 0);
	signal tag_invalidate_line_address : std_logic_vector(25 downto 0);

	signal cpu_command_is_not_a_clear_or_flush: boolean;

	signal tags_arrays_request_state: std_logic;
	signal tags_arrays_result_ready:  boolean;


	-- Added: in the multi-thread case, we need to ensure that lock is maintained.
	--        We will prevent fast path from getting in to the dcache if the lock
	--        is held by the slow path.
	signal slow_request_wants_lock, slow_request_has_lock, slow_request_selected: boolean;

	-- added: register the cache stall.
	signal CACHE_STALL_ENABLE_REG: std_logic_vector(0 downto 0);
	signal starting_new_memory_write,  invalidate_slot_return, DCACHE_STALL: boolean;
	signal free_invalidate_slot_count : integer range 0 to NUMBER_OF_INVALIDATE_SLOTS_PER_CORE-2;


	signal is_pure_mem_access_asi, is_mem_access_asi, is_mem_access_asi_reg : boolean;

	-- These are moved to global scope since they are used
	-- in multiple blocks.
	signal nc_tlb_match_base, nc_tlb_match: std_logic;
	signal access_tag_command: std_logic_vector(2 downto 0);
	signal lookup_acc: std_logic_vector(2 downto 0);

-- see comment above..
--##decl_synopsys_sync_set_reset##

begin
	-- once started, never finish!
	start_ack <= '1';
	fin_ack <= '0'; 
	tag_out <= tag_in;

	-- why the &^(%* is this getting lost..
	process(clk)
        begin
		if(clk'event and clk='1') then
			assert false report "Dcache State is " & StateToString(dcache_state)
					severity note;
		end if;
        end process;

	cpu_valid <= cpu_valid_fast or cpu_valid_slow;
	exec_cpu <= cpu_valid;
	exec_cpu_reg <= cpu_valid_reg;

	-- register the cache stall to cut combi path.
	process(clk,reset)
	begin
		if(clk'event and clk ='1') then 
			if(reset = '1') then
				CACHE_STALL_ENABLE_REG(0) <= '0';
			else
				CACHE_STALL_ENABLE_REG(0) <= CACHE_STALL_ENABLE(0);
			end if;
		end if;
	end process;

	-- Stall logic...  need to reserve an invalidation queue slot before
	--  starting a write operation.
    	NOBLOCK_INVALIDATE_SLOT_RETURN_pipe_read_req(0) <= '1';
	invalidate_slot_return <=
    		(NOBLOCK_INVALIDATE_SLOT_RETURN_pipe_read_ack(0) = '1') and
    			(NOBLOCK_INVALIDATE_SLOT_RETURN_pipe_read_data(0) = '1');
	starting_new_memory_write <=
		is_mem_access_asi and
			((is_memory_write(0) = '1') and ((is_thread_head(0) = '1') or (not DCACHE_TRAPPED)) and 
				(latch_cpu_commands or
					(cpu_bypass_command_available and cpu_bypass_command_accept)));

	process(clk, reset, starting_new_memory_write,
				invalidate_slot_return, CACHE_STALL_ENABLE_REG)
		variable next_free_invalidate_slot_count_var: 
			integer range 0 to NUMBER_OF_INVALIDATE_SLOTS_PER_CORE - 2 ;
		variable i1, d1: boolean;
	begin

		i1 := invalidate_slot_return;
		d1 := starting_new_memory_write;

		next_free_invalidate_slot_count_var := free_invalidate_slot_count;


		if(clk'event and (clk = '1')) then
			if((reset = '1') or (accept_cpu_reset and cpu_reset)) then 
				-- note: give up two slots for potential writes to
				--   page tables as part of mmu activity!
				free_invalidate_slot_count <= NUMBER_OF_INVALIDATE_SLOTS_PER_CORE - 2; 
			elsif (CACHE_STALL_ENABLE_REG(0) = '1') then
				if (i1 and (not d1)) then
					next_free_invalidate_slot_count_var :=
						next_free_invalidate_slot_count_var + 1;
				elsif ((not i1) and d1) then 
					next_free_invalidate_slot_count_var :=
						next_free_invalidate_slot_count_var - 1;
				end if;
				free_invalidate_slot_count <= next_free_invalidate_slot_count_var; 
			end if;
		end if;
		
	end process;
	DCACHE_STALL <= (free_invalidate_slot_count = 0);

			
	

	-----------------------------------------------------------------------------------------------
	--  invalidate logic..
	-----------------------------------------------------------------------------------------------
    	MMU_TO_DCACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_req(0) <= '1' when syn_inval_accept else '0';
	syn_inval_ready <= (MMU_TO_DCACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_ack(0) = '1');
	syn_inval_applicable <= syn_inval_ready and
					(MMU_TO_DCACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_data(26) = '1');
	syn_inval_accept <= (dcache_state = SYN_INVALIDATE);


    	NOBLOCK_MMU_TO_DCACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_req(0) <= 
			'1' when coherence_inval_accept else '0';
    	coherence_inval_ready <= (NOBLOCK_MMU_TO_DCACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_ack(0) = '1');
    	coherence_inval_applicable <= 
			coherence_inval_ready and 
			     (NOBLOCK_MMU_TO_DCACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_data(26) = '1');
	coherence_inval_accept <=  
		(not waiting_on_tags_arrays) and 
			(((cpu_valid(0) = '1') and cpu_command_is_not_a_clear_or_flush) 
						or ((cpu_valid(0) = '0') and (dcache_state = IDLE))); 

	tag_invalidate_apply(0) <= 
		'1' when ((syn_inval_accept and syn_inval_applicable) or 
				(coherence_inval_accept and coherence_inval_applicable))
											else '0'; 
	tag_invalidate_line_address
		<= MMU_TO_DCACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_data(25 downto 0)
				when (syn_inval_accept and syn_inval_applicable) else
					NOBLOCK_MMU_TO_DCACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_data(25 downto 0);
	
	cpu_command_is_not_a_clear_or_flush <=
			exec_tag_access_cpu and (dcache_needs_to_be_flushed(0) = '0');



	-------------------------------------------------------------------------------------------
	-- registers, muxes, parsing..
	-------------------------------------------------------------------------------------------
	beParse: parse_from_backend_Volatile 
			port map (
    					from_be  => from_backend ,
    					be_valid  => be_valid ,
    					be_counter  => be_counter ,
    					be_tag_command  => be_tag_command ,
    					be_array_command  => be_array_command ,
    					be_dword_id  => be_dword_id ,
    					be_last_dword  => be_last_dword ,
    					be_acc  => be_acc ,
    					be_cacheable  => be_cacheable ,
    					be_mae  => be_mae ,
    					be_access_error  => be_access_error ,
    					be_dword  => be_dword 
				);

	---------------------------------------------------------------------------------------
	-- slow request..  if slow_request_has_lock=true, then only slow requests will be
	-- 		permitted.  This is required to ensure sanctity of lock in the
	--		multi-threaded case
	---------------------------------------------------------------------------------------
	from_cpu_slow   <= cpu_slow_command;
	slow_request_selected <= (slow_request_has_lock and (from_cpu_slow(120) = '1'))
					or ((not slow_request_has_lock) and (from_cpu_slow(120) = '1') and
							(from_cpu_fast(120) = '0'));
	slow_request_wants_lock <= (from_cpu_fast(120) = '0') and (from_cpu_slow(120) = '1') and 
										(from_cpu_slow(118) = '1');

	process(clk, reset, slow_request_has_lock, slow_request_wants_lock, 
					latch_cpu_commands, slow_request_selected, 
					latch_cpu_commands, trap_dcache, untrap_dcache)
		variable slow_request_has_lock_var: boolean;
	begin
		slow_request_has_lock_var := slow_request_has_lock;
		if((latch_cpu_commands or cpu_bypass_command_available) and slow_request_selected) then
			-- modify only if not if this operation is trapped out...
			if (trap_dcache or (DCACHE_TRAPPED and (not untrap_dcache))) then
				slow_request_has_lock_var := false;
			else
				slow_request_has_lock_var := slow_request_wants_lock;
			end if;
		end if;

		if(clk'event and (clk = '1')) then
			-- coming out of reset or trap, clear the lock.
			if(reset = '1') then
				slow_request_has_lock <= false;
			else
				slow_request_has_lock <= slow_request_has_lock_var;
			end if;
		end if;
	end process;

	---------------------------------------------------------------------------------------
	-- fast request: suppressed when slow_request_has_lock = true  (line 1427).
	---------------------------------------------------------------------------------------
	from_cpu_fast <= cpu_fast_command;

	---------------------------------------------------------------------------------------
	-- registers.
	---------------------------------------------------------------------------------------
	process(clk,reset)
	begin
		if(clk'event and clk = '1') then
	   	   if reset = '1' then
			to_cpu_registered <= (others => '0');
			to_be_registered  <= (others => '0');

			latch_to_cpu_registered <= false;
			latch_to_be_registered <= false;

			cpu_valid_reg(0) <= '0';
			cpu_valid_fast_reg(0) <= '0';
			cpu_valid_slow_reg(0) <= '0';

			expect_be_response_reg <= false;

			dcache_in_trapped_state_reg <= (others => '0');
			cpu_req_type_reg <= (others => '0');
				
			fast_command_bypass_control_info_reg <= (others => '0');
			is_mem_access_asi_reg <= false;
		   else

			latch_to_cpu_registered <= latch_to_cpu;
			latch_to_be_registered <= latch_to_be;

			if(latch_cpu_commands) then

				skip_tag_lookup_slv_reg <= skip_tag_lookup_slv;

				cpu_valid_reg <= cpu_valid;
				cpu_valid_fast_reg <= cpu_valid_fast;
				cpu_valid_slow_reg <= cpu_valid_slow;

				cpu_req_type_reg <= cpu_req_type;
				cpu_asi_reg <= cpu_asi;
				is_mem_access_asi_reg <= is_mem_access_asi;

				cpu_byte_mask_reg <= cpu_byte_mask;
				cpu_addr_reg <= cpu_addr;
				cpu_write_data_reg <= cpu_write_data;

				lock_bus_reg <= lock_bus;
				is_flush_asi_reg <= is_flush_asi;
				is_mmu_ctrl_reg_write_reg <= is_mmu_ctrl_reg_write;
				flush_line_only_reg <= flush_line_only;
				is_supervisor_asi_reg <= is_supervisor_asi;
				is_mmu_access_asi_reg <= is_mmu_access_asi;
				is_memory_write_reg <= is_memory_write;
				is_memory_read_reg <= is_memory_read;
				is_mmu_fsr_write_reg <= is_mmu_fsr_write;
				is_stbar_reg <= is_stbar;
				is_ccu_request_reg <= is_ccu_request;

				dcache_in_trapped_state_reg <= dcache_in_trapped_state;

				fast_command_bypass_control_info_reg <= fast_command_bypass_control_info;
			
			elsif clear_cpu_commands then

				cpu_valid_reg(0) <= '0';
				cpu_valid_fast_reg(0) <= '0';
				cpu_valid_slow_reg(0) <= '0';

			end if;

			if(latch_to_cpu) then
				to_cpu_registered <= to_cpu;
			end if;

			if(latch_to_be) then
				to_be_registered <= to_be;
				expect_be_response_reg <= expect_be_response;
			end if;
                  end if;
		end if;
	end process;

	-------------------------------------------------------------------------------------------
	-- analyse commands.
	-------------------------------------------------------------------------------------------
	decodeCpu: merge_and_decode_from_cpu_VVD
		port map (from_cpu_fast => from_cpu_fast, from_cpu_slow => from_cpu_slow,
				is_thread_head => is_thread_head,
				lock_bus => lock_bus,
				cpu_valid_fast => cpu_valid_fast,
				cpu_valid_slow => cpu_valid_slow,
				cpu_req_type => cpu_req_type,
				cpu_asi => cpu_asi,
				cpu_byte_mask => cpu_byte_mask,
				cpu_addr => cpu_addr,
				cpu_write_data => cpu_write_data,
				is_flush_asi => is_flush_asi,
				is_mmu_ctrl_reg_write=> is_mmu_ctrl_reg_write,
				flush_line_only => flush_line_only,
				is_supervisor_asi => is_supervisor_asi,
				is_mmu_access_asi => is_mmu_access_asi,
				dcache_needs_to_be_flushed => dcache_needs_to_be_flushed,
				is_memory_read => is_memory_read,
				is_memory_write => is_memory_write,
				is_mmu_fsr_write => is_mmu_fsr_write,
				is_stbar => is_stbar,
				is_ccu_request => is_ccu_request);
	
	
	

	-------------------------------------------------------------------------------------------
	-- ACTIVE CPU FOR THIS REQUEST!
	-------------------------------------------------------------------------------------------
	cpu_thread_id <= cpu_req_type(5 downto 4);
	cpu_thread_id_registered <= cpu_req_type_reg(5 downto 4);
	active_cpu_thread_id <= cpu_thread_id when 
					(accept_cpu_commands and 
							(cpu_fast_command_valid or cpu_slow_command_valid))
								 else cpu_thread_id_registered;
	ACPU <= 0 when (active_cpu_thread_id = "00") else 1;

	
	-------------------------------------------------------------------------------------------
	-- DCACHE_TRAPPED is derived from dcache_trapped_vector
	-------------------------------------------------------------------------------------------
	process(dcache_trapped_vector, active_cpu_thread_id)
		variable tv : boolean;
	begin
		tv := true;
		if(active_cpu_thread_id = "00") then
			tv := (dcache_trapped_vector(0) = '1');
		elsif (active_cpu_thread_id = "01") then
			tv := (dcache_trapped_vector(1) = '1');
		end if;
		DCACHE_TRAPPED <= tv;
	end process;
	-------------------------------------------------------------------------------------------
			

	skip_tag_lookup_slv(0) <= '1' when skip_tag_lookup else '0';


        dcache_in_trapped_state(0) <= '1' when (DCACHE_TRAPPED and (is_thread_head(0) = '0')) else '0';


	idActions: identify_cpu_actions_VVD
			port map (
				-- inputs: note: except for is_a_hit, all
				-- are registered, because cpu-actions 
				-- are delayed by 1 cycle relative to the
				-- acceptance of the cpu-command (latch_command).
    				exec_cpu  => exec_cpu_reg ,
    				next_dcache_trapped  => dcache_in_trapped_state_reg,
    				is_ccu_request  => is_ccu_request_reg ,
    				is_a_hit  => is_a_hit ,
    				skip_tag_lookup  => skip_tag_lookup_slv_reg,
    				is_memory_write  => is_memory_write_reg,
    				is_memory_read  => is_memory_read_reg ,
    				is_flush_asi  => is_flush_asi_reg ,
    				is_stbar  => is_stbar_reg ,
    				is_mmu_access_asi  => is_mmu_access_asi_reg ,
    				is_mmu_fsr_write  => is_mmu_fsr_write_reg ,
				-- outputs..
    				write_dword_hit  => write_dword_hit ,
    				write_dword_miss  => write_dword_miss ,
    				read_dword_hit  => read_dword_hit ,
    				read_dword_miss  => read_dword_miss ,
    				finished_flush_or_nop  => finished_flush_or_nop ,
    				write_to_mmu_or_bypass  => write_to_mmu_or_bypass ,
    				read_from_mmu_or_bypass  => read_from_mmu_or_bypass ,
    				write_to_mmu_fsr  => write_to_mmu_fsr ,
    				send_to_be  => send_to_be ,
    				no_response_from_be  => no_response_from_be 
			);
	-------------------------------------------------------------------------------------------
	-- construct predicates/inputs
	-------------------------------------------------------------------------------------------
	is_a_hit <= is_hit  and cpu_permissions_ok;

	cpu_reset <= ((NOBLOCK_CPU_to_DCACHE_reset_pipe_read_ack(0) = '1') and 
				  (NOBLOCK_CPU_to_DCACHE_reset_pipe_read_data(0) = '1'));


	be_response_can_be_applied <= 
		(not waiting_on_tags_arrays) and  (be_valid(0) = '1') and 
			((dcache_state = RECV_WAIT_ON_BE_FIRST_DWORD)
				or
			  (dcache_state = RECV_WAIT_ON_BE_REMAINING_DWORDS));

	first_be_response_can_be_applied <= 
		(not waiting_on_tags_arrays) and
			(dcache_state = RECV_WAIT_ON_BE_FIRST_DWORD) and (be_valid(0) = '1'); 

	be_has_exception <= be_response_can_be_applied and ((be_mae(0) = '1') or (be_access_error(0) = '1'));
			
	be_response_available <= 
			((noblock_dcache_backend_to_frontend_command_pipe_read_ack(0) = '1') and 
				  (noblock_dcache_backend_to_frontend_command_pipe_read_data(83) = '1'));

	be_ready_for_command  <= (dcache_frontend_to_backend_pipe_write_ack(0) = '1');

	-- Two cases to consider
	--   fast valid 
	--   (not fast_valid) and slow_valid
	cpu_ready_for_response  <= 
			((cpu_valid_fast_reg(0) = '1') and (DCACHE_to_CPU_response_pipe_write_ack(0) = '1'))
				or
			((cpu_valid_fast_reg(0) = '0') and 
				(cpu_valid_slow_reg(0) = '1') and 
					(DCACHE_to_CPU_slow_response_pipe_write_ack(0) = '1'));


	-- exec cpu tag command every time a cpu command is latched!
	exec_tag_access_cpu <= (latch_cpu_commands and (cpu_valid(0) = '1'));


	-- 1 cycle after cpu-command is accepted..
	exec_be <= be_response_can_be_applied;

	be_is_needed <= (send_to_be(0) = '1');
	expect_be_response <= be_is_needed and (no_response_from_be(0) = '0');

	-- computed immediately when cpu-command is accepted.
	skip_tag_lookup <= ((is_flush_asi(0) = '1') or (is_mmu_access_asi(0) = '1') or
					(is_mmu_fsr_write(0) = '1') or
					(is_stbar(0) = '1'));
	do_tag_lookup <= (cpu_valid(0) = '1') and 
					(not skip_tag_lookup) and
					((is_memory_read(0) = '1') or (is_memory_write(0) = '1')) and
					((not trap_dcache) or (is_ccu_request(0) = '1'));
	---------------------------------------------------------------------------------------------
	-- control state machine
	---------------------------------------------------------------------------------------------
	process(clk, reset, dcache_state, 
			cpu_command_available,
			cpu_reset,
			be_ready_for_command,
			be_is_needed,
			expect_be_response,
			be_response_available,
			cpu_ready_for_response,
			be_has_exception,
			is_thread_head,
			dcache_trapped_vector,
			DCACHE_TRAPPED,
			ACPU,
			waiting_on_tags_arrays)
		variable next_dcache_state : DcacheState;
		variable accept_cpu_commands_var  : boolean;
		variable latch_cpu_commands_var  : boolean;
		variable clear_cpu_commands_var : boolean;
		variable latch_tag_results_var  : boolean;
		variable latch_be_info_var	: boolean;
		variable latch_to_be_var	: boolean;
		variable latch_to_cpu_var	: boolean;
		variable accept_be_response_var  : boolean;
		variable write_to_be_var	 : boolean;
		variable write_to_cpu_var	 : boolean;
		variable next_be_has_completed_var	 : boolean;
		variable next_dcache_trapped_vector_var: std_logic_vector(0 to 1);
		variable latch_expect_be_response_var : boolean;
		variable send_cpu_reset_ack_var : boolean;
		variable accept_cpu_reset_var : boolean;
	begin
		next_dcache_state := dcache_state;
		accept_cpu_commands_var := false;
		latch_cpu_commands_var  := false;
		clear_cpu_commands_var := false;
		accept_be_response_var  := false;
		latch_be_info_var := false;
		latch_to_be_var := false;
		latch_to_cpu_var := false;
		write_to_be_var	 := false;
		write_to_cpu_var	 := false;
		next_be_has_completed_var := false;
		latch_expect_be_response_var := false;
		send_cpu_reset_ack_var := false;
		accept_cpu_reset_var := false;

		-- inherit the trapped status.
		next_dcache_trapped_vector_var := dcache_trapped_vector;

		case dcache_state is 
			when IDLE => 
				-- Ready to accept..
			    accept_cpu_reset_var := true;

			    -- important: it is assumed that there is always room
			    -- for the reset ack to the cpu..
			    if ((not waiting_on_tags_arrays) and cpu_reset) then
				-- we will clear the tag valid bits..
				send_cpu_reset_ack_var := true;

				-- clear the trapped vector.
				next_dcache_trapped_vector_var := (others => '0');
			    elsif (not waiting_on_tags_arrays) then  
				accept_cpu_commands_var := true;
				if(cpu_command_available) then
					latch_cpu_commands_var := true;
					next_dcache_state := CHECK_HIT_OR_MISS;
					if(is_thread_head(0) = '1') then
						-- clear the trapped vector entry for ACPU.
						next_dcache_trapped_vector_var(ACPU) := '0';
					end if;
				end if;
			     end if;
			when CHECK_HIT_OR_MISS =>
				if (waiting_on_tags_arrays) then
					-- hang on..
					next_dcache_state := CHECK_HIT_OR_MISS;
				elsif (be_is_needed) then

					-- cpu command received in previous cycle and
					-- tags, arrays have been accessed.
					-- need to go to be with registered cpu information.
					write_to_be_var := true;
					if be_ready_for_command then
						-- be is accepting..
						if expect_be_response then
							-- be response is expected... go wait on it.
							if((write_dword_miss(0) = '1') or 
								(read_dword_miss(0) = '1')) then
								next_dcache_state := SYN_INVALIDATE;
							else
								next_dcache_state := RECV_WAIT_ON_BE_FIRST_DWORD;
							end if;
						else
							-- be response is not expected..
							-- can send response to CPU!
							write_to_cpu_var := true;
							if(cpu_ready_for_response) then
							   -- CPU has accepted.. see if it has a command..
							   -- provided stall is not asserted.
							        accept_cpu_commands_var := true;
								if(cpu_command_available) then
									latch_cpu_commands_var := true;
									if(is_thread_head(0) = '1') then
									  -- clear the trapped vector entry for ACPU.
										next_dcache_trapped_vector_var(ACPU) 
												:= '0';
									end if;
									-- stay in CHECK_HIT_OR_MISS.
								else
									clear_cpu_commands_var := true;
									next_dcache_state := IDLE;
								end if;
							else
								-- cpu not ready, never mind, but latch to_cpu!
								-- this is a write-through situation or a flush
								-- write to the mmu or a write-bypass... cpu
								-- return data value is not important.
								latch_to_cpu_var := true;
								next_dcache_state := SEND_WAIT_ON_CPU;	
							end if;
							-- be is trivially done...
							next_be_has_completed_var := true;
						end if;
					else
						-- be response is expected..  remember it.
						latch_expect_be_response_var := true;	

						-- be not ready to be receiver, latch to_be!
						latch_to_be_var := true;

						-- cpu will be responded to later... 
						--  so latch to_cpu.
						latch_to_cpu_var := true;
						next_dcache_state := SEND_WAIT_ON_BE;	
					end if;
				else -- be is not needed..
					next_be_has_completed_var := true;
					-- try to write to cpu...
					write_to_cpu_var := true;
					if cpu_ready_for_response then 
					   -- cpu write is on! only if no stall...
						accept_cpu_commands_var := true;
						if cpu_command_available then
							-- and new command is available!!
							latch_cpu_commands_var := true;
							if(is_thread_head(0) = '1') then
							        -- clear the trapped vector entry for ACPU.
								next_dcache_trapped_vector_var(ACPU) := '0';
							end if;
							-- stay in CHECK_HIT_OR_MISS.
						else
							-- no new command.. clear command info.
							clear_cpu_commands_var := true;
							next_dcache_state := IDLE;
						end if;
					else
						-- cpu not ready to receive response..
						-- delayed response to CPU.. latch to_cpu.
						latch_to_cpu_var := true;
						next_dcache_state := SEND_WAIT_ON_CPU;	
					end if;
				end if;
			when SYN_INVALIDATE =>
				if(syn_inval_ready) then
					next_dcache_state := RECV_WAIT_ON_BE_FIRST_DWORD;	
				end if;
			when SEND_WAIT_ON_BE =>
				write_to_be_var := true;
				if be_ready_for_command then
					if(expect_be_response_reg) then
						if((write_dword_miss(0) = '1') or 
							(read_dword_miss(0) = '1')) then
							next_dcache_state := SYN_INVALIDATE;
						else
							next_dcache_state := RECV_WAIT_ON_BE_FIRST_DWORD;
						end if;
					else
						-- No response is expected from the backend..
						-- we can send the response to CPU!
						write_to_cpu_var := true;
						if(cpu_ready_for_response) then
						-- CPU has accepted.. see if it has a command..
						-- but ensure no stall!
			    				accept_cpu_reset_var := true;
							if(cpu_reset) then
								send_cpu_reset_ack_var := true;
								-- clear the trapped vector.
								next_dcache_trapped_vector_var := 
										(others => '0');
								next_dcache_state := IDLE;
							else
								accept_cpu_commands_var := true;
								if(cpu_command_available) then
									latch_cpu_commands_var := true;
									if(is_thread_head(0) = '1') then
										-- clear trapped for ACPU
										next_dcache_trapped_vector_var(ACPU) 
												:= '0';
									end if;
									next_dcache_state := CHECK_HIT_OR_MISS;
								else
									clear_cpu_commands_var := true;
									next_dcache_state := IDLE;
								end if;
							end if;
						else
							-- cpu not ready for response..
						        -- to_cpu_reg has already been updated.	
							next_dcache_state := SEND_WAIT_ON_CPU;	
						end if;

						-- no response needed from be, ergo
						-- be has completed.
						next_be_has_completed_var := true;
					end if;
				end if;
			when RECV_WAIT_ON_BE_FIRST_DWORD =>

			    if(not waiting_on_tags_arrays) then 
				-- word from BE will be returned to the CPU
				-- and possible written into the cache array.
				accept_be_response_var := true;
				if (be_response_available) then

					-- cpu will get the response in the
					-- next cycle..
					next_dcache_state := SEND_WAIT_ON_CPU;
					latch_be_info_var := true;

					-- to_cpu will be computed in this
					-- state but used in the next.
					latch_to_cpu_var := true;

					if (be_has_exception) then
						-- mark that the ACPU thread has an exception.
						-- Note that the other thread will continue normal
						-- execution..
						next_dcache_trapped_vector_var(ACPU) := '1';
					end if;
					if(be_last_dword(0) = '1') then
						next_be_has_completed_var := true;
					end if;
				end if;
 	                     end if;
			when SEND_WAIT_ON_CPU =>
				-- in the previous state, we have probably accessed tags/arrays.
				-- ensure that these are done....
				if(waiting_on_tags_arrays) then
					next_be_has_completed_var := be_has_completed;
				else
				  write_to_cpu_var := true;
				  if cpu_ready_for_response then
				     if(be_has_completed) then
			    		accept_cpu_reset_var := true;
					if(cpu_reset) then
						send_cpu_reset_ack_var := true;
						next_dcache_trapped_vector_var := (others => '0');
						next_dcache_state := IDLE;
					else
						accept_cpu_commands_var := true;
						if (cpu_command_available) then
							latch_cpu_commands_var := true;
							if(is_thread_head(0) = '1') then
								-- clear the trapped state for ACPU.
								next_dcache_trapped_vector_var(ACPU) := '0';
							end if;
							next_dcache_state := CHECK_HIT_OR_MISS;
						else 
							clear_cpu_commands_var := true;
							next_dcache_state := IDLE;
						end if;
					end if;
				     else
					next_dcache_state := RECV_WAIT_ON_BE_REMAINING_DWORDS;
				     end if;
				  else
					-- if be has completed, it stays completed
					-- while we wait for the cpu.
					next_be_has_completed_var := be_has_completed;
				  end if;
				end if;
			when RECV_WAIT_ON_BE_REMAINING_DWORDS =>
				-- Technically, in this state, we should ensure that
				-- the tags/arrays are not pending..
				if(waiting_on_tags_arrays) then 
				  next_be_has_completed_var := be_has_completed; 
				else
				  accept_be_response_var := true;
				  if (be_response_available) then
					if(be_last_dword(0) = '1') then
						next_be_has_completed_var := true;
						clear_cpu_commands_var := true;
						next_dcache_state := IDLE;
					end if;
				  end if;
				end if;
		end case;

		accept_cpu_commands <= accept_cpu_commands_var;
		latch_cpu_commands <= latch_cpu_commands_var;
		clear_cpu_commands <= clear_cpu_commands_var;
		latch_be_info  <= latch_be_info_var;
		latch_to_be  <= latch_to_be_var;
		latch_to_cpu  <= latch_to_cpu_var;
		accept_be_response <= accept_be_response_var;
		write_to_be	   <= write_to_be_var;
		write_to_cpu	   <= write_to_cpu_var;

		untrap_dcache <= (DCACHE_TRAPPED and (next_dcache_trapped_vector_var(ACPU) = '0'));
		trap_dcache <= (next_dcache_trapped_vector_var(ACPU) = '1');

		send_cpu_reset_ack <= send_cpu_reset_ack_var;
		accept_cpu_reset <= accept_cpu_reset_var;
		

		if clk'event and clk = '1' then
			if reset = '1' then	
				dcache_state <= IDLE;
				be_has_completed <= false;
				dcache_trapped_vector <= (others => '0');
			else
				dcache_state <= next_dcache_state;
				be_has_completed <= next_be_has_completed_var;
				dcache_trapped_vector <= next_dcache_trapped_vector_var;
			end if;
		end if;	
	end process;

	------------------------------------------------------------------------------------------------------
	-- accessDcache
	------------------------------------------------------------------------------------------------------
	arrays_start_req  <= '1' when (send_cpu_reset_ack or latch_cpu_commands or be_response_can_be_applied) else '0';
	tags_start_req  <= arrays_start_req or tag_invalidate_apply(0);

	tags_arrays_trigger <= tags_start_req or arrays_start_req;

	

	init_flag  <= '1' when send_cpu_reset_ack else '0';
	access_mae <= be_mae(0) when be_response_can_be_applied else '0';
	access_tags_acc <= be_acc when be_response_can_be_applied  else (others => '0');

	-- note that when the BE command is executed, we use the registered supervisor bit from the cpu.
	access_S <= is_supervisor_asi_reg(0) when be_response_can_be_applied else is_supervisor_asi(0);

	-- note that when the BE command is executed, we use the registered address/byte-mask from the cpu.
	--
	-- Careful here... the byte mask to be used for the write to the array is the following..
	--    when cpu write is being performed .. cpu_byte_mask,  else 0xff.
	--
	access_byte_mask <=  cpu_byte_mask when latch_cpu_commands else byte_mask_ff;
	access_is_read <= '0' when be_response_can_be_applied else is_memory_read(0);
	access_is_ifetch <= '0';

	-- cpu_tag_command
	process(dcache_needs_to_be_flushed, flush_line_only, do_tag_lookup, trap_dcache, init_flag)
	begin
		if(init_flag = '1') then
			cpu_tag_command <= CACHE_TAG_CLEAR_ALL;
		elsif(trap_dcache and (is_ccu_request(0) = '0')) then
			cpu_tag_command <= CACHE_TAG_NOP;
		elsif(dcache_needs_to_be_flushed(0) = '1') then
			if(flush_line_only(0) = '1') then
				cpu_tag_command <= CACHE_TAG_CLEAR_LINE;
			else
				cpu_tag_command <= CACHE_TAG_CLEAR_ALL;
			end if;
		elsif do_tag_lookup then
			cpu_tag_command <= CACHE_TAG_LOOKUP;
		else
			cpu_tag_command <= CACHE_TAG_NOP;
		end if;
	end process;
			
	------------------------------------------------------------------------------------------------------

	TagsAndArraysBlock: block
    		signal access_tag_lookup, access_tag_insert, 
				access_tag_clear_line,
				access_tag_clear_all : std_logic;
    		signal access_tag_addr : std_logic_vector(31 downto 0);
    		signal tag_in: std_logic_vector(0 downto 0);
    		signal tag_out: std_logic_vector(0 downto 0);
    		signal access_array_command, cpu_array_command : std_logic_vector(2 downto 0);
    		signal access_array_addr : std_logic_vector(31 downto 0);
    		signal access_dword : std_logic_vector((8*(2**LOG2_DATA_WIDTH_IN_BYTES))-1 downto 0);
	begin
	   tag_in (0) <= '0';


	   -------------------  Tag side ---------------------------------------------------------------
	   --
	   -- NOTE: In the "be" case, tags are modified only in the first fetch.
	   --          In subsequent fetches, tags will be cleared if there is
	   --          an error or mae.
	   --       
	   access_tag_command <=  CACHE_TAG_CLEAR_LINE when (exec_be and ((be_mae(0) = '1') or (be_access_error(0) = '1')))
					 else be_tag_command when (exec_be and first_be_response_can_be_applied)
						 else cpu_tag_command when  exec_tag_access_cpu else CACHE_TAG_NOP;

	

	-- note that when the BE command is executed, we use the registered address/byte-mask from the cpu.
	   access_tag_addr <= cpu_addr_reg when exec_be else cpu_addr;
	
	

	--
	-- TODO: split access_tag_command into lookup, clear-line, clear-all, insert.   
	-- 	  The insert can only be from the BE side and the lookup can only be
	--	  from the CPU side.  Currently, the two are being smeared into 
	--        the same signal access_tag_command, which results in a false 
	--	  critical path being flagged!
	--	
	--
	   -----------------------------------------------------------------------------------------------
	
	   -------------------  Array side ---------------------------------------------------------------
	    -- cpu_array_command
	   cpu_array_command <= CACHE_ARRAY_NOP when ((trap_dcache and (is_ccu_request(0) = '0')) or 
					skip_tag_lookup or (init_flag = '1'))
				else CACHE_ARRAY_READ_DWORD when (is_memory_read(0) = '1') 
				else CACHE_ARRAY_WRITE_DWORD  when (is_memory_write(0) = '1') 
				else CACHE_ARRAY_NOP;

	   -----------------------------------------------------------------------------------
	   -- control logic
	   -----------------------------------------------------------------------------------
	   -- if dword being written has an exception/error, do not update the cache array.
	   access_array_command <= 	
			CACHE_ARRAY_NOP when 
				(exec_be and ((be_mae(0) = '1')  or (be_access_error(0) = '1')))
						else be_array_command when exec_be
						else cpu_array_command when exec_tag_access_cpu
						else CACHE_ARRAY_NOP;
	   access_array_addr <= (cpu_addr_reg(31 downto 6) & be_dword_id & "000") when exec_be else cpu_addr;
	   access_dword      <= be_dword when exec_be else cpu_write_data;


	 
	   -- merged tags and arrays into one....
           directMappedGen: if (LOG_DCACHE_SET_ASSOCIATIVITY = 0) generate 
	      tagsArraysInst: 
		GenericDcacheTagsArraysWithInvalidate
                        generic map (name => "dcache-tags-arrays",
                                        log2_number_of_blocks => LOG2_NUMBER_OF_BLOCKS, -- 9  
                                        log2_block_size_in_bytes => LOG2_BLOCK_SIZE_IN_BYTES, -- 6
                                        address_width => 32,
                                        log2_data_width_in_bytes => 3)
			port map (
					trigger => tags_arrays_trigger,	
					done => tags_arrays_done,	
					init_flag => init_flag,
					access_mae => access_mae,
					access_S => access_S,
					access_is_read => access_is_read,
					access_is_ifetch => access_is_ifetch,
					access_acc => access_tags_acc,
					access_tag_command => access_tag_command,
					access_tag_addr => access_tag_addr,
					invalidate => tag_invalidate_apply,
					invalidate_line_address => tag_invalidate_line_address,
					is_hit => is_hit,
					permissions_ok => cpu_permissions_ok,
    					access_array_command  => access_array_command ,
    					access_byte_mask  => access_byte_mask ,
    					access_array_addr  => access_array_addr ,
    					access_dword  => access_dword ,
    					dword_out  => dword_out ,
    					clk => clk,
					reset => reset
				);

			-- in direct mapped case, the tags/arrays are guaranteed to respond
			--  in one clock cycle..
			waiting_on_tags_arrays <= false;
		end generate directMappedGen;


    		setAssociativeGen: if (LOG_DCACHE_SET_ASSOCIATIVITY > 0) generate 
	   
			-- note that lookup is only from cpu side and insert is only from the
	   		-- be side.  This prevents a false path from being flagged.
	   		access_tag_lookup <= '1' when (exec_tag_access_cpu and (cpu_tag_command = CACHE_TAG_LOOKUP))
							else '0';
	   		access_tag_insert <= '1' when (exec_be and first_be_response_can_be_applied and
									(be_tag_command = CACHE_TAG_INSERT))
							else '0';
	   		access_tag_clear_line <= '1' when (access_tag_command = CACHE_TAG_CLEAR_LINE) else '0';
	   		access_tag_clear_all <= '1' when (access_tag_command = CACHE_TAG_CLEAR_ALL) else '0';

	   	   tagsArraysInst: 
			GenericSetAssociativeCacheTagsArraysWithInvalidate
                             generic map (name => "dcache-tags-arrays",
                                        log2_number_of_blocks => LOG2_NUMBER_OF_BLOCKS, 	-- 9  
                                        log2_block_size_in_bytes => LOG2_BLOCK_SIZE_IN_BYTES, 	-- 6
					log2_associativity => LOG_DCACHE_SET_ASSOCIATIVITY, 	-- 4-way set associative
                                        address_width => 32,
                                        log2_data_width_in_bytes => 3)
		 	     port map (
					trigger => tags_arrays_trigger,	
					done => tags_arrays_done,	
					init_flag => init_flag,
					access_mae => access_mae,
					access_S => access_S,
					access_is_read => access_is_read,
					access_is_ifetch => access_is_ifetch,
					access_acc => access_tags_acc,
					access_tag_lookup => access_tag_lookup,
					access_tag_insert => access_tag_insert,
					access_tag_clear_line => access_tag_clear_line,
					access_tag_clear_all => access_tag_clear_all,
    					access_array_command  => access_array_command ,
					access_addr => access_array_addr,
    					access_byte_mask  => access_byte_mask ,
    					access_dword  => access_dword ,
					-- invalidation...
					invalidate => tag_invalidate_apply,
					invalidate_line_address => tag_invalidate_line_address,
					-- outputs.
					is_hit => is_hit,
					permissions_ok => cpu_permissions_ok,
					lookup_acc => lookup_acc,
    					dword_out  => dword_out ,
    					clk => clk,
					-- clock, reset.
					reset => reset
				);

			-- in set associative case, tags/arrays may need more than
			--    one clock cycle...
			process(clk, reset, tags_arrays_trigger, tags_arrays_done)
			begin
				if(clk'event and (clk = '1')) then
					if(reset = '1') then
						wait_on_tags_arrays <= false;
					else
						if(tags_arrays_trigger = '1')  then
							wait_on_tags_arrays <= true;
						elsif (wait_on_tags_arrays and (tags_arrays_done = '1')) then
							wait_on_tags_arrays <= false;
						end if;
					end if;
				end if;
			end process;
			waiting_on_tags_arrays <= wait_on_tags_arrays and (tags_arrays_done = '0');

		end generate setAssociativeGen;
	end block tagsAndArraysBlock;


	--------------------------------------------------------------------------------------------------
	-- pipe-connections
	--------------------------------------------------------------------------------------------------
	data_to_cpu <= 
		dword_out when  (dcache_state = CHECK_HIT_OR_MISS) and (is_memory_read_reg(0) = '1') 
			else be_dword when (first_be_response_can_be_applied  and (is_memory_read_reg(0) = '1')) 
					else ZERO_64;
	is_a_hit_to_cpu(0) <= is_a_hit(0) when (dcache_state = CHECK_HIT_OR_MISS)  else '0';
	mae_to_cpu(0)   <= be_mae(0) when first_be_response_can_be_applied else '0';
	access_error_to_cpu(0)  <= be_access_error(0) when first_be_response_can_be_applied else '0';
	mae_8_to_cpu <= (ZERO_5 & is_a_hit_to_cpu & access_error_to_cpu & mae_to_cpu);

	-- to_cpu itself will be registered if necessary.
	to_cpu <= (mae_8_to_cpu & data_to_cpu);

	-- no need to use registered values unless mentioned.. to_be itself will be registered
	-- if necessary.
	to_be <= (no_response_from_be  &
				lock_bus_reg &  -- note: registered value!
				read_dword_miss &
				write_dword_miss &
				write_dword_hit &
				read_from_mmu_or_bypass &
				write_to_mmu_or_bypass &
				write_to_mmu_fsr &
				cpu_asi_reg	 &
				cpu_byte_mask_reg &
				cpu_addr_reg &
				cpu_write_data_reg);

	NOBLOCK_CPU_to_DCACHE_reset_pipe_read_req (0) <= '1' when accept_cpu_reset else '0';
			
	NOBLOCK_CPU_to_DCACHE_command_pipe_read_req (0) <= '1' when 
				(not slow_request_has_lock)
					and
				accept_cpu_commands 
					and
				((normal_case and (cpu_valid_fast(0) = '1')) 
					or
				  (cpu_bypass_command_accept and bypass_case and (cpu_valid_fast(0) = '1')))
				 else '0';
	NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_req (0) <= '1' when 
				(accept_cpu_commands and
					(normal_case or 
						(cpu_bypass_command_accept and bypass_case)))
				and (cpu_valid_fast(0) = '0') and (cpu_valid_slow(0) = '1') else '0';

					
	--
	-- Added: do not consider fast valid if slow request has
	--         lock.
	cpu_fast_command_valid <= (NOBLOCK_CPU_to_DCACHE_command_pipe_read_data (142) = '1') 
					and 
					(NOBLOCK_CPU_to_DCACHE_command_pipe_read_ack (0) = '1')
					and 
					(not slow_request_has_lock);

	cpu_slow_command_valid <= (NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_data (120) = '1') 
					and 
					(NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_ack (0) = '1');

	cpu_fast_command <= 
		NOBLOCK_CPU_to_DCACHE_command_pipe_read_data(142 downto 142) & NOBLOCK_CPU_to_DCACHE_command_pipe_read_data (119 downto 0)
						when cpu_fast_command_valid
									else (others => '0');
	fast_command_bypass_control_info <=
		NOBLOCK_CPU_to_DCACHE_command_pipe_read_data (141 downto 120)
						when cpu_fast_command_valid
									else (others => '0');

	cpu_slow_command <=  NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_data when cpu_slow_command_valid
						else (others => '0');

	noblock_dcache_backend_to_frontend_command_pipe_read_req (0) <= 
				'1' when (accept_be_response or accept_be_bypass_response) else '0';
	from_backend <= noblock_dcache_backend_to_frontend_command_pipe_read_data when
				noblock_dcache_backend_to_frontend_command_pipe_read_ack(0) = '1' else
					(others => '0');

	dcache_frontend_to_backend_pipe_write_req (0) <= '1' when 
					(write_to_be or write_to_be_from_bypass) else '0';
	dcache_frontend_to_backend_pipe_write_data  <= 
			to_be_from_bypass when write_to_be_from_bypass else
				to_be_registered when (dcache_state = SEND_WAIT_ON_BE) else to_be;

	DCACHE_to_CPU_response_pipe_write_req(0) <= 
			'1' when write_bypass_to_cpu_fast or 
				((cpu_valid_fast_reg(0) = '1') and write_to_cpu) else '0';
	DCACHE_to_CPU_response_pipe_write_data <= 
			bypass_response_to_cpu when write_bypass_to_cpu_fast else
				to_cpu when (dcache_state = CHECK_HIT_OR_MISS) else to_cpu_registered;

	DCACHE_to_CPU_slow_response_pipe_write_req(0) <= 
			'1' when 
				write_bypass_to_cpu_slow or
					((cpu_valid_fast_reg(0) = '0') and
							(cpu_valid_slow_reg(0) = '1') and write_to_cpu)
							 else '0';

	DCACHE_to_CPU_slow_response_pipe_write_data <= 
			bypass_response_to_cpu when write_bypass_to_cpu_slow else
				to_cpu when (dcache_state = CHECK_HIT_OR_MISS) else to_cpu_registered;

	DCACHE_to_CPU_reset_ack_pipe_write_req(0) <= '1' when send_cpu_reset_ack  else '0';
	DCACHE_to_CPU_reset_ack_pipe_write_data(0) <= '1';

	-----------------------------------------------------------------------------------------------
	-- bypass controller
	-----------------------------------------------------------------------------------------------
	is_bypass_asi    <= (cpu_asi(7 downto 4) = "0010");
	is_pure_mem_access_asi <= ((cpu_asi(3 downto 0) = "1000") or
				(cpu_asi(3 downto 0) = "1001") or
				(cpu_asi(3 downto 0) = "1010") or
				(cpu_asi(3 downto 0) = "1011"));
	is_mem_access_asi <= is_pure_mem_access_asi or is_bypass_asi;
				
	
	--
	-- on dcache trapped, do not bypass, unless its a memory read.
	--  Note: if it is an nc tlb match, then do not treat the operation as a bypass in any case.
	--
	bypass_case      <= ((nc_tlb_match = '1') or is_bypass_asi) and  (not DCACHE_STALL) and 
					((is_bypass_asi and (is_memory_read(0) = '1')) or (not DCACHE_TRAPPED)) 
						and (not cpu_reset);

	normal_case      <= (not bypass_case) and (not bypass_response_pending) and (not DCACHE_STALL);

	cpu_command_available <= 
		(cpu_fast_command_valid or cpu_slow_command_valid) and normal_case;

	-- start the bypass only when the main FSM is accepting new commands.
	cpu_bypass_command_available <= 
		(cpu_fast_command_valid or cpu_slow_command_valid) and bypass_case and accept_cpu_commands;

	cpu_fast_ready_for_bypass_response <= (DCACHE_to_CPU_response_pipe_write_ack(0) = '1');
	cpu_slow_ready_for_bypass_response <= (DCACHE_to_CPU_slow_response_pipe_write_ack(0) = '1');

	bc: DcacheBypassController
		port map (clk => clk, reset => reset,
				cpu_bypass_command_available => cpu_bypass_command_available,	
				cpu_bypass_command_accept => cpu_bypass_command_accept,
				cpu_fast_valid => cpu_valid_fast(0),
				cpu_slow_valid => cpu_valid_slow(0),
				is_memory_write => is_memory_write(0),
				locked_access => lock_bus(0),
				cpu_asi => cpu_asi,
				cpu_byte_mask => cpu_byte_mask,
				cpu_address => cpu_addr,
				cpu_write_data => cpu_write_data,
				cpu_slow_ready_for_bypass_response => cpu_slow_ready_for_bypass_response,
				cpu_fast_ready_for_bypass_response => cpu_fast_ready_for_bypass_response,
				write_to_cpu_slow => write_bypass_to_cpu_slow,
				write_to_cpu_fast => write_bypass_to_cpu_fast,
				response_to_cpu => bypass_response_to_cpu,
				be_ready_for_request => be_ready_for_command,
				be_write => write_to_be_from_bypass,
				to_be_from_bypass => to_be_from_bypass,
				be_response_ready => be_response_available,
				be_read => accept_be_bypass_response,
				be_dword => be_dword,
				bypass_response_pending => bypass_response_pending);

	------------------------------------------------------------------------------------------
	-- Non-cacheable logic.
	------------------------------------------------------------------------------------------
	ncGen: if (TREAT_NONCACHEABLE_AS_BYPASS = 1) generate
	  gB: block
		signal nc_tlb_clear, nc_tlb_insert: std_logic;
		signal nc_tlb_lookup_supervisor, nc_tlb_lookup_read, nc_tlb_lookup_ifetch: std_logic;
		signal nc_tlb_insert_acc: std_logic_vector(2 downto 0);

		signal write_dword_miss_reg, read_dword_miss_reg: std_logic_vector(0 downto 0);
	  begin

		-- some local registers
		process(clk, reset)
		begin
			if(clk'event and (clk = '1')) then
				if(reset = '1') then
					write_dword_miss_reg(0) <= '0';
					read_dword_miss_reg(0) <= '0';
				else
					if(dcache_state = CHECK_HIT_OR_MISS) then
						write_dword_miss_reg <= write_dword_miss;
						read_dword_miss_reg  <= read_dword_miss;
					end if;

				end if;
			end if;
		end process;

		-- on a miss, insert into the nc tlb if the backend returned status as non-cacheable 
		nc_tlb_insert <= '1' when
				(first_be_response_can_be_applied 
						and 
						(be_cacheable(0) = '0') 
						and 
						(be_mae(0) = '0') 
						and 
						((write_dword_miss_reg(0) = '1') or (read_dword_miss_reg(0) = '1'))
						and
						(be_tag_command /= CACHE_TAG_INSERT))
					else '0';
		nc_tlb_insert_acc <= be_acc;
	
		nc_tlb_clear <= '1' when 
				((tags_start_req = '1') and (access_tag_command = CACHE_TAG_CLEAR_ALL)) 
					else '0';

		nc_tlb_lookup_ifetch <= '0';
		nc_tlb_lookup_read <= is_memory_read(0);
		nc_tlb_lookup_supervisor <= is_supervisor_asi(0);


		nc_tlb: nonCacheablePageTlb
			generic map (number_of_entries => 4)
			port map (lookup_virtual_address => cpu_addr,
					lookup_supervisor => nc_tlb_lookup_supervisor,
					lookup_read => nc_tlb_lookup_read,
					lookup_ifetch => nc_tlb_lookup_ifetch,
					insert_virtual_address => cpu_addr_reg,
					insert_acc => nc_tlb_insert_acc, 
					match => nc_tlb_match_base,
					insert => nc_tlb_insert,
					clear => nc_tlb_clear,	
					clk => clk, reset => reset);

		-- NC TLB match only applicable to pure memory accesses!
		nc_tlb_match <= nc_tlb_match_base when is_pure_mem_access_asi  else '0';
	  end block;
	end generate ncGen;

	noNcGen: if (TREAT_NONCACHEABLE_AS_BYPASS = 0) generate
		nc_tlb_match <= '0';
	end generate noNcGen;

	-- the control information is in this form..
	--  valid thread-id stream-id slot-id do-not-bypass  rd to-iu to-fp to-cp
	--   1     4         2         6       1              5    1    1       1 =  22
	--
	-- The bypass signal has the following format..
	-- valid cpu-id thread-id stream-id slot-id signed-type byte-mask   rd  rdata
	--   1     2      4         2         6        1          8         5   64  = 92
	process(dcache_state, 
			is_a_hit, 
			dword_out,
			cpu_byte_mask_reg,
			fast_command_bypass_control_info_reg, 
			tags_arrays_done,
			cpu_valid_fast_reg,
			cpu_thread_id_registered)
		variable to_iu : std_logic_vector (92 downto 0);
		variable to_fu : std_logic_vector (92 downto 0);
		variable valid, signed_type : std_logic;
	begin
		valid := fast_command_bypass_control_info_reg(21);
		signed_type := fast_command_bypass_control_info_reg(8);

		to_iu(92) := (valid and fast_command_bypass_control_info_reg(2));
		to_fu(92) := (valid and fast_command_bypass_control_info_reg(1));

		to_iu(91 downto 90) := cpu_thread_id_registered;
		to_fu(91 downto 90) := cpu_thread_id_registered;
	
		-- thread stream slot
		to_iu(89 downto 78) := fast_command_bypass_control_info_reg(20 downto 9);
		to_fu(89 downto 78) := fast_command_bypass_control_info_reg(20 downto 9);

		to_iu(77) := signed_type;
		to_fu(77) := signed_type;

		-- byte-mask
		to_iu(76 downto 69) := cpu_byte_mask_reg;
		to_fu(76 downto 69) := cpu_byte_mask_reg;

		-- rd
		to_iu(68 downto 64) := fast_command_bypass_control_info_reg(7 downto 3);
		to_fu(68 downto 64) := fast_command_bypass_control_info_reg(7 downto 3);

		-- rdata 
		to_iu(63 downto 0) := dword_out;
		to_fu(63 downto 0) := dword_out;

		if ((valid = '1') and
				(cpu_valid_fast_reg(0) = '1') and 
				(tags_arrays_done = '1') and
				(dcache_state = CHECK_HIT_OR_MISS) and 
				(is_a_hit(0) = '1')) then

			NOBLOCK_DCACHE_TO_CPU_IU_BYPASS_pipe_write_data <= to_iu;	
			NOBLOCK_DCACHE_TO_CPU_IU_BYPASS_pipe_write_req(0) <= to_iu(92);

			NOBLOCK_DCACHE_TO_CPU_FU_BYPASS_pipe_write_data <= to_fu;	
			NOBLOCK_DCACHE_TO_CPU_FU_BYPASS_pipe_write_req(0) <= to_fu(92);
		else
			NOBLOCK_DCACHE_TO_CPU_IU_BYPASS_pipe_write_data <= (others => '0');	
			NOBLOCK_DCACHE_TO_CPU_IU_BYPASS_pipe_write_req(0) <= '0';

			NOBLOCK_DCACHE_TO_CPU_FU_BYPASS_pipe_write_data <= (others => '0');	
			NOBLOCK_DCACHE_TO_CPU_FU_BYPASS_pipe_write_req(0) <= '0';
		end if;
	end process;

end DcacheFrontendCoreDaemon_arch;
--
-- This is a shell which includes 1-cycle of buffering at the
-- CPU request side in order to reduce the critical path. If this
-- is specified.
--
--
library std;
use std.standard.all;

library ieee;
use ieee.std_logic_1164.all;

library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;

library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;

library AjitCustom;
use AjitCustom.AjitGlobalConfigurationPackage.all;
use AjitCustom.AjitCoreConfigurationPackage.all;
use AjitCustom.AjitCustomComponents.all;
use AjitCustom.CachePackage.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

entity DcacheFrontendWithStallDaemon is -- 
  generic (tag_length : integer := 1); 
  port ( -- 
    NOBLOCK_CPU_to_DCACHE_command_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_command_pipe_read_data : in   std_logic_vector(142 downto 0);
    NOBLOCK_CPU_to_DCACHE_reset_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_reset_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_reset_pipe_read_data : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_data : in   std_logic_vector(120 downto 0);
    noblock_dcache_backend_to_frontend_command_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_dcache_backend_to_frontend_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_dcache_backend_to_frontend_command_pipe_read_data : in   std_logic_vector(83 downto 0);
    -----------------------------------------------------------------------------------------------
    NOBLOCK_DCACHE_TO_CPU_IU_BYPASS_pipe_write_req: out std_logic_vector(0 downto 0);
    NOBLOCK_DCACHE_TO_CPU_IU_BYPASS_pipe_write_ack: in std_logic_vector(0 downto 0);
    NOBLOCK_DCACHE_TO_CPU_IU_BYPASS_pipe_write_data: out std_logic_vector(92 downto 0);
    -----------------------------------------------------------------------------------------------
    NOBLOCK_DCACHE_TO_CPU_FU_BYPASS_pipe_write_req:  out std_logic_vector(0 downto 0);
    NOBLOCK_DCACHE_TO_CPU_FU_BYPASS_pipe_write_ack:  in std_logic_vector(0 downto 0);
    NOBLOCK_DCACHE_TO_CPU_FU_BYPASS_pipe_write_data: out std_logic_vector(92 downto 0);
    -----------------------------------------------------------------------------------------------
    DCACHE_to_CPU_reset_ack_pipe_write_req : out  std_logic_vector(0 downto 0);
    DCACHE_to_CPU_reset_ack_pipe_write_ack : in   std_logic_vector(0 downto 0);
    DCACHE_to_CPU_reset_ack_pipe_write_data : out  std_logic_vector(0 downto 0);
    DCACHE_to_CPU_response_pipe_write_req : out  std_logic_vector(0 downto 0);
    DCACHE_to_CPU_response_pipe_write_ack : in   std_logic_vector(0 downto 0);
    DCACHE_to_CPU_response_pipe_write_data : out  std_logic_vector(71 downto 0);
    DCACHE_to_CPU_slow_response_pipe_write_req : out  std_logic_vector(0 downto 0);
    DCACHE_to_CPU_slow_response_pipe_write_ack : in   std_logic_vector(0 downto 0);
    DCACHE_to_CPU_slow_response_pipe_write_data : out  std_logic_vector(71 downto 0);
    MMU_TO_DCACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_req: out std_logic_vector(0 downto 0);
    MMU_TO_DCACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_ack: in std_logic_vector(0 downto 0);
    MMU_TO_DCACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_data: in std_logic_vector(26 downto 0);
    NOBLOCK_MMU_TO_DCACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_req: out std_logic_vector(0 downto 0);
    NOBLOCK_MMU_TO_DCACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_ack: in std_logic_vector(0 downto 0);
    NOBLOCK_MMU_TO_DCACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_data: in std_logic_vector(26 downto 0);
    CACHE_STALL_ENABLE: in std_logic_vector(0 downto 0);
    NOBLOCK_INVALIDATE_SLOT_RETURN_pipe_read_req : out std_logic_vector(0 downto 0);
    NOBLOCK_INVALIDATE_SLOT_RETURN_pipe_read_ack : in std_logic_vector(0 downto 0);
    NOBLOCK_INVALIDATE_SLOT_RETURN_pipe_read_data: in std_logic_vector(0 downto 0);
    dcache_frontend_to_backend_pipe_write_req : out  std_logic_vector(0 downto 0);
    dcache_frontend_to_backend_pipe_write_ack : in   std_logic_vector(0 downto 0);
    dcache_frontend_to_backend_pipe_write_data : out  std_logic_vector(119 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity DcacheFrontendWithStallDaemon;
architecture DcacheFrontendDaemon_arch of DcacheFrontendWithStallDaemon is -- 

    signal NOBLOCK_BUFFERED_CPU_to_DCACHE_command_pipe_read_req : std_logic_vector(0 downto 0);
    signal NOBLOCK_BUFFERED_CPU_to_DCACHE_command_pipe_read_ack : std_logic_vector(0 downto 0);
    signal NOBLOCK_BUFFERED_CPU_to_DCACHE_command_pipe_read_data : std_logic_vector(142 downto 0);

    signal NOBLOCK_BUFFERED_CPU_to_DCACHE_slow_command_pipe_read_req : std_logic_vector(0 downto 0);
    signal NOBLOCK_BUFFERED_CPU_to_DCACHE_slow_command_pipe_read_ack : std_logic_vector(0 downto 0);
    signal NOBLOCK_BUFFERED_CPU_to_DCACHE_slow_command_pipe_read_data : std_logic_vector(120 downto 0);
begin

	ifBuffer: if (DCACHE_BUFFER_REQUEST > 0) generate
		qBuf: QueueBase
			generic map (name => "DcacheRequestQueue", queue_depth => 2,
						data_width => 143, save_one_slot => false)
			port map (
				clk => clk,
				reset => reset,
				data_in => NOBLOCK_CPU_to_DCACHE_command_pipe_read_data,
				push_req => NOBLOCK_CPU_to_DCACHE_command_pipe_read_ack(0),
				push_ack => NOBLOCK_CPU_to_DCACHE_command_pipe_read_req(0),
				data_out => NOBLOCK_BUFFERED_CPU_to_DCACHE_command_pipe_read_data,
				pop_req =>  NOBLOCK_BUFFERED_CPU_to_DCACHE_command_pipe_read_req(0),
				pop_ack =>  NOBLOCK_BUFFERED_CPU_to_DCACHE_command_pipe_read_ack(0)
			);
		qBufSlow: QueueBase
			generic map (name => "DcacheSlowRequestQueue", queue_depth => 2,
						data_width => 121, save_one_slot => false)
			port map (
				clk => clk,
				reset => reset,
				data_in => NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_data,
				push_req => NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_ack(0),
				push_ack => NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_req(0),
				data_out => NOBLOCK_BUFFERED_CPU_to_DCACHE_slow_command_pipe_read_data,
				pop_req =>  NOBLOCK_BUFFERED_CPU_to_DCACHE_slow_command_pipe_read_req(0),
				pop_ack =>  NOBLOCK_BUFFERED_CPU_to_DCACHE_slow_command_pipe_read_ack(0)
			);
	end generate ifBuffer;

	ifNoBuffer: if (DCACHE_BUFFER_REQUEST = 0) generate

		NOBLOCK_CPU_to_DCACHE_command_pipe_read_req <= NOBLOCK_BUFFERED_CPU_to_DCACHE_command_pipe_read_req;
    		NOBLOCK_BUFFERED_CPU_to_DCACHE_command_pipe_read_ack <= NOBLOCK_CPU_to_DCACHE_command_pipe_read_ack;
    		NOBLOCK_BUFFERED_CPU_to_DCACHE_command_pipe_read_data <= NOBLOCK_CPU_to_DCACHE_command_pipe_read_data;

		NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_req <= NOBLOCK_BUFFERED_CPU_to_DCACHE_slow_command_pipe_read_req;
    		NOBLOCK_BUFFERED_CPU_to_DCACHE_slow_command_pipe_read_ack <= NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_ack;
    		NOBLOCK_BUFFERED_CPU_to_DCACHE_slow_command_pipe_read_data <= NOBLOCK_CPU_to_DCACHE_slow_command_pipe_read_data;

	end generate ifNoBuffer;

	coreInst: DcacheFrontendWithStallCoreDaemon
			generic map (tag_length => tag_length)
			port map (
    				NOBLOCK_BUFFERED_CPU_to_DCACHE_command_pipe_read_req,
    				NOBLOCK_BUFFERED_CPU_to_DCACHE_command_pipe_read_ack,
    				NOBLOCK_BUFFERED_CPU_to_DCACHE_command_pipe_read_data,
    				NOBLOCK_CPU_to_DCACHE_reset_pipe_read_req,
    				NOBLOCK_CPU_to_DCACHE_reset_pipe_read_ack,
    				NOBLOCK_CPU_to_DCACHE_reset_pipe_read_data,
    				NOBLOCK_BUFFERED_CPU_to_DCACHE_slow_command_pipe_read_req,
    				NOBLOCK_BUFFERED_CPU_to_DCACHE_slow_command_pipe_read_ack,
    				NOBLOCK_BUFFERED_CPU_to_DCACHE_slow_command_pipe_read_data,
    				noblock_dcache_backend_to_frontend_command_pipe_read_req,
    				noblock_dcache_backend_to_frontend_command_pipe_read_ack,
    				noblock_dcache_backend_to_frontend_command_pipe_read_data,
    				-----------------------------------------------------------------------------------------------
    				NOBLOCK_DCACHE_TO_CPU_IU_BYPASS_pipe_write_req,
    				NOBLOCK_DCACHE_TO_CPU_IU_BYPASS_pipe_write_ack,
    				NOBLOCK_DCACHE_TO_CPU_IU_BYPASS_pipe_write_data,
    				-----------------------------------------------------------------------------------------------
    				NOBLOCK_DCACHE_TO_CPU_FU_BYPASS_pipe_write_req,
    				NOBLOCK_DCACHE_TO_CPU_FU_BYPASS_pipe_write_ack,
    				NOBLOCK_DCACHE_TO_CPU_FU_BYPASS_pipe_write_data,
    				-----------------------------------------------------------------------------------------------
    				DCACHE_to_CPU_reset_ack_pipe_write_req,
    				DCACHE_to_CPU_reset_ack_pipe_write_ack,
    				DCACHE_to_CPU_reset_ack_pipe_write_data,
    				DCACHE_to_CPU_response_pipe_write_req,
    				DCACHE_to_CPU_response_pipe_write_ack,
    				DCACHE_to_CPU_response_pipe_write_data,
    				DCACHE_to_CPU_slow_response_pipe_write_req,
    				DCACHE_to_CPU_slow_response_pipe_write_ack,
    				DCACHE_to_CPU_slow_response_pipe_write_data,
    				MMU_TO_DCACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_req,
    				MMU_TO_DCACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_ack,
    				MMU_TO_DCACHE_SYNONYM_INVALIDATE_PIPE_pipe_read_data,
    				NOBLOCK_MMU_TO_DCACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_req, 
    				NOBLOCK_MMU_TO_DCACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_ack, 
    				NOBLOCK_MMU_TO_DCACHE_COHERENCE_INVALIDATE_PIPE_pipe_read_data,
    				CACHE_STALL_ENABLE, 
    				NOBLOCK_INVALIDATE_SLOT_RETURN_pipe_read_req ,
    				NOBLOCK_INVALIDATE_SLOT_RETURN_pipe_read_ack ,
    				NOBLOCK_INVALIDATE_SLOT_RETURN_pipe_read_data,
    				dcache_frontend_to_backend_pipe_write_req ,
    				dcache_frontend_to_backend_pipe_write_ack ,
    				dcache_frontend_to_backend_pipe_write_data ,
    				tag_in,
    				tag_out,
    				clk ,
    				reset ,
    				start_req ,
    				start_ack ,
    				fin_req ,
    				fin_ack 
				);
end DcacheFrontendDaemon_arch;
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.Types.all;
use ahir.Subprograms.all;

entity nonCacheablePageTlb is
	generic (number_of_entries: integer := 4);
	port (
		lookup_virtual_address: in std_logic_vector(31 downto 0);
		lookup_supervisor, lookup_read, lookup_ifetch: in std_logic;

		insert_virtual_address: in std_logic_vector(31 downto 0);
		insert_acc: in std_logic_vector (2 downto 0);

		match: out std_logic;
		insert: in std_logic;
		clear : in std_logic;
		clk, reset:  in std_logic
	);
end entity;

architecture Behavioural of nonCacheablePageTlb is
	-- page ids.
	type TlbArray is array (natural range <>) of std_logic_vector(22 downto 0);
	signal tlb_array: TlbArray (number_of_entries-1 downto 0);
	signal valids: std_logic_vector(number_of_entries-1 downto 0);
	signal last_inserted_pointer: integer range 0 to number_of_entries-1;
	signal match_sig: std_logic;
	signal insert_match_sig: boolean;
	signal insert_match_pointer: integer range 0 to number_of_entries-1;

	function IncrementPointer(x: integer) return integer is
		variable ret_val: integer range 0 to number_of_entries-1;
	begin
		if(x = number_of_entries-1) then
			ret_val := 0;
		else
			ret_val := x + 1;
		end if;

		return(ret_val);
	end function;

	function nonCacheablePageTlbPermissionsOk (supervisor, read, ifetch: std_logic; acc: std_logic_vector(2 downto 0))
		return boolean is
		variable ret_var : boolean;
	begin
		ret_var := false;
		case acc is 
				      -- user : supervisor...
			when "000" => -- read : read
				ret_var := (ifetch = '0') and (read = '1');
			when "001" => -- read/write: read/write
				ret_var := (ifetch = '0');
			when "010" => -- read/exec : read/exec
				ret_var := ((read = '1') or (ifetch = '1'));
			when "011" => -- read/write/exec: read/write/exec
				ret_var := true;
			when "100" => -- exec : exec
				ret_var := (ifetch = '1');
			when "101" => -- read : read/write
				ret_var := (ifetch = '0') and
						((supervisor = '1') or (read = '1'));
			when "110" =>  -- none : read/exec
				ret_var := ((supervisor = '1') and 
						((read = '1') or (ifetch = '1')));
			when "111" => -- none : read/write/exec.
				ret_var := (supervisor = '1');
			when others  =>
				ret_var := false;
		end case;
		return ret_var;
	end function;

begin
	-- match process
	process(tlb_array, valids, lookup_virtual_address, lookup_supervisor, lookup_read, lookup_ifetch,
				insert, insert_acc, insert_virtual_address)

		variable match_var: std_logic_vector(number_of_entries-1 downto 0);
		variable tlb_entry : std_logic_vector(22 downto 0);
		variable acc_flags : std_logic_vector(2 downto 0);
		variable tlb_va : std_logic_vector(19 downto 0);
		variable acc_ok, insert_match, local_match,  lookup_match: boolean;
		variable insert_match_pointer_var: integer range 0 to number_of_entries-1;
	
	begin

		match_var := (others => '0');
		insert_match := false;
		local_match := false;
		insert_match_pointer_var := 0;
		
		for I in 0 to number_of_entries-1 loop
			tlb_entry := tlb_array(I);
			acc_flags := tlb_entry (22 downto 20);
			tlb_va    := tlb_entry (19 downto 0);

			acc_ok := 
				nonCacheablePageTlbPermissionsOk(lookup_supervisor, lookup_read, 
										lookup_ifetch, acc_flags);
			local_match     := ((insert = '1') and 
						    ((tlb_va = insert_virtual_address(31 downto 12))
							and (acc_flags = insert_acc)));
			if(local_match) then
				insert_match_pointer_var := I;
			end if;

			insert_match := insert_match or local_match;
			lookup_match     := (insert = '0') and acc_ok and
						(tlb_va = lookup_virtual_address(31 downto 12));
			if(lookup_match) then
				match_var(I) := valids(I);
			end if;
		end loop;

		match_sig <= OrReduce(match_var);
		insert_match_sig <= insert_match;
		insert_match_pointer <= insert_match_pointer_var;
	end process;
	match <= match_sig;


	-- management process
	process(clk, reset, valids, insert_acc, 
			insert_virtual_address, tlb_array, insert_match_sig, insert_match_pointer, last_inserted_pointer) 
		variable insert_pointer_var : integer range 0 to number_of_entries-1;
	begin
		if(insert_match_sig) then
			insert_pointer_var := insert_match_pointer;
		else
			insert_pointer_var := IncrementPointer (last_inserted_pointer);
		end if;

		if(clk'event and clk = '1') then
			if((reset = '1') or (clear = '1')) then
				valids <= (others => '0');
				last_inserted_pointer <= 0;
			elsif (insert = '1') then
				valids(insert_pointer_var) <= '1';
				tlb_array(insert_pointer_var) <= 
					insert_acc & insert_virtual_address(31 downto 12);
				last_inserted_pointer <= insert_pointer_var;
			end if;
		end if;
	end process;

end Behavioural;

--
-- THIS MUST BE IN SYNCH WITH fpunit/exec/fpu_module/merge_outs.aa
-- a simple mux.. fast-pipe is always read. If the top-bit of
-- fast-pipe is '0', then slow-pipe is read and forwarded.
-- Else fast-pipe itself is forwarded.
--
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
entity fpunit_exec_pipe_merge_daemon is -- 
  generic (tag_length: integer);
  port ( -- 
    fpunit_exec_to_writeback_fast_pipe_read_req : out  std_logic_vector(0 downto 0);
    fpunit_exec_to_writeback_fast_pipe_read_ack : in   std_logic_vector(0 downto 0);
    fpunit_exec_to_writeback_fast_pipe_read_data : in   std_logic_vector(96-1 downto 0);
    fpunit_exec_to_writeback_slow_pipe_read_req : out  std_logic_vector(0 downto 0);
    fpunit_exec_to_writeback_slow_pipe_read_ack : in   std_logic_vector(0 downto 0);
    fpunit_exec_to_writeback_slow_pipe_read_data : in   std_logic_vector(96-1 downto 0);
    fpunit_exec_to_writeback_pipe_write_req : out  std_logic_vector(0 downto 0);
    fpunit_exec_to_writeback_pipe_write_ack : in   std_logic_vector(0 downto 0);
    fpunit_exec_to_writeback_pipe_write_data : out  std_logic_vector(96-1 downto 0);
    clk : in std_logic;
    reset : in std_logic;
    start_req: in std_logic;
    start_ack: out std_logic;
    fin_req: in std_logic;
    fin_ack: out std_logic;
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0)
  );
  -- 
end entity fpunit_exec_pipe_merge_daemon;

architecture very_simple of fpunit_exec_pipe_merge_daemon is
	signal fpunit_exec_to_writeback_slow_pipe_needed: boolean;
	signal write_to_out : boolean;
begin
	start_ack <= '1';
	fin_ack <= '0';
	tag_out <= (others => '0');

	fpunit_exec_to_writeback_slow_pipe_needed <= 
		(fpunit_exec_to_writeback_fast_pipe_read_ack(0) = '1') and (fpunit_exec_to_writeback_fast_pipe_read_data(96-1) = '0');
	
	fpunit_exec_to_writeback_pipe_write_data <= 
		fpunit_exec_to_writeback_slow_pipe_read_data 
			when fpunit_exec_to_writeback_slow_pipe_needed 
				else fpunit_exec_to_writeback_fast_pipe_read_data;
	write_to_out <= ((fpunit_exec_to_writeback_fast_pipe_read_ack(0) = '1') and (not fpunit_exec_to_writeback_slow_pipe_needed))
				 or
			((fpunit_exec_to_writeback_slow_pipe_read_ack(0) = '1') and fpunit_exec_to_writeback_slow_pipe_needed);

	fpunit_exec_to_writeback_fast_pipe_read_req(0) <= fpunit_exec_to_writeback_pipe_write_ack(0)  when write_to_out else '0';
	fpunit_exec_to_writeback_slow_pipe_read_req(0) <= fpunit_exec_to_writeback_pipe_write_ack(0)  
						when (fpunit_exec_to_writeback_slow_pipe_needed and write_to_out) else '0';

	fpunit_exec_to_writeback_pipe_write_req(0) <= '1' when write_to_out else '0';
end very_simple;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;

library AjitCustom;
use AjitCustom.AjitCustomComponents.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

entity mul24_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    L : in  std_logic_vector(23 downto 0);
    R : in  std_logic_vector(23 downto 0);
    RESULT : out  std_logic_vector(47 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity mul24_Operator;
architecture mul24_Operator_arch of mul24_Operator is -- 
   signal start_req, start_ack, fin_req, fin_ack: std_logic;
   signal tag_in, tag_out: std_logic_vector(0 downto 0);
   signal umul_out, umul_out_reg: std_logic_vector(47 downto 0);
   signal update_ack_sig: boolean;

-- see comment above..
--##decl_synopsys_sync_set_reset##

begin
   tag_in(0) <= '0';
   update_ack <= update_ack_sig;

   p2l: Sample_Pulse_To_Level_Translate_Entity
		generic map(name => "mul24_Operator_p2l")
		port map (rL => sample_req, rR => start_req,
				aL => sample_ack, aR => start_ack,
					clk => clk, reset => reset);
   l2p: Level_To_Pulse_Translate_Entity
		generic map(name => "mul24_Operator_l2p")
		port map (rL => fin_req, rR => update_req,
				aL => fin_ack, aR => update_ack_sig, clk => clk, reset => reset);
				
   mul_inst: mul24
		generic map(tag_length => 1)
		port map( L => L, R => R,
				RESULT => umul_out,
				clk => clk, reset => reset,
				tag_in => tag_in , tag_out => tag_out,
				start_req => start_req, fin_req => fin_req,
				start_ack => start_ack, fin_ack => fin_ack);

   rrr: BypassRegister 
		generic map(data_width => umul_out'length, bypass => true)
		port map (clk => clk, reset => reset, din => umul_out, enable => update_ack_sig, q => RESULT);
			
end mul24_Operator_arch;


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library ahir;
use ahir.BaseComponents.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

entity mul24 is -- 
    generic (tag_length : integer);
    port ( -- 
      L : in  std_logic_vector(23 downto 0);
      R : in  std_logic_vector(23 downto 0);
      RESULT : out  std_logic_vector(47 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
end entity mul24;

architecture Struct of mul24 is
	signal uL : unsigned (23 downto 0);
	signal uR : unsigned (23 downto 0);	
	signal uRESULT: unsigned(47 downto 0);

	signal enable: std_logic;
	signal fin_ack_sig: bit;
-- see comment above..
--##decl_synopsys_sync_set_reset##
begin

   	fin_ack <= '1' when fin_ack_sig = '1' else '0';
	start_ack <= enable;

	uL <= to_unsigned(L);
	uR <= to_unsigned(R);
	uRESULT <= uL*uR;

	process(clk,reset)
	begin
		if(clk'event and clk = '1') then
		    if(enable = '1') then
			RESULT <= To_SLV(uRESULT);
		    end if;
		end if;
	end process;

	process(clk,reset, fin_req, start_req, fin_ack_sig)
		variable next_fin_ack_sig: bit;
		variable enable_var : std_logic;
	begin
		next_fin_ack_sig := fin_ack_sig;
		enable_var := '0';

		case fin_ack_sig is
			when '0' =>
				if(start_req = '1') then
					enable_var := '1';
					next_fin_ack_sig := '1';
				end if;
			when '1' =>
				if((fin_req = '1') and (start_req  = '1')) then
					enable_var := '1';
				elsif (fin_req = '1') then
					next_fin_ack_sig := '0';
				end if;
			when others => 
				null;
		end case;

		enable <= enable_var;

		if(clk'event and clk = '1') then
			if(reset = '1') then
				fin_ack_sig <= '0';
			else
				fin_ack_sig <= next_fin_ack_sig;
				if(enable_var = '1') then
					tag_out <= tag_in;
				end if;
			end if;
		end if;

	end process;
end Struct;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library ahir;
use ahir.BaseComponents.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

entity mul24_deterministic_pipeline_operator is -- 
    port ( -- 
      L : in  std_logic_vector(23 downto 0);
      R : in  std_logic_vector(23 downto 0);
      RESULT : out  std_logic_vector(47 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      enable: in std_logic;
      stall : in std_logic_vector(1 to 1)
    );
end entity mul24_deterministic_pipeline_operator;

architecture Struct of mul24_deterministic_pipeline_operator is
	signal uL : unsigned (23 downto 0);
	signal uR : unsigned (23 downto 0);	
	signal uRESULT: unsigned(47 downto 0);
-- see comment above..
--##decl_synopsys_sync_set_reset##
begin
	uL <= to_unsigned(L);
	uR <= to_unsigned(R);
	uRESULT <= uL*uR;

	process(clk,reset)
	begin
		if(clk'event and clk = '1') then
		    if ((enable = '1') and (stall(1) = '0')) then
			RESULT <= To_SLV(uRESULT);
		    end if;
		end if;
	end process;
end Struct;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;

library AjitCustom;
use AjitCustom.AjitCustomComponents.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

entity mul53_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    L : in  std_logic_vector(52 downto 0);
    R : in  std_logic_vector(52 downto 0);
    RESULT : out  std_logic_vector(105 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity mul53_Operator;
architecture mul53_Operator_arch of mul53_Operator is -- 
   signal start_req, start_ack, fin_req, fin_ack: std_logic;
   signal tag_in, tag_out: std_logic_vector(0 downto 0);
   signal umul_out, umul_out_reg: std_logic_vector(105 downto 0);
   signal update_ack_sig: boolean;

-- see comment above..
--##decl_synopsys_sync_set_reset##

begin
   tag_in(0) <= '0';
   update_ack <= update_ack_sig;

   p2l: Sample_Pulse_To_Level_Translate_Entity
		generic map(name => "mul53_Operator_p2l")
		port map (rL => sample_req, rR => start_req,
				aL => sample_ack, aR => start_ack,
					clk => clk, reset => reset);
   l2p: Level_To_Pulse_Translate_Entity
		generic map(name => "mul53_Operator_l2p")
		port map (rL => fin_req, rR => update_req,
				aL => fin_ack, aR => update_ack_sig, clk => clk, reset => reset);
				
   mul_inst: mul53
		generic map(tag_length => 1)
		port map( L => L, R => R,
				RESULT => umul_out,
				clk => clk, reset => reset,
				tag_in => tag_in , tag_out => tag_out,
				start_req => start_req, fin_req => fin_req,
				start_ack => start_ack, fin_ack => fin_ack);

   rrr: BypassRegister 
		generic map(data_width => umul_out'length, bypass => true)
		port map (clk => clk, reset => reset, din => umul_out, enable => update_ack_sig, q => RESULT);
			
end mul53_Operator_arch;


library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library ahir;
use ahir.BaseComponents.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

entity mul53 is -- 
    generic (tag_length : integer);
    port ( -- 
      L : in  std_logic_vector(52 downto 0);
      R : in  std_logic_vector(52 downto 0);
      RESULT : out  std_logic_vector(105 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
end entity mul53;

architecture Struct of mul53 is
	signal uL : unsigned (52 downto 0);
	signal uR : unsigned (52 downto 0);	
	signal uRESULT: unsigned(105 downto 0);

	signal enable: std_logic;
	signal fin_ack_sig: bit;
-- see comment above..
--##decl_synopsys_sync_set_reset##
begin

   	fin_ack <= '1' when fin_ack_sig = '1' else '0';
	start_ack <= enable;

	uL <= to_unsigned(L);
	uR <= to_unsigned(R);
	uRESULT <= uL*uR;

	process(clk,reset)
	begin
		if(clk'event and clk = '1') then
		    if(enable = '1') then
			RESULT <= To_SLV(uRESULT);
		    end if;
		end if;
	end process;

	process(clk,reset, fin_req, start_req, fin_ack_sig)
		variable next_fin_ack_sig: bit;
		variable enable_var : std_logic;
	begin
		next_fin_ack_sig := fin_ack_sig;
		enable_var := '0';

		case fin_ack_sig is
			when '0' =>
				if(start_req = '1') then
					enable_var := '1';
					next_fin_ack_sig := '1';
				end if;
			when '1' =>
				if((fin_req = '1') and (start_req  = '1')) then
					enable_var := '1';
				elsif (fin_req = '1') then
					next_fin_ack_sig := '0';
				end if;
			when others => 
				null;
		end case;

		enable <= enable_var;

		if(clk'event and clk = '1') then
			if(reset = '1') then
				fin_ack_sig <= '0';
			else
				fin_ack_sig <= next_fin_ack_sig;
				if(enable_var = '1') then
					tag_out <= tag_in;
				end if;
			end if;
		end if;

	end process;
end Struct;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library ahir;
use ahir.BaseComponents.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

entity mul53_deterministic_pipeline_operator is -- 
    port ( -- 
      L : in  std_logic_vector(52 downto 0);
      R : in  std_logic_vector(52 downto 0);
      RESULT : out  std_logic_vector(105 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      enable: in std_logic;
      stall : in std_logic_vector(1 to 1)
    );
end entity mul53_deterministic_pipeline_operator;

architecture Struct of mul53_deterministic_pipeline_operator is
	signal uL : unsigned (52 downto 0);
	signal uR : unsigned (52 downto 0);	
	signal uRESULT: unsigned(105 downto 0);
-- see comment above..
--##decl_synopsys_sync_set_reset##
begin
	uL <= to_unsigned(L);
	uR <= to_unsigned(R);
	uRESULT <= uL*uR;

	process(clk,reset)
	begin
		if(clk'event and clk = '1') then
		    if ((enable = '1') and (stall(1) = '0')) then
			RESULT <= To_SLV(uRESULT);
		    end if;
		end if;
	end process;
end Struct;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##

entity interrupt_stub_daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    INTR_LEVEL : in std_logic_vector(3 downto 0);
    ENV_to_CPU_irl_pipe_write_req : out  std_logic_vector(0 downto 0);
    ENV_to_CPU_irl_pipe_write_ack : in   std_logic_vector(0 downto 0);
    ENV_to_CPU_irl_pipe_write_data : out  std_logic_vector(7 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity interrupt_stub_daemon;
architecture interrupt_stub_daemon_arch of interrupt_stub_daemon is -- 
	signal INTR_LEVEL_d, INTR_LEVEL_dd : std_logic_vector(3 downto 0);
	signal counter: unsigned (1 downto 0);
	constant ZZZ4 : std_logic_vector(3 downto 0) := "0000";
-- see comment above..
--##decl_synopsys_sync_set_reset##
begin

	tag_out <= tag_in;

	start_ack <= '1';
	fin_ack <= '0';

	ENV_to_CPU_irl_pipe_write_data <=  ZZZ4 & INTR_LEVEL_dd;

	
	process(clk, reset)
	begin
		if(clk'event and clk = '1') then
			if(reset = '1') then
				ENV_to_CPU_irl_pipe_write_req(0) <= '0'; 
				counter <= (others => '0');
			else 
				ENV_to_CPU_irl_pipe_write_req(0) <= '1'; 
				counter <= counter + 1;
			end if;
		end if;
	end process;

	process(clk, reset, counter)
	begin
		if(clk'event and clk = '1') then
		   if(reset = '1') then
			INTR_LEVEL_d <= ZZZ4;
			INTR_LEVEL_dd <= ZZZ4;
		   elsif (counter = "11") then
			INTR_LEVEL_d <= INTR_LEVEL;
			INTR_LEVEL_dd <= INTR_LEVEL_d;
		   end if;
		end if;
	end process;

end interrupt_stub_daemon_arch;
-- IN NO EVENT SHALL THE CONTRIBUTORS OR COPYRIGHT HOLDERS BE LIABLE FOR
-- ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN ACTION OF CONTRACT,
-- TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN CONNECTION WITH THE
-- SOFTWARE OR THE USE OR OTHER DEALINGS WITH THE SOFTWARE.
------------------------------------------------------------------------------------------------
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.BaseComponents.all;

library AjitCustom;
use AjitCustom.AjitCustomComponents.all;

entity iu_umul32_Operator is -- 
    port ( -- 
      L : in  std_logic_vector(31 downto 0);
      R : in  std_logic_vector(31 downto 0);
      ret_val_x_x : out  std_logic_vector(63 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      sample_req : in Boolean;
      sample_ack : out Boolean;
      update_req : in Boolean;
      update_ack   : out Boolean
    );
end entity iu_umul32_Operator;

architecture Struct of iu_umul32_Operator is
   signal start_req, start_ack, fin_req, fin_ack: std_logic;
   signal tag_in, tag_out: std_logic_vector(0 downto 0);
   signal umul_out, umul_out_reg: std_logic_vector(63 downto 0);
   signal update_ack_sig: boolean;
begin
   tag_in(0) <= '0';
   update_ack <= update_ack_sig;

   p2l: Sample_Pulse_To_Level_Translate_Entity
		generic map(name => "iu_umul32_Operator_p2l")
		port map (rL => sample_req, rR => start_req,
				aL => sample_ack, aR => start_ack,
					clk => clk, reset => reset);
   l2p: Level_To_Pulse_Translate_Entity
		generic map(name => "iu_umul32_Operator_l2p")
		port map (rL => fin_req, rR => update_req,
				aL => fin_ack, aR => update_ack_sig, clk => clk, reset => reset);
				
   mul_inst: iu_umul32
		generic map(tag_length => 1)
		port map( L => L, R => R,
				RESULT => umul_out,
				clk => clk, reset => reset,
				tag_in => tag_in , tag_out => tag_out,
				start_req => start_req, fin_req => fin_req,
				start_ack => start_ack, fin_ack => fin_ack);

   rrr: BypassRegister 
		generic map(data_width => umul_out'length, bypass => true)
		port map (clk => clk, reset => reset, din => umul_out, enable => update_ack_sig, q => ret_val_x_x);
			
end Struct;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.BaseComponents.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;

entity iu_umul32 is -- 
    generic (tag_length : integer);
    port ( -- 
      L : in  std_logic_vector(31 downto 0);
      R : in  std_logic_vector(31 downto 0);
      RESULT : out  std_logic_vector(63 downto 0);
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic;
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) -- 
    );
end entity iu_umul32;

architecture Struct of iu_umul32 is
	signal uL : unsigned (31 downto 0);
	signal uR : unsigned (31 downto 0);	
	signal uRESULT: unsigned(63 downto 0);

	signal enable: std_logic;
	signal fin_ack_sig: bit;
begin

   	fin_ack <= '1' when fin_ack_sig = '1' else '0';
	start_ack <= enable;

	uL <= to_unsigned(L);
	uR <= to_unsigned(R);
	uRESULT <= uL*uR;

	process(clk,reset)
	begin
		if(clk'event and clk = '1') then
		    if(enable = '1') then
			RESULT <= To_SLV(uRESULT);
		    end if;
		end if;
	end process;

	process(clk,reset, fin_req, start_req, fin_ack_sig)
		variable next_fin_ack_sig: bit;
		variable enable_var : std_logic;
	begin
		next_fin_ack_sig := fin_ack_sig;
		enable_var := '0';

		case fin_ack_sig is
			when '0' =>
				if(start_req = '1') then
					enable_var := '1';
					next_fin_ack_sig := '1';
				end if;
			when '1' =>
				if((fin_req = '1') and (start_req  = '1')) then
					enable_var := '1';
				elsif (fin_req = '1') then
					next_fin_ack_sig := '0';
				end if;
			when others => 
				null;
		end case;

		enable <= enable_var;

		if(clk'event and clk = '1') then
			if(reset = '1') then
				fin_ack_sig <= '0';
			else
				fin_ack_sig <= next_fin_ack_sig;
				if(enable_var = '1') then
					tag_out <= tag_in;
				end if;
			end if;
		end if;

	end process;
end Struct;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.BaseComponents.all;
use ahir.Subprograms.all;
use ahir.Utilities.all;

entity iu_umul32_Volatile is -- 
    port ( -- 
      L : in  std_logic_vector(31 downto 0);
      R : in  std_logic_vector(31 downto 0);
      ret_val_x_x : out  std_logic_vector(63 downto 0)
    );
end entity iu_umul32_Volatile;

architecture Struct of iu_umul32_Volatile is
	signal uL : unsigned (31 downto 0);
	signal uR : unsigned (31 downto 0);	
	signal uRESULT: unsigned(63 downto 0);
begin
	uL <= to_unsigned(L);
	uR <= to_unsigned(R);
	uRESULT <= uL*uR;
	ret_val_x_x <= To_SLV(uRESULT);
end Struct;

library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
entity analyze_dcache_response_VVP is -- 
  port ( -- 
    addr : in  std_logic_vector(31 downto 0);
    dcache_response : in  std_logic_vector(71 downto 0);
    is_load : in  std_logic_vector(0 downto 0);
    is_store : in  std_logic_vector(0 downto 0);
    signed_type : in  std_logic_vector(0 downto 0);
    unsigned_type : in  std_logic_vector(0 downto 0);
    byte : in  std_logic_vector(0 downto 0);
    half_word : in  std_logic_vector(0 downto 0);
    word : in  std_logic_vector(0 downto 0);
    double_word : in  std_logic_vector(0 downto 0);
    dout_h : out  std_logic_vector(31 downto 0);
    dout_l : out  std_logic_vector(31 downto 0);
    data_access_exception : out  std_logic_vector(0 downto 0);
    data_access_error : out  std_logic_vector(0 downto 0);
    dcache_hit : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity analyze_dcache_response_VVP;
architecture analyze_dcache_response_VVP_arch of analyze_dcache_response_VVP is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(112-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal addr_buffer :  std_logic_vector(31 downto 0);
  signal dcache_response_buffer :  std_logic_vector(71 downto 0);
  signal is_load_buffer :  std_logic_vector(0 downto 0);
  signal is_store_buffer :  std_logic_vector(0 downto 0);
  signal signed_type_buffer :  std_logic_vector(0 downto 0);
  signal unsigned_type_buffer :  std_logic_vector(0 downto 0);
  signal byte_buffer :  std_logic_vector(0 downto 0);
  signal half_word_buffer :  std_logic_vector(0 downto 0);
  signal word_buffer :  std_logic_vector(0 downto 0);
  signal double_word_buffer :  std_logic_vector(0 downto 0);
  -- output port buffer signals
  signal dout_h_buffer :  std_logic_vector(31 downto 0);
  signal dout_l_buffer :  std_logic_vector(31 downto 0);
  signal data_access_exception_buffer :  std_logic_vector(0 downto 0);
  signal data_access_error_buffer :  std_logic_vector(0 downto 0);
  signal dcache_hit_buffer :  std_logic_vector(0 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  addr_buffer <= addr;
  dcache_response_buffer <= dcache_response;
  is_load_buffer <= is_load;
  is_store_buffer <= is_store;
  signed_type_buffer <= signed_type;
  unsigned_type_buffer <= unsigned_type;
  byte_buffer <= byte;
  half_word_buffer <= half_word;
  word_buffer <= word;
  double_word_buffer <= double_word;
  -- output handling  -------------------------------------------------------
  dout_h <= dout_h_buffer;
  dout_l <= dout_l_buffer;
  data_access_exception <= data_access_exception_buffer;
  data_access_error <= data_access_error_buffer;
  dcache_hit <= dcache_hit_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u32_u1_1216_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1226_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1233_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1241_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1248_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1259_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_1266_wire : std_logic_vector(0 downto 0);
    signal MUX_1230_wire : std_logic_vector(7 downto 0);
    signal MUX_1237_wire : std_logic_vector(7 downto 0);
    signal MUX_1245_wire : std_logic_vector(7 downto 0);
    signal MUX_1252_wire : std_logic_vector(7 downto 0);
    signal MUX_1263_wire : std_logic_vector(15 downto 0);
    signal MUX_1270_wire : std_logic_vector(15 downto 0);
    signal MUX_1287_wire : std_logic_vector(31 downto 0);
    signal MUX_1289_wire : std_logic_vector(31 downto 0);
    signal MUX_1299_wire : std_logic_vector(31 downto 0);
    signal MUX_1301_wire : std_logic_vector(31 downto 0);
    signal MUX_1308_wire : std_logic_vector(31 downto 0);
    signal OR_u1_u1_1217_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1305_wire : std_logic_vector(0 downto 0);
    signal OR_u32_u32_1302_wire : std_logic_vector(31 downto 0);
    signal OR_u8_u8_1238_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_1253_wire : std_logic_vector(7 downto 0);
    signal a10_1207 : std_logic_vector(1 downto 0);
    signal dcache_mae_1184 : std_logic_vector(7 downto 0);
    signal ext_byte_1255 : std_logic_vector(7 downto 0);
    signal ext_half_word_1272 : std_logic_vector(15 downto 0);
    signal konst_1191_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1196_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1201_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1215_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1225_wire_constant : std_logic_vector(1 downto 0);
    signal konst_1229_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1232_wire_constant : std_logic_vector(1 downto 0);
    signal konst_1236_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1240_wire_constant : std_logic_vector(1 downto 0);
    signal konst_1244_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1247_wire_constant : std_logic_vector(1 downto 0);
    signal konst_1251_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1258_wire_constant : std_logic_vector(1 downto 0);
    signal konst_1262_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1265_wire_constant : std_logic_vector(1 downto 0);
    signal konst_1269_wire_constant : std_logic_vector(15 downto 0);
    signal konst_1288_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1300_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1307_wire_constant : std_logic_vector(31 downto 0);
    signal loaded_high_word_1211 : std_logic_vector(31 downto 0);
    signal loaded_low_word_1222 : std_logic_vector(31 downto 0);
    signal loaded_word_1188 : std_logic_vector(63 downto 0);
    signal slice_1219_wire : std_logic_vector(31 downto 0);
    signal slice_1228_wire : std_logic_vector(7 downto 0);
    signal slice_1235_wire : std_logic_vector(7 downto 0);
    signal slice_1243_wire : std_logic_vector(7 downto 0);
    signal slice_1250_wire : std_logic_vector(7 downto 0);
    signal slice_1261_wire : std_logic_vector(15 downto 0);
    signal slice_1268_wire : std_logic_vector(15 downto 0);
    signal type_cast_1282_wire : std_logic_vector(7 downto 0);
    signal type_cast_1283_wire : std_logic_vector(31 downto 0);
    signal type_cast_1284_wire : std_logic_vector(31 downto 0);
    signal type_cast_1286_wire : std_logic_vector(31 downto 0);
    signal type_cast_1294_wire : std_logic_vector(15 downto 0);
    signal type_cast_1295_wire : std_logic_vector(31 downto 0);
    signal type_cast_1296_wire : std_logic_vector(31 downto 0);
    signal type_cast_1298_wire : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    konst_1191_wire_constant <= "00000000";
    konst_1196_wire_constant <= "00000001";
    konst_1201_wire_constant <= "00000010";
    konst_1215_wire_constant <= "00000000000000000000000000000010";
    konst_1225_wire_constant <= "00";
    konst_1229_wire_constant <= "00000000";
    konst_1232_wire_constant <= "01";
    konst_1236_wire_constant <= "00000000";
    konst_1240_wire_constant <= "10";
    konst_1244_wire_constant <= "00000000";
    konst_1247_wire_constant <= "11";
    konst_1251_wire_constant <= "00000000";
    konst_1258_wire_constant <= "00";
    konst_1262_wire_constant <= "0000000000000000";
    konst_1265_wire_constant <= "10";
    konst_1269_wire_constant <= "0000000000000000";
    konst_1288_wire_constant <= "00000000000000000000000000000000";
    konst_1300_wire_constant <= "00000000000000000000000000000000";
    konst_1307_wire_constant <= "00000000000000000000000000000000";
    -- flow-through select operator MUX_1221_inst
    loaded_low_word_1222 <= slice_1219_wire when (OR_u1_u1_1217_wire(0) /=  '0') else loaded_high_word_1211;
    -- flow-through select operator MUX_1230_inst
    MUX_1230_wire <= slice_1228_wire when (EQ_u2_u1_1226_wire(0) /=  '0') else konst_1229_wire_constant;
    -- flow-through select operator MUX_1237_inst
    MUX_1237_wire <= slice_1235_wire when (EQ_u2_u1_1233_wire(0) /=  '0') else konst_1236_wire_constant;
    -- flow-through select operator MUX_1245_inst
    MUX_1245_wire <= slice_1243_wire when (EQ_u2_u1_1241_wire(0) /=  '0') else konst_1244_wire_constant;
    -- flow-through select operator MUX_1252_inst
    MUX_1252_wire <= slice_1250_wire when (EQ_u2_u1_1248_wire(0) /=  '0') else konst_1251_wire_constant;
    -- flow-through select operator MUX_1263_inst
    MUX_1263_wire <= slice_1261_wire when (EQ_u2_u1_1259_wire(0) /=  '0') else konst_1262_wire_constant;
    -- flow-through select operator MUX_1270_inst
    MUX_1270_wire <= slice_1268_wire when (EQ_u2_u1_1266_wire(0) /=  '0') else konst_1269_wire_constant;
    -- flow-through select operator MUX_1287_inst
    MUX_1287_wire <= type_cast_1284_wire when (signed_type_buffer(0) /=  '0') else type_cast_1286_wire;
    -- flow-through select operator MUX_1289_inst
    MUX_1289_wire <= MUX_1287_wire when (byte_buffer(0) /=  '0') else konst_1288_wire_constant;
    -- flow-through select operator MUX_1299_inst
    MUX_1299_wire <= type_cast_1296_wire when (signed_type_buffer(0) /=  '0') else type_cast_1298_wire;
    -- flow-through select operator MUX_1301_inst
    MUX_1301_wire <= MUX_1299_wire when (half_word_buffer(0) /=  '0') else konst_1300_wire_constant;
    -- flow-through select operator MUX_1308_inst
    MUX_1308_wire <= loaded_low_word_1222 when (OR_u1_u1_1305_wire(0) /=  '0') else konst_1307_wire_constant;
    -- flow-through slice operator slice_1183_inst
    dcache_mae_1184 <= dcache_response_buffer(71 downto 64);
    -- flow-through slice operator slice_1187_inst
    loaded_word_1188 <= dcache_response_buffer(63 downto 0);
    -- flow-through slice operator slice_1206_inst
    a10_1207 <= addr_buffer(1 downto 0);
    -- flow-through slice operator slice_1210_inst
    loaded_high_word_1211 <= loaded_word_1188(63 downto 32);
    -- flow-through slice operator slice_1219_inst
    slice_1219_wire <= loaded_word_1188(31 downto 0);
    -- flow-through slice operator slice_1228_inst
    slice_1228_wire <= loaded_low_word_1222(31 downto 24);
    -- flow-through slice operator slice_1235_inst
    slice_1235_wire <= loaded_low_word_1222(23 downto 16);
    -- flow-through slice operator slice_1243_inst
    slice_1243_wire <= loaded_low_word_1222(15 downto 8);
    -- flow-through slice operator slice_1250_inst
    slice_1250_wire <= loaded_low_word_1222(7 downto 0);
    -- flow-through slice operator slice_1261_inst
    slice_1261_wire <= loaded_low_word_1222(31 downto 16);
    -- flow-through slice operator slice_1268_inst
    slice_1268_wire <= loaded_low_word_1222(15 downto 0);
    -- interlock W_dout_h_1273_inst
    process(loaded_high_word_1211) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := loaded_high_word_1211(31 downto 0);
      dout_h_buffer <= tmp_var; -- 
    end process;
    -- interlock type_cast_1282_inst
    process(ext_byte_1255) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ext_byte_1255(7 downto 0);
      type_cast_1282_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1284_inst
    process(type_cast_1283_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := type_cast_1283_wire(31 downto 0);
      type_cast_1284_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1286_inst
    process(ext_byte_1255) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := ext_byte_1255(7 downto 0);
      type_cast_1286_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1294_inst
    process(ext_half_word_1272) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := ext_half_word_1272(15 downto 0);
      type_cast_1294_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1296_inst
    process(type_cast_1295_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := type_cast_1295_wire(31 downto 0);
      type_cast_1296_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1298_inst
    process(ext_half_word_1272) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 15 downto 0) := ext_half_word_1272(15 downto 0);
      type_cast_1298_wire <= tmp_var; -- 
    end process;
    -- binary operator BITSEL_u32_u1_1216_inst
    process(addr_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(addr_buffer, konst_1215_wire_constant, tmp_var);
      BITSEL_u32_u1_1216_wire <= tmp_var; --
    end process;
    -- binary operator BITSEL_u8_u1_1192_inst
    process(dcache_mae_1184) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(dcache_mae_1184, konst_1191_wire_constant, tmp_var);
      data_access_exception_buffer <= tmp_var; --
    end process;
    -- binary operator BITSEL_u8_u1_1197_inst
    process(dcache_mae_1184) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(dcache_mae_1184, konst_1196_wire_constant, tmp_var);
      data_access_error_buffer <= tmp_var; --
    end process;
    -- binary operator BITSEL_u8_u1_1202_inst
    process(dcache_mae_1184) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(dcache_mae_1184, konst_1201_wire_constant, tmp_var);
      dcache_hit_buffer <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1226_inst
    process(a10_1207) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(a10_1207, konst_1225_wire_constant, tmp_var);
      EQ_u2_u1_1226_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1233_inst
    process(a10_1207) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(a10_1207, konst_1232_wire_constant, tmp_var);
      EQ_u2_u1_1233_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1241_inst
    process(a10_1207) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(a10_1207, konst_1240_wire_constant, tmp_var);
      EQ_u2_u1_1241_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1248_inst
    process(a10_1207) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(a10_1207, konst_1247_wire_constant, tmp_var);
      EQ_u2_u1_1248_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1259_inst
    process(a10_1207) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(a10_1207, konst_1258_wire_constant, tmp_var);
      EQ_u2_u1_1259_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_1266_inst
    process(a10_1207) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(a10_1207, konst_1265_wire_constant, tmp_var);
      EQ_u2_u1_1266_wire <= tmp_var; --
    end process;
    -- binary operator OR_u16_u16_1271_inst
    process(MUX_1263_wire, MUX_1270_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1263_wire, MUX_1270_wire, tmp_var);
      ext_half_word_1272 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1217_inst
    process(double_word_buffer, BITSEL_u32_u1_1216_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(double_word_buffer, BITSEL_u32_u1_1216_wire, tmp_var);
      OR_u1_u1_1217_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1305_inst
    process(word_buffer, double_word_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(word_buffer, double_word_buffer, tmp_var);
      OR_u1_u1_1305_wire <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1302_inst
    process(MUX_1289_wire, MUX_1301_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1289_wire, MUX_1301_wire, tmp_var);
      OR_u32_u32_1302_wire <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_1309_inst
    process(OR_u32_u32_1302_wire, MUX_1308_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u32_u32_1302_wire, MUX_1308_wire, tmp_var);
      dout_l_buffer <= tmp_var; --
    end process;
    -- binary operator OR_u8_u8_1238_inst
    process(MUX_1230_wire, MUX_1237_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1230_wire, MUX_1237_wire, tmp_var);
      OR_u8_u8_1238_wire <= tmp_var; --
    end process;
    -- binary operator OR_u8_u8_1253_inst
    process(MUX_1245_wire, MUX_1252_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1245_wire, MUX_1252_wire, tmp_var);
      OR_u8_u8_1253_wire <= tmp_var; --
    end process;
    -- binary operator OR_u8_u8_1254_inst
    process(OR_u8_u8_1238_wire, OR_u8_u8_1253_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u8_u8_1238_wire, OR_u8_u8_1253_wire, tmp_var);
      ext_byte_1255 <= tmp_var; --
    end process;
    -- unary operator type_cast_1283_inst
    process(type_cast_1282_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", type_cast_1282_wire, tmp_var);
      type_cast_1283_wire <= tmp_var; -- 
    end process;
    -- unary operator type_cast_1295_inst
    process(type_cast_1294_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntToApIntSigned", type_cast_1294_wire, tmp_var);
      type_cast_1295_wire <= tmp_var; -- 
    end process;
    -- 
  end Block; -- data_path
  -- 
end analyze_dcache_response_VVP_arch;

library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
entity decode_routing_control_info_VVP is -- 
  port ( -- 
    control_info : in  std_logic_vector(96 downto 0);
    read_simple : out  std_logic_vector(0 downto 0);
    read_messy : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity decode_routing_control_info_VVP;
architecture decode_routing_control_info_VVP_arch of decode_routing_control_info_VVP is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(97-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal control_info_buffer :  std_logic_vector(96 downto 0);
  -- output port buffer signals
  signal read_simple_buffer :  std_logic_vector(0 downto 0);
  signal read_messy_buffer :  std_logic_vector(0 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  control_info_buffer <= control_info;
  -- output handling  -------------------------------------------------------
  read_simple <= read_simple_buffer;
  read_messy <= read_messy_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal addr_4166 : std_logic_vector(31 downto 0);
    signal byte_4134 : std_logic_vector(0 downto 0);
    signal dbg_wp_read_hit_4154 : std_logic_vector(0 downto 0);
    signal dbg_wp_reg_id_4150 : std_logic_vector(1 downto 0);
    signal dbg_wp_write_hit_4158 : std_logic_vector(0 downto 0);
    signal double_word_4146 : std_logic_vector(0 downto 0);
    signal early_ls_traps_4114 : std_logic_vector(2 downto 0);
    signal half_word_4138 : std_logic_vector(0 downto 0);
    signal is_load_4118 : std_logic_vector(0 downto 0);
    signal is_store_4122 : std_logic_vector(0 downto 0);
    signal signed_type_4126 : std_logic_vector(0 downto 0);
    signal simple_store_signature_4162 : std_logic_vector(31 downto 0);
    signal slot_id_4086 : std_logic_vector(5 downto 0);
    signal stream_id_4082 : std_logic_vector(1 downto 0);
    signal thread_id_4078 : std_logic_vector(3 downto 0);
    signal to_cu_4098 : std_logic_vector(0 downto 0);
    signal to_fu_4094 : std_logic_vector(0 downto 0);
    signal to_iu_4090 : std_logic_vector(0 downto 0);
    signal to_retire_4102 : std_logic_vector(0 downto 0);
    signal unsigned_type_4130 : std_logic_vector(0 downto 0);
    signal word_4142 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    -- flow-through slice operator slice_4077_inst
    thread_id_4078 <= control_info_buffer(96 downto 93);
    -- flow-through slice operator slice_4081_inst
    stream_id_4082 <= control_info_buffer(92 downto 91);
    -- flow-through slice operator slice_4085_inst
    slot_id_4086 <= control_info_buffer(90 downto 85);
    -- flow-through slice operator slice_4089_inst
    to_iu_4090 <= control_info_buffer(84 downto 84);
    -- flow-through slice operator slice_4093_inst
    to_fu_4094 <= control_info_buffer(83 downto 83);
    -- flow-through slice operator slice_4097_inst
    to_cu_4098 <= control_info_buffer(82 downto 82);
    -- flow-through slice operator slice_4101_inst
    to_retire_4102 <= control_info_buffer(81 downto 81);
    -- flow-through slice operator slice_4105_inst
    read_messy_buffer <= control_info_buffer(80 downto 80);
    -- flow-through slice operator slice_4109_inst
    read_simple_buffer <= control_info_buffer(79 downto 79);
    -- flow-through slice operator slice_4113_inst
    early_ls_traps_4114 <= control_info_buffer(78 downto 76);
    -- flow-through slice operator slice_4117_inst
    is_load_4118 <= control_info_buffer(75 downto 75);
    -- flow-through slice operator slice_4121_inst
    is_store_4122 <= control_info_buffer(74 downto 74);
    -- flow-through slice operator slice_4125_inst
    signed_type_4126 <= control_info_buffer(73 downto 73);
    -- flow-through slice operator slice_4129_inst
    unsigned_type_4130 <= control_info_buffer(72 downto 72);
    -- flow-through slice operator slice_4133_inst
    byte_4134 <= control_info_buffer(71 downto 71);
    -- flow-through slice operator slice_4137_inst
    half_word_4138 <= control_info_buffer(70 downto 70);
    -- flow-through slice operator slice_4141_inst
    word_4142 <= control_info_buffer(69 downto 69);
    -- flow-through slice operator slice_4145_inst
    double_word_4146 <= control_info_buffer(68 downto 68);
    -- flow-through slice operator slice_4149_inst
    dbg_wp_reg_id_4150 <= control_info_buffer(67 downto 66);
    -- flow-through slice operator slice_4153_inst
    dbg_wp_read_hit_4154 <= control_info_buffer(65 downto 65);
    -- flow-through slice operator slice_4157_inst
    dbg_wp_write_hit_4158 <= control_info_buffer(64 downto 64);
    -- flow-through slice operator slice_4161_inst
    simple_store_signature_4162 <= control_info_buffer(63 downto 32);
    -- flow-through slice operator slice_4165_inst
    addr_4166 <= control_info_buffer(31 downto 0);
    -- 
  end Block; -- data_path
  -- 
end decode_routing_control_info_VVP_arch;


library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
entity loadstore_router_core_VVP is -- 
  port ( -- 
    control_info : in  std_logic_vector(96 downto 0);
    simple_info : in  std_logic_vector(71 downto 0);
    messy_info : in  std_logic_vector(97 downto 0);
    to_iu : out  std_logic_vector(0 downto 0);
    to_fu : out  std_logic_vector(0 downto 0);
    to_cu : out  std_logic_vector(0 downto 0);
    to_retire : out  std_logic_vector(0 downto 0);
    to_iu_fu_data : out  std_logic_vector(77 downto 0);
    to_cu_data : out  std_logic_vector(13 downto 0);
    data_to_iretire : out  std_logic_vector(53 downto 0)-- 
  );
  -- 
end entity loadstore_router_core_VVP;
architecture loadstore_router_core_VVP_arch of loadstore_router_core_VVP is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(267-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal control_info_buffer :  std_logic_vector(96 downto 0);
  signal simple_info_buffer :  std_logic_vector(71 downto 0);
  signal messy_info_buffer :  std_logic_vector(97 downto 0);
  -- output port buffer signals
  signal to_iu_buffer :  std_logic_vector(0 downto 0);
  signal to_fu_buffer :  std_logic_vector(0 downto 0);
  signal to_cu_buffer :  std_logic_vector(0 downto 0);
  signal to_retire_buffer :  std_logic_vector(0 downto 0);
  signal to_iu_fu_data_buffer :  std_logic_vector(77 downto 0);
  signal to_cu_data_buffer :  std_logic_vector(13 downto 0);
  signal data_to_iretire_buffer :  std_logic_vector(53 downto 0);
  -- volatile/operator module components. 
  component analyze_dcache_response_VVP is -- 
    port ( -- 
      addr : in  std_logic_vector(31 downto 0);
      dcache_response : in  std_logic_vector(71 downto 0);
      is_load : in  std_logic_vector(0 downto 0);
      is_store : in  std_logic_vector(0 downto 0);
      signed_type : in  std_logic_vector(0 downto 0);
      unsigned_type : in  std_logic_vector(0 downto 0);
      byte : in  std_logic_vector(0 downto 0);
      half_word : in  std_logic_vector(0 downto 0);
      word : in  std_logic_vector(0 downto 0);
      double_word : in  std_logic_vector(0 downto 0);
      dout_h : out  std_logic_vector(31 downto 0);
      dout_l : out  std_logic_vector(31 downto 0);
      data_access_exception : out  std_logic_vector(0 downto 0);
      data_access_error : out  std_logic_vector(0 downto 0);
      dcache_hit : out  std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component; 
  -- 
begin --  
  -- input handling ------------------------------------------------
  control_info_buffer <= control_info;
  simple_info_buffer <= simple_info;
  messy_info_buffer <= messy_info;
  -- output handling  -------------------------------------------------------
  to_iu <= to_iu_buffer;
  to_fu <= to_fu_buffer;
  to_cu <= to_cu_buffer;
  to_retire <= to_retire_buffer;
  to_iu_fu_data <= to_iu_fu_data_buffer;
  to_cu_data <= to_cu_data_buffer;
  data_to_iretire <= data_to_iretire_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_9626_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_9629_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_9635_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_9638_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u13_u16_9771_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u1_u2_9700_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_9768_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_9774_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_9779_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u33_9687_wire : std_logic_vector(32 downto 0);
    signal CONCAT_u2_u34_9781_wire : std_logic_vector(33 downto 0);
    signal CONCAT_u2_u3_9746_wire : std_logic_vector(2 downto 0);
    signal CONCAT_u2_u3_9770_wire : std_logic_vector(2 downto 0);
    signal CONCAT_u2_u4_9776_wire : std_logic_vector(3 downto 0);
    signal CONCAT_u33_u65_9689_wire : std_logic_vector(64 downto 0);
    signal CONCAT_u3_u32_9749_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u4_u38_9782_wire : std_logic_vector(37 downto 0);
    signal CONCAT_u4_u6_9680_wire : std_logic_vector(5 downto 0);
    signal CONCAT_u4_u6_9695_wire : std_logic_vector(5 downto 0);
    signal CONCAT_u4_u6_9761_wire : std_logic_vector(5 downto 0);
    signal CONCAT_u6_u12_9697_wire : std_logic_vector(11 downto 0);
    signal CONCAT_u6_u13_9684_wire : std_logic_vector(12 downto 0);
    signal CONCAT_u6_u13_9765_wire : std_logic_vector(12 downto 0);
    signal CONCAT_u6_u7_9683_wire : std_logic_vector(6 downto 0);
    signal CONCAT_u6_u7_9764_wire : std_logic_vector(6 downto 0);
    signal MUX_9659_wire : std_logic_vector(31 downto 0);
    signal MUX_9663_wire : std_logic_vector(31 downto 0);
    signal MUX_9670_wire : std_logic_vector(31 downto 0);
    signal MUX_9674_wire : std_logic_vector(31 downto 0);
    signal MUX_9751_wire : std_logic_vector(31 downto 0);
    signal MUX_9755_wire : std_logic_vector(31 downto 0);
    signal NEQ_u3_u1_9644_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_9646_wire : std_logic_vector(0 downto 0);
    signal addr_9579 : std_logic_vector(31 downto 0);
    signal byte_9547 : std_logic_vector(0 downto 0);
    signal data_access_error_9640 : std_logic_vector(0 downto 0);
    signal data_access_exception_9631 : std_logic_vector(0 downto 0);
    signal dbg_wp_hit_9654 : std_logic_vector(0 downto 0);
    signal dbg_wp_read_hit_9567 : std_logic_vector(0 downto 0);
    signal dbg_wp_reg_id_9563 : std_logic_vector(1 downto 0);
    signal dbg_wp_write_hit_9571 : std_logic_vector(0 downto 0);
    signal double_word_9559 : std_logic_vector(0 downto 0);
    signal dout_h_9665 : std_logic_vector(31 downto 0);
    signal dout_l_9676 : std_logic_vector(31 downto 0);
    signal early_ls_traps_9527 : std_logic_vector(2 downto 0);
    signal half_word_9551 : std_logic_vector(0 downto 0);
    signal illegal_instr_trap_9736 : std_logic_vector(0 downto 0);
    signal is_load_9531 : std_logic_vector(0 downto 0);
    signal is_store_9535 : std_logic_vector(0 downto 0);
    signal konst_9643_wire_constant : std_logic_vector(2 downto 0);
    signal konst_9658_wire_constant : std_logic_vector(31 downto 0);
    signal konst_9662_wire_constant : std_logic_vector(31 downto 0);
    signal konst_9669_wire_constant : std_logic_vector(31 downto 0);
    signal konst_9673_wire_constant : std_logic_vector(31 downto 0);
    signal konst_9750_wire_constant : std_logic_vector(31 downto 0);
    signal konst_9754_wire_constant : std_logic_vector(31 downto 0);
    signal late_load_store_trap_9649 : std_logic_vector(0 downto 0);
    signal mem_address_not_aligned_trap_9740 : std_logic_vector(0 downto 0);
    signal messy_dout_h_9595 : std_logic_vector(31 downto 0);
    signal messy_dout_l_9599 : std_logic_vector(31 downto 0);
    signal messy_error_9587 : std_logic_vector(0 downto 0);
    signal messy_store_signature_9591 : std_logic_vector(31 downto 0);
    signal messy_trap_9583 : std_logic_vector(0 downto 0);
    signal privileged_instr_trap_9732 : std_logic_vector(0 downto 0);
    signal read_messy_9519 : std_logic_vector(0 downto 0);
    signal read_simple_9523 : std_logic_vector(0 downto 0);
    signal signed_type_9539 : std_logic_vector(0 downto 0);
    signal simple_data_access_error_9615 : std_logic_vector(0 downto 0);
    signal simple_data_access_exception_9615 : std_logic_vector(0 downto 0);
    signal simple_dcache_hit_9615 : std_logic_vector(0 downto 0);
    signal simple_dout_h_9615 : std_logic_vector(31 downto 0);
    signal simple_dout_l_9615 : std_logic_vector(31 downto 0);
    signal simple_store_signature_9575 : std_logic_vector(31 downto 0);
    signal slice_9744_wire : std_logic_vector(1 downto 0);
    signal slice_9748_wire : std_logic_vector(28 downto 0);
    signal slot_id_9499 : std_logic_vector(5 downto 0);
    signal store_signature_9757 : std_logic_vector(31 downto 0);
    signal stream_id_9495 : std_logic_vector(1 downto 0);
    signal thread_id_9491 : std_logic_vector(3 downto 0);
    signal unsigned_type_9543 : std_logic_vector(0 downto 0);
    signal word_9555 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    konst_9643_wire_constant <= "000";
    konst_9658_wire_constant <= "00000000000000000000000000000000";
    konst_9662_wire_constant <= "00000000000000000000000000000000";
    konst_9669_wire_constant <= "00000000000000000000000000000000";
    konst_9673_wire_constant <= "00000000000000000000000000000000";
    konst_9750_wire_constant <= "00000000000000000000000000000000";
    konst_9754_wire_constant <= "00000000000000000000000000000000";
    -- flow-through select operator MUX_9659_inst
    MUX_9659_wire <= simple_dout_h_9615 when (read_simple_9523(0) /=  '0') else konst_9658_wire_constant;
    -- flow-through select operator MUX_9663_inst
    MUX_9663_wire <= messy_dout_h_9595 when (read_messy_9519(0) /=  '0') else konst_9662_wire_constant;
    -- flow-through select operator MUX_9670_inst
    MUX_9670_wire <= simple_dout_l_9615 when (read_simple_9523(0) /=  '0') else konst_9669_wire_constant;
    -- flow-through select operator MUX_9674_inst
    MUX_9674_wire <= messy_dout_l_9599 when (read_messy_9519(0) /=  '0') else konst_9673_wire_constant;
    -- flow-through select operator MUX_9751_inst
    MUX_9751_wire <= CONCAT_u3_u32_9749_wire when (read_simple_9523(0) /=  '0') else konst_9750_wire_constant;
    -- flow-through select operator MUX_9755_inst
    MUX_9755_wire <= messy_store_signature_9591 when (read_messy_9519(0) /=  '0') else konst_9754_wire_constant;
    -- flow-through slice operator slice_9490_inst
    thread_id_9491 <= control_info_buffer(96 downto 93);
    -- flow-through slice operator slice_9494_inst
    stream_id_9495 <= control_info_buffer(92 downto 91);
    -- flow-through slice operator slice_9498_inst
    slot_id_9499 <= control_info_buffer(90 downto 85);
    -- flow-through slice operator slice_9502_inst
    to_iu_buffer <= control_info_buffer(84 downto 84);
    -- flow-through slice operator slice_9506_inst
    to_fu_buffer <= control_info_buffer(83 downto 83);
    -- flow-through slice operator slice_9510_inst
    to_cu_buffer <= control_info_buffer(82 downto 82);
    -- flow-through slice operator slice_9514_inst
    to_retire_buffer <= control_info_buffer(81 downto 81);
    -- flow-through slice operator slice_9518_inst
    read_messy_9519 <= control_info_buffer(80 downto 80);
    -- flow-through slice operator slice_9522_inst
    read_simple_9523 <= control_info_buffer(79 downto 79);
    -- flow-through slice operator slice_9526_inst
    early_ls_traps_9527 <= control_info_buffer(78 downto 76);
    -- flow-through slice operator slice_9530_inst
    is_load_9531 <= control_info_buffer(75 downto 75);
    -- flow-through slice operator slice_9534_inst
    is_store_9535 <= control_info_buffer(74 downto 74);
    -- flow-through slice operator slice_9538_inst
    signed_type_9539 <= control_info_buffer(73 downto 73);
    -- flow-through slice operator slice_9542_inst
    unsigned_type_9543 <= control_info_buffer(72 downto 72);
    -- flow-through slice operator slice_9546_inst
    byte_9547 <= control_info_buffer(71 downto 71);
    -- flow-through slice operator slice_9550_inst
    half_word_9551 <= control_info_buffer(70 downto 70);
    -- flow-through slice operator slice_9554_inst
    word_9555 <= control_info_buffer(69 downto 69);
    -- flow-through slice operator slice_9558_inst
    double_word_9559 <= control_info_buffer(68 downto 68);
    -- flow-through slice operator slice_9562_inst
    dbg_wp_reg_id_9563 <= control_info_buffer(67 downto 66);
    -- flow-through slice operator slice_9566_inst
    dbg_wp_read_hit_9567 <= control_info_buffer(65 downto 65);
    -- flow-through slice operator slice_9570_inst
    dbg_wp_write_hit_9571 <= control_info_buffer(64 downto 64);
    -- flow-through slice operator slice_9574_inst
    simple_store_signature_9575 <= control_info_buffer(63 downto 32);
    -- flow-through slice operator slice_9578_inst
    addr_9579 <= control_info_buffer(31 downto 0);
    -- flow-through slice operator slice_9582_inst
    messy_trap_9583 <= messy_info_buffer(97 downto 97);
    -- flow-through slice operator slice_9586_inst
    messy_error_9587 <= messy_info_buffer(96 downto 96);
    -- flow-through slice operator slice_9590_inst
    messy_store_signature_9591 <= messy_info_buffer(95 downto 64);
    -- flow-through slice operator slice_9594_inst
    messy_dout_h_9595 <= messy_info_buffer(63 downto 32);
    -- flow-through slice operator slice_9598_inst
    messy_dout_l_9599 <= messy_info_buffer(31 downto 0);
    -- flow-through slice operator slice_9731_inst
    privileged_instr_trap_9732 <= early_ls_traps_9527(2 downto 2);
    -- flow-through slice operator slice_9735_inst
    illegal_instr_trap_9736 <= early_ls_traps_9527(1 downto 1);
    -- flow-through slice operator slice_9739_inst
    mem_address_not_aligned_trap_9740 <= early_ls_traps_9527(0 downto 0);
    -- flow-through slice operator slice_9744_inst
    slice_9744_wire <= simple_store_signature_9575(31 downto 30);
    -- flow-through slice operator slice_9748_inst
    slice_9748_wire <= simple_store_signature_9575(28 downto 0);
    -- binary operator AND_u1_u1_9626_inst
    process(read_simple_9523, simple_data_access_exception_9615) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(read_simple_9523, simple_data_access_exception_9615, tmp_var);
      AND_u1_u1_9626_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_9629_inst
    process(read_messy_9519, messy_trap_9583) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(read_messy_9519, messy_trap_9583, tmp_var);
      AND_u1_u1_9629_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_9635_inst
    process(read_simple_9523, simple_data_access_error_9615) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(read_simple_9523, simple_data_access_error_9615, tmp_var);
      AND_u1_u1_9635_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_9638_inst
    process(read_messy_9519, messy_error_9587) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(read_messy_9519, messy_error_9587, tmp_var);
      AND_u1_u1_9638_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u12_u14_9701_inst
    process(CONCAT_u6_u12_9697_wire, CONCAT_u1_u2_9700_wire) -- 
      variable tmp_var : std_logic_vector(13 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u6_u12_9697_wire, CONCAT_u1_u2_9700_wire, tmp_var);
      to_cu_data_buffer <= tmp_var; --
    end process;
    -- binary operator CONCAT_u13_u16_9771_inst
    process(CONCAT_u6_u13_9765_wire, CONCAT_u2_u3_9770_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u6_u13_9765_wire, CONCAT_u2_u3_9770_wire, tmp_var);
      CONCAT_u13_u16_9771_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u13_u78_9690_inst
    process(CONCAT_u6_u13_9684_wire, CONCAT_u33_u65_9689_wire) -- 
      variable tmp_var : std_logic_vector(77 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u6_u13_9684_wire, CONCAT_u33_u65_9689_wire, tmp_var);
      to_iu_fu_data_buffer <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u54_9783_inst
    process(CONCAT_u13_u16_9771_wire, CONCAT_u4_u38_9782_wire) -- 
      variable tmp_var : std_logic_vector(53 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u13_u16_9771_wire, CONCAT_u4_u38_9782_wire, tmp_var);
      data_to_iretire_buffer <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_9700_inst
    process(dbg_wp_hit_9654, late_load_store_trap_9649) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(dbg_wp_hit_9654, late_load_store_trap_9649, tmp_var);
      CONCAT_u1_u2_9700_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_9768_inst
    process(illegal_instr_trap_9736, privileged_instr_trap_9732) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(illegal_instr_trap_9736, privileged_instr_trap_9732, tmp_var);
      CONCAT_u1_u2_9768_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_9774_inst
    process(mem_address_not_aligned_trap_9740, data_access_error_9640) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(mem_address_not_aligned_trap_9740, data_access_error_9640, tmp_var);
      CONCAT_u1_u2_9774_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_9779_inst
    process(dbg_wp_read_hit_9567, dbg_wp_write_hit_9571) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(dbg_wp_read_hit_9567, dbg_wp_write_hit_9571, tmp_var);
      CONCAT_u1_u2_9779_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u33_9687_inst
    process(late_load_store_trap_9649, dout_h_9665) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(late_load_store_trap_9649, dout_h_9665, tmp_var);
      CONCAT_u1_u33_9687_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u2_u34_9781_inst
    process(CONCAT_u1_u2_9779_wire, store_signature_9757) -- 
      variable tmp_var : std_logic_vector(33 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_9779_wire, store_signature_9757, tmp_var);
      CONCAT_u2_u34_9781_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u2_u3_9746_inst
    process(slice_9744_wire, simple_dcache_hit_9615) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_9744_wire, simple_dcache_hit_9615, tmp_var);
      CONCAT_u2_u3_9746_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u2_u3_9770_inst
    process(CONCAT_u1_u2_9768_wire, data_access_exception_9631) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_9768_wire, data_access_exception_9631, tmp_var);
      CONCAT_u2_u3_9770_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u2_u4_9776_inst
    process(CONCAT_u1_u2_9774_wire, dbg_wp_reg_id_9563) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_9774_wire, dbg_wp_reg_id_9563, tmp_var);
      CONCAT_u2_u4_9776_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u33_u65_9689_inst
    process(CONCAT_u1_u33_9687_wire, dout_l_9676) -- 
      variable tmp_var : std_logic_vector(64 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u33_9687_wire, dout_l_9676, tmp_var);
      CONCAT_u33_u65_9689_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u3_u32_9749_inst
    process(CONCAT_u2_u3_9746_wire, slice_9748_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u2_u3_9746_wire, slice_9748_wire, tmp_var);
      CONCAT_u3_u32_9749_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u4_u38_9782_inst
    process(CONCAT_u2_u4_9776_wire, CONCAT_u2_u34_9781_wire) -- 
      variable tmp_var : std_logic_vector(37 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u2_u4_9776_wire, CONCAT_u2_u34_9781_wire, tmp_var);
      CONCAT_u4_u38_9782_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u4_u6_9680_inst
    process(thread_id_9491, stream_id_9495) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApConcat_proc(thread_id_9491, stream_id_9495, tmp_var);
      CONCAT_u4_u6_9680_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u4_u6_9695_inst
    process(thread_id_9491, stream_id_9495) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApConcat_proc(thread_id_9491, stream_id_9495, tmp_var);
      CONCAT_u4_u6_9695_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u4_u6_9761_inst
    process(thread_id_9491, stream_id_9495) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApConcat_proc(thread_id_9491, stream_id_9495, tmp_var);
      CONCAT_u4_u6_9761_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u6_u12_9697_inst
    process(CONCAT_u4_u6_9695_wire, slot_id_9499) -- 
      variable tmp_var : std_logic_vector(11 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u4_u6_9695_wire, slot_id_9499, tmp_var);
      CONCAT_u6_u12_9697_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u6_u13_9684_inst
    process(CONCAT_u4_u6_9680_wire, CONCAT_u6_u7_9683_wire) -- 
      variable tmp_var : std_logic_vector(12 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u4_u6_9680_wire, CONCAT_u6_u7_9683_wire, tmp_var);
      CONCAT_u6_u13_9684_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u6_u13_9765_inst
    process(CONCAT_u4_u6_9761_wire, CONCAT_u6_u7_9764_wire) -- 
      variable tmp_var : std_logic_vector(12 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u4_u6_9761_wire, CONCAT_u6_u7_9764_wire, tmp_var);
      CONCAT_u6_u13_9765_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u6_u7_9683_inst
    process(slot_id_9499, dbg_wp_hit_9654) -- 
      variable tmp_var : std_logic_vector(6 downto 0); -- 
    begin -- 
      ApConcat_proc(slot_id_9499, dbg_wp_hit_9654, tmp_var);
      CONCAT_u6_u7_9683_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u6_u7_9764_inst
    process(slot_id_9499, late_load_store_trap_9649) -- 
      variable tmp_var : std_logic_vector(6 downto 0); -- 
    begin -- 
      ApConcat_proc(slot_id_9499, late_load_store_trap_9649, tmp_var);
      CONCAT_u6_u7_9764_wire <= tmp_var; --
    end process;
    -- binary operator NEQ_u3_u1_9644_inst
    process(early_ls_traps_9527) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(early_ls_traps_9527, konst_9643_wire_constant, tmp_var);
      NEQ_u3_u1_9644_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_9630_inst
    process(AND_u1_u1_9626_wire, AND_u1_u1_9629_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_9626_wire, AND_u1_u1_9629_wire, tmp_var);
      data_access_exception_9631 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_9639_inst
    process(AND_u1_u1_9635_wire, AND_u1_u1_9638_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_9635_wire, AND_u1_u1_9638_wire, tmp_var);
      data_access_error_9640 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_9646_inst
    process(NEQ_u3_u1_9644_wire, data_access_exception_9631) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NEQ_u3_u1_9644_wire, data_access_exception_9631, tmp_var);
      OR_u1_u1_9646_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_9648_inst
    process(OR_u1_u1_9646_wire, data_access_error_9640) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_9646_wire, data_access_error_9640, tmp_var);
      late_load_store_trap_9649 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_9653_inst
    process(dbg_wp_read_hit_9567, dbg_wp_write_hit_9571) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(dbg_wp_read_hit_9567, dbg_wp_write_hit_9571, tmp_var);
      dbg_wp_hit_9654 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_9664_inst
    process(MUX_9659_wire, MUX_9663_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_9659_wire, MUX_9663_wire, tmp_var);
      dout_h_9665 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_9675_inst
    process(MUX_9670_wire, MUX_9674_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_9670_wire, MUX_9674_wire, tmp_var);
      dout_l_9676 <= tmp_var; --
    end process;
    -- binary operator OR_u32_u32_9756_inst
    process(MUX_9751_wire, MUX_9755_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_9751_wire, MUX_9755_wire, tmp_var);
      store_signature_9757 <= tmp_var; --
    end process;
    volatile_operator_analyze_dcache_response_8445: analyze_dcache_response_VVP port map(addr => addr_9579, dcache_response => simple_info_buffer, is_load => is_load_9531, is_store => is_store_9535, signed_type => signed_type_9539, unsigned_type => unsigned_type_9543, byte => byte_9547, half_word => half_word_9551, word => word_9555, double_word => double_word_9559, dout_h => simple_dout_h_9615, dout_l => simple_dout_l_9615, data_access_exception => simple_data_access_exception_9615, data_access_error => simple_data_access_error_9615, dcache_hit => simple_dcache_hit_9615); 
    -- 
  end Block; -- data_path
  -- 
end loadstore_router_core_VVP_arch;

library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
entity load_store_router_daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    DCACHE_to_CPU_response_pipe_read_req : out  std_logic_vector(0 downto 0);
    DCACHE_to_CPU_response_pipe_read_ack : in   std_logic_vector(0 downto 0);
    DCACHE_to_CPU_response_pipe_read_data : in   std_logic_vector(71 downto 0);
    load_store_messy_to_router_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    load_store_messy_to_router_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    load_store_messy_to_router_pipe_pipe_read_data : in   std_logic_vector(97 downto 0);
    load_store_router_control_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    load_store_router_control_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    load_store_router_control_pipe_pipe_read_data : in   std_logic_vector(96 downto 0);
    teu_loadstore_to_fpunit_pipe_write_req : out  std_logic_vector(0 downto 0);
    teu_loadstore_to_fpunit_pipe_write_ack : in   std_logic_vector(0 downto 0);
    teu_loadstore_to_fpunit_pipe_write_data : out  std_logic_vector(77 downto 0);
    teu_loadstore_to_iretire_pipe_write_req : out  std_logic_vector(0 downto 0);
    teu_loadstore_to_iretire_pipe_write_ack : in   std_logic_vector(0 downto 0);
    teu_loadstore_to_iretire_pipe_write_data : out  std_logic_vector(53 downto 0);
    teu_loadstore_to_iunit_pipe_write_req : out  std_logic_vector(0 downto 0);
    teu_loadstore_to_iunit_pipe_write_ack : in   std_logic_vector(0 downto 0);
    teu_loadstore_to_iunit_pipe_write_data : out  std_logic_vector(77 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity load_store_router_daemon;
architecture load_store_router_daemon_arch of load_store_router_daemon is -- 
  -- volatile/operator module components. 
  component decode_routing_control_info_VVP is -- 
    port ( -- 
      control_info : in  std_logic_vector(96 downto 0);
      read_simple : out  std_logic_vector(0 downto 0);
      read_messy : out  std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component; 
  component loadstore_router_core_VVP is -- 
    port ( -- 
      control_info : in  std_logic_vector(96 downto 0);
      simple_info : in  std_logic_vector(71 downto 0);
      messy_info : in  std_logic_vector(97 downto 0);
      to_iu : out  std_logic_vector(0 downto 0);
      to_fu : out  std_logic_vector(0 downto 0);
      to_cu : out  std_logic_vector(0 downto 0);
      to_retire : out  std_logic_vector(0 downto 0);
      to_iu_fu_data : out  std_logic_vector(77 downto 0);
      to_cu_data : out  std_logic_vector(13 downto 0);
      data_to_iretire : out  std_logic_vector(53 downto 0)-- 
    );
    -- 
  end component; 
  
  signal do_transfer: boolean;
  signal read_simple, read_messy: std_logic_vector(0 downto 0);

  signal to_iu, to_fu, to_cu, to_retire: std_logic_vector(0 downto 0);
  signal to_iu_fu_data : std_logic_vector(77 downto 0);
  signal to_cu_data : std_logic_vector(13 downto 0);
  signal data_to_iretire : std_logic_vector(53 downto 0);

  signal dcache_rdy, messy_rdy, iu_rdy, fu_rdy, retire_rdy, ctrl_rdy: boolean;

  signal pop_req_to_ctrl, pop_ack_from_ctrl: std_logic;
  signal pop_req_to_messy, pop_ack_from_messy: std_logic;
  signal pop_req_to_dcache, pop_ack_from_dcache: std_logic;

  signal data_from_dcache : std_logic_vector(71 downto 0);
  signal data_from_ctrl: std_logic_vector(96 downto 0);
  signal data_from_messy : std_logic_vector(97 downto 0);
begin --  
    tag_out <= (others => '0');
    start_ack <= '1';
    fin_ack <= '0';

    --      Input Queues!
    qCtrl: QueueBase
		generic map (name => "ls_router_qCtrl",
				queue_depth => 2, data_width => 97)
		port map (clk => clk, reset => reset,
				data_in => load_store_router_control_pipe_pipe_read_data,
				 push_req => load_store_router_control_pipe_pipe_read_ack(0),
				 push_ack => load_store_router_control_pipe_pipe_read_req(0),
				data_out => data_from_ctrl, 
				 pop_req => pop_req_to_ctrl,
				 pop_ack => pop_ack_from_ctrl);

    qMessy: QueueBase
		generic map (name => "ls_router_qMessy",
				queue_depth => 2, data_width => 98)
		port map (clk => clk, reset => reset,
				data_in => load_store_messy_to_router_pipe_pipe_read_data,
				 push_req => load_store_messy_to_router_pipe_pipe_read_ack(0),
				 push_ack => load_store_messy_to_router_pipe_pipe_read_req(0),
				data_out => data_from_messy, 
				 pop_req => pop_req_to_messy,
				 pop_ack => pop_ack_from_messy);

    -- dcache bypassed into iunit/fpunit..  This seems to be an issue
    -- in the ASIC, since delays are a bit large..
    qDcache: QueueWithBypass
		generic map (name => "ls_router_qDcache",
				queue_depth => 2, data_width => 72)
		port map (clk => clk, reset => reset,
				data_in => DCACHE_to_CPU_response_pipe_read_data,
				 push_req => DCACHE_to_CPU_response_pipe_read_ack(0),
				 push_ack => DCACHE_to_CPU_response_pipe_read_req(0),
				data_out => data_from_dcache, 
				 pop_req => pop_req_to_dcache,
				 pop_ack => pop_ack_from_dcache);

    -- decode incoming!
    decRtr: decode_routing_control_info_VVP
		port map (control_info => data_from_ctrl,
					read_simple => read_simple, read_messy => read_messy);
    coreInst: loadstore_router_core_VVP
			port map (control_info => data_from_ctrl,
					simple_info => data_from_dcache,
					   messy_info => data_from_messy,
					     to_iu => to_iu, to_fu => to_fu, to_cu => to_cu, to_retire => to_retire,
						to_iu_fu_data => to_iu_fu_data, to_cu_data => to_cu_data, data_to_iretire => data_to_iretire);

    -- determine if transfer should go ahead.
    ctrl_rdy   <=   (pop_ack_from_ctrl = '1');
    dcache_rdy <=   ((read_simple(0) = '0') or  (pop_ack_from_dcache = '1'));
    messy_rdy  <=   ((read_messy(0) = '0') or (pop_ack_from_messy = '1'));
    iu_rdy     <=   ((to_iu(0) = '0') or (teu_loadstore_to_iunit_pipe_write_ack(0) = '1'));
    fu_rdy     <=   ((to_fu(0) = '0') or (teu_loadstore_to_fpunit_pipe_write_ack(0) = '1'));
    retire_rdy <=   ((to_retire(0) = '0') or (teu_loadstore_to_iretire_pipe_write_ack(0) = '1'));

    do_transfer <= ctrl_rdy
			and dcache_rdy
			and messy_rdy
			and iu_rdy
			and fu_rdy
			and retire_rdy;

    -- writes to targets.
    teu_loadstore_to_iunit_pipe_write_data <= to_iu_fu_data; 
    teu_loadstore_to_iunit_pipe_write_req(0) <= '1' when do_transfer and (to_iu(0) = '1') else '0';

    teu_loadstore_to_fpunit_pipe_write_data <= to_iu_fu_data; 
    teu_loadstore_to_fpunit_pipe_write_req(0) <= '1' when do_transfer and (to_fu(0) = '1') else '0';


    teu_loadstore_to_iretire_pipe_write_data <= data_to_iretire; 
    teu_loadstore_to_iretire_pipe_write_req(0) <= '1' when do_transfer and (to_retire(0) = '1') else '0';

    -- reqs to sources.
    pop_req_to_ctrl <= '1' when do_transfer else '0';
    pop_req_to_messy <= '1' when do_transfer and (read_messy(0) = '1') else '0';
    pop_req_to_dcache <= '1' when do_transfer and (read_simple(0) = '1') else '0';

end load_store_router_daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
entity needSignalFromRetire_VVV is -- 
  port ( -- 
    msg_from_sc : in  std_logic_vector(147 downto 0);
    sc_valid : out  std_logic_vector(0 downto 0);
    wait_on_iretire : out  std_logic_vector(0 downto 0)-- 
  );
  -- 
end entity needSignalFromRetire_VVV;
architecture needSignalFromRetire_VVV_arch of needSignalFromRetire_VVV is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(148-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal msg_from_sc_buffer :  std_logic_vector(147 downto 0);
  -- output port buffer signals
  signal sc_valid_buffer :  std_logic_vector(0 downto 0);
  signal wait_on_iretire_buffer :  std_logic_vector(0 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  msg_from_sc_buffer <= msg_from_sc;
  -- output handling  -------------------------------------------------------
  sc_valid <= sc_valid_buffer;
  wait_on_iretire <= wait_on_iretire_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal w_9142 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    -- flow-through slice operator slice_9137_inst
    sc_valid_buffer <= msg_from_sc_buffer(147 downto 147);
    -- flow-through slice operator slice_9141_inst
    w_9142 <= msg_from_sc_buffer(134 downto 134);
    -- binary operator AND_u1_u1_9146_inst
    process(sc_valid_buffer, w_9142) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      -- ApIntAnd_proc(sc_valid_buffer, w_9142, tmp_var);
      tmp_var := sc_valid_buffer and w_9142;
      wait_on_iretire_buffer <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end needSignalFromRetire_VVV_arch;

library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.types.all;
use ahir.BaseComponents.all;

entity sc_iretire_join_daemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    noblock_teu_stream_corrector_to_idispatch_pipe_read_req : out  std_logic_vector(0 downto 0);
    noblock_teu_stream_corrector_to_idispatch_pipe_read_ack : in   std_logic_vector(0 downto 0);
    noblock_teu_stream_corrector_to_idispatch_pipe_read_data : in   std_logic_vector(147 downto 0);
    teu_iretire_to_idispatch_pipe_read_req : out  std_logic_vector(0 downto 0);
    teu_iretire_to_idispatch_pipe_read_ack : in   std_logic_vector(0 downto 0);
    teu_iretire_to_idispatch_pipe_read_data : in   std_logic_vector(0 downto 0);
    noblock_joined_iretire_sc_to_idispatch_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_joined_iretire_sc_to_idispatch_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_joined_iretire_sc_to_idispatch_pipe_write_data : out  std_logic_vector(147 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity sc_iretire_join_daemon;
architecture sc_iretire_join_daemon_arch of sc_iretire_join_daemon is -- 
  -- volatile/operator module components. 
  component needSignalFromRetire_VVV is -- 
    port ( -- 
      msg_from_sc : in  std_logic_vector(147 downto 0);
      sc_valid : out  std_logic_vector(0 downto 0);
      wait_on_iretire : out  std_logic_vector(0 downto 0)-- 
    );
    -- 
  end component; 

  signal msg_from_sc : std_logic_vector(147 downto 0);
  signal wait_on_iretire, sc_valid: std_logic_vector(0 downto 0);
 
  signal sc_ok, iretire_ok, dest_ready: boolean;
  signal write_to_dest_valid, need_iretire: boolean;
  
  signal pop_req_to_sc, pop_ack_from_sc: std_logic;
  signal data_from_sc: std_logic_vector(147 downto 0);

begin --  
	start_ack <= '1';
	fin_ack <= '0';
	tag_out <= tag_in;

        -- receive the data in a queue.
	qbSC: QueueBase
		generic map (name => "sc_iretire_join_qbSC",
				queue_depth => 1, data_width => 148)
		port map (clk => clk, reset => reset,
				data_in => noblock_teu_stream_corrector_to_idispatch_pipe_read_data ,
				 push_req => noblock_teu_stream_corrector_to_idispatch_pipe_read_ack(0),
				 push_ack => noblock_teu_stream_corrector_to_idispatch_pipe_read_req(0),
				 data_out => data_from_sc, 
				 pop_req => pop_req_to_sc,
				 pop_ack => pop_ack_from_sc);


	-- raw message from sc.. forwarded.
	noblock_joined_iretire_sc_to_idispatch_pipe_write_data <= data_from_sc;

	-- writers ok?
	sc_ok <= pop_ack_from_sc = '1';
        iretire_ok <= teu_iretire_to_idispatch_pipe_read_ack(0) = '1';

	-- destination ready?
	dest_ready <= noblock_joined_iretire_sc_to_idispatch_pipe_write_ack(0) = '1'; 

	-- needs to join iretire?
	need_iretire <= sc_ok and (sc_valid(0) = '1') and (wait_on_iretire(0) = '1');

	-- can write to dest?  if sc-ok and iretire ok..
	write_to_dest_valid <= sc_ok and (sc_valid(0) = '1') and ((not need_iretire) or iretire_ok);


	-- write request if writers are available.
	noblock_joined_iretire_sc_to_idispatch_pipe_write_req(0) <= '1' when write_to_dest_valid else '0';

	-- requests go out if transfer possible.
	pop_req_to_sc <= '1' when (write_to_dest_valid and dest_ready) else '0';

	-- iretire to idispatch.
	teu_iretire_to_idispatch_pipe_read_req (0) <= 
				'1' when (write_to_dest_valid and need_iretire and dest_ready) 
								else '0';

  	decInst: needSignalFromRetire_VVV
			port map (msg_from_sc => data_from_sc, wait_on_iretire => wait_on_iretire,
								sc_valid => sc_valid);



end sc_iretire_join_daemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##
library ahir;
use ahir.basecomponents.all;

entity stream_corrector_in_mux_daemon_v2 is -- 
  generic (tag_length : integer := 1); 
  port ( -- 
    teu_idispatch_to_stream_corrector_pipe_read_req : out  std_logic_vector(0 downto 0);
    teu_idispatch_to_stream_corrector_pipe_read_ack : in   std_logic_vector(0 downto 0);
    teu_idispatch_to_stream_corrector_pipe_read_data : in   std_logic_vector(204 downto 0);
    teu_fpunit_cc_to_stream_corrector_pipe_read_req : out  std_logic_vector(0 downto 0);
    teu_fpunit_cc_to_stream_corrector_pipe_read_ack : in   std_logic_vector(0 downto 0);
    teu_fpunit_cc_to_stream_corrector_pipe_read_data : in   std_logic_vector(14 downto 0);
    teu_iunit_cc_to_stream_corrector_pipe_read_req : out  std_logic_vector(0 downto 0);
    teu_iunit_cc_to_stream_corrector_pipe_read_ack : in   std_logic_vector(0 downto 0);
    teu_iunit_cc_to_stream_corrector_pipe_read_data : in   std_logic_vector(16 downto 0);
    teu_iunit_rs1_to_stream_corrector_pipe_read_req : out  std_logic_vector(0 downto 0);
    teu_iunit_rs1_to_stream_corrector_pipe_read_ack : in   std_logic_vector(0 downto 0);
    teu_iunit_rs1_to_stream_corrector_pipe_read_data : in   std_logic_vector(31 downto 0);
    teu_iunit_to_stream_corrector_pipe_read_req : out  std_logic_vector(0 downto 0);
    teu_iunit_to_stream_corrector_pipe_read_ack : in   std_logic_vector(0 downto 0);
    teu_iunit_to_stream_corrector_pipe_read_data : in   std_logic_vector(89 downto 0);
    noblock_stream_corrector_in_args_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_stream_corrector_in_args_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_stream_corrector_in_args_pipe_write_data : out  std_logic_vector(359 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity stream_corrector_in_mux_daemon_v2;
architecture stream_corrector_in_mux_daemon_arch of stream_corrector_in_mux_daemon_v2 is -- 

   signal pop_req_to_dispatch, pop_ack_from_dispatch : std_logic;
   signal data_from_dispatch:  std_logic_vector(204 downto 0);

   signal other_data: std_logic_vector(153 downto 0);

   signal pop_req_to_iu_cc, pop_ack_from_iu_cc : std_logic;
   signal data_from_iu_cc : std_logic_vector(16 downto 0);

   signal pop_req_to_iu_rs1, pop_ack_from_iu_rs1 : std_logic;
   signal data_from_iu_rs1 : std_logic_vector(31 downto 0);

   signal pop_req_to_fp_cc, pop_ack_from_fp_cc : std_logic;
   signal data_from_fp_cc : std_logic_vector(14 downto 0);

   signal pop_req_to_iu, pop_ack_from_iu : std_logic;
   signal data_from_iu : std_logic_vector(89 downto 0);


   signal dispatch_valid, read_iu, read_iu_cc, read_iu_rs1, read_fp_cc: boolean;
   signal dest_rdy, iu_cc_rdy, iu_rs1_rdy, iu_rdy, fp_cc_rdy : boolean;

   signal write_to_dest, do_transfer : boolean;

   signal const_one_sig: std_logic_vector(0 downto 0);
   constant debug_print_flag: boolean := false;

-- see comment above..
--##decl_synopsys_sync_set_reset##


begin --  

	-- stubbing.
	start_ack <= '1';
	fin_ack   <= '0';
	tag_out   <= tag_in;
	const_one_sig(0) <= '1';

	dispatch_valid <= (pop_ack_from_dispatch = '1');

	read_iu_cc <= dispatch_valid and (data_from_dispatch(137) = '1');
	iu_cc_rdy     <= (not read_iu_cc) or (pop_ack_from_iu_cc = '1');

	read_fp_cc <= dispatch_valid and (data_from_dispatch(136) = '1');
	fp_cc_rdy     <= (not read_fp_cc) or (pop_ack_from_fp_cc = '1');

	read_iu_rs1 <= dispatch_valid and (data_from_dispatch(135) = '1');
	iu_rs1_rdy     <= (not read_iu_rs1) or (pop_ack_from_iu_rs1 = '1');

	read_iu    <= dispatch_valid and (data_from_dispatch(134) = '1');
	iu_rdy     <= (not read_iu) or (pop_ack_from_iu = '1');

	-- qualified other data
	process (data_from_iu_cc, 
			data_from_iu_rs1, 
			data_from_iu, 
			data_from_fp_cc,
			read_iu_cc, 
			read_iu_rs1, 
			read_iu, 
			read_fp_cc)
		variable data_from_iu_cc_var: std_logic_vector(16 downto 0);
		variable data_from_iu_rs1_var: std_logic_vector(31 downto 0);
		variable data_from_fp_cc_var: std_logic_vector(14 downto 0);
		variable data_from_iu_var: std_logic_vector(89 downto 0);

	begin
		if(read_iu_cc) then
			data_from_iu_cc_var := data_from_iu_cc;
		else	
			data_from_iu_cc_var := (others => '0');
		end if;
		if(read_iu_rs1) then
			data_from_iu_rs1_var := data_from_iu_rs1;
		else	
			data_from_iu_rs1_var := (others => '0');
		end if;
		if(read_fp_cc) then
			data_from_fp_cc_var := data_from_fp_cc;
		else	
			data_from_fp_cc_var := (others => '0');
		end if;
		if(read_iu) then
			data_from_iu_var := data_from_iu;
		else	
			data_from_iu_var := (others => '0');
		end if;

		other_data <= data_from_iu_cc_var & data_from_iu_rs1_var & data_from_iu_var & data_from_fp_cc_var;

	end process;

	-- Need to cut the long path...
	qbDispatch: QueueBase
		generic map (name => "sc_in_mux_qbDispatch", queue_depth => 2, data_width => 205)
		port map (
			clk => clk, reset => reset,
			data_in => teu_idispatch_to_stream_corrector_pipe_read_data,
			push_req => teu_idispatch_to_stream_corrector_pipe_read_ack(0),
			push_ack => teu_idispatch_to_stream_corrector_pipe_read_req(0),
			data_out => data_from_dispatch,
			pop_req  => pop_req_to_dispatch,
			pop_ack  => pop_ack_from_dispatch);

	-- bypass..  registered downstream..
	qbIUCC: QueueWithBypass
		generic map (name => "sc_in_mux_qbIUCC", queue_depth => 2, data_width => 17)
		port map (
			clk => clk, reset => reset,
			data_in => teu_iunit_cc_to_stream_corrector_pipe_read_data,
			push_req => teu_iunit_cc_to_stream_corrector_pipe_read_ack(0),
			push_ack => teu_iunit_cc_to_stream_corrector_pipe_read_req(0),
			data_out => data_from_iu_cc,
			pop_req  => pop_req_to_iu_cc,
			pop_ack  => pop_ack_from_iu_cc);

	qbIURS1: QueueWithBypass
		generic map (name => "sc_in_mux_qbIURS1", queue_depth => 2, data_width => 32)
		port map (
			clk => clk, reset => reset,
			data_in => teu_iunit_rs1_to_stream_corrector_pipe_read_data,
			push_req => teu_iunit_rs1_to_stream_corrector_pipe_read_ack(0),
			push_ack => teu_iunit_rs1_to_stream_corrector_pipe_read_req(0),
			data_out => data_from_iu_rs1,
			pop_req  => pop_req_to_iu_rs1,
			pop_ack  => pop_ack_from_iu_rs1);


	-- not critical...
	qbIU: QueueBase
		generic map (name => "sc_in_mux_qbIU", queue_depth => 1, data_width => 90)
		port map (
			clk => clk, reset => reset,
			data_in => teu_iunit_to_stream_corrector_pipe_read_data,
			push_req => teu_iunit_to_stream_corrector_pipe_read_ack(0),
			push_ack => teu_iunit_to_stream_corrector_pipe_read_req(0),
			data_out => data_from_iu,
			pop_req  => pop_req_to_iu,
			pop_ack  => pop_ack_from_iu);

	qbFPCC: QueueWithBypass
		generic map (name => "sc_in_mux_qbFPCC", queue_depth => 2, data_width => 15)
		port map (
			clk => clk, reset => reset,
			data_in => teu_fpunit_cc_to_stream_corrector_pipe_read_data,
			push_req => teu_fpunit_cc_to_stream_corrector_pipe_read_ack(0),
			push_ack => teu_fpunit_cc_to_stream_corrector_pipe_read_req(0),
			data_out => data_from_fp_cc,
			pop_req  => pop_req_to_fp_cc,
			pop_ack  => pop_ack_from_fp_cc);

	-- destination side..
	dest_rdy   <= (noblock_stream_corrector_in_args_pipe_write_ack(0) = '1'); 


	-- do transfer.
	do_transfer <= dest_rdy and 
				dispatch_valid and 
				iu_cc_rdy and 
				iu_rs1_rdy and
				iu_rdy and
				fp_cc_rdy;

	-- pops!
	pop_req_to_dispatch <= '1' when do_transfer else '0';
	pop_req_to_iu_cc <= '1' when (do_transfer and read_iu_cc) else '0';
	pop_req_to_iu_rs1 <= '1' when (do_transfer and read_iu_rs1) else '0';
	pop_req_to_iu     <= '1' when (do_transfer and read_iu) else '0';
	pop_req_to_fp_cc     <= '1' when (do_transfer and read_fp_cc) else '0';

	


	write_to_dest <= do_transfer;
	noblock_stream_corrector_in_args_pipe_write_req(0) <= '1' when write_to_dest else '0';
	noblock_stream_corrector_in_args_pipe_write_data <= (const_one_sig & data_from_dispatch & other_data);

end stream_corrector_in_mux_daemon_arch;

library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
-- Synopsys DC ($^^$@!)  needs you to declare an attribute
-- to infer a synchronous set/reset ... unbelievable.
--##decl_synopsys_attribute_lib##
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
entity stream_corrector_in_mux_daemon is -- 
  generic (tag_length : integer := 1); 
  port ( -- 
    teu_idispatch_to_stream_corrector_pipe_read_req : out  std_logic_vector(0 downto 0);
    teu_idispatch_to_stream_corrector_pipe_read_ack : in   std_logic_vector(0 downto 0);
    teu_idispatch_to_stream_corrector_pipe_read_data : in   std_logic_vector(203 downto 0);
    teu_fpunit_cc_to_stream_corrector_pipe_read_req : out  std_logic_vector(0 downto 0);
    teu_fpunit_cc_to_stream_corrector_pipe_read_ack : in   std_logic_vector(0 downto 0);
    teu_fpunit_cc_to_stream_corrector_pipe_read_data : in   std_logic_vector(14 downto 0);
    teu_iunit_cc_to_stream_corrector_pipe_read_req : out  std_logic_vector(0 downto 0);
    teu_iunit_cc_to_stream_corrector_pipe_read_ack : in   std_logic_vector(0 downto 0);
    teu_iunit_cc_to_stream_corrector_pipe_read_data : in   std_logic_vector(16 downto 0);
    teu_iunit_to_stream_corrector_pipe_read_req : out  std_logic_vector(0 downto 0);
    teu_iunit_to_stream_corrector_pipe_read_ack : in   std_logic_vector(0 downto 0);
    teu_iunit_to_stream_corrector_pipe_read_data : in   std_logic_vector(89 downto 0);
    noblock_stream_corrector_in_args_pipe_write_req : out  std_logic_vector(0 downto 0);
    noblock_stream_corrector_in_args_pipe_write_ack : in   std_logic_vector(0 downto 0);
    noblock_stream_corrector_in_args_pipe_write_data : out  std_logic_vector(326 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity stream_corrector_in_mux_daemon;
architecture stream_corrector_in_mux_daemon_arch of stream_corrector_in_mux_daemon is -- 

   signal pop_req_to_dispatch, pop_ack_from_dispatch : std_logic;
   signal data_from_dispatch, data_from_dispatch_reg: std_logic_vector(203 downto 0);


   signal other_data_reg, other_data: std_logic_vector(121 downto 0);


   signal pop_req_to_iu_cc, pop_ack_from_iu_cc : std_logic;
   signal data_from_iu_cc : std_logic_vector(16 downto 0);

   signal pop_req_to_fp_cc, pop_ack_from_fp_cc : std_logic;
   signal data_from_fp_cc : std_logic_vector(14 downto 0);

   signal pop_req_to_iu, pop_ack_from_iu : std_logic;
   signal data_from_iu : std_logic_vector(89 downto 0);


   signal dispatch_valid, read_iu, read_iu_cc, read_fp_cc: boolean;
   signal dest_rdy, iu_cc_rdy, iu_rdy, fp_cc_rdy : boolean;

   signal write_to_dest : boolean;

   type FsmState is (Idle, WaitOnInputs, WaitOnDestination);
   signal fsm_state: FsmState;

   -- from FSM.
   signal read_iu_cc_reg, read_fp_cc_reg, read_iu_reg: boolean;

   signal latch_dispatch_data, latch_other_data: boolean;
   signal clear_dispatch_data, clear_other_data: boolean;


   signal const_one_sig: std_logic_vector(0 downto 0);

   constant debug_print_flag: boolean := false;

-- see comment above..
--##decl_synopsys_sync_set_reset##


begin --  

	-- stubbing.
	start_ack <= '1';
	fin_ack   <= '0';
	tag_out   <= tag_in;
	const_one_sig(0) <= '1';

	dispatch_valid <= (pop_ack_from_dispatch = '1');

	read_iu_cc <= dispatch_valid and (data_from_dispatch(136) = '1');
	iu_cc_rdy     <= (pop_ack_from_iu_cc = '1');

	read_fp_cc <= dispatch_valid and (data_from_dispatch(135) = '1');
	fp_cc_rdy     <= (pop_ack_from_fp_cc = '1');

	read_iu    <= dispatch_valid and (data_from_dispatch(134) = '1');
	iu_rdy     <= (pop_ack_from_iu = '1');

        dbgGen: if debug_print_flag generate

	  process(clk, reset)
	  begin
		if(clk'event and clk = '1') then
			if(reset = '0') then
				assert (not ((read_iu_cc and read_iu) or
						(read_iu_cc and read_fp_cc)))
					report "Error: in stream_corrector_in_mux_daemon:  two inputs selected" 
						severity error;
			end if;
		end if;
	  end process;

        end generate dbgGen;


	process(clk, fsm_state, dispatch_valid, read_iu_cc, read_fp_cc, read_iu, 
					iu_cc_rdy, fp_cc_rdy, iu_rdy, dest_rdy,
					read_iu_cc, read_iu, read_fp_cc,
					read_iu_cc_reg, read_iu_reg, read_fp_cc_reg)
		variable next_read_iu_cc_reg_var, next_read_fp_cc_reg_var, next_read_iu_reg_var: boolean;
		variable next_fsm_state_var: FsmState;

		variable latch_dispatch_data_var, latch_other_data_var: boolean;
		variable clear_dispatch_data_var, clear_other_data_var: boolean;

		variable iu_cc_value_var: std_logic_vector(16 downto 0);
		variable fp_cc_value_var: std_logic_vector(14 downto 0);
		variable iu_value_var: std_logic_vector(89 downto 0);

		variable write_to_dest_var: boolean;
   		variable pop_req_to_dispatch_var,
				pop_req_to_iu_var, pop_req_to_iu_cc_var, pop_req_to_fp_cc_var: std_logic;

	begin
		next_fsm_state_var := fsm_state;

		latch_dispatch_data_var := false;
		clear_dispatch_data_var := false;

		latch_other_data_var := false;
		clear_other_data_var := false;

		write_to_dest_var := false;

		-- remember what we are doing..
		next_read_iu_cc_reg_var := read_iu_cc_reg;
		next_read_fp_cc_reg_var := read_fp_cc_reg;
		next_read_iu_reg_var    := read_iu_reg;

		pop_req_to_dispatch_var := '0';
		pop_req_to_iu_var := '0';
		pop_req_to_iu_cc_var := '0';
		pop_req_to_fp_cc_var := '0';

		case fsm_state is
			when Idle =>

				-- ready to pick up data from dispatch
				pop_req_to_dispatch_var := '1';
				if(dispatch_valid) then

					-- dispatch is valid, latch the data from dispatch.
					latch_dispatch_data_var := true;
					-- clear stale old data.			
					clear_other_data_var:= true;

					-- remember the read-flags.
					next_read_iu_cc_reg_var :=  read_iu_cc;
					next_read_fp_cc_reg_var :=  read_fp_cc;
					next_read_iu_reg_var    :=  read_iu;

					next_fsm_state_var := WaitOnInputs;

				end if;

			when WaitOnInputs =>

				--
				-- set up the pops... exactly one of these
				-- will be acked.
				--
				if(read_iu_cc_reg) then
					pop_req_to_iu_cc_var := '1';
				end if;
				if(read_iu_reg) then
					pop_req_to_iu_var := '1';
				end if;
				if(read_fp_cc_reg) then
					pop_req_to_fp_cc_var := '1';
				end if;

				if (((not read_iu_cc_reg) or iu_cc_rdy) and
					((not read_iu_reg) or iu_rdy) and
					((not read_fp_cc_reg) or fp_cc_rdy)) then

					-- all pops are acked?  send response
					write_to_dest_var := true;

					if dest_rdy then
					-- destination is accepting the response..

						-- check if dispatch has something for us.
						pop_req_to_dispatch_var := '1';

						if(dispatch_valid) then
						-- yes it does... 
	
							-- latch the dispatch-data.	
							latch_dispatch_data_var := true;

							-- clear the old-data
							clear_other_data_var:= true;

							-- register the read flags.
							next_read_iu_cc_reg_var :=  read_iu_cc;
							next_read_fp_cc_reg_var :=  read_fp_cc;
							next_read_iu_reg_var    :=  read_iu;

							-- stay in this state.

						else
							next_fsm_state_var := Idle;
							
							next_read_iu_cc_reg_var :=  false;
							next_read_fp_cc_reg_var :=  false;
							next_read_iu_reg_var :=  false;

							clear_other_data_var:= true;
						end if;
					 else
						-- other data is ready but destination is not.
						next_fsm_state_var := WaitOnDestination;

						-- remember other data.
						latch_other_data_var := true;
					 end if;
				end if;
					
			when WaitOnDestination =>
				write_to_dest_var := true;
				if dest_rdy then
					-- same logic as before..
					pop_req_to_dispatch_var := '1';
					clear_other_data_var:= true;

					if(dispatch_valid) then

						latch_dispatch_data_var := true;

						next_read_iu_cc_reg_var :=  read_iu_cc;
						next_read_fp_cc_reg_var :=  read_fp_cc;
						next_read_iu_reg_var    :=  read_iu;

						next_fsm_state_var := WaitOnInputs;
					else
						next_fsm_state_var := Idle;
							
						next_read_iu_cc_reg_var :=  false;
						next_read_fp_cc_reg_var :=  false;
						next_read_iu_reg_var :=  false;
					end if;
				end if;
		end case;

		latch_dispatch_data <= latch_dispatch_data_var;
		clear_dispatch_data <= clear_dispatch_data_var;

		latch_other_data <= latch_other_data_var;
		clear_other_data <= clear_other_data_var;

		write_to_dest <= write_to_dest_var;

		pop_req_to_dispatch <= pop_req_to_dispatch_var;
		pop_req_to_iu_cc <= pop_req_to_iu_cc_var;
		pop_req_to_iu    <= pop_req_to_iu_var;
		pop_req_to_fp_cc <= pop_req_to_fp_cc_var;

		if(clk'event and clk = '1') then
			if(reset = '1') then
				fsm_state <= Idle;
				read_iu_cc_reg <= false;
				read_fp_cc_reg <= false;
				read_iu_reg <= false;
			else
				fsm_state <= next_fsm_state_var;
				read_iu_cc_reg <= next_read_iu_cc_reg_var;
				read_fp_cc_reg <= next_read_fp_cc_reg_var;
				read_iu_reg <= next_read_iu_reg_var;
			end if;
		end if;
	end process;


	-- qualified other data
	process (data_from_iu_cc, data_from_iu, data_from_fp_cc,
			read_iu_cc, read_iu, read_fp_cc,
			read_iu_cc_reg, read_iu_reg, read_fp_cc_reg)
		variable data_from_iu_cc_var: std_logic_vector(16 downto 0);
		variable data_from_fp_cc_var: std_logic_vector(14 downto 0);
		variable data_from_iu_var: std_logic_vector(89 downto 0);

	begin
		if(read_iu_cc_reg) then
			data_from_iu_cc_var := data_from_iu_cc;
		else	
			data_from_iu_cc_var := (others => '0');
		end if;
		if(read_fp_cc_reg) then
			data_from_fp_cc_var := data_from_fp_cc;
		else	
			data_from_fp_cc_var := (others => '0');
		end if;
		if(read_iu_reg) then
			data_from_iu_var := data_from_iu;
		else	
			data_from_iu_var := (others => '0');
		end if;

		other_data <= data_from_iu_cc_var & data_from_iu_var & data_from_fp_cc_var;

	end process;


	-- registers.
	process (clk)
	begin
		if(clk'event and (clk = '1') ) then
			if(latch_dispatch_data ) then
				data_from_dispatch_reg <= data_from_dispatch;
			elsif (clear_dispatch_data) then
				data_from_dispatch_reg <= (others => '0');
			end if;
			if(latch_other_data) then
				other_data_reg <= other_data;
			elsif (clear_other_data) then
				other_data_reg <= (others => '0');
			end if;
		end if;
	end process;

	-- Zero delay works well.  Need to confirm with synth.
	qbDispatch: QueueBase
		generic map (name => "sc_in_mux_qbDispatch", queue_depth => 0, data_width => 204)
		port map (
			clk => clk, reset => reset,
			data_in => teu_idispatch_to_stream_corrector_pipe_read_data,
			push_req => teu_idispatch_to_stream_corrector_pipe_read_ack(0),
			push_ack => teu_idispatch_to_stream_corrector_pipe_read_req(0),
			data_out => data_from_dispatch,
			pop_req  => pop_req_to_dispatch,
			pop_ack  => pop_ack_from_dispatch);

	-- bypass..  registered downstream..
	qbIUCC: QueueWithBypass
		generic map (name => "sc_in_mux_qbIUCC", queue_depth => 2, data_width => 17)
		port map (
			clk => clk, reset => reset,
			data_in => teu_iunit_cc_to_stream_corrector_pipe_read_data,
			push_req => teu_iunit_cc_to_stream_corrector_pipe_read_ack(0),
			push_ack => teu_iunit_cc_to_stream_corrector_pipe_read_req(0),
			data_out => data_from_iu_cc,
			pop_req  => pop_req_to_iu_cc,
			pop_ack  => pop_ack_from_iu_cc);

	-- bypass, registered down-stream
	qbIU: QueueWithBypass
		generic map (name => "sc_in_mux_qbIU", queue_depth => 1, data_width => 90)
		port map (
			clk => clk, reset => reset,
			data_in => teu_iunit_to_stream_corrector_pipe_read_data,
			push_req => teu_iunit_to_stream_corrector_pipe_read_ack(0),
			push_ack => teu_iunit_to_stream_corrector_pipe_read_req(0),
			data_out => data_from_iu,
			pop_req  => pop_req_to_iu,
			pop_ack  => pop_ack_from_iu);

	-- bypass, registered downstream.
	qbFPCC: QueueWithBypass
		generic map (name => "sc_in_mux_qbFPCC", queue_depth => 2, data_width => 15)
		port map (
			clk => clk, reset => reset,
			data_in => teu_fpunit_cc_to_stream_corrector_pipe_read_data,
			push_req => teu_fpunit_cc_to_stream_corrector_pipe_read_ack(0),
			push_ack => teu_fpunit_cc_to_stream_corrector_pipe_read_req(0),
			data_out => data_from_fp_cc,
			pop_req  => pop_req_to_fp_cc,
			pop_ack  => pop_ack_from_fp_cc);

	-- destination side..
	dest_rdy   <= (noblock_stream_corrector_in_args_pipe_write_ack(0) = '1'); 
	noblock_stream_corrector_in_args_pipe_write_req(0) <= '1' when write_to_dest else '0';
	noblock_stream_corrector_in_args_pipe_write_data <= 
		(const_one_sig & data_from_dispatch_reg & other_data_reg) when (fsm_state = WaitOnDestination) 
			else (const_one_sig & data_from_dispatch_reg & other_data);

end stream_corrector_in_mux_daemon_arch;

-- VHDL global package produced by vc2vhdl from virtual circuit (vc) description 
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library ahir;
use ahir.BaseComponents.all;
use ahir.mem_component_pack.all;

library AjitCustom;

entity bpbV2_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    bpb_init : in  std_logic_vector(0 downto 0);
    add_entry : in  std_logic_vector(0 downto 0);
    add_pc : in  std_logic_vector(31 downto 0);
    add_nnpc : in  std_logic_vector(31 downto 0);
    lookup_pc : in  std_logic_vector(31 downto 0);
    bpb_result : out  std_logic_vector(32 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity bpbV2_Operator;
architecture bpbV2_Operator_arch of bpbV2_Operator is -- 

    signal mem_write_address: std_logic_vector(7 downto 0);
    signal mem_write_data, ignore_data_0: std_logic_vector(51 downto 0);
    signal mem_write_enable, mem_write_enable_bar: std_logic;

    signal mem_read_address: std_logic_vector(7 downto 0);
    signal mem_read_address_delayed: std_logic_vector(7 downto 0);
    signal mem_read_data, zero_data_1: std_logic_vector(51 downto 0);
    signal mem_read_enable: std_logic;

    signal valids: std_logic_vector(255 downto 0);

    signal joined_sig: Boolean;
    signal trigger: std_logic;

    signal lookup_pc_tag: std_logic_vector(21 downto 0);
    signal trigger_reg  : std_logic;


    signal const_one : std_logic;
  
    signal bpb_result_prereg, bpb_result_reg : std_logic_vector(32 downto 0);
    signal write_read_clash, write_read_clash_reg : boolean;

begin --  
    zero_data_1 <= (others => '0');
    const_one <= '1';


    trigger <= '1' when joined_sig else '0';

    trig_join: join2 generic map (name => "bpbV2:trig-join", bypass => true)
			port map (pred0 => sample_req, pred1 => update_req,
					symbol_out => joined_sig, clk => clk, reset => reset);
   
    sample_ack <= joined_sig;

    process(clk, reset)
    begin
	if(clk'event and clk='1') then
		if(reset = '1') then
			update_ack <= false;
			trigger_reg <= '0';
			write_read_clash_reg <= false;
		else

			mem_read_address_delayed <= mem_read_address;

			lookup_pc_tag <= lookup_pc(31 downto 10);
			update_ack <= joined_sig;
	
			trigger_reg <= trigger;
			write_read_clash_reg <= write_read_clash;
		end if;
	end if;
    end process;

    mem_write_address <= add_pc (9 downto 2);
    mem_write_data    <= add_pc (31 downto 10) & add_nnpc (31 downto 2);
    mem_write_enable  <= (not bpb_init(0)) and trigger and add_entry(0);
    mem_write_enable_bar <= not mem_write_enable;

    mem_read_address  <= lookup_pc (9 downto 2);
    mem_read_enable   <= (not bpb_init(0)) and trigger;

    write_read_clash <= joined_sig and (mem_write_address = mem_read_address);

    process(clk, reset)
    begin
        if(clk'event and (clk='1')) then
		if((reset = '1') or ((trigger = '1') and (bpb_init(0) = '1'))) then
			valids <= (others => '0');
		else
			if ((trigger = '1') and (add_entry(0) = '1')) then
				valids(to_integer(unsigned(mem_write_address))) <= '1';
			end if;
		end if;
	end if;
    end process;
     
    dpram: base_bank_dual_port
		generic map (name =>  "bpbV2:dpram",
				g_addr_width => 8,
					g_data_width => 52)
		port map (
			datain_0 => mem_write_data,
			dataout_0 => ignore_data_0,
			addrin_0 => mem_write_address,
			enable_0 => mem_write_enable,
			writebar_0 => mem_write_enable_bar,
			datain_1 => zero_data_1,
			dataout_1 => mem_read_data,
			addrin_1 => mem_read_address,
			enable_1   => mem_read_enable,
			writebar_1 => const_one,
			clk => clk , reset => reset);
			

	process(valids, trigger_reg, mem_read_address_delayed, mem_read_data, lookup_pc_tag)
		variable result_var: std_logic_vector(32 downto 0);
	begin
		result_var := (others => '0');
		if((valids(to_integer(unsigned(mem_read_address_delayed))) = '1') and
			(mem_read_data(51 downto 30) = lookup_pc_tag) and (not write_read_clash_reg)) then
			result_var(32) := trigger_reg;
		else
			result_var(32) := '0';
		end if;
		result_var(31 downto 2) := mem_read_data(29 downto 0);

		bpb_result_prereg <= result_var;
	end process;

	-- Important: need to maintain the bpb result until the next trigger..
	process(clk, reset)
	begin
		if(clk'event and clk = '1') then
			if(reset = '1') then
				bpb_result_reg <= (others => '0');
			elsif (trigger_reg = '1') then
				bpb_result_reg <= bpb_result_prereg;
			end if;
		end if;
	end process;
	bpb_result <= bpb_result_prereg when (trigger_reg = '1') else bpb_result_reg;

end bpbV2_Operator_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


library ahir;
use ahir.mem_component_pack.all;
use ahir.basecomponents.all;

entity bpbV3_dual_port_mem_Operator is -- 
  port ( -- 
    init : in  std_logic_vector(0 downto 0);
    enable_0 : in  std_logic_vector(0 downto 0);
    addr_0 : in  std_logic_vector(7 downto 0);
    enable_1 : in  std_logic_vector(0 downto 0);
    write_bar_1 : in  std_logic_vector(0 downto 0);
    addr_1 : in  std_logic_vector(7 downto 0);
    write_data_1 : in  std_logic_vector(53 downto 0);
    read_data : out  std_logic_vector(109 downto 0);
    clk : in std_logic;
    reset : in std_logic;
    sample_req : in Boolean;
    sample_ack : out Boolean;
    update_req : in Boolean;
    update_ack   : out Boolean-- 
  );
  -- 
end entity bpbV3_dual_port_mem_Operator;

architecture bpbV3_dual_port_mem_arch of bpbV3_dual_port_mem_Operator is -- 
    signal valids: std_logic_vector(255 downto 0);
    signal Z54, read_data_0, read_data_1 : std_logic_vector(53 downto 0);

    signal joined_sig: Boolean;
    signal trigger, trigger_reg: Boolean;

    signal One1: std_logic_vector(0 downto 0);
    signal valid_0, valid_1: std_logic_vector(0 downto 0);
    signal read_data_prereg, read_data_reg : std_logic_vector(109 downto 0);

begin --  

    One1(0)  <= '1';

    Z54 <= (others => '0');

    trigger <= joined_sig;

    trig_join: join2 generic map (name => "bpbV2:trig-join", bypass => true)
			port map (pred0 => sample_req, pred1 => update_req,
					symbol_out => joined_sig, clk => clk, reset => reset);
   
    sample_ack <= joined_sig;

    process(clk, reset)
    begin
	if(clk'event and clk='1') then
		if(reset = '1') then
			update_ack <= false;
			trigger_reg <= false;
		else
			update_ack <= joined_sig;
			trigger_reg <= trigger;
		end if;
	end if;
    end process;

    -- valids extraction..
    process(clk, reset)
    begin
	if(clk'event and clk='1') then
		if((reset = '1')  or (init(0) = '1')) then
			valid_0(0) <= '0';
			valid_1(0) <= '0';
			valids <= (others => '0');
		else

			if(trigger and (enable_0(0) = '1')) then
				valid_0(0) <= valids (to_integer(unsigned(addr_0)));
			end if;
		
			if(trigger and (enable_1(0) = '1')) then
			    if (write_bar_1(0) = '0') then
				valids(to_integer(unsigned(addr_1))) <= '1';
			    else 
			        valid_1(0) <= valids (to_integer(unsigned(addr_1)));
			    end if;
			end if;
		end if;
	end if;
    end process;

    -- dual port mem.
    dpram: base_bank_dual_port
		generic map (name =>  "bpbV3:dpram",
				g_addr_width => 8,
					g_data_width => 54)
		port map (
			datain_0 => Z54,
			dataout_0 => read_data_0,
			addrin_0 => addr_0,
			enable_0 => enable_0(0),
			writebar_0 => One1(0),
			datain_1 => write_data_1,
			dataout_1 => read_data_1,
			addrin_1 => addr_1,
			enable_1   => enable_1(0),
			writebar_1 => write_bar_1(0),
			clk => clk , reset => reset);
			

   read_data_prereg <= valid_0 & read_data_0 & valid_1 & read_data_1;
   process(clk, reset)
   begin
	if(clk'event and clk = '1') then
		if(trigger_reg) then
			read_data_reg <= read_data_prereg;
		end if;
	end if;
   end process;
   read_data <= read_data_prereg when trigger_reg else read_data_reg;

end bpbV3_dual_port_mem_arch;
-- VHDL global package produced by vc2vhdl from virtual circuit (vc) description 
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library ahir;
use ahir.BaseComponents.all;
use ahir.mem_component_pack.all;

library AjitCustom;
use AjitCustom.AjitCoreConfigurationPackage.all; 

entity ibuf_cache_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    ibuf_cache_init : in  std_logic_vector(0 downto 0);
    add_entry : in  std_logic_vector(0 downto 0);
    add_pc : in  std_logic_vector(31 downto 0);
    add_acc : in  std_logic_vector(2 downto 0);
    add_ipair : in  std_logic_vector(63 downto 0);
    lookup_S : in  std_logic_vector(0 downto 0);
    lookup_pc : in  std_logic_vector(31 downto 0);
    ibuf_cache_result : out  std_logic_vector(64 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity ibuf_cache_Operator;
architecture ibuf_cache_Operator_arch of ibuf_cache_Operator is -- 

    constant data_width: integer := IBUF_CACHE_TAG_WIDTH + 67;

    function ibufPermissionsOk (S: std_logic; acc: std_logic_vector(2 downto 0)) 
	return boolean is
	variable ret_var: boolean;
	variable acc_int: integer range 0 to 7;
    begin
	acc_int := to_integer (unsigned(acc));
	ret_var := ((acc_int > 2) and (acc_int < 5)) or
			((S = '1') and (acc_int > 5));
	return(ret_var);
    end function;

    signal mem_write_address: std_logic_vector(LOG_IBUF_CACHE_SIZE-1 downto 0);
    signal mem_write_data, ignore_data_0: std_logic_vector(data_width-1 downto 0);
    signal mem_write_enable, mem_write_enable_bar: std_logic;

    signal mem_read_address: std_logic_vector(LOG_IBUF_CACHE_SIZE-1 downto 0);
    signal mem_read_address_delayed: std_logic_vector(LOG_IBUF_CACHE_SIZE-1 downto 0);
    signal mem_read_data, zero_data_1: std_logic_vector(data_width-1 downto 0);
    signal mem_read_enable: std_logic;

    signal valids: std_logic_vector(IBUF_CACHE_SIZE-1 downto 0);

    signal joined_sig: Boolean;
    signal trigger: std_logic;

    signal lookup_pc_tag: std_logic_vector(IBUF_CACHE_TAG_WIDTH-1 downto 0);
    signal trigger_reg  : std_logic;


    signal const_one : std_logic;
  
    signal ibuf_cache_result_prereg, ibuf_cache_result_reg : std_logic_vector(64 downto 0);
    signal write_read_clash, write_read_clash_reg : boolean;

begin --  
    zero_data_1 <= (others => '0');
    const_one <= '1';


    trigger <= '1' when joined_sig else '0';

    trig_join: join2 generic map (name => "ibuf_cache:trig-join", bypass => true)
			port map (pred0 => sample_req, pred1 => update_req,
					symbol_out => joined_sig, clk => clk, reset => reset);
   
    sample_ack <= joined_sig;

    process(clk, reset)
    begin
	if(clk'event and clk='1') then
		if(reset = '1') then
			update_ack <= false;
			trigger_reg <= '0';
			write_read_clash_reg <= false;
		else

			mem_read_address_delayed <= mem_read_address;

			lookup_pc_tag <= lookup_pc(31 downto (3 + LOG_IBUF_CACHE_SIZE));
			update_ack <= joined_sig;
	
			trigger_reg <= trigger;
			write_read_clash_reg <= write_read_clash;
		end if;
	end if;
    end process;

    -- index into memory..
    mem_write_address <= add_pc ((3 + LOG_IBUF_CACHE_SIZE -1) downto 3);

    -- tag acc ipair.
    mem_write_data    <= add_pc (31 downto (3 + LOG_IBUF_CACHE_SIZE)) & add_acc & add_ipair;
    mem_write_enable  <= (not ibuf_cache_init(0)) and trigger and add_entry(0);
    mem_write_enable_bar <= not mem_write_enable;

    -- index into memory..
    mem_read_address  <= lookup_pc ((3 + LOG_IBUF_CACHE_SIZE -1) downto 3);
    mem_read_enable   <= (not ibuf_cache_init(0)) and trigger;

    write_read_clash <= joined_sig and (mem_write_address = mem_read_address);

    process(clk, reset)
    begin
        if(clk'event and (clk='1')) then
		if((reset = '1') or ((trigger = '1') and (ibuf_cache_init(0) = '1'))) then
			valids <= (others => '0');
		else
			if ((trigger = '1') and (add_entry(0) = '1')) then
				valids(to_integer(unsigned(mem_write_address))) <= '1';
			end if;
		end if;
	end if;
    end process;
     
    dpram: base_bank_dual_port
		generic map (name =>  "ibuf_cache:dpram",
				g_addr_width => LOG_IBUF_CACHE_SIZE,
					g_data_width => data_width)
		port map (
			datain_0 => mem_write_data,
			dataout_0 => ignore_data_0,
			addrin_0 => mem_write_address,
			enable_0 => mem_write_enable,
			writebar_0 => mem_write_enable_bar,
			datain_1 => zero_data_1,
			dataout_1 => mem_read_data,
			addrin_1 => mem_read_address,
			enable_1   => mem_read_enable,
			writebar_1 => const_one,
			clk => clk , reset => reset);
			

	process(valids, trigger_reg, mem_read_address_delayed, mem_read_data, lookup_pc_tag)
		variable result_var: std_logic_vector(64 downto 0);
	begin
		result_var := (others => '0');
		if((valids(to_integer(unsigned(mem_read_address_delayed))) = '1') and
			(mem_read_data((IBUF_CACHE_TAG_WIDTH + 66) downto 67) = lookup_pc_tag) and (not write_read_clash_reg)
				and ibufPermissionsOk (lookup_S(0), mem_read_data (66 downto 64))) then
			result_var(64) := trigger_reg;
		else
			result_var(64) := '0';
		end if;
		result_var(63 downto 0) := mem_read_data(63 downto 0);

		ibuf_cache_result_prereg <= result_var;
	end process;

	-- Important: need to maintain the ibuf_cache result until the next trigger..
	process(clk, reset)
	begin
		if(clk'event and clk = '1') then
			if(reset = '1') then
				ibuf_cache_result_reg <= (others => '0');
			elsif (trigger_reg = '1') then
				ibuf_cache_result_reg <= ibuf_cache_result_prereg;
			end if;
		end if;
	end process;
	ibuf_cache_result <= ibuf_cache_result_prereg when (trigger_reg = '1') else ibuf_cache_result_reg;

end ibuf_cache_Operator_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library ahir;
use ahir.mem_component_pack.all;
library AjitCustom;
use AjitCustom.AjitCoreConfigurationPackage.all;
entity ras_daemon is -- 
  generic (tag_length : integer := 1); 
  port ( -- 
    teu_ras_access_pipe_pipe_read_req : out  std_logic_vector(0 downto 0);
    teu_ras_access_pipe_pipe_read_ack : in   std_logic_vector(0 downto 0);
    teu_ras_access_pipe_pipe_read_data : in   std_logic_vector(32 downto 0);
    teu_ras_top_of_stack_pipe_write_req : out  std_logic_vector(0 downto 0);
    teu_ras_top_of_stack_pipe_write_ack : in   std_logic_vector(0 downto 0);
    teu_ras_top_of_stack_pipe_write_data : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity ras_daemon;
architecture ras_daemon_arch of ras_daemon is -- 

	signal push, pop, flush, command_available, command_available_reg, valid_bit: std_logic;
	signal valids: std_logic_vector (RAS_DEPTH-1 downto 0);
	
	signal mem_address: std_logic_vector (LOG_RAS_DEPTH-1 downto 0);
	signal mem_enable, mem_enable_reg: std_logic;
	signal mem_write_bar, mem_write_bar_reg : std_logic;
	signal mem_write_data, mem_read_data, mem_read_data_reg: std_logic_vector(29 downto 0);


	-- maintains the top of the stack..
	signal top_of_stack_pointer: unsigned(LOG_RAS_DEPTH-1 downto 0);
	
    	signal pop_data_qualified, push_data_qualified : std_logic_vector(31 downto 0);

	signal last_is_pop, last_is_push, last_is_flush: std_logic;
	signal command_reg: std_logic_vector(32 downto 0);
	constant ZZ: unsigned(LOG_RAS_DEPTH-1 downto 0) := (others => '0');
	constant OO: unsigned(LOG_RAS_DEPTH-1 downto 0) := (others => '1');
begin --  

	tag_out <= (others => '0');
	start_ack <= '1';
	fin_ack <= '0';

	command_available <= teu_ras_access_pipe_pipe_read_ack(0);

	-- always ready to read!
	teu_ras_access_pipe_pipe_read_req(0) <= '1';
	
	-- commands.	
	push <= command_available and teu_ras_access_pipe_pipe_read_data(32);
	pop  <= command_available and teu_ras_access_pipe_pipe_read_data(31);
	flush  <= command_available and teu_ras_access_pipe_pipe_read_data(30);

	-- mem written from access command.
	mem_write_data <= teu_ras_access_pipe_pipe_read_data(29 downto 0);
	mem_enable <= (not flush) and (push or pop);
	mem_write_bar <= (flush or (not push));

	
	process(clk, reset, command_available, valids, valid_bit,
			top_of_stack_pointer,
			push, pop, flush, teu_ras_access_pipe_pipe_read_data,
			mem_enable,mem_write_bar, mem_enable_reg, mem_write_bar_reg,
			mem_read_data) 
		variable next_last_is_push, next_last_is_pop, next_last_is_flush: std_logic;
		variable next_top_of_stack_pointer : unsigned(LOG_RAS_DEPTH-1 downto 0);
		variable next_valids: std_logic_vector (RAS_DEPTH-1 downto 0);
		variable next_valid_bit: std_logic;
		variable mem_address_var: std_logic_vector (LOG_RAS_DEPTH-1 downto 0);
	begin
		next_last_is_push := last_is_push;
		next_last_is_pop := last_is_pop;
		next_last_is_flush := last_is_flush;
		next_top_of_stack_pointer := top_of_stack_pointer;
		next_valids := valids;
		next_valid_bit := valid_bit;
		mem_address_var := (others => '0');
				
		if(flush = '1') then
			next_valids := (others => '0');
			next_top_of_stack_pointer := OO;
			next_last_is_push := '0';
			next_last_is_pop  := '0';
			next_last_is_flush := '1';
			next_valid_bit := '0';
		elsif(push = '1') then
			next_last_is_push := '1';
			next_last_is_pop  := '0';
			next_last_is_flush := '0';
			next_valid_bit := '1';

			-- increment top of stack..
			if(top_of_stack_pointer = OO) then
				next_top_of_stack_pointer := ZZ;
			else 
				next_top_of_stack_pointer := top_of_stack_pointer + 1;
			end if;

			-- write to incremented slot.
			next_valids(to_integer(next_top_of_stack_pointer)) := '1';
			mem_address_var := std_logic_vector(next_top_of_stack_pointer);

		elsif (pop = '1') then

			next_last_is_push := '0';
			next_last_is_pop  := '1';
			next_last_is_flush := '0';

			-- clear the valid for the top of stack...
			next_valids(to_integer(top_of_stack_pointer)) := '0';

			-- decrement top of stack..
			if(top_of_stack_pointer = ZZ) then
				next_top_of_stack_pointer := OO;
			else 
				next_top_of_stack_pointer := top_of_stack_pointer - 1;
			end if;

			-- capture validity of new top of stack?
			next_valid_bit := valids(to_integer(next_top_of_stack_pointer));
	
			--
			-- new top of stack data read using address as  decremented top of stack
			--
			mem_address_var := std_logic_vector(next_top_of_stack_pointer);
		end if;


		mem_address <= mem_address_var;
		if(clk'event and clk = '1') then
			if(reset = '1') then
				valids <= (others => '0');

				last_is_pop <= '0';
				last_is_push <= '0';
				last_is_flush <= '1';

				command_available_reg <= '0';
				valid_bit <= '0';

				top_of_stack_pointer <= ZZ;

				mem_enable_reg <='0';
				mem_write_bar_reg <= '1';
			else
				mem_enable_reg <= mem_enable;
				mem_write_bar_reg <= mem_write_bar;

				valids <= next_valids;
				valid_bit <= next_valid_bit;

				command_available_reg <= command_available;

				last_is_pop <= next_last_is_pop;
				last_is_push <= next_last_is_push;
				last_is_flush <= next_last_is_flush;

				if(command_available = '1') then 
					command_reg <= teu_ras_access_pipe_pipe_read_data;
				end if;

				top_of_stack_pointer <= next_top_of_stack_pointer;

				if((mem_enable_reg = '1') and (mem_write_bar_reg = '1')) then
					mem_read_data_reg <= mem_read_data;
				end if;
			end if;
		end if;
	end process;

	bb: base_bank
		generic map (name => "RAS-BB", g_addr_width => LOG_RAS_DEPTH, g_data_width => 30)
		port map (clk => clk, reset => reset,
					datain => mem_write_data,
					dataout => mem_read_data,
					addrin => mem_address,
					enable => mem_enable,
					writebar => mem_write_bar);
		
	-- hold for one cycle, when memory access has completed.
	teu_ras_top_of_stack_pipe_write_req(0) <= last_is_push or last_is_pop or last_is_flush; 	
	teu_ras_top_of_stack_pipe_write_data 	
				<= push_data_qualified when (last_is_push = '1')
					 else pop_data_qualified when (last_is_pop = '1')  else (others => '0');

	-- push data.. from command, but with valid bit attached.
	push_data_qualified(31 downto 2) <= command_reg (29 downto 0);
	push_data_qualified(1) <= '0';
	push_data_qualified(0) <= valid_bit;


	-- pop data.. from memory, with valid bit attached.
	pop_data_qualified(31 downto 2) <= 
		mem_read_data(29 downto 0) when ((mem_enable_reg = '1') and (mem_write_bar_reg = '1')) 
									else mem_read_data_reg(29 downto 0);
	pop_data_qualified(1) <= '0';
	pop_data_qualified(0) <= valid_bit;


end ras_daemon_arch;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity ahb_splitter is -- 
    -- address range is specified for upper memory and for lower
    -- memory.  Address is not modified on the way out.  Addresses
    -- that do not fall in either range are just ignored.
    generic (
		UPPER_ADDRESS_LOWER_BOUND, UPPER_ADDRESS_UPPER_BOUND: integer;
		LOWER_ADDRESS_LOWER_BOUND, LOWER_ADDRESS_UPPER_BOUND: integer);
    port( -- 

  -- main input.. will be split..
      main_HADDR : in std_logic_vector(31 downto 0);
  -- ignored.
      main_HMASTLOCK : in std_logic;
  -- ignored.
      main_HPROT : in std_logic_vector(3 downto 0); 
  -- ignored.
      main_HBURST : in std_logic_vector(2 downto 0); 
  -- ignored.. all accesses are 32-bits wide.
      main_HSIZE : in std_logic_vector(2 downto 0);
   -- should be NONSEQ or SEQ to indicate transfer
      main_HTRANS : in std_logic_vector(1 downto 0);
  -- write data
      main_HWDATA : in std_logic_vector(31 downto 0); 
  -- "1" implies write
      main_HWRITE : in std_logic;
  -- read data
      main_HRDATA : out std_logic_vector(31 downto 0); 
  -- always "1".
      main_HREADY : out std_logic;
  -- response.
      main_HRESP : out std_logic_vector(1 downto 0); -- always "00"

  -- upper addr..
      upper_HADDR : out std_logic_vector(31 downto 0);
  -- ignored.
      upper_HMASTLOCK : out std_logic;
  -- ignored.
      upper_HPROT : out std_logic_vector(3 downto 0); 
  -- ignored.
      upper_HBURST : out std_logic_vector(2 downto 0); 
  -- ignored.. all accesses are 32-bits wide.
      upper_HSIZE : out std_logic_vector(2 downto 0);
   -- should be NONSEQ or SEQ to indicate transfer
      upper_HTRANS : out std_logic_vector(1 downto 0);
  -- write data
      upper_HWDATA : out std_logic_vector(31 downto 0); 
  -- "1" implies write
      upper_HWRITE : out std_logic;
  -- read data
      upper_HRDATA : in std_logic_vector(31 downto 0); 
  -- always "1".
      upper_HREADY : in std_logic;
  -- response.
      upper_HRESP : in std_logic_vector(1 downto 0); -- always "00"

  -- lower addr..
      lower_HADDR : out std_logic_vector(31 downto 0);
  -- ignored.
      lower_HMASTLOCK : out std_logic;
  -- ignored.
      lower_HPROT : out std_logic_vector(3 downto 0); 
  -- ignored.
      lower_HBURST : out std_logic_vector(2 downto 0); 
  -- ignored.. all accesses are 32-bits wide.
      lower_HSIZE : out std_logic_vector(2 downto 0);
   -- should be NONSEQ or SEQ to indicate transfer
      lower_HTRANS : out std_logic_vector(1 downto 0);
  -- write data
      lower_HWDATA : out std_logic_vector(31 downto 0); 
  -- "1" implies write
      lower_HWRITE : out std_logic;
  -- read data
      lower_HRDATA : in std_logic_vector(31 downto 0); 
  -- always "1".
      lower_HREADY : in std_logic;
  -- response.
      lower_HRESP : in std_logic_vector(1 downto 0); -- always "00"
  -- positive edge of clock is used, reset is active high.
      clk, reset: in std_logic 
    );
end entity;


--
-- a simple interface.. serves single/burst requests..
--   it is assumed that the host never goes into a busy cycle.
--
architecture Mixed of ahb_splitter is

  constant HTRANS_IDLE : std_logic_vector(1 downto 0) := "00";
  constant HTRANS_BUSY : std_logic_vector(1 downto 0) := "01";
  constant HTRANS_NONSEQ : std_logic_vector(1 downto 0) := "10";
  constant HTRANS_SEQ : std_logic_vector(1 downto 0) := "11";
  constant HSIZE_1   : std_logic_vector(2 downto 0)  := "000"; -- 1-byte transfer
  constant HSIZE_2   : std_logic_vector(2 downto 0)  := "001"; -- 2-byte transfer
  constant HSIZE_4   : std_logic_vector(2 downto 0)  := "010"; -- 4-byte transfer
  constant HSIZE_8   : std_logic_vector(2 downto 0)  := "011"; -- 8-byte transfer

  constant HBURST_SINGLE   : std_logic_vector(2 downto 0)  := "000"; -- 8-byte transfer
  constant SLAVE_RESPONSE_OK   : std_logic_vector(1 downto 0)  := "00"; -- OK
  constant SLAVE_RESPONSE_ERROR   : std_logic_vector(1 downto 0)  := "01"; -- Error
    
  type FsmState is (LatchRequestState, RequestState, RequestSentState);
  signal fsm_state: FsmState;

  signal upper_half_selected: std_logic;
  signal upper_half_selected_reg: std_logic;

  signal lower_half_selected: std_logic;
  signal lower_half_selected_reg: std_logic;

  signal latch_request, latch_hwdata: std_logic;
      
   -- registered main request.
  signal HADDR_reg :  std_logic_vector(31 downto 0);
  signal HMASTLOCK_reg : std_logic;
  signal HPROT_reg : std_logic_vector(3 downto 0); 
  signal HBURST_reg : std_logic_vector(2 downto 0); 
  signal HSIZE_reg : std_logic_vector(2 downto 0);
  signal HTRANS_reg : std_logic_vector(1 downto 0);
  signal HWDATA_reg : std_logic_vector(31 downto 0); 
  signal HWRITE_reg : std_logic;

begin 
  upper_half_selected <= '1' when  
      (to_integer(unsigned(main_HADDR)) >=  UPPER_ADDRESS_LOWER_BOUND) and
      (to_integer(unsigned(main_HADDR)) <=  UPPER_ADDRESS_UPPER_BOUND) 
        else '0';
  lower_half_selected <= '1' when  
      (to_integer(unsigned(main_HADDR)) >=  LOWER_ADDRESS_LOWER_BOUND) and
      (to_integer(unsigned(main_HADDR)) <=  LOWER_ADDRESS_UPPER_BOUND) 
	else '0';

  -- registers
  process(clk, reset)
  begin
    if (clk'event and (clk='1')) then
	if (reset = '1') then
		upper_half_selected_reg <= '0';	
		lower_half_selected_reg <= '0';	
	elsif latch_request = '1' then
  		HADDR_reg  <= main_HADDR;
        	HMASTLOCK_reg <= main_HMASTLOCK;
        	HPROT_reg <= main_HPROT;
        	HBURST_reg <= main_HBURST;
        	HSIZE_reg <= main_HSIZE;
        	HTRANS_reg <= main_HTRANS;
        	HWRITE_reg <= main_HWRITE;

		upper_half_selected_reg <= upper_half_selected;
		lower_half_selected_reg <= lower_half_selected;
	end if;

	if latch_hwdata = '1' then
		HWDATA_reg <= main_HWDATA;
	end if;
    end if;
  end process;


  -- state machine.
  process(clk, reset, 
	    -- fsm state.
	    fsm_state,  
	    -- main side request
            main_HADDR,
            main_HMASTLOCK,
            main_HPROT,
            main_HBURST,
            main_HSIZE,
            main_HTRANS,
            main_HWDATA,
            main_HWRITE,
            -- upper side responses
            upper_HRDATA,
            upper_HREADY,
            upper_HRESP,
            -- lower side responses
            lower_HRDATA,
            lower_HREADY,
            lower_HRESP,
	    -- which half is active?
     	    upper_half_selected, 
	    upper_half_selected_reg,
     	    lower_half_selected, 
	    lower_half_selected_reg
	)

    variable next_fsm_state : FsmState;
    variable latch_request_var: std_logic;
  
    variable upper_HADDR_var :  std_logic_vector(31 downto 0);
    variable upper_HMASTLOCK_var : std_logic;
    variable upper_HPROT_var : std_logic_vector(3 downto 0); 
    variable upper_HBURST_var : std_logic_vector(2 downto 0); 
    variable upper_HSIZE_var : std_logic_vector(2 downto 0);
    variable upper_HTRANS_var : std_logic_vector(1 downto 0);
    variable upper_HWDATA_var : std_logic_vector(31 downto 0); 
    variable upper_HWRITE_var : std_logic;

    variable lower_HADDR_var :  std_logic_vector(31 downto 0);
    variable lower_HMASTLOCK_var : std_logic;
    variable lower_HPROT_var : std_logic_vector(3 downto 0); 
    variable lower_HBURST_var : std_logic_vector(2 downto 0); 
    variable lower_HSIZE_var : std_logic_vector(2 downto 0);
    variable lower_HTRANS_var : std_logic_vector(1 downto 0);
    variable lower_HWDATA_var : std_logic_vector(31 downto 0); 
    variable lower_HWRITE_var : std_logic;

    variable main_HRESP_var  : std_logic_vector(1 downto 0);
    variable main_HREADY_var : std_logic;
    variable main_HRDATA_var : std_logic_vector(31 downto 0);

    variable slave_response_ready_var : boolean;
    variable slave_is_ready_var : boolean;

    variable next_latch_hwdata_var: std_logic;

  begin
    next_fsm_state := fsm_state;

    latch_request_var := '0';
    next_latch_hwdata_var  := '0';

    slave_response_ready_var := false;
    slave_is_ready_var := false;

    main_HREADY_var  := '0';
    main_HRESP_var := SLAVE_RESPONSE_OK;
    main_HRDATA_var := (others => '0');

    upper_HTRANS_var := HTRANS_IDLE;
    upper_HMASTLOCK_var :=  '0';
    upper_HSIZE_var := HSIZE_4;
    upper_HBURST_var := HBURST_SINGLE;
    upper_HPROT_var  := (others => '0');
    upper_HWDATA_var  := (others => '0');
    upper_HWRITE_var  := '0';
    upper_HADDR_var := (others => '0');

    lower_HTRANS_var := HTRANS_IDLE;
    lower_HMASTLOCK_var :=  '0';
    lower_HSIZE_var := HSIZE_4;
    lower_HBURST_var := HBURST_SINGLE;
    lower_HPROT_var  := (others => '0');
    lower_HWDATA_var  := (others => '0');
    lower_HWRITE_var  := '0';
    lower_HADDR_var := (others => '0');


    case fsm_state is 
      when LatchRequestState =>
	main_HREADY_var := '1';
        -- if main request is valid then register the request.
	--   Note: only nonseq requests are entertained.
	--   Note: this is a dead state which reduces the throughput.
        if(main_HTRANS = HTRANS_NONSEQ) then
	  latch_request_var := '1';
	  next_latch_hwdata_var := '1';
	  next_fsm_state := RequestState;
	end if;
      when RequestState =>

          if (upper_half_selected_reg = '1') then
            upper_HTRANS_var := HTRANS_reg;
            upper_HWRITE_var := HWRITE_reg;
            upper_HSIZE_var  := HSIZE_reg;
            upper_HMASTLOCK_var := HMASTLOCK_reg;
	    upper_HADDR_var := HADDR_REG;
            if(upper_HREADY = '1') then
               slave_is_ready_var := true;
            end if;
          elsif (lower_half_selected_reg = '1') then
            lower_HTRANS_var := HTRANS_reg;
            lower_HWRITE_var := HWRITE_reg;
            lower_HSIZE_var  := HSIZE_reg;
            lower_HMASTLOCK_var := HMASTLOCK_reg;
	    lower_HADDR_var := HADDR_REG;
            if(lower_HREADY = '1') then
               slave_is_ready_var := true;
            end if;
	  else
               slave_is_ready_var := true;
          end if;

	  if slave_is_ready_var then
	     next_fsm_state := RequestSentState;
	     next_latch_hwdata_var := '1';
          end if;
      when RequestSentState => 
        if (upper_half_selected_reg = '1') then

          upper_HMASTLOCK_var := HMASTLOCK_reg;
          upper_HWDATA_var := HWDATA_reg;
	  upper_HADDR_var := HADDR_reg;

          main_HRESP_var   := upper_HRESP;
          main_HRDATA_var  := upper_HRDATA;

          if(upper_HREADY = '1') then
            slave_response_ready_var := true;
          end if;

        elsif (lower_half_selected_reg = '1') then

          lower_HMASTLOCK_var := HMASTLOCK_reg;
          lower_HWDATA_var := HWDATA_reg;
	  lower_HADDR_var := HADDR_reg;

          main_HRESP_var   := lower_HRESP;
          main_HRDATA_var  := lower_HRDATA;

          if(lower_HREADY = '1') then
            slave_response_ready_var := true;
          end if;
        else
            slave_response_ready_var := true;
        end if;

        if(slave_response_ready_var) then

	  main_HREADY_var := '1';

          if(main_HTRANS = HTRANS_NONSEQ) then
		latch_request_var := '1';
	  	next_latch_hwdata_var := '1';
		next_fsm_state := RequestState;
	  else
	  	next_fsm_state := LatchRequestState;
	  end if;

        end if;
    end case;

    upper_HTRANS <= upper_HTRANS_var;
    upper_HADDR <= upper_HADDR_var;
    upper_HWRITE <= upper_HWRITE_var;
    upper_HMASTLOCK <= upper_HMASTLOCK_var;
    upper_HSIZE <= upper_HSIZE_var;
    upper_HBURST <= upper_HBURST_var;
    upper_HPROT <= upper_HPROT_var;
    upper_HWDATA <= upper_HWDATA_var;

    lower_HTRANS <= lower_HTRANS_var;
    lower_HADDR <= lower_HADDR_var;
    lower_HWRITE <= lower_HWRITE_var;
    lower_HMASTLOCK <= lower_HMASTLOCK_var;
    lower_HSIZE <= lower_HSIZE_var;
    lower_HBURST <= lower_HBURST_var;
    lower_HPROT <= lower_HPROT_var;
    lower_HWDATA <= lower_HWDATA_var;
          
    main_HREADY <= main_HREADY_var;
    main_HRESP  <= main_HRESP_var;
    main_HRDATA <= main_HRDATA_var;

    latch_request <= latch_request_var;

    if(clk'event and clk = '1') then
      if(reset = '1') then
        fsm_state <= LatchRequestState;
    	latch_hwdata  <= '0';
      else
        fsm_state <= next_fsm_state;
    	latch_hwdata  <= next_latch_hwdata_var;
      end if;
    end if;
  end process;



end Mixed;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
entity memAccessRequestMergeDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    fast_mem_access_and_send_response_command_pipe_read_req : out  std_logic_vector(0 downto 0);
    fast_mem_access_and_send_response_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
    fast_mem_access_and_send_response_command_pipe_read_data : in   std_logic_vector(124 downto 0);
    slow_mem_access_and_send_response_command_pipe_read_req : out  std_logic_vector(0 downto 0);
    slow_mem_access_and_send_response_command_pipe_read_ack : in   std_logic_vector(0 downto 0);
    slow_mem_access_and_send_response_command_pipe_read_data : in   std_logic_vector(209 downto 0);
    mem_access_and_send_response_command_pipe_write_req : out  std_logic_vector(0 downto 0);
    mem_access_and_send_response_command_pipe_write_ack : in   std_logic_vector(0 downto 0);
    mem_access_and_send_response_command_pipe_write_data : out  std_logic_vector(207 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity memAccessRequestMergeDaemon;
architecture memAccessRequestMergeDaemon_arch of memAccessRequestMergeDaemon is -- 
  component mergeCommands_VVV is -- 
    port ( -- 
      fast_cmd : in  std_logic_vector(124 downto 0);
      slow_cmd : in  std_logic_vector(207 downto 0);
      merged_cmd : out  std_logic_vector(207 downto 0)-- 
    );
    -- 
  end component; 

  signal fast_valid, slow_needed, all_ready, slow_valid, rx_ready: boolean;
  signal merged_command: std_logic_vector(207 downto 0);
  signal command_counter : std_logic_vector(1 downto 0);
begin --  

	start_ack <= '1';
	fin_ack   <= '0';
	tag_out   <= (others => '0');

	command_counter <= slow_mem_access_and_send_response_command_pipe_read_data(209 downto 208);

	mc: mergeCommands_VVV
		port map (fast_cmd =>fast_mem_access_and_send_response_command_pipe_read_data ,
				slow_cmd => slow_mem_access_and_send_response_command_pipe_read_data(207 downto 0),
				 merged_cmd => merged_command);

	mem_access_and_send_response_command_pipe_write_data <=  merged_command;

	fast_valid  <= (fast_mem_access_and_send_response_command_pipe_read_ack(0) = '1');
	slow_needed <= fast_valid and (fast_mem_access_and_send_response_command_pipe_read_data(124) = '1');
	slow_valid  <= (slow_mem_access_and_send_response_command_pipe_read_ack(0) = '1');

	rx_ready  <= (mem_access_and_send_response_command_pipe_write_ack(0) = '1');
	all_ready <= (fast_valid and rx_ready and ((not slow_needed) or slow_valid));

	fast_mem_access_and_send_response_command_pipe_read_req(0) <= '1' when all_ready  else '0';
	slow_mem_access_and_send_response_command_pipe_read_req(0)  <= '1' when (slow_valid and all_ready) else '0';
	mem_access_and_send_response_command_pipe_write_req(0) <= '1' when all_ready else '0';
			
end memAccessRequestMergeDaemon_arch;

library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;

entity mergeCommands_VVV is -- 
  port ( -- 
    fast_cmd : in  std_logic_vector(124 downto 0);
    slow_cmd : in  std_logic_vector(207 downto 0);
    merged_cmd : out  std_logic_vector(207 downto 0)-- 
  );
  -- 
end entity mergeCommands_VVV;
architecture mergeCommands_VVV_arch of mergeCommands_VVV is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(333-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal fast_cmd_buffer :  std_logic_vector(124 downto 0);
  signal slow_cmd_buffer :  std_logic_vector(207 downto 0);
  -- output port buffer signals
  signal merged_cmd_buffer :  std_logic_vector(207 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  fast_cmd_buffer <= fast_cmd;
  slow_cmd_buffer <= slow_cmd;
  -- output handling  -------------------------------------------------------
  merged_cmd <= merged_cmd_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u12_u95_4802_wire : std_logic_vector(94 downto 0);
    signal CONCAT_u1_u2_4783_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_4806_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_4809_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u9_4788_wire : std_logic_vector(8 downto 0);
    signal CONCAT_u1_u9_4813_wire : std_logic_vector(8 downto 0);
    signal CONCAT_u2_u3_4785_wire : std_logic_vector(2 downto 0);
    signal CONCAT_u2_u4_4810_wire : std_logic_vector(3 downto 0);
    signal CONCAT_u33_u83_4800_wire_constant : std_logic_vector(82 downto 0);
    signal CONCAT_u36_u100_4816_wire : std_logic_vector(99 downto 0);
    signal CONCAT_u3_u12_4789_wire : std_logic_vector(11 downto 0);
    signal CONCAT_u4_u113_4818_wire : std_logic_vector(112 downto 0);
    signal CONCAT_u9_u109_4817_wire : std_logic_vector(108 downto 0);
    signal byte_mask_4771 : std_logic_vector(7 downto 0);
    signal default_cacheable_bit_4743 : std_logic_vector(0 downto 0);
    signal flags_4767 : std_logic_vector(7 downto 0);
    signal is_read_dword_4759 : std_logic_vector(0 downto 0);
    signal is_read_line_4763 : std_logic_vector(0 downto 0);
    signal is_write_dword_4755 : std_logic_vector(0 downto 0);
    signal lock_bus_4735 : std_logic_vector(0 downto 0);
    signal mmu_enabled_4739 : std_logic_vector(0 downto 0);
    signal physical_addr_to_mem_4775 : std_logic_vector(35 downto 0);
    signal reconstructed_fast_cmd_4820 : std_logic_vector(207 downto 0);
    signal send_response_4751 : std_logic_vector(0 downto 0);
    signal to_dcache_4747 : std_logic_vector(0 downto 0);
    signal type_cast_4804_wire_constant : std_logic_vector(0 downto 0);
    signal use_slow_4731 : std_logic_vector(0 downto 0);
    signal write_data_4779 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    CONCAT_u33_u83_4800_wire_constant <= "00000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    type_cast_4804_wire_constant <= "0";
    -- flow-through select operator MUX_4825_inst
    merged_cmd_buffer <= slow_cmd_buffer when (use_slow_4731(0) /=  '0') else reconstructed_fast_cmd_4820;
    -- flow-through slice operator slice_4730_inst
    use_slow_4731 <= fast_cmd_buffer(124 downto 124);
    -- flow-through slice operator slice_4734_inst
    lock_bus_4735 <= fast_cmd_buffer(123 downto 123);
    -- flow-through slice operator slice_4738_inst
    mmu_enabled_4739 <= fast_cmd_buffer(122 downto 122);
    -- flow-through slice operator slice_4742_inst
    default_cacheable_bit_4743 <= fast_cmd_buffer(121 downto 121);
    -- flow-through slice operator slice_4746_inst
    to_dcache_4747 <= fast_cmd_buffer(120 downto 120);
    -- flow-through slice operator slice_4750_inst
    send_response_4751 <= fast_cmd_buffer(119 downto 119);
    -- flow-through slice operator slice_4754_inst
    is_write_dword_4755 <= fast_cmd_buffer(118 downto 118);
    -- flow-through slice operator slice_4758_inst
    is_read_dword_4759 <= fast_cmd_buffer(117 downto 117);
    -- flow-through slice operator slice_4762_inst
    is_read_line_4763 <= fast_cmd_buffer(116 downto 116);
    -- flow-through slice operator slice_4766_inst
    flags_4767 <= fast_cmd_buffer(115 downto 108);
    -- flow-through slice operator slice_4770_inst
    byte_mask_4771 <= fast_cmd_buffer(107 downto 100);
    -- flow-through slice operator slice_4774_inst
    physical_addr_to_mem_4775 <= fast_cmd_buffer(99 downto 64);
    -- flow-through slice operator slice_4778_inst
    write_data_4779 <= fast_cmd_buffer(63 downto 0);
    -- binary operator CONCAT_u12_u95_4802_inst
    process(CONCAT_u3_u12_4789_wire) -- 
      variable tmp_var : std_logic_vector(94 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u3_u12_4789_wire, CONCAT_u33_u83_4800_wire_constant, tmp_var);
      CONCAT_u12_u95_4802_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_4783_inst
    process(mmu_enabled_4739, default_cacheable_bit_4743) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(mmu_enabled_4739, default_cacheable_bit_4743, tmp_var);
      CONCAT_u1_u2_4783_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_4806_inst
    process(type_cast_4804_wire_constant, lock_bus_4735) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_4804_wire_constant, lock_bus_4735, tmp_var);
      CONCAT_u1_u2_4806_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_4809_inst
    process(is_write_dword_4755, is_read_dword_4759) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(is_write_dword_4755, is_read_dword_4759, tmp_var);
      CONCAT_u1_u2_4809_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u9_4788_inst
    process(to_dcache_4747, flags_4767) -- 
      variable tmp_var : std_logic_vector(8 downto 0); -- 
    begin -- 
      ApConcat_proc(to_dcache_4747, flags_4767, tmp_var);
      CONCAT_u1_u9_4788_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u9_4813_inst
    process(is_read_line_4763, byte_mask_4771) -- 
      variable tmp_var : std_logic_vector(8 downto 0); -- 
    begin -- 
      ApConcat_proc(is_read_line_4763, byte_mask_4771, tmp_var);
      CONCAT_u1_u9_4813_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u2_u3_4785_inst
    process(CONCAT_u1_u2_4783_wire, send_response_4751) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_4783_wire, send_response_4751, tmp_var);
      CONCAT_u2_u3_4785_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u2_u4_4810_inst
    process(CONCAT_u1_u2_4806_wire, CONCAT_u1_u2_4809_wire) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_4806_wire, CONCAT_u1_u2_4809_wire, tmp_var);
      CONCAT_u2_u4_4810_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u36_u100_4816_inst
    process(physical_addr_to_mem_4775, write_data_4779) -- 
      variable tmp_var : std_logic_vector(99 downto 0); -- 
    begin -- 
      ApConcat_proc(physical_addr_to_mem_4775, write_data_4779, tmp_var);
      CONCAT_u36_u100_4816_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u3_u12_4789_inst
    process(CONCAT_u2_u3_4785_wire, CONCAT_u1_u9_4788_wire) -- 
      variable tmp_var : std_logic_vector(11 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u2_u3_4785_wire, CONCAT_u1_u9_4788_wire, tmp_var);
      CONCAT_u3_u12_4789_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u4_u113_4818_inst
    process(CONCAT_u2_u4_4810_wire, CONCAT_u9_u109_4817_wire) -- 
      variable tmp_var : std_logic_vector(112 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u2_u4_4810_wire, CONCAT_u9_u109_4817_wire, tmp_var);
      CONCAT_u4_u113_4818_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u95_u208_4819_inst
    process(CONCAT_u12_u95_4802_wire, CONCAT_u4_u113_4818_wire) -- 
      variable tmp_var : std_logic_vector(207 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u12_u95_4802_wire, CONCAT_u4_u113_4818_wire, tmp_var);
      reconstructed_fast_cmd_4820 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u9_u109_4817_inst
    process(CONCAT_u1_u9_4813_wire, CONCAT_u36_u100_4816_wire) -- 
      variable tmp_var : std_logic_vector(108 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u9_4813_wire, CONCAT_u36_u100_4816_wire, tmp_var);
      CONCAT_u9_u109_4817_wire <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end mergeCommands_VVV_arch;
-- VHDL global package produced by vc2vhdl from virtual circuit (vc) description 
library ieee;
use ieee.std_logic_1164.all;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
entity constructDcacheMmuRequest_VVV is -- 
  port ( -- 
    from_dcache : in  std_logic_vector(119 downto 0);
    to_mmu : out  std_logic_vector(121 downto 0)-- 
  );
  -- 
end entity constructDcacheMmuRequest_VVV;
architecture constructDcacheMmuRequest_VVV_arch of constructDcacheMmuRequest_VVV is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(120-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal from_dcache_buffer :  std_logic_vector(119 downto 0);
  -- output port buffer signals
  signal to_mmu_buffer :  std_logic_vector(121 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  from_dcache_buffer <= from_dcache;
  -- output handling  -------------------------------------------------------
  to_mmu <= to_mmu_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u16_u56_92_wire : std_logic_vector(55 downto 0);
    signal CONCAT_u64_u65_96_wire : std_logic_vector(64 downto 0);
    signal CONCAT_u65_u66_99_wire : std_logic_vector(65 downto 0);
    signal CONCAT_u8_u16_88_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u40_91_wire : std_logic_vector(39 downto 0);
    signal addr_80 : std_logic_vector(31 downto 0);
    signal asi_68 : std_logic_vector(7 downto 0);
    signal byte_mask_72 : std_logic_vector(7 downto 0);
    signal request_type_76 : std_logic_vector(7 downto 0);
    signal type_cast_95_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_98_wire_constant : std_logic_vector(0 downto 0);
    signal write_data_84 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    type_cast_95_wire_constant <= "1";
    type_cast_98_wire_constant <= "1";
    -- flow-through slice operator slice_67_inst
    asi_68 <= from_dcache_buffer(119 downto 112);
    -- flow-through slice operator slice_71_inst
    byte_mask_72 <= from_dcache_buffer(111 downto 104);
    -- flow-through slice operator slice_75_inst
    request_type_76 <= from_dcache_buffer(103 downto 96);
    -- flow-through slice operator slice_79_inst
    addr_80 <= from_dcache_buffer(95 downto 64);
    -- flow-through slice operator slice_83_inst
    write_data_84 <= from_dcache_buffer(63 downto 0);
    -- binary operator CONCAT_u16_u56_92_inst
    process(CONCAT_u8_u16_88_wire, CONCAT_u8_u40_91_wire) -- 
      variable tmp_var : std_logic_vector(55 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_88_wire, CONCAT_u8_u40_91_wire, tmp_var);
      CONCAT_u16_u56_92_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u56_u122_100_inst
    process(CONCAT_u16_u56_92_wire, CONCAT_u65_u66_99_wire) -- 
      variable tmp_var : std_logic_vector(121 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u16_u56_92_wire, CONCAT_u65_u66_99_wire, tmp_var);
      to_mmu_buffer <= tmp_var; --
    end process;
    -- binary operator CONCAT_u64_u65_96_inst
    process(write_data_84) -- 
      variable tmp_var : std_logic_vector(64 downto 0); -- 
    begin -- 
      ApConcat_proc(write_data_84, type_cast_95_wire_constant, tmp_var);
      CONCAT_u64_u65_96_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u65_u66_99_inst
    process(CONCAT_u64_u65_96_wire) -- 
      variable tmp_var : std_logic_vector(65 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u64_u65_96_wire, type_cast_98_wire_constant, tmp_var);
      CONCAT_u65_u66_99_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u16_88_inst
    process(asi_68, request_type_76) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(asi_68, request_type_76, tmp_var);
      CONCAT_u8_u16_88_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u40_91_inst
    process(byte_mask_72, addr_80) -- 
      variable tmp_var : std_logic_vector(39 downto 0); -- 
    begin -- 
      ApConcat_proc(byte_mask_72, addr_80, tmp_var);
      CONCAT_u8_u40_91_wire <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end constructDcacheMmuRequest_VVV_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
entity constructIcacheMmuRequest_VVV is -- 
  port ( -- 
    from_icache : in  std_logic_vector(47 downto 0);
    to_mmu : out  std_logic_vector(121 downto 0)-- 
  );
  -- 
end entity constructIcacheMmuRequest_VVV;
architecture constructIcacheMmuRequest_VVV_arch of constructIcacheMmuRequest_VVV is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(48-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal from_icache_buffer :  std_logic_vector(47 downto 0);
  -- output port buffer signals
  signal to_mmu_buffer :  std_logic_vector(121 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  from_icache_buffer <= from_icache;
  -- output handling  -------------------------------------------------------
  to_mmu <= to_mmu_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u16_u56_127_wire : std_logic_vector(55 downto 0);
    signal CONCAT_u65_u66_136_wire_constant : std_logic_vector(65 downto 0);
    signal CONCAT_u8_u16_121_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u40_126_wire : std_logic_vector(39 downto 0);
    signal NOT_u8_u8_124_wire_constant : std_logic_vector(7 downto 0);
    signal addr_117 : std_logic_vector(31 downto 0);
    signal asi_109 : std_logic_vector(7 downto 0);
    signal request_type_113 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    CONCAT_u65_u66_136_wire_constant <= "000000000000000000000000000000000000000000000000000000000000000001";
    NOT_u8_u8_124_wire_constant <= "11111111";
    -- flow-through slice operator slice_108_inst
    asi_109 <= from_icache_buffer(47 downto 40);
    -- flow-through slice operator slice_112_inst
    request_type_113 <= from_icache_buffer(39 downto 32);
    -- flow-through slice operator slice_116_inst
    addr_117 <= from_icache_buffer(31 downto 0);
    -- binary operator CONCAT_u16_u56_127_inst
    process(CONCAT_u8_u16_121_wire, CONCAT_u8_u40_126_wire) -- 
      variable tmp_var : std_logic_vector(55 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_121_wire, CONCAT_u8_u40_126_wire, tmp_var);
      CONCAT_u16_u56_127_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u56_u122_138_inst
    process(CONCAT_u16_u56_127_wire) -- 
      variable tmp_var : std_logic_vector(121 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u16_u56_127_wire, CONCAT_u65_u66_136_wire_constant, tmp_var);
      to_mmu_buffer <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u16_121_inst
    process(asi_109, request_type_113) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(asi_109, request_type_113, tmp_var);
      CONCAT_u8_u16_121_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u40_126_inst
    process(NOT_u8_u8_124_wire_constant, addr_117) -- 
      variable tmp_var : std_logic_vector(39 downto 0); -- 
    begin -- 
      ApConcat_proc(NOT_u8_u8_124_wire_constant, addr_117, tmp_var);
      CONCAT_u8_u40_126_wire <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end constructIcacheMmuRequest_VVV_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
entity mmuDcacheServiceDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    DCACHE_to_MMU_request_pipe_read_req : out  std_logic_vector(0 downto 0);
    DCACHE_to_MMU_request_pipe_read_ack : in   std_logic_vector(0 downto 0);
    DCACHE_to_MMU_request_pipe_read_data : in   std_logic_vector(119 downto 0);
    NOBLOCK_DCACHE_TO_MMU_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_DCACHE_TO_MMU_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_DCACHE_TO_MMU_REQUEST_pipe_write_data : out  std_logic_vector(121 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity mmuDcacheServiceDaemon;
architecture mmuDcacheServiceDaemon_arch of mmuDcacheServiceDaemon is -- 
  -- volatile/operator module components. 
  component constructDcacheMmuRequest_VVV is -- 
    port ( -- 
      from_dcache : in  std_logic_vector(119 downto 0);
      to_mmu : out  std_logic_vector(121 downto 0)-- 
    );
  end component; 
begin --  
	tag_out <= tag_in;
	start_ack <= '1';
	fin_ack <= '0';
	
    	NOBLOCK_DCACHE_TO_MMU_REQUEST_pipe_write_req <= DCACHE_to_MMU_request_pipe_read_ack;
	DCACHE_to_MMU_request_pipe_read_req <= NOBLOCK_DCACHE_TO_MMU_REQUEST_pipe_write_ack;

	gR: constructDcacheMmuRequest_VVV 
			port map (from_dcache => DCACHE_to_MMU_request_pipe_read_data,
					to_mmu => NOBLOCK_DCACHE_TO_MMU_REQUEST_pipe_write_data);

end mmuDcacheServiceDaemon_arch;


library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
entity mmuIcacheServiceDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    ICACHE_to_MMU_request_pipe_read_req : out  std_logic_vector(0 downto 0);
    ICACHE_to_MMU_request_pipe_read_ack : in   std_logic_vector(0 downto 0);
    ICACHE_to_MMU_request_pipe_read_data : in   std_logic_vector(47 downto 0);
    NOBLOCK_ICACHE_TO_MMU_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_ICACHE_TO_MMU_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_ICACHE_TO_MMU_REQUEST_pipe_write_data : out  std_logic_vector(121 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity mmuIcacheServiceDaemon;
architecture mmuIcacheServiceDaemon_arch of mmuIcacheServiceDaemon is -- 
  component constructIcacheMmuRequest_VVV is -- 
    port ( -- 
      from_icache : in  std_logic_vector(47 downto 0);
      to_mmu : out  std_logic_vector(121 downto 0)-- 
    );
    -- 
  end component; 
begin --  
	start_ack <= '1';
	fin_ack <= '0';
	tag_out <= tag_in;
	
    	NOBLOCK_ICACHE_TO_MMU_REQUEST_pipe_write_req <= ICACHE_to_MMU_request_pipe_read_ack;
	ICACHE_to_MMU_request_pipe_read_req <= NOBLOCK_ICACHE_TO_MMU_REQUEST_pipe_write_ack;

	gR: constructIcacheMmuRequest_VVV 
			port map (from_icache => ICACHE_to_MMU_request_pipe_read_data,
					to_mmu => NOBLOCK_ICACHE_TO_MMU_REQUEST_pipe_write_data);

end mmuIcacheServiceDaemon_arch;

library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
entity mmuMuxDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    NOBLOCK_DCACHE_TO_MMU_REQUEST_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_DCACHE_TO_MMU_REQUEST_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_DCACHE_TO_MMU_REQUEST_pipe_read_data : in   std_logic_vector(121 downto 0);
    NOBLOCK_ICACHE_TO_MMU_REQUEST_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_ICACHE_TO_MMU_REQUEST_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_ICACHE_TO_MMU_REQUEST_pipe_read_data : in   std_logic_vector(121 downto 0);
    NOBLOCK_CACHE_TO_MMU_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_CACHE_TO_MMU_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_CACHE_TO_MMU_REQUEST_pipe_write_data : out  std_logic_vector(121 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity mmuMuxDaemon;
architecture mmuMuxDaemon_arch of mmuMuxDaemon is -- 
	signal icache_has_priority: boolean;

	signal icache_is_valid: boolean;
	signal dcache_is_valid: boolean;

	signal select_icache, select_dcache, send_something: std_logic;

	signal send_to_mmu, mmu_ready: std_logic;

	type FsmState is (IDLE, WAIT_ON_MMU);
	signal fsm_state: FsmState;

	signal ack_icache, ack_dcache: std_logic;

	signal dcache_queue_data_out : std_logic_vector(121 downto 0);
	signal dcache_queue_pop_req,  dcache_queue_pop_ack: std_logic;

	signal dcache_wants_lock, dcache_has_lock: boolean;
	
begin --  
	start_ack <= '1';
	fin_ack  <= '0';
	tag_out <= tag_in;

	-- a little bit of queueing on the dcache side which generates
	-- lots of write through requests to the mmu..  But note the bypass.
	qb: QueueWithBypass
		generic map (name => "mmu_mux_dcache_request_queue",
				queue_depth => 2, data_width => dcache_queue_data_out'length)
		port map (
			clk => clk, reset => reset,
			data_in  => NOBLOCK_DCACHE_TO_MMU_REQUEST_pipe_read_data,
			push_req => NOBLOCK_DCACHE_TO_MMU_REQUEST_pipe_read_ack(0), 
			push_ack => NOBLOCK_DCACHE_TO_MMU_REQUEST_pipe_read_req(0), 
			data_out => dcache_queue_data_out,
			pop_req  => dcache_queue_pop_req,
			pop_ack  => dcache_queue_pop_ack);

	icache_is_valid <= (NOBLOCK_ICACHE_TO_MMU_REQUEST_pipe_read_ack(0) = '1') and
					(NOBLOCK_ICACHE_TO_MMU_REQUEST_pipe_read_data(0) = '1'); 
	dcache_is_valid <= (dcache_queue_pop_ack = '1') and (dcache_queue_data_out(0) = '1'); 

	-- dcache lock is bit 6 of request
	--    asi [121:114]
	--    request [113:106], so [112]
	dcache_wants_lock <=  (dcache_is_valid and (dcache_queue_data_out(112) = '1'));


	select_icache <= '1' when (icache_is_valid and (not dcache_has_lock) and 
					((not dcache_is_valid) or icache_has_priority)) else '0';
	select_dcache <= '1' when (dcache_is_valid and
					(dcache_has_lock or 
						(not icache_is_valid) or (not icache_has_priority))) else '0';
				
	send_something <= (select_icache or select_dcache);
	

	process(clk, reset, fsm_state, mmu_ready, select_icache, select_dcache, send_something,
				icache_has_priority, dcache_wants_lock, dcache_has_lock)
		variable next_fsm_state_var : FsmState;
		variable send_to_mmu_var: std_logic;
		variable ack_icache_var, ack_dcache_var: std_logic;
		variable next_icache_has_priority_var: boolean;
		variable next_dcache_has_lock_var: boolean;
	begin
		next_fsm_state_var := fsm_state;
		send_to_mmu_var    := '0';
		next_icache_has_priority_var := icache_has_priority;
		ack_icache_var := '0';
		ack_dcache_var := '0';

		next_dcache_has_lock_var := dcache_has_lock;

		case fsm_state is
			when IDLE => 
				if(send_something = '1') then
					send_to_mmu_var := '1';
					if(mmu_ready = '1') then
						ack_icache_var := select_icache;
						ack_dcache_var := select_dcache;
						next_icache_has_priority_var := not icache_has_priority;
					else 
						next_fsm_state_var := WAIT_ON_MMU;
					end if;
				end if;
			when WAIT_ON_MMU => 
				send_to_mmu_var := '1';
				if(mmu_ready = '1') then
					next_icache_has_priority_var := not icache_has_priority;
					ack_icache_var := select_icache;
					ack_dcache_var := select_dcache;
					next_fsm_state_var := IDLE;
				end if;
		end case;	


		if(select_dcache = '1') then
			if(dcache_wants_lock) then
				next_dcache_has_lock_var := true;
			else
				next_dcache_has_lock_var := false;
			end if;
		end if;

		ack_icache <= ack_icache_var;
		ack_dcache <= ack_dcache_var;
		send_to_mmu <= send_to_mmu_var;

		if(clk'event and (clk = '1')) then
			if(reset = '1') then
				fsm_state <= IDLE;
				dcache_has_lock <= false;
			else
				fsm_state <= next_fsm_state_var;
				icache_has_priority <= next_icache_has_priority_var;
				dcache_has_lock <= next_dcache_has_lock_var;
			end if;
		end if;
	end process;

    	NOBLOCK_CACHE_TO_MMU_REQUEST_pipe_write_req(0) <= send_to_mmu;
    	mmu_ready <= NOBLOCK_CACHE_TO_MMU_REQUEST_pipe_write_ack(0);

    	NOBLOCK_CACHE_TO_MMU_REQUEST_pipe_write_data <= 
			NOBLOCK_ICACHE_TO_MMU_REQUEST_pipe_read_data when (select_icache = '1') 
					else dcache_queue_data_out when (select_dcache = '1') else
						(others => '0'); 
		
    	dcache_queue_pop_req <= ack_dcache;
    	NOBLOCK_ICACHE_TO_MMU_REQUEST_pipe_read_req(0) <= ack_icache;

end mmuMuxDaemon_arch;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.mem_component_pack.all;


-- a generic fully associative memory for use in the MMU TLB.
entity genericFullyAssociativeMemory is
	generic (tag_width: integer := 8;
			data_width: integer := 32;
			log_number_of_entries: integer := 6;
			ignore_collisions: boolean := true;
			use_mem_cuts: boolean:= true);
	port (  start_req: in std_logic;
		start_ack: out std_logic;
		fin_req: in std_logic;
		fin_ack: out std_logic;

		-- clear all valids.
		clear_flag: in std_logic_vector(0 downto 0);

		-- add entry
		erase_flag: in std_logic_vector(0 downto 0);
		write_flag: in std_logic_vector(0 downto 0);
		write_data: in std_logic_vector(data_width-1 downto 0);
		write_tag : in std_logic_vector(tag_width-1 downto 0);

		-- lookup entry
		lookup_flag: in std_logic_vector(0 downto 0);
		lookup_tag : in std_logic_vector(tag_width-1 downto 0);
		lookup_valid: out std_logic_vector(0 downto 0);
		lookup_data: out std_logic_vector(data_width-1 downto 0);

		clk,reset: in std_logic);

end entity genericFullyAssociativeMemory;


-- read and then write.
architecture genericFullyAssociativeMemoryArch of genericFullyAssociativeMemory is


	-- tags for all entries in a set are maintained in a single word.
	signal last_written_index, update_index: integer range 0 to (2**log_number_of_entries);

	signal valids_vector : std_logic_vector((2**log_number_of_entries)-1 downto 0);
	signal tags_vector   : std_logic_vector((2**log_number_of_entries)*tag_width-1 downto 0);

	signal collision_flag_reg : std_logic;
	signal erase_collision_flag_reg : std_logic;

	subtype TagWord is std_logic_vector(tag_width-1 downto 0);
	type TagWordArray is array (natural range <> ) of TagWord;
	function tagArrayToVector (x: TagWordArray) 
		return std_logic_vector is
		alias twa : TagWordArray((2**log_number_of_entries)-1 downto 0) is x;
		variable ret_var : std_logic_vector((2**log_number_of_entries)*tag_width -1 downto 0);
	begin
		for I in 0 to (2**log_number_of_entries)-1 loop
			ret_var(((I+1)*tag_width)-1 downto (I*tag_width)) := twa(I);
		end loop;
		return(ret_var);
	end function;
	function tagVectorToArray (x: std_logic_vector) return TagWordArray is
		alias tx : std_logic_vector((2**log_number_of_entries)*tag_width - 1 downto 0) is x;
		variable ret_var: TagWordArray((2**log_number_of_entries-1) downto 0);
	begin
		for I in 0 to (2**log_number_of_entries)-1 loop
			 ret_var(I) := tx(((I+1)*tag_width)-1 downto (I*tag_width));
		end loop;
		return(ret_var);
	end function;
		
	-- data memory access signals
	signal data_mem_write_data, data_mem_read_data: std_logic_vector(data_width-1 downto 0);
	signal data_mem_address: std_logic_vector(log_number_of_entries-1 downto 0);
	signal data_mem_enable, data_mem_write_bar: std_logic;

	type FsmState is (IDLE, WRITE_STATE);
	signal fsm_state: FsmState;
	signal done_reg: std_logic;

	signal lookup_match_index, write_match_index, write_match_index_reg: integer range 0 to (2**log_number_of_entries);

	signal lookup_flag_reg: std_logic_vector(0 downto 0);
	signal lookup_valid_reg: std_logic;
		
	signal write_flag_reg	: std_logic_vector(0 downto 0);
	signal write_data_reg	: std_logic_vector(data_width-1 downto 0);
	signal write_tag_reg 	: std_logic_vector(tag_width-1 downto 0);

	signal sample_write_inputs: boolean;

	function matchTag (tags: std_logic_vector; ltag: std_logic_vector; valids: std_logic_vector; W: integer) 
		return integer is
		variable ret_var: integer;

		alias ltags: std_logic_vector((W*tag_width)-1 downto 0) is tags;
		alias lltag: std_logic_vector(tag_width-1 downto 0) is ltag;
		alias lvalids: std_logic_vector(W-1 downto 0) is valids;
		variable lret_var, rret_var: integer;
	begin
		ret_var := -1;

		if(W = 1) then
			if((lvalids(0) = '1') and (ltags = lltag)) then
				ret_var := 0;
			end if;
		else 
			rret_var := matchTag(ltags((W*tag_width)-1 downto (W/2)*tag_width), ltag, 
								lvalids (W-1 downto W/2), W - (W/2));
			lret_var := matchTag(ltags(((W/2)*tag_width)-1 downto 0), ltag, 
								lvalids ((W/2)-1 downto 0), W/2);
			if(rret_var >= 0) then
				ret_var := rret_var + W - (W/2);
			elsif (lret_var >= 0) then
				ret_var := lret_var;
			end if;
		end if;
		return ret_var;
	end matchTag;

	function findMatchIndex (tags: std_logic_vector; valids: std_logic_vector; search_tag: std_logic_vector)
		return integer is
		variable ret_var: integer range 0 to (2**log_number_of_entries);
		variable T: integer;
		alias ltags: std_logic_vector((tag_width*(2**log_number_of_entries))-1 downto 0) is tags;
		alias lvalids: std_logic_vector((2**log_number_of_entries)-1 downto 0) is valids;
		alias llookup_tag: std_logic_vector(tag_width-1 downto 0) is search_tag;
	begin
		ret_var := (2**log_number_of_entries);
		--T := matchTag(ltags, llookup_tag, lvalids, valids'length);
		--if(T >= 0) then
			--ret_var := T;
		--end if;
		--return (ret_var);
		for I in 0 to  (2**log_number_of_entries)-1 loop
			if(lvalids(I) = '1') then
				if(ltags(((I+1)*tag_width)-1 downto (I*tag_width)) = search_tag) then
					ret_var := I;
					exit;
				end if;
			end if;
		end loop;
		return ret_var;
	end function;

						
	function IncrementWrittenIndex(last_windex: integer) 
		return integer is
		variable ret_var: integer range 0 to (2**log_number_of_entries);
	begin

		if(last_windex >= ((2**log_number_of_entries)-1)) then
			ret_var := 0;
		else
			ret_var := last_windex + 1;
		end if;	

		return (ret_var);
	end function;

begin

   lookup_match_index  <= findMatchIndex (tags_vector, valids_vector, lookup_tag);
   write_match_index   <= findMatchIndex (tags_vector, valids_vector, write_tag);
   
   process(fsm_state, clear_flag, 
			erase_flag, 
			lookup_flag, 
			write_flag, 
			lookup_match_index, 
			write_match_index,
			start_req, fin_req, 
			done_reg,
			collision_flag_reg,
			erase_collision_flag_reg,
			clk, reset)
	variable next_fsm_state_var : FsmState;
	variable next_valids_var : std_logic_vector((2**log_number_of_entries)-1 downto 0);
	variable next_tags_var: TagWordArray((2**log_number_of_entries-1) downto 0);
	variable next_lookup_valid_var: std_logic;
	variable data_mem_write_data_var: std_logic_vector(data_width-1 downto 0);
	variable data_mem_address_var: std_logic_vector(log_number_of_entries-1 downto 0);
	variable data_mem_enable_var, data_mem_write_bar_var: std_logic;
	variable sample_write_inputs_var : boolean;
	variable next_last_written_index_var: integer range 0 to (2**log_number_of_entries);
	variable update_index_var: integer range 0 to (2**log_number_of_entries);
	variable start_ack_var, fin_ack_var: std_logic;
	variable next_lookup_flag_reg_var: std_logic_vector(0 downto 0);
	variable next_done_var : std_logic;
	variable collision_var : std_logic;
	variable erase_collision_var : std_logic;
   begin
	next_fsm_state_var := fsm_state;
	next_valids_var    := valids_vector;
	next_lookup_valid_var := lookup_valid_reg;
	next_lookup_flag_reg_var := lookup_flag_reg;
	next_done_var := done_reg;
	collision_var := collision_flag_reg;
	erase_collision_var := erase_collision_flag_reg;


	next_tags_var := tagVectorToArray(tags_vector);
	next_last_written_index_var := last_written_index;

	sample_write_inputs_var := false;

	data_mem_write_data_var := (others => '0');
	data_mem_address_var := (others => '0');
	data_mem_enable_var := '0';
	data_mem_write_bar_var := '1';

	fin_ack_var := '0';
	start_ack_var := '0';


	case fsm_state is 
		when IDLE =>
			fin_ack_var := done_reg;
			if((done_reg = '0') or (fin_req = '1'))  then 
				next_done_var := '0';

				-- can start again
			  	start_ack_var := '1';
			  	if(start_req = '1') then  

				  	sample_write_inputs_var := true;
				  	next_lookup_flag_reg_var := lookup_flag;

					-- by default we are done in one step 
					-- except as indicated below.
					next_done_var := '1';

					erase_collision_var := '0';
					collision_var := '0';

					if ((not ignore_collisions) and
						(lookup_flag(0) = '1') and
						(clear_flag(0) = '0') and 
						((write_flag(0) = '1') or
							(erase_flag(0) = '1'))
						and (lookup_tag = write_tag)) then

						collision_var := '1';

						-- erase and collision means invalid.
						if(erase_flag(0) = '1') then
							erase_collision_var := '1';
						end if;
					end if;

		
					-- must clear it!  Not clearing it was a bug.
					next_lookup_valid_var := '0';

				  	-- clear flag: clear all valids.
				  	if(clear_flag(0) = '1') then
						next_valids_var := (others => '0');
				  	end if;
	
				  	-- erase flag: clear the write tag entry.
				  	if(erase_flag(0) = '1') then
					  	if(write_match_index < (2**log_number_of_entries)) then
							next_valids_var(write_match_index) := '0';
					  	end if;
				  	end if;
	
				  	-- lookup?  read the data if there is a match.
  				  	if(lookup_flag(0) = '1') then

					  	if(lookup_match_index < (2**log_number_of_entries)) then
						    -- need to read only if there is no collision.
						    if(collision_var = '0') then
						  	data_mem_address_var := 
						      		std_logic_vector(to_unsigned(lookup_match_index, 
											log_number_of_entries));
						  	data_mem_enable_var  := '1';
						  	data_mem_write_bar_var := '1';
                                                    end if;

						    -- erase collision?   invalid lookup
						    if(erase_collision_var = '0') then
						    	next_lookup_valid_var := '1';
						    end if;

					  	end if;
	
					  	if(write_flag(0) = '1') then
						  	next_fsm_state_var := WRITE_STATE;

							-- next done.. make it '0' because you need
							-- to do the write in the next cycle.
							next_done_var := '0';
					  	end if;

				  	elsif(write_flag(0) = '1') then
						-- write in a new entry.
						if(write_match_index < (2**log_number_of_entries)) then
							update_index_var := write_match_index;
						else 
					  		next_last_written_index_var := 
									IncrementWrittenIndex(last_written_index);
							update_index_var := next_last_written_index_var;
						end if;
					  	data_mem_write_data_var := write_data;
					  	data_mem_address_var := 
						  	std_logic_vector(to_unsigned(update_index_var, 
											log_number_of_entries));
					  	data_mem_enable_var  := '1';
					  	data_mem_write_bar_var := '0';
					  	next_valids_var(update_index_var) := '1';
					  	next_tags_var(update_index_var) := write_tag;
							
						-- next_done_var stays '1'.
						-- stay in IDLE.
				  	end if;
			  	end if;
			end if;

		when WRITE_STATE =>

			-- done_reg is '0' when you enter this state.

			if(write_match_index_reg < (2**log_number_of_entries))then
				update_index_var := write_match_index_reg;
			else 
				next_last_written_index_var := IncrementWrittenIndex(last_written_index);
				update_index_var := next_last_written_index_var;
			end if;

			data_mem_write_data_var := write_data_reg;
			data_mem_address_var := 
				std_logic_vector(to_unsigned(update_index_var,log_number_of_entries));
			data_mem_enable_var  := '1';
			data_mem_write_bar_var := '0';
			next_valids_var(update_index_var) := '1';
			next_tags_var(update_index_var) := write_tag_reg;

			next_fsm_state_var := IDLE;
			next_done_var := '1';
	end case;

	data_mem_write_data <= data_mem_write_data_var;
	data_mem_address <= data_mem_address_var;
	data_mem_enable  <= data_mem_enable_var;
	data_mem_write_bar <= data_mem_write_bar_var;

	start_ack <= start_ack_var;
	fin_ack   <= done_reg;

	if(clk'event and (clk = '1')) then
		if(reset = '1') then
			fsm_state <= IDLE;
			valids_vector <= (others => '0');
			tags_vector <= (others => '0');
			last_written_index <= (2**log_number_of_entries);
			lookup_valid_reg <= '0';
			lookup_flag_reg(0) <= '0';
			done_reg <= '0';
			collision_flag_reg <= '0';
			erase_collision_flag_reg <= '0';
		else
			fsm_state <= next_fsm_state_var;
			lookup_valid_reg <= next_lookup_valid_var;
			valids_vector <= next_valids_var;
			tags_vector   <= tagArrayToVector(next_tags_var);
			last_written_index <= next_last_written_index_var;
			lookup_flag_reg <= next_lookup_flag_reg_var;
			

			done_reg <= next_done_var;
			collision_flag_reg <= collision_var;
			erase_collision_flag_reg <= erase_collision_var;

			if(sample_write_inputs_var) then
				write_flag_reg	<= write_flag;
				write_data_reg	<= write_data;
				write_tag_reg 	<= write_tag;
				write_match_index_reg <= write_match_index;
			end if;
		end if;
	end if;
   end process;
  

   	
   memCutBB: if use_mem_cuts generate 
   	data_bb: base_bank 
		generic map  (name => "genericFullyAssociativeMemory:data_base_bank", 
						g_addr_width => log_number_of_entries,
						g_data_width => data_width)
		port map (
				datain => data_mem_write_data,
				addrin => data_mem_address,
				dataout => data_mem_read_data,
				enable => data_mem_enable,
				writebar => data_mem_write_bar,
				clk => clk, reset => reset
			);
   end generate memCutBB;
   regBB: if not use_mem_cuts generate 
   	data_bb: base_bank_with_registers
		generic map  (name => "genericFullyAssociativeMemory:data_base_bank", 
						g_addr_width => log_number_of_entries,
						g_data_width => data_width)
		port map (
				datain => data_mem_write_data,
				addrin => data_mem_address,
				dataout => data_mem_read_data,
				enable => data_mem_enable,
				writebar => data_mem_write_bar,
				clk => clk, reset => reset);
   end generate regBB;

   lookup_valid(0) <= lookup_valid_reg or (collision_flag_reg and (not erase_collision_flag_reg));
   lookup_data     <= write_data_reg when (collision_flag_reg = '1')  
				else data_mem_read_data 
					when ((lookup_valid_reg = '1') and (lookup_flag_reg(0) = '1')) 
							else (others => '0');

end genericFullyAssociativeMemoryArch;

		
	
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.BaseComponents.all;

library AjitCustom;
use AjitCustom.AjitCustomComponents.all;


-- a generic fully associative memory for use in the MMU TLB.
entity genericFullyAssociativeMemory_Operator is
	generic (tag_width: integer := 8;
			data_width: integer := 32;
			log_number_of_entries: integer := 6;
			ignore_collisions: boolean := true;
			use_mem_cuts: boolean:= true);
	port (  sample_req: in boolean;
		sample_ack: out boolean;
		update_req: in boolean;
		update_ack: out boolean;

		-- clear all valids.
		clear_flag: in std_logic_vector(0 downto 0);

		-- add entry
		erase_flag: in std_logic_vector(0 downto 0);
		write_flag: in std_logic_vector(0 downto 0);
		write_data: in std_logic_vector(data_width-1 downto 0);
		write_tag : in std_logic_vector(tag_width-1 downto 0);

		-- lookup entry
		lookup_flag: in std_logic_vector(0 downto 0);
		lookup_tag : in std_logic_vector(tag_width-1 downto 0);
		lookup_valid: out std_logic_vector(0 downto 0);
		lookup_data: out std_logic_vector(data_width-1 downto 0);

		clk,reset: in std_logic);

end entity genericFullyAssociativeMemory_Operator;


architecture simpleTon of genericFullyAssociativeMemory_Operator is
	signal start_req, start_ack: std_logic;
	signal fin_req, fin_ack: std_logic;

	signal br_lookup_data: std_logic_vector(data_width-1 downto 0);
	signal br_lookup_valid: std_logic_vector(0 downto 0);
	signal br_data_in, br_data_out: std_logic_vector(data_width downto 0);

   	signal update_ack_sig: boolean;

begin

   p2l: Sample_Pulse_To_Level_Translate_Entity
                generic map(name => "genericFullyAssociativeMemory-Operator-p2l")
                port map (rL => sample_req, rR => start_req,
                                aL => sample_ack, aR => start_ack,
                                        clk => clk, reset => reset);
   l2p: Level_To_Pulse_Translate_Entity
		generic map(name => "genericFullyAssociativeMemory-Operator-l2p")
		port map (rL => fin_req, rR => update_req,
				aL => fin_ack, aR => update_ack_sig, clk => clk, reset => reset);


   update_ack <= update_ack_sig;

   br_data_in <= br_lookup_valid & br_lookup_data;


   br: BypassRegister 
		generic map(data_width => data_width+1, bypass => true)
		port map (clk => clk, reset => reset, din => br_data_in, enable => update_ack_sig, 
					q => br_data_out);

   lookup_valid(0) <= br_data_out(data_width);
   lookup_data <= br_data_out(data_width-1 downto 0);

   bmem: genericFullyAssociativeMemory
			generic map (tag_width => tag_width,
					log_number_of_entries => log_number_of_entries,
					data_width => data_width,
					ignore_collisions => ignore_collisions,
					use_mem_cuts => use_mem_cuts)
			port map (
				start_req => start_req,
				start_ack => start_ack,
				fin_req =>   fin_req,
				fin_ack =>   fin_ack,
    				clear_flag => clear_flag,
    				write_flag => write_flag,
    				write_data => write_data,
				write_tag => write_tag,
				erase_flag => erase_flag,
				lookup_flag => lookup_flag,
				lookup_tag => lookup_tag,
    				lookup_valid => br_lookup_valid,
    				lookup_data =>  br_lookup_data,
    				clk => clk, reset => reset);

end simpleTon;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.mem_component_pack.all;


-- a generic fully associative memory for use in the MMU TLB.
entity genericFullyAssociativeMemoryNoData is
	generic (tag_width: integer := 8; log_number_of_entries: integer := 6; ignore_collisions: boolean := true);
	port (  start_req: in std_logic;
		start_ack: out std_logic;
		fin_req: in std_logic;
		fin_ack: out std_logic;

		-- clear all valids.
		clear_flag: in std_logic_vector(0 downto 0);

		-- add entry
		erase_flag: in std_logic_vector(0 downto 0);
		write_flag: in std_logic_vector(0 downto 0);
		write_tag : in std_logic_vector(tag_width-1 downto 0);

		-- lookup entry
		lookup_flag: in std_logic_vector(0 downto 0);
		lookup_tag : in std_logic_vector(tag_width-1 downto 0);
		lookup_valid: out std_logic_vector(0 downto 0);

		clk,reset: in std_logic);

end entity genericFullyAssociativeMemoryNoData;


-- read and then write.
architecture genericFullyAssociativeMemoryNoDataArch of genericFullyAssociativeMemoryNoData is


	-- tags for all entries in a set are maintained in a single word.
	signal last_written_index: integer range 0 to (2**log_number_of_entries);

	signal valids_vector : std_logic_vector((2**log_number_of_entries)-1 downto 0);
	signal tags_vector   : std_logic_vector((2**log_number_of_entries)*tag_width-1 downto 0);

	subtype TagWord is std_logic_vector(tag_width-1 downto 0);
	type TagWordArray is array (natural range <> ) of TagWord;
	function tagArrayToVector (x: TagWordArray) 
		return std_logic_vector is
		alias twa : TagWordArray((2**log_number_of_entries)-1 downto 0) is x;
		variable ret_var : std_logic_vector((2**log_number_of_entries)*tag_width -1 downto 0);
	begin
		for I in 0 to (2**log_number_of_entries)-1 loop
			ret_var(((I+1)*tag_width)-1 downto (I*tag_width)) := twa(I);
		end loop;
		return(ret_var);
	end function;
	function tagVectorToArray (x: std_logic_vector) return TagWordArray is
		alias tx : std_logic_vector((2**log_number_of_entries)*tag_width - 1 downto 0) is x;
		variable ret_var: TagWordArray((2**log_number_of_entries-1) downto 0);
	begin
		for I in 0 to (2**log_number_of_entries)-1 loop
			 ret_var(I) := tx(((I+1)*tag_width)-1 downto (I*tag_width));
		end loop;
		return(ret_var);
	end function;
		

	type FsmState is (IDLE, DONE_WAIT);
	signal fsm_state: FsmState;

	signal lookup_match_index, write_match_index: integer range 0 to (2**log_number_of_entries);
	signal lookup_valid_reg: std_logic;

	function matchTag (tags: std_logic_vector; ltag: std_logic_vector; valids: std_logic_vector; W: integer) 
		return integer is
		variable ret_var: integer;

		alias ltags: std_logic_vector((W*tag_width)-1 downto 0) is tags;
		alias lltag: std_logic_vector(tag_width-1 downto 0) is ltag;
		alias lvalids: std_logic_vector(W-1 downto 0) is valids;
		variable lret_var, rret_var: integer;
	begin
		ret_var := -1;

		if(W = 1) then
			if((lvalids(0) = '1') and (ltags = lltag)) then
				ret_var := 0;
			end if;
		else 
			rret_var := matchTag(ltags((W*tag_width)-1 downto (W/2)*tag_width), ltag, 
								lvalids (W-1 downto W/2), W - (W/2));
			lret_var := matchTag(ltags(((W/2)*tag_width)-1 downto 0), ltag, 
								lvalids ((W/2)-1 downto 0), W/2);
			if(rret_var >= 0) then
				ret_var := rret_var + W - (W/2);
			elsif (lret_var >= 0) then
				ret_var := lret_var;
			end if;
		end if;
		return ret_var;
	end matchTag;

	function findMatchIndex (tags: std_logic_vector; valids: std_logic_vector; search_tag: std_logic_vector)
		return integer is
		variable ret_var: integer range 0 to (2**log_number_of_entries);
		variable T: integer;
		alias ltags: std_logic_vector((tag_width*(2**log_number_of_entries))-1 downto 0) is tags;
		alias lvalids: std_logic_vector((2**log_number_of_entries)-1 downto 0) is valids;
		alias llookup_tag: std_logic_vector(tag_width-1 downto 0) is search_tag;
	begin
		ret_var := (2**log_number_of_entries);
		--T := matchTag(ltags, llookup_tag, lvalids, valids'length);
		--if(T >= 0) then
			--ret_var := T;
		--end if;
		--return (ret_var);
		for I in 0 to  (2**log_number_of_entries)-1 loop
			if(lvalids(I) = '1') then
				if(ltags(((I+1)*tag_width)-1 downto (I*tag_width)) = search_tag) then
					ret_var := I;
					exit;
				end if;
			end if;
		end loop;
		return ret_var;
	end function;

						
	function IncrementWriteIndex(last_windex: integer) 
		return integer is
		variable ret_var: integer range 0 to (2**log_number_of_entries);
	begin

		if(last_windex >= ((2**log_number_of_entries) - 1)) then
			ret_var := 0;
		else
			ret_var := last_windex + 1;
		end if;	
		return (ret_var);

	end function;

begin

   lookup_match_index  <= findMatchIndex (tags_vector, valids_vector, lookup_tag);
   write_match_index   <= findMatchIndex (tags_vector, valids_vector, write_tag);
   
   process(fsm_state, clear_flag, 
			erase_flag, 
			lookup_flag, 
			write_flag, 
			lookup_match_index, 
			write_match_index,
			start_req, fin_req, 
			clk, reset)
	variable next_fsm_state_var : FsmState;
	variable next_valids_var : std_logic_vector((2**log_number_of_entries)-1 downto 0);
	variable next_tags_var: TagWordArray((2**log_number_of_entries-1) downto 0);
	variable next_lookup_valid_var: std_logic;
	variable sample_write_inputs_var : boolean;
	variable next_last_written_index_var: integer range 0 to (2**log_number_of_entries);
	variable start_ack_var, fin_ack_var: std_logic;
	variable collision_var: std_logic;
   begin
	next_fsm_state_var := fsm_state;
	next_valids_var    := valids_vector;
	next_lookup_valid_var := lookup_valid_reg;

	next_tags_var := tagVectorToArray(tags_vector);
	next_last_written_index_var := last_written_index;

	sample_write_inputs_var := false;

	collision_var := '0';


	fin_ack_var := '0';
	start_ack_var := '0';


	if(fsm_state = DONE_WAIT) then
		fin_ack_var := '1';
	end if;

	if((fsm_state = IDLE) or (fin_req = '1'))  then 

		-- can start again
	  	start_ack_var := '1';
	  	if(start_req = '1') then  
			next_lookup_valid_var := '0';
			if((not ignore_collisions) and
				(clear_flag(0) = '0') and ((write_flag(0)  = '1') or (erase_flag(0) = '1'))
					and (lookup_flag(0) = '1') and
						(write_tag = lookup_tag)) then
				collision_var := '1';
			end if;

		  	-- clear flag: clear all valids.
		  	if(clear_flag(0) = '1') then
				next_valids_var := (others => '0');
		  	end if;
	
		  	-- erase flag: clear the write tag entry.
		  	if(erase_flag(0) = '1') then
			  	if(write_match_index < (2**log_number_of_entries)) then
					next_valids_var(write_match_index) := '0';
			  	end if;
		  	end if;
	
		  	-- lookup?  read the data if there is a match.
  		  	if(lookup_flag(0) = '1') then
			  	if(lookup_match_index < (2**log_number_of_entries)) then
					if ((collision_var = '0') or (erase_flag(0) = '0')) then
				  		next_lookup_valid_var := '1';
					end if;
				elsif ((collision_var = '1') and (erase_flag(0) = '0')) then
				  	next_lookup_valid_var := '1';
			  	end if;
			end if;

		  	if((write_flag(0) = '1') and (write_match_index >= (2**log_number_of_entries))) then
				-- write in a new entry.
			  	next_last_written_index_var := IncrementWriteIndex(last_written_index);
			  	next_valids_var(next_last_written_index_var) := '1';
			  	next_tags_var(next_last_written_index_var) := write_tag;
		  	end if;
			next_fsm_state_var := DONE_WAIT;

	  	else -- if (start_req = '0')
			-- could have started again, but no start_req present.
			next_fsm_state_var := IDLE;
	  	end if;
	else 
		-- (fsm_state = DONE) and (fin_req = '0')
		next_fsm_state_var := DONE_WAIT;
	end if;

	start_ack <= start_ack_var;
	fin_ack   <= fin_ack_var;

	if(clk'event and (clk = '1')) then
		if(reset = '1') then
			fsm_state <= IDLE;
			valids_vector <= (others => '0');
			tags_vector <= (others => '0');
			last_written_index <= (2**log_number_of_entries);
			lookup_valid_reg <= '0';
		else
			fsm_state <= next_fsm_state_var;
			lookup_valid_reg <= next_lookup_valid_var;
			valids_vector <= next_valids_var;
			tags_vector   <= tagArrayToVector(next_tags_var);
			last_written_index <= next_last_written_index_var;
		end if;
	end if;
   end process;

   lookup_valid(0) <= lookup_valid_reg;

end genericFullyAssociativeMemoryNoDataArch;

		
	
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.BaseComponents.all;

library AjitCustom;
use AjitCustom.AjitCustomComponents.all;


-- a generic fully associative memory for use in the MMU TLB.
entity genericFullyAssociativeMemoryNoData_Operator is
	generic (tag_width: integer := 8; log_number_of_entries: integer := 6; ignore_collisions: boolean := true);
	port (  sample_req: in boolean;
		sample_ack: out boolean;
		update_req: in boolean;
		update_ack: out boolean;

		-- clear all valids.
		clear_flag: in std_logic_vector(0 downto 0);

		-- add entry
		erase_flag: in std_logic_vector(0 downto 0);
		write_flag: in std_logic_vector(0 downto 0);
		write_tag : in std_logic_vector(tag_width-1 downto 0);

		-- lookup entry
		lookup_flag: in std_logic_vector(0 downto 0);
		lookup_tag : in std_logic_vector(tag_width-1 downto 0);
		lookup_valid: out std_logic_vector(0 downto 0);

		clk,reset: in std_logic);

end entity genericFullyAssociativeMemoryNoData_Operator;


architecture simpleTon of genericFullyAssociativeMemoryNoData_Operator is
	signal start_req, start_ack: std_logic;
	signal fin_req, fin_ack: std_logic;
	signal br_lookup_valid: std_logic_vector(0 downto 0);

   	signal update_ack_sig: boolean;

begin

   p2l: Sample_Pulse_To_Level_Translate_Entity
                generic map(name => "genericFullyAssociativeMemoryNoData-Operator-p2l")
                port map (rL => sample_req, rR => start_req,
                                aL => sample_ack, aR => start_ack,
                                        clk => clk, reset => reset);
   l2p: Level_To_Pulse_Translate_Entity
		generic map(name => "genericFullyAssociativeMemoryNoData-Operator-l2p")
		port map (rL => fin_req, rR => update_req,
				aL => fin_ack, aR => update_ack_sig, clk => clk, reset => reset);


   update_ack <= update_ack_sig;


   br: BypassRegister 
		generic map(data_width => 1, bypass => true)
		port map (clk => clk, reset => reset, din => br_lookup_valid, enable => update_ack_sig, 
					q => lookup_valid);

   bmem: genericFullyAssociativeMemoryNoData
			generic map (tag_width => tag_width, 
					log_number_of_entries => log_number_of_entries,
					ignore_collisions => ignore_collisions)
			port map (
				start_req => start_req,
				start_ack => start_ack,
				fin_req =>   fin_req,
				fin_ack =>   fin_ack,
    				clear_flag => clear_flag,
    				write_flag => write_flag,
				write_tag => write_tag,
				erase_flag => erase_flag,
				lookup_flag => lookup_flag,
				lookup_tag => lookup_tag,
    				lookup_valid => br_lookup_valid,
    				clk => clk, reset => reset);

end simpleTon;

library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.mem_component_pack.all;


-- a generic set associative memory for potential use in the MMU TLB.
--   This could probably be used in the caches as well..
entity genericSetAssociativeMemory is
	generic (
			-- width of tag.
			tag_width: integer := 8;
			-- width of data.
			data_width: integer := 32;
			-- size of the set associative memory is 2**log_number_of_entries
			log_number_of_entries: integer := 8;
			-- 0 means direct mapped.
			log_associativity: integer := 0;
			-- ignore write->lookup collisions?
			ignore_collisions: boolean := true;
			-- use memory cuts or registers?
			use_mem_cuts: boolean:= true;
			-- ignore data, behave like a set and not a map.
			g_ignore_data: boolean := false
		);
	port (  start_req: in std_logic;
		start_ack: out std_logic;
		fin_req: in std_logic;
		fin_ack: out std_logic;

		-- clear all valids.
		clear_flag: in std_logic_vector(0 downto 0);

		-- add/erase entry specified by write_* ports.
		erase_flag: in std_logic_vector(0 downto 0);
		write_flag: in std_logic_vector(0 downto 0);
		
		-- write data 
		write_data: in std_logic_vector(data_width-1 downto 0);
		-- write tag (computed by environment)
		write_tag : in std_logic_vector(tag_width-1 downto 0);
		-- write set id (specified by environment)
		write_set_id: in std_logic_vector((log_number_of_entries-log_associativity)-1 downto 0);

		-- lookup entry
		lookup_flag: in std_logic_vector(0 downto 0);
		-- lookup tag.
		lookup_tag : in std_logic_vector(tag_width-1 downto 0);
		-- lookup set id.
		lookup_set_id: in std_logic_vector((log_number_of_entries-log_associativity)-1 downto 0);
		-- lookup is valid.. hit.
		lookup_valid: out std_logic_vector(0 downto 0);
		-- lookup data.
		lookup_data: out std_logic_vector(data_width-1 downto 0);
		clk,reset: in std_logic);

end entity genericSetAssociativeMemory;


-- read and then write.
architecture genericSetAssociativeMemoryArch of genericSetAssociativeMemory is


	constant number_of_entries: integer := (2**log_number_of_entries);
	constant number_of_elements_in_set: integer := (2**log_associativity);
	constant number_of_sets: integer := (2**(log_number_of_entries - log_associativity));

	-- tags for all entries in a set are maintained in a single word.

	-- tags for the set, prefixed by most-recently-updated index.
	constant set_tag_word_length: integer := (log_associativity + (number_of_elements_in_set*tag_width));

	-- data for all entries in a set is maintained in a single word.
	constant set_data_word_length: integer := (number_of_elements_in_set*data_width);

	-- number of address bits to identify set.
	constant n_set_address_bits: integer := (log_number_of_entries - log_associativity);

	-- separate valids vector for ease of clearing.
	signal valids : std_logic_vector(number_of_entries-1 downto 0);
		
	-- write information.
	signal erase_flag_reg: std_logic_vector(0 downto 0);
	signal write_flag_reg: std_logic_vector(0 downto 0);
	signal write_data_reg: std_logic_vector(data_width-1 downto 0);
	signal write_tag_reg : std_logic_vector(tag_width-1 downto 0);
	signal write_set_id_reg: std_logic_vector((log_number_of_entries-log_associativity)-1 downto 0);

	-- lookup information.
	signal lookup_flag_reg: std_logic_vector(0 downto 0);
	signal lookup_tag_reg : std_logic_vector(tag_width-1 downto 0);
	signal lookup_set_id_reg: std_logic_vector((log_number_of_entries-log_associativity)-1 downto 0);


	signal lookup_recorded_valid, lookup_recorded_valid_reg : std_logic;

	-- tag word is last-written-id  (tag)* .  This is stored in tag memory..
	subtype TagRecord is 
		std_logic_vector(set_tag_word_length-1 downto 0);
	type TagArray is array (natural range <>) of std_logic_vector(tag_width-1 downto 0);

	function tagArrayToVector (x: TagArray) 
		return std_logic_vector is
		alias twa : TagArray(number_of_elements_in_set-1 downto 0) is x;
		variable ret_var : std_logic_vector(number_of_elements_in_set*tag_width -1 downto 0);
	begin
		for I in 0 to number_of_elements_in_set-1 loop
			ret_var(((I+1)*tag_width)-1 downto (I*tag_width)) := twa(I);
		end loop;
		return(ret_var);
	end function;
	function tagVectorToArray (x: std_logic_vector) return TagArray is
		alias tx : std_logic_vector(number_of_elements_in_set*tag_width - 1 downto 0) is x;
		variable ret_var: TagArray(number_of_elements_in_set-1 downto 0);
	begin
		for I in 0 to number_of_elements_in_set-1 loop
			 ret_var(I) := tx(((I+1)*tag_width)-1 downto (I*tag_width));
		end loop;
		return(ret_var);
	end function;
		


	subtype DataRecord is 
		std_logic_vector(set_data_word_length-1 downto 0);
	type DataArray is array (natural range <>) of std_logic_vector(data_width-1 downto 0);
	function dataArrayToVector (x: DataArray) 
		return std_logic_vector is
		alias twa : DataArray(number_of_elements_in_set-1 downto 0) is x;
		variable ret_var : std_logic_vector(number_of_elements_in_set*data_width -1 downto 0);
	begin
		for I in 0 to number_of_elements_in_set-1 loop
			ret_var(((I+1)*data_width)-1 downto (I*data_width)) := twa(I);
		end loop;
		return(ret_var);
	end function;
	function dataVectorToArray (x: std_logic_vector) return DataArray is
		alias tx : std_logic_vector(number_of_elements_in_set*data_width - 1 downto 0) is x;
		variable ret_var: DataArray(number_of_elements_in_set-1 downto 0);
	begin
		for I in 0 to number_of_elements_in_set-1 loop
			 ret_var(I) := tx(((I+1)*data_width)-1 downto (I*data_width));
		end loop;
		return(ret_var);
	end function;
	

	-- tag memory access signals.
	signal tag_mem_write_data, tag_mem_read_data, tag_mem_read_data_reg, tag_mem_lookup_data: TagRecord;
	signal tag_mem_address: std_logic_vector(((log_number_of_entries-log_associativity)-1) downto 0);
	signal tag_mem_enable, tag_mem_write_bar: std_logic;

	-- data memory access signals
	signal data_mem_write_data, data_mem_read_data, data_mem_read_data_reg, data_mem_lookup_data: DataRecord;
	signal data_mem_address: std_logic_vector((log_number_of_entries-log_associativity)-1 downto 0);
	signal data_mem_enable, data_mem_write_bar: std_logic;

	-- FSM state
	type sFsmState is (INIT_STATE, IDLE, READ_FOR_WRITE, WRITE_STATE);
	signal fsm_state : sFsmState;

	-- flag used to indicate when tag lookup read data is to be sampled.
	signal record_lookup_outputs: boolean;

	-- index of lookup information in the set.
	--   note the invalid value 2**log_associativity.
	signal lookup_index_in_set: integer range 0 to number_of_elements_in_set;
	signal lookup_set_id_int : integer range 0 to number_of_sets-1;
	signal index_in_set : integer range 0 to number_of_elements_in_set;

	signal collision_flag_reg, erase_collision_flag_reg: std_logic;

	function extractLastWrittenIndex(x: TagRecord) 
			return integer is
		variable ret_var: integer range 0 to number_of_elements_in_set-1;
	begin
		ret_var := to_integer(unsigned(x(set_tag_word_length-1 downto 
								(number_of_elements_in_set*tag_width))));
		return(ret_var);
	end function;

	function findMatchingIndexInSet(tag_data: std_logic_vector;
					 svalids: std_logic_vector;
					 tag: std_logic_vector) return
			integer is
		alias ltag_mem_lookup_data: std_logic_vector(tag_data'length-1 downto 0) is tag_data;
		alias ltag: std_logic_vector(tag'length-1 downto 0) is tag;
		alias lsvalids: std_logic_vector(number_of_elements_in_set-1 downto 0) is svalids;

		variable ret_var: integer range 0 to number_of_elements_in_set;
	begin
		ret_var := number_of_elements_in_set;
		for I in 0 to number_of_elements_in_set-1 loop
			if(ltag_mem_lookup_data(((I+1)*tag_width)-1 downto (I*tag_width)) = ltag) then
				if(lsvalids(I) = '1') then
					ret_var := I;
					exit;
				end if;
			end if;
		end loop;
		return(ret_var);
	end function;

	function findInsertIndexInSet (tag_record: TagRecord;
					set_id_var: integer;
					v: std_logic_vector;
					wtag: std_logic_vector)
		return integer is
		alias ltag_mem_read_data: std_logic_vector(tag_record'length-1 downto 0) is tag_record;
		alias lwrite_tag: std_logic_vector(wtag'length-1 downto 0) is wtag;
		alias lvalids: std_logic_vector(number_of_entries-1 downto 0) is v;

		variable ret_var,t_var: integer range 0 to number_of_elements_in_set-1;
		variable found_flag: boolean;
	begin
		ret_var := 0;
		found_flag := false;
		for I in 0 to number_of_elements_in_set-1 loop
			if(ltag_mem_read_data(((I+1)*tag_width)-1 downto (I*tag_width)) = lwrite_tag) 
				and (lvalids((set_id_var*number_of_elements_in_set)+I) = '1') then
				ret_var := I;
				found_flag := true;
				exit;
			end if;
		end loop;
		if(not found_flag) then
			t_var := extractLastWrittenIndex(ltag_mem_read_data);
			if(t_var >= number_of_elements_in_set-1) then
				ret_var := 0;
			else
				ret_var := (t_var + 1);
			end if;
		end if;
		return(ret_var);
	end function;

						
	function insertDataItem(x_vec: std_logic_vector;
				 index: integer; 
				  x: std_logic_vector) return std_logic_vector is
		alias lx_vec: std_logic_vector(x_vec'length-1 downto 0) is x_vec;
		alias lx : std_logic_vector(x'length-1 downto 0) is x;
		variable ret_var: std_logic_vector(number_of_elements_in_set*data_width-1 downto 0);
		variable dwa : DataArray(number_of_elements_in_set-1 downto 0);
	begin
		dwa := dataVectorToArray(lx_vec);
		dwa(index) := lx;
		ret_var := dataArrayToVector(dwa);

		return(ret_var);
	end function;

	function insertTagItem(x_vec: std_logic_vector;
				 index: integer; 
				  x: std_logic_vector) return std_logic_vector is
		alias lx_vec: std_logic_vector(number_of_elements_in_set*tag_width-1 downto 0) is x_vec;
		alias lx : std_logic_vector(tag_width-1 downto 0) is x;
		variable ret_var: std_logic_vector(number_of_elements_in_set*tag_width-1 downto 0);
		variable twa : TagArray(number_of_elements_in_set-1 downto 0);
	begin

		twa := tagVectorToArray(lx_vec);
		twa(index) := lx;
		ret_var := tagArrayToVector(twa);

		return(ret_var);
	end function;

	function determineValidity(v: std_logic_vector; set_id: integer; idx_in_set: integer)
		return std_logic is
		variable ret_var: std_logic;
	begin
		ret_var := '0';
		if(idx_in_set < number_of_elements_in_set) then
			if(v((set_id*number_of_elements_in_set)+idx_in_set) = '1') then
				ret_var := '1';
			end if;
		end if;
		return(ret_var);
	end function;

	function extractDataFromSet (r: std_logic_vector; index: integer)
		return std_logic_vector is
		variable ret_var: std_logic_vector(data_width-1 downto 0);

		alias lr: std_logic_vector(r'length-1 downto 0) is r;
		variable dwa : DataArray(number_of_elements_in_set-1 downto 0);
	begin
		dwa := dataVectorToArray(lr);
		ret_var := (others => '0');

		if(index < number_of_elements_in_set) then
			ret_var := dwa(index);
		end if;

		return(ret_var);
	end function;

	function updateValids(nv: std_logic_vector; sid: integer; iid: integer; vval: std_logic)
		return std_logic_vector is
		alias lnv : std_logic_vector(nv'length-1 downto 0) is nv;
		variable ret_var: std_logic_vector(nv'length-1 downto 0);
	begin
		ret_var := lnv;
		ret_var((sid*number_of_elements_in_set) + iid) := vval;
		return ret_var;
	end function;

	signal reset_counter: integer range 0 to number_of_sets-1;

	signal done_reg: std_logic;
	signal ignore_collision_generic_sig: boolean;
begin

	ignore_collision_generic_sig <= ignore_collisions;


				
	--
	-- state machine.
	--    For lookups, the sequence is 
	--		IDLE -> IDLE
	--                 (lookup-read)
	--	      or IDLE -> IDLE
	--                 (lookup-read)
	--
	--    For lookups and simultaneous writes the
	--	sequence is
	--		IDLE  ->  READ_FOR_WRITE  -> WRITE     ->    IDLE
	--                (lookup-read)      (read-for-write)  (write) 
	--
	--    For writes, the squence is
	--		IDLE ->              WRITE   -> 	 IDLE
	--                (read-for-write)         (write)
	--    
	process(clk, reset, fsm_state, start_req, fin_req, clear_flag, write_flag, erase_flag, lookup_flag,
				valids, tag_mem_read_data, data_mem_read_data,
				write_data, write_data_reg, lookup_tag, lookup_tag_reg,
				write_set_id, write_set_id_reg,
				lookup_set_id, lookup_set_id_reg, done_reg, collision_flag_reg,
				erase_collision_flag_reg)
		variable next_fsm_state_var: sFsmState;
		variable tag_mem_enable_var, tag_mem_write_bar_var: std_logic;
		variable data_mem_enable_var, data_mem_write_bar_var: std_logic;
		variable start_ack_var: std_logic;
		variable latch_inputs_var: std_logic;
		variable collision_var : std_logic;
		variable erase_collision_var : std_logic;

		variable next_valids_var: std_logic_vector(number_of_entries-1 downto 0);
		variable next_done_var: std_logic;

		variable tag_mem_address_var: std_logic_vector((log_number_of_entries-log_associativity)-1 downto 0);
		variable data_mem_address_var: std_logic_vector((log_number_of_entries-log_associativity)-1 downto 0);

		variable tag_mem_write_data_var: TagRecord;
		variable data_mem_write_data_var: DataRecord;


		variable next_record_lookup_outputs_var: boolean;
		variable set_id_var : integer range 0 to number_of_sets-1;
		variable index_in_set_var : integer range 0 to number_of_elements_in_set;
	
		variable next_reset_counter_var: 
				integer range 0 to number_of_sets-1;
		variable valid_value_var: std_logic;

	begin

		collision_var := collision_flag_reg;
		erase_collision_var := erase_collision_flag_reg;
		valid_value_var := '0';

		next_done_var := done_reg;
		next_reset_counter_var := reset_counter;
		set_id_var := 0;
		next_record_lookup_outputs_var := false;

		index_in_set_var := 0;

		tag_mem_write_bar_var := '1';
		tag_mem_enable_var := '0';

		tag_mem_address_var := (others => '0');
		data_mem_address_var := (others => '0');

		tag_mem_write_data_var := (others => '0');
		data_mem_write_data_var := (others => '0');

		data_mem_write_bar_var := '1';
		data_mem_enable_var := '0';

		next_fsm_state_var := fsm_state;

		start_ack_var := '0';

		latch_inputs_var := '0';
		next_valids_var := valids;

		case fsm_state is
			when INIT_STATE => 
				tag_mem_enable_var := '1';
				tag_mem_write_bar_var := '0';
				tag_mem_write_data_var := (others => '0');
				tag_mem_address_var := 	
					std_logic_vector(to_unsigned(reset_counter,n_set_address_bits));
				if(reset_counter = number_of_sets-1) then
					next_fsm_state_var := IDLE;
				else
					next_reset_counter_var := reset_counter + 1;
				end if;
			when IDLE =>
				if((done_reg = '0') or (fin_req = '1')) then
					next_done_var := '0';

					-- can start again..
					start_ack_var := '1';
					if (start_req = '1') then
						collision_var := '0';
						erase_collision_var := '0';

						if ((not ignore_collisions) and 
						      (lookup_flag(0) = '1') and
							(clear_flag(0) = '0') and 
								((write_flag(0) = '1') or
									(erase_flag(0) = '1'))
								and (lookup_tag = write_tag) and
									(lookup_set_id = write_set_id)) then
							collision_var := '1';
							if(erase_flag(0) = '1') then
								erase_collision_var := '1';
							end if;
						end if;

						-- latch for read-for-write
						latch_inputs_var := '1';

						-- if init, then all valids are cleared.
						if(clear_flag(0) = '1') then
							next_valids_var := (others => '0');
						end if;
	
						-- Note: both lookup and write could be active
						if(lookup_flag(0) = '1') then
							-- read the set tag using the lookup address.
							tag_mem_enable_var := '1';
							tag_mem_address_var := 	lookup_set_id;
							-- read the data using the lookup address.
							data_mem_enable_var := '1';
							data_mem_address_var := lookup_set_id;
		
							-- in the next cycle, record the lookup outputs.
							next_record_lookup_outputs_var := true;

							if((write_flag(0) = '1')  or (erase_flag(0) = '1')) then
								-- need to read entry for write.
								next_fsm_state_var := READ_FOR_WRITE;
							else
								-- no write, done. stay in IDLE, set done_reg.
								next_done_var := '1';
							end if;
						elsif ((write_flag(0) = '1') or (erase_flag(0) = '1')) then
							-- read the tag using the write address.
							tag_mem_enable_var := '1';
							tag_mem_address_var := 	write_set_id;
							if(write_flag(0) = '1') then
								-- read the data using the write address.
								data_mem_enable_var := '1';
								data_mem_address_var :=	write_set_id;
							end if;
							next_fsm_state_var := WRITE_STATE;
						else
							-- stay in IDLE, and set done_reg
							next_done_var := '1';
						end if;
					end if;
				end if;
			when READ_FOR_WRITE => 
				-- read the set tag using the registered write address.
				tag_mem_enable_var := '1';
				tag_mem_address_var := 	write_set_id_reg;
				-- read the data using the registered write address.
				data_mem_enable_var := '1';
				data_mem_address_var :=	write_set_id_reg;
				next_fsm_state_var := WRITE_STATE;

				-- one more cycle!
				next_done_var := '0';

			when WRITE_STATE =>

				-- index of the set.
				set_id_var := to_integer(unsigned(write_set_id_reg));

				-- index in set at which word is written... return either a 
				-- matching index, or a free index, or an NMRU replacement index.
				-- 	 the set, and then find the index within the set.
				index_in_set_var := 
					findInsertIndexInSet(
								-- result of tag mem read.
								tag_mem_read_data, 
								-- set id.
								set_id_var,
								-- use set_id to extract the
								-- valids for the set.
								valids, 
								-- write tag to look for slot.
								write_tag_reg);

				if(erase_flag_reg(0) = '0') then 
					-- write the tag using the registered write information.
					tag_mem_enable_var := '1';
					tag_mem_write_bar_var  := '0';
					tag_mem_address_var := 	write_set_id_reg;

					-- tag mem entry.
					tag_mem_write_data_var((number_of_elements_in_set*tag_width)-1 downto 0) :=
					    insertTagItem(
 					       tag_mem_read_data((number_of_elements_in_set*tag_width)-1 downto 0),
								index_in_set_var, write_tag_reg);
					tag_mem_write_data_var(tag_mem_write_data'high downto 
   						   				number_of_elements_in_set*tag_width)
							:= std_logic_vector(to_unsigned(index_in_set_var, 
											log_associativity));

					-- write the data using the registered write information.
					data_mem_enable_var := '1';
					data_mem_write_bar_var  := '0';
					data_mem_address_var := write_set_id_reg;
					data_mem_write_data_var :=
						insertDataItem(data_mem_read_data, index_in_set_var, write_data_reg);
				end if;
	
				-- next valids..
				valid_value_var := (not erase_flag_reg(0));
				next_valids_var := 
					updateValids(next_valids_var, set_id_var, index_in_set_var, valid_value_var);

				-- go to IDLE...
				next_fsm_state_var := IDLE;
				next_done_var := '1';
		end case;

		tag_mem_write_data <= tag_mem_write_data_var;
		tag_mem_enable <= tag_mem_enable_var;
		tag_mem_write_bar <= tag_mem_write_bar_var;
		tag_mem_address <= tag_mem_address_var;

		data_mem_write_data 
				   <= data_mem_write_data_var;
		data_mem_enable    <= data_mem_enable_var;
		data_mem_write_bar <= data_mem_write_bar_var;
		data_mem_address   <= data_mem_address_var;

		index_in_set <= index_in_set_var;

		fin_ack <= done_reg;
		start_ack <= start_ack_Var;
		

		if(clk'event and clk = '1') then
			if(reset = '1') then
				fsm_state <= INIT_STATE;
				valids <= (others => '0');
				reset_counter <= 0;
				collision_flag_reg <= '0';
				erase_collision_flag_reg <= '0';
				done_reg <= '0';
			else
				fsm_state <= next_fsm_state_var;
				valids    <= next_valids_var;

				record_lookup_outputs <= next_record_lookup_outputs_var;
				collision_flag_reg  <= collision_var;
				erase_collision_flag_reg  <= erase_collision_var;

				done_reg <= next_done_var;

				if(latch_inputs_var = '1') then

					write_flag_reg <= write_flag;
					write_data_reg <= write_data;
					write_tag_reg  <= write_tag;
					write_set_id_reg <= write_set_id;

					lookup_flag_reg <= lookup_flag;
					lookup_tag_reg  <= lookup_tag;
					lookup_set_id_reg <= lookup_set_id;

					erase_flag_reg <= erase_flag;

				end if;

				reset_counter <= next_reset_counter_var;
			end if;
		end if;
	end process;

		
	-- record lookup values at the point they are available.
	process(clk, record_lookup_outputs, reset, tag_mem_read_data, data_mem_read_data)
	begin
		
		if(clk'event and clk = '1') then
			if (reset = '1') then 
				tag_mem_read_data_reg     <= (others => '0');
			elsif(record_lookup_outputs) then
				tag_mem_read_data_reg     <= tag_mem_read_data;
				data_mem_read_data_reg    <= data_mem_read_data;
			end if;
		end if;
	end process;
				
	tag_mem_lookup_data <= tag_mem_read_data when record_lookup_outputs 
					else tag_mem_read_data_reg when (lookup_flag_reg(0) = '1') 
						else (others => '0');
	data_mem_lookup_data <= data_mem_read_data when record_lookup_outputs 
					else data_mem_read_data_reg when (lookup_flag_reg(0) = '1') 
						else (others => '0');

	lookup_set_id_int       <= to_integer(unsigned(lookup_set_id_reg));

	-- will return (2**log_associativity if none found).
	process(tag_mem_lookup_data, lookup_set_id_int, lookup_tag_reg)
           variable sel_var: std_logic_vector(number_of_elements_in_set-1 downto 0);
        begin
	   for I in 0 to number_of_elements_in_set-1 loop
	   	sel_var(I) := valids((lookup_set_id_int*number_of_elements_in_set)+I);
	   end loop;
	   lookup_index_in_set <=  findMatchingIndexInSet(tag_mem_lookup_data, sel_var, lookup_tag_reg);
	end process;

	-- if in bounds, validity determined by looking at index.
	--  	Note: there was a bug here earlier.  The lookup valid value must be
	--		sampled at the correct point, since in the lookup + write
	--		case, the valids can get modified by the write and clobber
	--		the state for the lookup.
	lookup_recorded_valid     
		<=  lookup_flag_reg(0) and  (not erase_collision_flag_reg) and 
					(collision_flag_reg  or 
					    determineValidity(valids, lookup_set_id_int, lookup_index_in_set));
	process(clk, reset, record_lookup_outputs, lookup_set_id_int, lookup_index_in_set, valids)
	begin
		if(clk'event and (clk = '1')) then
			if(reset = '1') then	
				lookup_recorded_valid_reg <= '0';
			else
				if(record_lookup_outputs) then
					lookup_recorded_valid_reg <= lookup_recorded_valid;
				end if;
			end if;
		end if;
	end process;
	lookup_valid(0) <= lookup_recorded_valid when record_lookup_outputs else lookup_recorded_valid_reg;
	
	-- if in bounds, extract..
	lookup_data         <=  write_data_reg when (collision_flag_reg = '1')  else 
						extractDataFromSet (data_mem_lookup_data, lookup_index_in_set);


	
   memCutBB: if use_mem_cuts generate 
   	tag_bb: base_bank 
		generic map  (name => "genericSetAssociativeMemory:tag_base_bank", 
						g_addr_width => log_number_of_entries - log_associativity,
						g_data_width => set_tag_word_length)
		port map (
				datain => tag_mem_write_data,
				addrin => tag_mem_address,
				dataout => tag_mem_read_data,
				enable => tag_mem_enable,
				writebar => tag_mem_write_bar,
				clk => clk, reset => reset
			);
        UseDataGen: if (not g_ignore_data) generate 
   	  data_bb: base_bank 
		generic map  (name => "genericSetAssociativeMemory:data_base_bank", 
						g_addr_width => log_number_of_entries - log_associativity,
						g_data_width => set_data_word_length)
		port map (
				datain => data_mem_write_data,
				addrin => data_mem_address,
				dataout => data_mem_read_data,
				enable => data_mem_enable,
				writebar => data_mem_write_bar,
				clk => clk, reset => reset
			);
         end generate UseDataGen;

	IgnDataGen: if g_ignore_data generate
		data_mem_read_data <= (others => '0');
	end generate IgnDataGen;

   end generate memCutBB;
   regBB: if not use_mem_cuts generate 
   	tag_bb: base_bank_with_registers
		generic map  (name => "genericSetAssociativeMemory:tag_base_bank", 
						g_addr_width => log_number_of_entries - log_associativity,
						g_data_width => set_tag_word_length)
		port map (
				datain => tag_mem_write_data,
				addrin => tag_mem_address,
				dataout => tag_mem_read_data,
				enable => tag_mem_enable,
				writebar => tag_mem_write_bar,
				clk => clk, reset => reset
			);
        UseDataGen: if not g_ignore_data generate
   	  data_bb: base_bank_with_registers
		generic map  (name => "genericSetAssociativeMemory:data_base_bank", 
						g_addr_width => log_number_of_entries - log_associativity,
						g_data_width => set_data_word_length)
		port map (
				datain => data_mem_write_data,
				addrin => data_mem_address,
				dataout => data_mem_read_data,
				enable => data_mem_enable,
				writebar => data_mem_write_bar,
				clk => clk, reset => reset);
         end generate UseDataGen;

	IgnDataGen: if g_ignore_data generate
		data_mem_read_data <= (others => '0');
	end generate IgnDataGen;
   end generate regBB;
 

end genericSetAssociativeMemoryArch;

		
	
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.BaseComponents.all;

library AjitCustom;
use AjitCustom.AjitCustomComponents.all;


-- operator form of generic set associative memory for potential use in the MMU TLB.
--   This could probably be used in the caches as well..
entity genericSetAssociativeMemory_Operator is
	generic (
			-- width of tag.
			tag_width: integer := 8;
			-- width of data.
			data_width: integer := 32;
			-- size of the set associative memory is 2**log_number_of_entries
			log_number_of_entries: integer := 8;
			-- 0 means direct mapped.
			log_associativity: integer := 0;
			-- ignore write->lookup collisions?
			ignore_collisions: boolean := true;
			-- use memory cuts or registers?
			use_mem_cuts: boolean:= true;
			-- ignore data, behave like a set and not a map.
			g_ignore_data: boolean := false);
	port (  sample_req: in boolean;
		sample_ack: out boolean;
		update_req: in boolean;
		update_ack: out boolean;

		-- clear all valids.
		clear_flag: in std_logic_vector(0 downto 0);

		-- add/erase entry specified by write_* ports.
		erase_flag: in std_logic_vector(0 downto 0);
		write_flag: in std_logic_vector(0 downto 0);
		
		-- write data 
		write_data: in std_logic_vector(data_width-1 downto 0);
		-- write tag (computed by environment)
		write_tag : in std_logic_vector(tag_width-1 downto 0);
		-- write set id (specified by environment)
		write_set_id: in std_logic_vector((log_number_of_entries-log_associativity)-1 downto 0);

		-- lookup entry
		lookup_flag: in std_logic_vector(0 downto 0);
		-- lookup tag.
		lookup_tag : in std_logic_vector(tag_width-1 downto 0);
		-- lookup set id.
		lookup_set_id: in std_logic_vector((log_number_of_entries-log_associativity)-1 downto 0);
		-- lookup is valid.. hit.
		lookup_valid: out std_logic_vector(0 downto 0);
		-- lookup data.
		lookup_data: out std_logic_vector(data_width-1 downto 0);
		clk,reset: in std_logic);

end entity genericSetAssociativeMemory_Operator;


architecture SimpleTon of genericSetAssociativeMemory_Operator is
	signal start_req, start_ack: std_logic;
	signal fin_req, fin_ack: std_logic;

	signal br_lookup_data: std_logic_vector(data_width-1 downto 0);
	signal br_lookup_valid: std_logic_vector(0 downto 0);
	signal br_data_in, br_data_out: std_logic_vector(data_width downto 0);

   	signal update_ack_sig: boolean;
begin

   p2l: Sample_Pulse_To_Level_Translate_Entity
                generic map(name => "genericSetAssociativeMemory-Operator-p2l")
                port map (rL => sample_req, rR => start_req,
                                aL => sample_ack, aR => start_ack,
                                        clk => clk, reset => reset);

   l2p: Level_To_Pulse_Translate_Entity
		generic map(name => "genericSetAssociativeMemory-Operator-l2p")
		port map (rL => fin_req, rR => update_req,
				aL => fin_ack, aR => update_ack_sig, clk => clk, reset => reset);

   update_ack <= update_ack_sig;

   br_data_in <= br_lookup_valid & br_lookup_data;


   br: BypassRegister 
		generic map(data_width => data_width+1, bypass => true)
		port map (clk => clk, reset => reset, din => br_data_in, enable => update_ack_sig, 
					q => br_data_out);

   lookup_valid(0) <= br_data_out(data_width);
   lookup_data <= br_data_out(data_width-1 downto 0);

   bmem: genericSetAssociativeMemory 
		generic map (
				tag_width => tag_width,
				data_width => data_width,
				log_number_of_entries => log_number_of_entries,
				log_associativity => log_associativity,
				ignore_collisions => ignore_collisions,
				use_mem_cuts => use_mem_cuts,
				g_ignore_data => g_ignore_data)
		port map (
		  	start_req => start_req,
		  	start_ack => start_ack,
		  	fin_req => fin_req,
	   	  	fin_ack => fin_ack,
		  	clear_flag => clear_flag,
		  	erase_flag => erase_flag,
		  	write_flag => write_flag,
		  	write_data => write_data,
		  	write_tag  => write_tag ,
		  	write_set_id => write_set_id,
		  	lookup_flag => lookup_flag,
		  	lookup_tag  => lookup_tag ,
		  	lookup_set_id => lookup_set_id,
		  	lookup_valid => br_lookup_valid,
		  	lookup_data => br_lookup_data,
		  	clk => clk,
		  	reset => reset);

end SimpleTon;

-- VHDL global package produced by vc2vhdl from virtual circuit (vc) description 
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library ahir;
use ahir.BaseComponents.all;
use ahir.mem_component_pack.all;

library AjitCustom;

entity genericDirectMappedAssociativeMemory is -- 
  generic (tag_width: integer := 32;
		data_width: integer := 67;
		log2_number_of_entries : integer := 8);
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    init_flag : in  std_logic_vector(0 downto 0);
    insert_flag : in  std_logic_vector(0 downto 0);
    insert_tag : in  std_logic_vector(tag_width-1 downto 0);
    insert_data : in  std_logic_vector(data_width-1 downto 0);
    lookup_flag : in  std_logic_vector(0 downto 0);
    lookup_tag : in  std_logic_vector(tag_width-1 downto 0);
    lookup_match : out  std_logic_vector(0 downto 0);
    lookup_data : out  std_logic_vector(data_width-1 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity genericDirectMappedAssociativeMemory;
architecture dm_Operator_arch of genericDirectMappedAssociativeMemory is -- 

    constant number_of_entries: integer := (2**log2_number_of_entries);
    constant reduced_tag_width : integer := (tag_width - log2_number_of_entries);
    constant augmented_data_width : integer := (data_width + reduced_tag_width);

    signal mem_write_address: std_logic_vector(log2_number_of_entries-1 downto 0);
    signal mem_write_data, ignore_data_0: std_logic_vector(augmented_data_width-1 downto 0);
    signal mem_write_enable, mem_write_enable_bar: std_logic;

    signal mem_read_address: std_logic_vector(log2_number_of_entries-1 downto 0);
    signal mem_read_address_delayed: std_logic_vector(log2_number_of_entries-1 downto 0);
    signal mem_read_data, zero_data_1: std_logic_vector(augmented_data_width-1 downto 0);
    signal mem_read_enable: std_logic;

    signal valids: std_logic_vector(number_of_entries-1 downto 0);

    signal joined_sig: Boolean;
    signal trigger: std_logic;

    signal insert_tag_reduced, 
		lookup_tag_reduced: std_logic_vector((tag_width-log2_number_of_entries)-1 downto 0);
    signal trigger_reg  : std_logic;


    signal const_one : std_logic;
  
    signal aggr_result, aggr_result_prereg, aggr_result_reg : std_logic_vector(data_width downto 0);
    signal write_read_clash, write_read_clash_reg : boolean;

    signal tag_in_mem_read_data: std_logic_vector(reduced_tag_width-1 downto 0);
    signal lookup_tag_match: boolean;
    
    signal init_flag_reg : std_logic_vector(0 downto 0);

begin --  

    insert_tag_reduced <= insert_tag(tag_width-1 downto log2_number_of_entries);

    zero_data_1 <= (others => '0');
    const_one <= '1';


    trigger <= '1' when joined_sig else '0';

    trig_join: join2 generic map (name => "bpbV2:trig-join", bypass => true)
			port map (pred0 => sample_req, pred1 => update_req,
					symbol_out => joined_sig, clk => clk, reset => reset);
   
    sample_ack <= joined_sig;

    process(clk, reset)
    begin
	if(clk'event and clk='1') then
		if(reset = '1') then
			update_ack <= false;
			trigger_reg <= '0';
			write_read_clash_reg <= false;
			init_flag_reg(0) <= '0';
		else

			mem_read_address_delayed <= mem_read_address;
    		        lookup_tag_reduced <= lookup_tag(tag_width-1 downto log2_number_of_entries);
			update_ack <= joined_sig;
	
			trigger_reg <= trigger;
			write_read_clash_reg <= write_read_clash;
			if(trigger  = '1') then
				init_flag_reg(0) <= init_flag(0);
			end if;

		end if;
	end if;
    end process;

    mem_write_address <= insert_tag (log2_number_of_entries-1 downto 0);
    mem_write_data    <= insert_tag_reduced & insert_data;

    mem_write_enable  <= (not init_flag(0)) and trigger and insert_flag(0);
    mem_write_enable_bar <= not mem_write_enable;

    mem_read_address  <= lookup_tag (log2_number_of_entries-1 downto 0);
    mem_read_enable   <= (not init_flag(0)) and trigger;

    write_read_clash <= joined_sig and (mem_write_address = mem_read_address);

    process(clk, reset)
    begin
        if(clk'event and (clk='1')) then
		if((reset = '1') or ((trigger = '1') and (init_flag(0) = '1'))) then
			valids <= (others => '0');
		else
			if ((trigger = '1') and (insert_flag(0) = '1')) then
				valids(to_integer(unsigned(mem_write_address))) <= '1';
			end if;
		end if;
	end if;
    end process;
     
    dpram: base_bank_dual_port
		generic map (name =>  "bpbV2:dpram",
				g_addr_width => log2_number_of_entries,
					g_data_width => augmented_data_width)
		port map (
			datain_0 => mem_write_data,
			dataout_0 => ignore_data_0,
			addrin_0 => mem_write_address,
			enable_0 => mem_write_enable,
			writebar_0 => mem_write_enable_bar,
			datain_1 => zero_data_1,
			dataout_1 => mem_read_data,
			addrin_1 => mem_read_address,
			enable_1   => mem_read_enable,
			writebar_1 => const_one,
			clk => clk , reset => reset);
			

	process(valids, trigger_reg, lookup_tag_match, mem_read_data)
		variable result_var: std_logic_vector(data_width downto 0);
	begin
		result_var := (others => '0');
		if(lookup_tag_match) then 
			result_var(data_width) := trigger_reg;
		else
			result_var(data_width) := '0';
		end if;

		result_var(data_width-1 downto 0) := mem_read_data(data_width-1 downto 0);

		aggr_result_prereg <= result_var;
	end process;

	lookup_tag_match <= 
		((init_flag_reg(0) = '0') and
			(valids(to_integer(unsigned(mem_read_address_delayed))) = '1') and
			(mem_read_data(augmented_data_width-1  downto data_width) = 
						lookup_tag_reduced) and (not write_read_clash_reg));

	-- Important: need to maintain the bpb result until the next trigger..
	process(clk, reset)
	begin
		if(clk'event and clk = '1') then
			if(reset = '1') then
				aggr_result_reg <= (others => '0');
			elsif (trigger_reg = '1') then
				aggr_result_reg <= aggr_result_prereg;
			end if;
		end if;
	end process;
	aggr_result <= aggr_result_prereg when (trigger_reg = '1') else aggr_result_reg;

	lookup_match(0) <= aggr_result(data_width);
	lookup_data  <= aggr_result(data_width-1 downto 0);

end dm_Operator_arch;
library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.mem_component_pack.all;
use ahir.BaseComponents.all;

entity genericSinglePortMemory_Operator is

	generic ( data_width: integer := 32; address_width: integer := 32);
	port (sample_req: in boolean;
		sample_ack: out boolean;
		update_req: in boolean;
		update_ack: out boolean;

		enable: in std_logic_vector(0 downto 0);	
		write_bar: in std_logic_vector(0 downto 0);	
		write_data: in std_logic_vector(data_width-1 downto 0);
		read_data: out std_logic_vector(data_width-1 downto 0);
		address: in std_logic_vector(address_width-1 downto 0);

		clk,reset: in std_logic);

end entity genericSinglePortMemory_Operator;


architecture SimpleBehavioural of genericSinglePortMemory_Operator is
	signal jsig: boolean;
	signal enable_sig: std_logic;
begin
	ji: join2 generic map (bypass => true, name => "genericSinglePortMemory:join2")
		port map (pred0 => sample_req, pred1 => update_req, symbol_out => jsig,
					clk => clk, reset => reset);

	enable_sig <= '1' when jsig else '0';

	sample_ack <= jsig;

	process(clk, reset)
	begin
		if(clk'event and (clk = '1')) then
			if(reset = '1') then
				update_ack <= false;
			else
				update_ack <= jsig;
			end if;
		end if;
	end process;

	bb: base_bank
		generic map (name => "genericSinglePortMemory:bb", g_addr_width => address_width,
					g_data_width => data_width)
		port map(
				datain => write_data,
				dataout => read_data,
				enable => enable_sig,
				writebar => write_bar(0),
				addrin => address,
				clk => clk, reset => reset);

end SimpleBehavioural;

library ieee;
use ieee.std_logic_1164.all;

library ahir;
use ahir.mem_component_pack.all;
use ahir.BaseComponents.all;

entity genericDualPortMemory_Operator is

	generic ( data_width: integer := 32; address_width: integer := 32);
	port (sample_req: in boolean;
		sample_ack: out boolean;
		update_req: in boolean;
		update_ack: out boolean;

		enable_0: in std_logic_vector(0 downto 0);	
		write_bar_0: in std_logic_vector(0 downto 0);	
		write_data_0: in std_logic_vector(data_width-1 downto 0);
		read_data_0: out std_logic_vector(data_width-1 downto 0);
		address_0: in std_logic_vector(address_width-1 downto 0);

		enable_1: in std_logic_vector(0 downto 0);	
		write_bar_1: in std_logic_vector(0 downto 0);	
		write_data_1: in std_logic_vector(data_width-1 downto 0);
		read_data_1: out std_logic_vector(data_width-1 downto 0);
		address_1: in std_logic_vector(address_width-1 downto 0);

		clk,reset: in std_logic);

end entity genericDualPortMemory_Operator;


architecture SimpleBehavioural of genericDualPortMemory_Operator is
	signal jsig: boolean;
	signal enable_sig: std_logic;
	signal enable_sig_0, enable_sig_1: std_logic;
begin
	ji: join2 generic map (bypass => true, name =>  "genericDualPortMemory:join2")
		port map (pred0 => sample_req, pred1 => update_req, symbol_out => jsig,
					clk => clk, reset => reset);

	enable_sig <= '1' when jsig else '0';
	enable_sig_0 <= enable_sig and enable_0(0);
	enable_sig_1 <= enable_sig and enable_1(0);

	sample_ack <= jsig;

	process(clk, reset)
	begin
		if(clk'event and (clk = '1')) then
			if(reset = '1') then
				update_ack <= false;
			else
				update_ack <= jsig;
			end if;
		end if;
	end process;

	bb: base_bank_dual_port
		generic map (name => ":genericDualPortMemory:bb", g_addr_width => address_width,
					g_data_width => data_width)
		port map(
				datain_0 => write_data_0,
				dataout_0 => read_data_0,
				enable_0 => enable_sig_0,
				writebar_0 => write_bar_0(0),
				addrin_0 => address_0,

				datain_1 => write_data_1,
				dataout_1 => read_data_1,
				enable_1 => enable_sig_1,
				writebar_1 => write_bar_1(0),
				addrin_1 => address_1,

				clk => clk, reset => reset);

end SimpleBehavioural;

library ieee;
use ieee.std_logic_1164.all;

library AjitCustom;
use AjitCustom.AjitCoreConfigurationPackage.all;
use AjitCustom.AjitGlobalConfigurationPackage.all;
use AjitCustom.AjitCustomComponents.all;

entity accessRlutBase_Operator is -- 
  generic (
		g_LOG_BASE_PAGE_SIZE: integer;
		g_LOG_CACHE_LINE_SIZE: integer;
		g_CACHE_WAY_SIZE: integer;
		g_RLUT_TAG_WIDTH : integer;
		g_RLUT_REDUCED_DATA_WIDTH: integer;
		g_RLUT_LOG_N_SETS: integer;
		g_RLUT_LOG_MEMORY_SIZE: integer;
		g_RLUT_LOG_SET_SIZE: integer
	);
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    lookup : in  std_logic_vector(0 downto 0);
    update : in  std_logic_vector(0 downto 0);
    clear : in  std_logic_vector(0 downto 0);
    physical_addr_of_line : in  std_logic_vector(29 downto 0);
    virtual_addr_of_line : in  std_logic_vector(25 downto 0);
    syn_invalidate_word : out  std_logic_vector(26 downto 0);
    clk, reset: in std_logic
    -- 
  );
end entity;

architecture SimpleStruct of accessRlutBase_Operator  is
	signal zero_sig: std_logic_vector(0 downto 0);
	signal write_tag: std_logic_vector(g_RLUT_TAG_WIDTH-1 downto 0);
	signal set_id: std_logic_vector(g_RLUT_LOG_N_SETS-1 downto 0);
	signal sample_ack_sig: boolean;

	signal hit: std_logic_vector(0 downto 0);
	signal hit_va: std_logic_vector(25 downto 0);
	signal pa_reg: std_logic_vector((g_LOG_BASE_PAGE_SIZE - g_LOG_CACHE_LINE_SIZE)-1 downto 0);

	constant ZZSIZE : integer := 
		(26 - (g_RLUT_REDUCED_DATA_WIDTH + (g_LOG_BASE_PAGE_SIZE - g_LOG_CACHE_LINE_SIZE)));

	constant c_triv_threshold : integer := (2 ** (g_LOG_BASE_PAGE_SIZE - g_LOG_CACHE_LINE_SIZE));

begin
	write_tag <= physical_addr_of_line (29 downto g_RLUT_LOG_N_SETS);
	set_id    <= physical_addr_of_line (g_RLUT_LOG_N_SETS-1 downto 0);

	zero_sig(0) <= '0';
	sample_ack <= sample_ack_sig;

	process(clk, reset, sample_ack_sig)
	begin
  	  if(clk'event and clk = '1') then
		if(sample_ack_sig) then
			pa_reg <= 
				physical_addr_of_line((g_LOG_BASE_PAGE_SIZE - g_LOG_CACHE_LINE_SIZE)-1 downto 0);
		end if;
	  end if;
	end process;

    NonTrivGen:  if (g_CACHE_WAY_SIZE > c_triv_threshold) generate
     bb: block 
	signal hit_va_reduced, va_reduced: std_logic_vector(g_RLUT_REDUCED_DATA_WIDTH-1 downto 0);
	signal zz_fill: std_logic_vector(ZZSIZE -1  downto 0);
     begin

	zz_fill <= (others => '0');

	-- need to keep only 3-bits for 32KB cache.
	va_reduced <= virtual_addr_of_line 
		((g_RLUT_REDUCED_DATA_WIDTH + g_LOG_BASE_PAGE_SIZE - g_LOG_CACHE_LINE_SIZE)-1 downto
					(g_LOG_BASE_PAGE_SIZE - g_LOG_CACHE_LINE_SIZE));

	basemem:genericSetAssociativeMemory_Operator
			generic map(
					tag_width => g_RLUT_TAG_WIDTH,
					data_width => g_RLUT_REDUCED_DATA_WIDTH,
					log_number_of_entries => g_RLUT_LOG_MEMORY_SIZE,
					log_associativity     => g_RLUT_LOG_SET_SIZE,
					ignore_collisions => true,
					use_mem_cuts => true,
					g_ignore_data => false -- use as a map.
				    )
			port map(
					sample_req => sample_req,
					sample_ack => sample_ack_sig,
					update_req => update_req,
					update_ack => update_ack,
					clear_flag => clear,
					erase_flag => zero_sig,
					write_flag => update,
					write_data => va_reduced,
					write_tag =>  write_tag,
					write_set_id => set_id,
					lookup_flag => lookup,
					lookup_tag => write_tag,
					lookup_set_id => set_id,
					lookup_valid => hit,
					lookup_data => hit_va_reduced,
					clk => clk, reset => reset);
	
        hit_va <= zz_fill & hit_va_reduced & pa_reg;
	syn_invalidate_word <= hit & hit_va;

      end block bb;
    end generate NonTrivGen;

	-- The trivial case,   hit needs to be calculated but
	-- The bits PA[11:6] are sent as the matching VA for invalidation.
    TrivGen:  if (g_CACHE_WAY_SIZE <= c_triv_threshold) generate
      bb: block
	signal hit_va_reduced, va_reduced: std_logic_vector(0 downto 0);
      begin
	-- 1-bit data, sacrificial..
	va_reduced(0) <= '0';

	basemem:genericSetAssociativeMemory_Operator
			generic map(
					tag_width => g_RLUT_TAG_WIDTH,
					data_width => 1,
					log_number_of_entries => g_RLUT_LOG_MEMORY_SIZE,
					log_associativity     => g_RLUT_LOG_SET_SIZE,
					ignore_collisions => true,
					use_mem_cuts => true,
					g_ignore_data => true -- use a set, not as a map
				    )
			port map(
					sample_req => sample_req,
					sample_ack => sample_ack_sig,
					update_req => update_req,
					update_ack => update_ack,
					clear_flag => clear,
					erase_flag => zero_sig,
					write_flag => update,
					write_data => va_reduced,
					write_tag =>  write_tag,
					write_set_id => set_id,
					lookup_flag => lookup,
					lookup_tag => write_tag,
					lookup_set_id => set_id,
					lookup_valid => hit,
					lookup_data => hit_va_reduced,
					clk => clk, reset => reset);
	
	-- in the trivial case, pa_reg is forwarded
	-- as the set id..
        process(hit, pa_reg)
           variable siw: std_logic_vector (26 downto 0);
        begin
	   siw := (others => '0');
	   siw (26) := hit(0);
           siw (pa_reg'length-1 downto 0) := pa_reg;

	   syn_invalidate_word <= siw;
        end process;
      end block bb;
    end generate TrivGen;

end SimpleStruct;

library ieee;
use ieee.std_logic_1164.all;

library AjitCustom;
use AjitCustom.AjitCoreConfigurationPackage.all;
use AjitCustom.AjitGlobalConfigurationPackage.all;
use AjitCustom.AjitCustomComponents.all;

entity accessIcacheRlut_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    lookup : in  std_logic_vector(0 downto 0);
    update : in  std_logic_vector(0 downto 0);
    clear : in  std_logic_vector(0 downto 0);
    physical_addr_of_line : in  std_logic_vector(29 downto 0);
    virtual_addr_of_line : in  std_logic_vector(25 downto 0);
    syn_invalidate_word : out  std_logic_vector(26 downto 0);
    clk, reset: in std_logic
    -- 
  );
end entity;
architecture SimpleStruct of accessIcacheRlut_Operator  is
begin
	baseInst: accessRlutBase_Operator
	  generic map 
		(
			g_LOG_BASE_PAGE_SIZE => LOG_BASE_PAGE_SIZE,
			g_LOG_CACHE_LINE_SIZE => LOG_CACHE_LINE_SIZE,
			g_CACHE_WAY_SIZE => ICACHE_WAY_SIZE,
			g_RLUT_TAG_WIDTH  => ICACHE_RLUT_TAG_WIDTH,
			g_RLUT_REDUCED_DATA_WIDTH => ICACHE_RLUT_REDUCED_DATA_WIDTH,
			g_RLUT_LOG_N_SETS => ICACHE_RLUT_LOG_N_SETS,
			g_RLUT_LOG_MEMORY_SIZE => ICACHE_RLUT_LOG_MEMORY_SIZE,
			g_RLUT_LOG_SET_SIZE => ICACHE_RLUT_LOG_SET_SIZE
		)
	  port map 
		(
			sample_req => sample_req,
			sample_ack => sample_ack,
			update_req => update_req,
			update_ack => update_ack,
			lookup => lookup,
			update => update,
			clear => clear,
			physical_addr_of_line => physical_addr_of_line,
			virtual_addr_of_line => virtual_addr_of_line,
    			syn_invalidate_word => syn_invalidate_word,
    			clk => clk, reset => reset
	        );
end SimpleStruct;

library ieee;
use ieee.std_logic_1164.all;

library AjitCustom;
use AjitCustom.AjitCoreConfigurationPackage.all;
use AjitCustom.AjitGlobalConfigurationPackage.all;
use AjitCustom.AjitCustomComponents.all;

entity accessDcacheRlut_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    lookup : in  std_logic_vector(0 downto 0);
    update : in  std_logic_vector(0 downto 0);
    clear : in  std_logic_vector(0 downto 0);
    physical_addr_of_line : in  std_logic_vector(29 downto 0);
    virtual_addr_of_line : in  std_logic_vector(25 downto 0);
    syn_invalidate_word : out  std_logic_vector(26 downto 0);
    clk, reset: in std_logic
    -- 
  );
end entity;
architecture SimpleStruct of accessDcacheRlut_Operator  is
begin
	baseInst: accessRlutBase_Operator
	  generic map 
		(
			g_LOG_BASE_PAGE_SIZE => LOG_BASE_PAGE_SIZE,
			g_LOG_CACHE_LINE_SIZE => LOG_CACHE_LINE_SIZE,
			g_CACHE_WAY_SIZE => DCACHE_WAY_SIZE,
			g_RLUT_TAG_WIDTH  => DCACHE_RLUT_TAG_WIDTH,
			g_RLUT_REDUCED_DATA_WIDTH => DCACHE_RLUT_REDUCED_DATA_WIDTH,
			g_RLUT_LOG_N_SETS => DCACHE_RLUT_LOG_N_SETS,
			g_RLUT_LOG_MEMORY_SIZE => DCACHE_RLUT_LOG_MEMORY_SIZE,
			g_RLUT_LOG_SET_SIZE => DCACHE_RLUT_LOG_SET_SIZE
		)
	  port map 
		(
			sample_req => sample_req,
			sample_ack => sample_ack,
			update_req => update_req,
			update_ack => update_ack,
			lookup => lookup,
			update => update,
			clear => clear,
			physical_addr_of_line => physical_addr_of_line,
			virtual_addr_of_line => virtual_addr_of_line,
    			syn_invalidate_word => syn_invalidate_word,
    			clk => clk, reset => reset
	        );
end SimpleStruct;

library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;

library AjitCustom;
use AjitCustom.AjitCustomComponents.all;

entity accessL2DataMemGeneric is -- 
  generic (LOG2_NUMBER_OF_LINES : integer := 11; 
		LINE_WIDTH_IN_BYTES: integer := 64);
  port ( -- 
    start_req: in std_logic;
    start_ack: out std_logic;
    fin_req: in std_logic;
    fin_ack: out std_logic;
    -- if true, read data line..
    read_data_line : in  std_logic_vector(0 downto 0);
    -- if true, write data word...
    data_write_dword : in  std_logic_vector(0 downto 0);
    -- if true, read data word (note: read_data_line will also be true in this case)
    data_read_dword : in  std_logic_vector(0 downto 0);
    -- write new line into data mem, (note: insert write dword if data_write_dword is true).
    data_write_new_line : in  std_logic_vector(0 downto 0);
    -- this is now redundant..  write_new_line is always the replaced line.
    do_write_replaced_line_to_mem : in  std_logic_vector(0 downto 0);
    -- byte mask for dword write.
    byte_mask : in  std_logic_vector(7 downto 0);
    -- address of line.
    line_id : in  std_logic_vector(LOG2_NUMBER_OF_LINES-1 downto 0);
    -- offset in line for write dword.
    pa_dword_id : in  std_logic_vector(2 downto 0);
    -- write dword.
    w_dword : in  std_logic_vector(63 downto 0);
    -- line to be written into memory..
    line_to_be_inserted : in  std_logic_vector((8*LINE_WIDTH_IN_BYTES)-1 downto 0);
    -- read data
    read_dword_from_data : out  std_logic_vector(63 downto 0);
    -- line that was read out of memory.. this line will be written eventually to main memory.
    writeback_line_from_data : out  std_logic_vector((8*LINE_WIDTH_IN_BYTES)-1 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity accessL2DataMemGeneric;
architecture accessL2DataMemGenericArch of accessL2DataMemGeneric is -- 

	constant LINE_WIDTH_IN_DWORDS : integer := LINE_WIDTH_IN_BYTES/8;
	constant MAX_DWORD_INDEX : integer := LINE_WIDTH_IN_DWORDS-1;

	type MemDataAggregate is array (natural range <>) of std_logic_vector(63 downto 0);
	signal mem_read_data, mem_write_data, line_from_mem_2D, line_from_mem_2D_reg: 
							MemDataAggregate (0 to LINE_WIDTH_IN_DWORDS-1);
	signal mem_enable, mem_write_bar: std_logic;
    	signal mem_address : std_logic_vector(LOG2_NUMBER_OF_LINES-1 downto 0);

	type ByteMaskAggregate is array (natural range <>) of std_logic_vector(7 downto 0);
	signal mem_byte_mask: ByteMaskAggregate (0 to LINE_WIDTH_IN_DWORDS-1);

	-- note:  These cases can occur.
	-- 
	--       read_data_line write_new_line read_dword write_dword
	--           1               1             1            0
	--        extract read dword out of the new line.
	--
	--           1               1             0            1
	--	  insert new dword into write-line
	--        read   data line.
	--
	--           1                0            x            x
	--        read out line for replacement.
	--
	--           0               0              1           0
	--	  read dword from memory
	--
	--           0               0              0           1
	--	  read dword from memory
	--
	type FsmState is (IDLE_STATE, WRITE_AFTER_READ_STATE);


	signal fsm_state: FsmState;
	signal done_reg: boolean;

	signal is_two_cycle_operation: boolean;
	signal is_read_operation : boolean;
	signal is_write_operation: boolean;

    	signal data_read_dword_reg, data_write_dword_reg: std_logic_vector(0 downto 0);
    	signal data_write_new_line_reg: std_logic_vector(0 downto 0);
    	signal do_write_replaced_line_to_mem_reg: std_logic_vector(0 downto 0);
    	signal line_id_reg: std_logic_vector(LOG2_NUMBER_OF_LINES-1 downto 0);
    	signal pa_dword_id_reg: std_logic_vector(2 downto 0);
    	signal byte_mask_reg:  std_logic_vector(7 downto 0);
    	signal w_dword_reg: std_logic_vector(63 downto 0);
    	signal line_to_be_inserted_reg : std_logic_vector((8*LINE_WIDTH_IN_BYTES)-1 downto 0);
		
	signal dword_index, dword_index_reg : integer range 0 to LINE_WIDTH_IN_DWORDS-1;

	signal fin_ack_sig: std_logic;
	signal latch_outputs: boolean;
    	signal writeback_line_from_data_pre_reg : std_logic_vector((8*64)-1 downto 0);
    	signal writeback_line_from_data_reg : std_logic_vector((8*64)-1 downto 0);
    	signal read_dword_from_data_pre_reg : std_logic_vector(63 downto 0);
    	signal read_dword_from_data_reg : std_logic_vector(63 downto 0);
							
	function calculateInsertDwordValue(ins_dword: std_logic_vector(63 downto 0); 
						byte_mask: std_logic_vector(7 downto 0);
						orig_dword: std_logic_vector(63 downto 0))
		return std_logic_vector is
			variable ret_dword: std_logic_vector(63 downto 0);
	begin
		for I in 7 downto 0 loop
			if(byte_mask(I) = '1') then
				ret_dword(((I+1)*8)-1 downto (I*8)) := 
						ins_dword(((I+1)*8)-1 downto (I*8));
			else
				ret_dword(((I+1)*8)-1 downto (I*8)) := 
						orig_dword(((I+1)*8)-1 downto (I*8));
			end if;
		end loop;
		return(ret_dword);
	end function;
begin --  
	-- note: we do not need to read if a new line is being written into the
	--       cache.  This is because the read data is extracted from the
	--       new line that is being written.
	is_read_operation <= 
		(((data_read_dword(0) = '1') and (data_write_new_line(0) = '0')) or 
								(read_data_line(0) = '1'));
	is_write_operation <= (data_write_dword(0) = '1') or (data_write_new_line(0) = '1');
	is_two_cycle_operation <= is_read_operation and is_write_operation;


	process(clk, reset, start_req, fin_req, fsm_state,done_reg,
			read_data_line, data_read_dword,
			data_write_dword, data_write_new_line,
			is_two_cycle_operation, is_read_operation, is_write_operation,
			line_id, line_id_reg, dword_index, dword_index_reg)
		variable next_fsm_state_var: FsmState;
		variable next_done_reg_var : boolean;
		variable start_ack_var, fin_ack_var: std_logic;
		variable latch_inputs_var: boolean;
		variable mem_enable_var, mem_write_bar_var: std_logic;
    		variable mem_address_var : std_logic_vector(LOG2_NUMBER_OF_LINES-1 downto 0);
		variable mem_byte_mask_var: ByteMaskAggregate (0 to LINE_WIDTH_IN_DWORDS-1);

	begin
		next_fsm_state_var := fsm_state;
		next_done_reg_var  := done_reg;
		start_ack_var := '0';
		fin_ack_var := '0';
		latch_inputs_var := false;
		mem_enable_var := '0';
		mem_write_bar_var := '1';
		mem_address_var := (others => '0');
		mem_byte_mask_var := (others => (others => '0'));

		case fsm_state is 
			when IDLE_STATE =>
				if(done_reg) then
					fin_ack_var := '1';
					if(fin_req = '1') then 
						next_done_reg_var := false;
					end if;
				end if;
				if(not next_done_reg_var) then
					start_ack_var := '1';
					if(start_req = '1') then

						latch_inputs_var := true;
						mem_address_var := line_id;

						-- first read then write for two cycle operation.
						if(is_two_cycle_operation or is_read_operation) then
							mem_enable_var := '1';
							mem_byte_mask_var := (others => (others => '1'));
						elsif (is_write_operation) then
							mem_enable_var := '1';
							mem_write_bar_var := '0';

							-- note: mem write data will be assembled
							--       in a separate process to avoid 
							--       clutter here.
							if(data_write_new_line(0) = '1')  then
								mem_byte_mask_var := (others => (others => '1'));
							else
								mem_byte_mask_var(dword_index) := byte_mask;
							end if;
						end if;

						if(is_two_cycle_operation) then
							next_fsm_state_var := WRITE_AFTER_READ_STATE;
						else 
							next_done_reg_var := true;
						end if;
					end if;
				end if; 
			when WRITE_AFTER_READ_STATE =>
				-- it has to be a write operation.
				--   either a write_line (with write_dword)
				--   or a plain write_dword.
				mem_enable_var := '1';
				mem_write_bar_var := '0';
				mem_address_var := line_id_reg;

				if(data_write_new_line_reg(0) = '1')  then
					mem_byte_mask_var := (others => (others => '1'));
				else
					mem_byte_mask_var(dword_index_reg) := byte_mask_reg;
				end if;

				next_done_reg_var := true;
				next_fsm_state_var := IDLE_STATE;
		end case;

		start_ack <= start_ack_var;
		fin_ack_sig   <= fin_ack_var;

		mem_enable <= mem_enable_var;
		mem_write_bar <= mem_write_bar_var;
		mem_address <= mem_address_var;
		mem_byte_mask <= mem_byte_mask_var;

		if(clk'event and (clk = '1')) then
			if(reset = '1') then
				fsm_state <= IDLE_STATE;
				done_reg <= false;
			else
				fsm_state <= next_fsm_state_var;
				done_reg <= next_done_reg_var;
    				if(latch_inputs_var) then
    					data_read_dword_reg  <= data_read_dword;
    					data_write_dword_reg  <= data_write_dword;
    					data_write_new_line_reg <= data_write_new_line;
    					do_write_replaced_line_to_mem_reg <= do_write_replaced_line_to_mem;
    					line_id_reg <= line_id;
    					pa_dword_id_reg <= pa_dword_id;
    					byte_mask_reg <= byte_mask;
    					w_dword_reg <= w_dword;
    					line_to_be_inserted_reg <= line_to_be_inserted;
				end if;
			end if;
		end if;
	end process;	
	fin_ack <= fin_ack_sig;

		
	dword_index <= to_integer(unsigned(pa_dword_id));
	dword_index_reg <= to_integer(unsigned(pa_dword_id_reg));

	genDwords: for D in 0 to LINE_WIDTH_IN_DWORDS-1 generate
	  bblk: block
		signal use_w_dword: boolean;
		signal use_w_dword_reg: boolean;

          begin
		-- reorganize the line being written into the memory..
		line_from_mem_2D_reg(D) <= 
			line_to_be_inserted_reg((((MAX_DWORD_INDEX-D)+1)*64)-1 downto ((MAX_DWORD_INDEX-D)*64));
					
		use_w_dword_reg <=  ((data_write_dword_reg(0) = '1') and (dword_index_reg = D));
		use_w_dword     <=  ((data_write_dword(0) = '1') and (dword_index = D));

		bb: generic_single_port_memory_with_byte_mask
			generic map (name => "accessL2Data:bb:" & Convert_To_String(D),
						g_addr_width => line_id'length, g_data_width => 64)
			port map (
					clk => clk, reset => reset,
					enable => mem_enable,
					writebar => mem_write_bar,
					bytemask => mem_byte_mask(D),
					datain => mem_write_data (D),
					dataout => mem_read_data (D),
					addrin  => mem_address
				);

		process(w_dword, w_dword_reg,  use_w_dword, use_w_dword_reg,
					 data_write_new_line, data_write_new_line_reg,
					 line_to_be_inserted, line_to_be_inserted_reg)
			variable inserted_dword_var: std_logic_vector(63 downto 0);
			variable line_dword_var: std_logic_vector(63 downto 0);
		begin
			inserted_dword_var := (others => '0');
			if(fsm_state = WRITE_AFTER_READ_STATE) then
				line_dword_var :=
					line_to_be_inserted_reg((((MAX_DWORD_INDEX-D)+1)*64)-1 downto 
									((MAX_DWORD_INDEX-D)*64));
				if(use_w_dword_reg) then 
					if(data_write_new_line_reg(0) = '1') then 
						-- insert dword into line dword and then
						-- write the full line!
						inserted_dword_var :=  
							calculateInsertDwordValue(w_dword_reg, 
											byte_mask_reg,
											line_dword_var);
					else
						inserted_dword_var :=  w_dword_reg;
					end if;
				elsif (data_write_new_line_reg(0) = '1') then 
					inserted_dword_var :=  line_dword_var;
				end if;
				mem_write_data(D) <= inserted_dword_var;
			else
				line_dword_var :=
					line_to_be_inserted((((MAX_DWORD_INDEX-D)+1)*64)-1 downto 
									((MAX_DWORD_INDEX-D)*64));
				if(use_w_dword) then 
					if(data_write_new_line(0) = '1') then 
						-- insert dword into line dword and then
						-- write the full line!
						inserted_dword_var :=  
							calculateInsertDwordValue(w_dword, 
											byte_mask,
											line_dword_var);
					else
						inserted_dword_var :=  w_dword;
					end if;
				elsif (data_write_new_line(0) = '1') then 
					inserted_dword_var :=  line_dword_var;
				end if;
			end if;
			mem_write_data(D) <= inserted_dword_var;
		end process;


		-- write back line is returned to the outside world.
		 writeback_line_from_data_pre_reg ((((MAX_DWORD_INDEX-D)+1)*64)-1 downto 
							((MAX_DWORD_INDEX-D)*64)) <= mem_read_data(D);
	  end block bblk;	
	end generate genDwords;

	-- here you have to be careful.. 
	-- read dword can come mem_read_data or from the replacing line.
    	read_dword_from_data_pre_reg <= 
		line_from_mem_2D_reg(dword_index_reg) when
			((data_write_new_line_reg(0) = '1') and (data_read_dword_reg(0) = '1')) 
				else mem_read_data(dword_index_reg);

	-- output stage: note the output goes to an UnloadBuffer which handles the
	--               update req/ack exchange with no races.
	writeback_line_from_data <= writeback_line_from_data_pre_reg;
	read_dword_from_data <= read_dword_from_data_pre_reg;

end accessL2DataMemGenericArch;
--------------------------------------------------------------------------------------------
--------------------------------------------------------------------------------------------
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;

library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
entity accessL2DataMemGeneric_Operator is -- 
  generic (     name: string;
		LOG2_NUMBER_OF_LINES: integer := 10;
		LINE_WIDTH_IN_BYTES: integer := 64
	);
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    -- if true, read data line..
    read_data_line : in  std_logic_vector(0 downto 0);
    -- if true, write data word...
    data_write_dword : in  std_logic_vector(0 downto 0);
    -- if true, read data word (note: read_data_line will also be true in this case)
    data_read_dword : in  std_logic_vector(0 downto 0);
    -- write new line into data mem, (note: insert write dword if data_write_dword is true).
    data_write_new_line : in  std_logic_vector(0 downto 0);
    -- this is now redundant..  write_new_line is always the replaced line.
    do_write_replaced_line_to_mem : in  std_logic_vector(0 downto 0);
    -- byte mask for dword write.
    byte_mask : in  std_logic_vector(7 downto 0);
    -- address of line.
    line_id : in  std_logic_vector(LOG2_NUMBER_OF_LINES-1 downto 0);
    -- offset in line for write dword.
    pa_dword_id : in  std_logic_vector(2 downto 0);
    -- write dword.
    w_dword : in  std_logic_vector(63 downto 0);
    -- line to be written into memory..
    line_to_be_inserted : in  std_logic_vector((8*LINE_WIDTH_IN_BYTES)-1 downto 0);
    -- read data
    read_dword_from_data : out  std_logic_vector(63 downto 0);
    -- line that was read out of memory.. this line will be written eventually to main memory.
    writeback_line_from_data : out  std_logic_vector((8*LINE_WIDTH_IN_BYTES)-1 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity accessL2DataMemGeneric_Operator;

architecture Trivial of accessL2DataMemGeneric_Operator is
	signal start_req, start_ack: std_logic;
	signal push_ack, push_req, pop_req, pop_ack: std_logic;
	signal push_data, pop_data: 
		std_logic_vector(writeback_line_from_data'length + read_dword_from_data'length -1
					downto 0);
			
    	signal read_dword_from_data_base : std_logic_vector(63 downto 0);
    	signal writeback_line_from_data_base : std_logic_vector((8*LINE_WIDTH_IN_BYTES)-1 downto 0);
	signal has_data: std_logic;

begin
	push_data <=  writeback_line_from_data_base & read_dword_from_data_base;

	writeback_line_from_data <= pop_data (pop_data'length-1 downto read_dword_from_data'length);
	read_dword_from_data <= pop_data (read_dword_from_data'length-1 downto 0);
	

	p2lInst:
		Sample_Pulse_To_Level_Translate_Entity
			generic map ("accessL2DataMem_P2L")
			port map 
				( rL => sample_req,
					rR => start_req,
					aL => sample_ack,
					aR => start_ack,
					clk => clk, reset => reset);	


	baseInst: accessL2DataMemGeneric
  		generic map(LOG2_NUMBER_OF_LINES => LOG2_NUMBER_OF_LINES, 
						LINE_WIDTH_IN_BYTES => LINE_WIDTH_IN_BYTES)
  		port map ( -- 
    				start_req => start_req,
    				start_ack => start_ack,
				-- This will push into the output queue.
    				fin_req => push_ack,
    				fin_ack => push_req,
    				read_data_line  => read_data_line ,
    				data_write_dword  => data_write_dword ,
    				data_read_dword  => data_read_dword ,
    				data_write_new_line  => data_write_new_line ,
    				do_write_replaced_line_to_mem  => do_write_replaced_line_to_mem ,
    				byte_mask  => byte_mask ,
    				line_id  => line_id ,
    				pa_dword_id  => pa_dword_id ,
    				w_dword  => w_dword ,
    				line_to_be_inserted  => line_to_be_inserted ,
    				read_dword_from_data  => read_dword_from_data_base ,
    				writeback_line_from_data  => writeback_line_from_data_base ,
    				clk => clk, reset => reset
  				);

	-- Unload buffer... for a coherent update req/ack connection.
	ub: UnloadBuffer
		generic map (name => "accessL2DataMem:ub",
				buffer_size => 2, 
				data_width => push_data'length,
				bypass_flag => true, 
				nonblocking_reaD_flag => false,
				use_unload_register => true)
		port map (clk => clk, reset => reset,
				write_req => push_req,
				write_ack => push_ack,
				write_data => push_data,
				unload_req  => update_req,
				unload_ack  => update_ack,
				read_data => pop_data,
				has_data => has_data);

end Trivial;
-------------------------------------------------------------------------------------------------------
-------------------------------------------------------------------------------------------------------
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;

library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
entity accessL2DataMemX1024X512_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    -- if true, read data line..
    read_data_line : in  std_logic_vector(0 downto 0);
    -- if true, write data word...
    data_write_dword : in  std_logic_vector(0 downto 0);
    -- if true, read data word (note: read_data_line will also be true in this case)
    data_read_dword : in  std_logic_vector(0 downto 0);
    -- write new line into data mem, (note: insert write dword if data_write_dword is true).
    data_write_new_line : in  std_logic_vector(0 downto 0);
    -- this is now redundant..  write_new_line is always the replaced line.
    do_write_replaced_line_to_mem : in  std_logic_vector(0 downto 0);
    -- byte mask for dword write.
    byte_mask : in  std_logic_vector(7 downto 0);
    -- address of line.
    line_id : in  std_logic_vector(9 downto 0);
    -- offset in line for write dword.
    pa_dword_id : in  std_logic_vector(2 downto 0);
    -- write dword.
    w_dword : in  std_logic_vector(63 downto 0);
    -- line to be written into memory..
    line_to_be_inserted : in  std_logic_vector((8*64)-1 downto 0);
    -- read data
    read_dword_from_data : out  std_logic_vector(63 downto 0);
    -- line that was read out of memory.. this line will be written eventually to main memory.
    writeback_line_from_data : out  std_logic_vector((8*64)-1 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity accessL2DataMemX1024X512_Operator;

architecture Trivial of accessL2DataMemX1024X512_Operator is

begin
	baseInst: accessL2DataMemGeneric_Operator
  		generic map(name => "accessL2DataMemX1024X512",
  				LOG2_NUMBER_OF_LINES => 10, LINE_WIDTH_IN_BYTES => 64)
  		port map ( -- 
    				sample_req => sample_req,
    				sample_ack => sample_ack,
    				update_req => update_req,
    				update_ack => update_ack,
    				read_data_line  => read_data_line ,
    				data_write_dword  => data_write_dword ,
    				data_read_dword  => data_read_dword ,
    				data_write_new_line  => data_write_new_line ,
    				do_write_replaced_line_to_mem  => do_write_replaced_line_to_mem ,
    				byte_mask  => byte_mask ,
    				line_id  => line_id ,
    				pa_dword_id  => pa_dword_id ,
    				w_dword  => w_dword ,
    				line_to_be_inserted  => line_to_be_inserted ,
    				read_dword_from_data  => read_dword_from_data ,
    				writeback_line_from_data  => writeback_line_from_data,
    				clk => clk, reset => reset
  				);

end Trivial;
-------------------------------------------------------------------------------------------------------
-------------------------------------------------------------------------------------------------------
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;

library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
entity accessL2DataMemX2048X512_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    -- if true, read data line..
    read_data_line : in  std_logic_vector(0 downto 0);
    -- if true, write data word...
    data_write_dword : in  std_logic_vector(0 downto 0);
    -- if true, read data word (note: read_data_line will also be true in this case)
    data_read_dword : in  std_logic_vector(0 downto 0);
    -- write new line into data mem, (note: insert write dword if data_write_dword is true).
    data_write_new_line : in  std_logic_vector(0 downto 0);
    -- this is now redundant..  write_new_line is always the replaced line.
    do_write_replaced_line_to_mem : in  std_logic_vector(0 downto 0);
    -- byte mask for dword write.
    byte_mask : in  std_logic_vector(7 downto 0);
    -- address of line.
    line_id : in  std_logic_vector(10 downto 0);
    -- offset in line for write dword.
    pa_dword_id : in  std_logic_vector(2 downto 0);
    -- write dword.
    w_dword : in  std_logic_vector(63 downto 0);
    -- line to be written into memory..
    line_to_be_inserted : in  std_logic_vector((8*64)-1 downto 0);
    -- read data
    read_dword_from_data : out  std_logic_vector(63 downto 0);
    -- line that was read out of memory.. this line will be written eventually to main memory.
    writeback_line_from_data : out  std_logic_vector((8*64)-1 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity accessL2DataMemX2048X512_Operator;

architecture Trivial of accessL2DataMemX2048X512_Operator is
begin
	baseInst: accessL2DataMemGeneric_Operator
  		generic map(name => "accessL2DataMemX2048X512",
				LOG2_NUMBER_OF_LINES => 11, LINE_WIDTH_IN_BYTES => 64)
  		port map ( -- 
    				sample_req => sample_req,
    				sample_ack => sample_ack,
    				update_req => update_req,
    				update_ack => update_ack,
    				read_data_line  => read_data_line ,
    				data_write_dword  => data_write_dword ,
    				data_read_dword  => data_read_dword ,
    				data_write_new_line  => data_write_new_line ,
    				do_write_replaced_line_to_mem  => do_write_replaced_line_to_mem ,
    				byte_mask  => byte_mask ,
    				line_id  => line_id ,
    				pa_dword_id  => pa_dword_id ,
    				w_dword  => w_dword ,
    				line_to_be_inserted  => line_to_be_inserted ,
    				read_dword_from_data  => read_dword_from_data,
    				writeback_line_from_data  => writeback_line_from_data,
    				clk => clk, reset => reset
  				);
end Trivial;
-------------------------------------------------------------------------------------------------------
-------------------------------------------------------------------------------------------------------
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;

library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
entity accessL2DataMemX4096X512_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    -- if true, read data line..
    read_data_line : in  std_logic_vector(0 downto 0);
    -- if true, write data word...
    data_write_dword : in  std_logic_vector(0 downto 0);
    -- if true, read data word (note: read_data_line will also be true in this case)
    data_read_dword : in  std_logic_vector(0 downto 0);
    -- write new line into data mem, (note: insert write dword if data_write_dword is true).
    data_write_new_line : in  std_logic_vector(0 downto 0);
    -- this is now redundant..  write_new_line is always the replaced line.
    do_write_replaced_line_to_mem : in  std_logic_vector(0 downto 0);
    -- byte mask for dword write.
    byte_mask : in  std_logic_vector(7 downto 0);
    -- address of line.
    line_id : in  std_logic_vector(11 downto 0);
    -- offset in line for write dword.
    pa_dword_id : in  std_logic_vector(2 downto 0);
    -- write dword.
    w_dword : in  std_logic_vector(63 downto 0);
    -- line to be written into memory..
    line_to_be_inserted : in  std_logic_vector((8*64)-1 downto 0);
    -- read data
    read_dword_from_data : out  std_logic_vector(63 downto 0);
    -- line that was read out of memory.. this line will be written eventually to main memory.
    writeback_line_from_data : out  std_logic_vector((8*64)-1 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity accessL2DataMemX4096X512_Operator;

architecture Trivial of accessL2DataMemX4096X512_Operator is
begin
	baseInst: accessL2DataMemGeneric_Operator
  		generic map(name => "accessL2DataMemX4096X512",
					LOG2_NUMBER_OF_LINES => 12, LINE_WIDTH_IN_BYTES => 64)
  		port map ( -- 
    				sample_req => sample_req,
    				sample_ack => sample_ack,
    				update_req => update_req,
    				update_ack => update_ack,
    				read_data_line  => read_data_line ,
    				data_write_dword  => data_write_dword ,
    				data_read_dword  => data_read_dword ,
    				data_write_new_line  => data_write_new_line ,
    				do_write_replaced_line_to_mem  => do_write_replaced_line_to_mem ,
    				byte_mask  => byte_mask ,
    				line_id  => line_id ,
    				pa_dword_id  => pa_dword_id ,
    				w_dword  => w_dword ,
    				line_to_be_inserted  => line_to_be_inserted ,
    				read_dword_from_data  => read_dword_from_data,
    				writeback_line_from_data  => writeback_line_from_data,
    				clk => clk, reset => reset
  				);
end Trivial;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.basecomponents.all;
use ahir.mem_component_pack.all;
use ahir.utilities.all;

library AjitCustom;
use AjitCustom.AjitGlobalConfigurationPackage.all;
use AjitCustom.AjitCustomComponents.all;

-- generic Tag memory model with configurable
--   number of lines, associativity, dwords-per-line and physical address width.
entity accessL2TagMemGeneric is -- 
  generic (
		LOG2_NUMBER_OF_LINES: integer := 12;
		LOG2_ASSOCIATIVITY: integer := 3;
		LOG2_DWORDS_PER_LINE: integer := 3;
		PA_ADDRESS_WIDTH: integer := 36
	  );
  port ( -- 
    start_req: in std_logic;
    start_ack: out std_logic;
    fin_req: in std_logic;
    fin_ack: out std_logic;
    init_flag : in  std_logic_vector(0 downto 0);
    tag_mem_read : in  std_logic_vector(0 downto 0);
    tag_mem_write : in  std_logic_vector(0 downto 0);
    read_set_id : in  std_logic_vector((LOG2_NUMBER_OF_LINES-LOG2_ASSOCIATIVITY)-1 downto 0);
    write_set_id : in  std_logic_vector((LOG2_NUMBER_OF_LINES-LOG2_ASSOCIATIVITY)-1 downto 0);
    tags_have_been_modified : in  std_logic_vector(0 downto 0);
    lwi_has_been_modified : in  std_logic_vector(0 downto 0);
    valids_have_been_modified : in  std_logic_vector(0 downto 0);
    dirty_bits_have_been_modified : in  std_logic_vector(0 downto 0);
    updated_set_tags : in  
	std_logic_vector(((2**LOG2_ASSOCIATIVITY)*(30-(LOG2_NUMBER_OF_LINES-LOG2_ASSOCIATIVITY)))-1 downto 0);
    updated_set_lwi : in  
	std_logic_vector(LOG2_ASSOCIATIVITY-1 downto 0);
    updated_set_valids : in  
	std_logic_vector((2**LOG2_ASSOCIATIVITY)-1 downto 0);
    updated_set_dirty_dword_masks : in  
	std_logic_vector(((2**LOG2_DWORDS_PER_LINE)*(2**LOG2_ASSOCIATIVITY))-1 downto 0);
    tag_mem_response : out  
	std_logic_vector(((2**LOG2_ASSOCIATIVITY)*(30-(LOG2_NUMBER_OF_LINES-LOG2_ASSOCIATIVITY))) +
			LOG2_ASSOCIATIVITY + (2**LOG2_ASSOCIATIVITY) + 
			((2**LOG2_DWORDS_PER_LINE)*(2**LOG2_ASSOCIATIVITY))-1  downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity accessL2TagMemGeneric;
architecture accessL2TagMemGeneric_arch of accessL2TagMemGeneric is -- 

	constant LOG2_NUMBER_OF_SETS : integer := (LOG2_NUMBER_OF_LINES - LOG2_ASSOCIATIVITY);
	constant NUMBER_OF_SETS: integer := (2**LOG2_NUMBER_OF_SETS);
	constant ASSOCIATIVITY : integer := (2**LOG2_ASSOCIATIVITY);
	constant DWORDS_PER_LINE: integer := (2**LOG2_DWORDS_PER_LINE);

	constant PA_LINE_ADDRESS_WIDTH: integer := (PA_ADDRESS_WIDTH - (LOG2_DWORDS_PER_LINE  + 3));
	constant PA_TAG_WIDTH : integer := (PA_LINE_ADDRESS_WIDTH - LOG2_NUMBER_OF_SETS);

	-- We will have two memories:
	--    a single ported memory for the pa_tags
	--    a dual ported memory for the dirty-bits, the last-written-indices and for the valids..
	--
	constant spmem_data_width : integer := PA_TAG_WIDTH*ASSOCIATIVITY;

	signal spmem_write_data: std_logic_vector(spmem_data_width-1 downto 0);
	signal spmem_read_data : std_logic_vector(spmem_data_width-1 downto 0);
	signal spmem_enable, spmem_write_bar: std_logic;
	signal spmem_address : std_logic_vector(LOG2_NUMBER_OF_SETS-1 downto 0);

	-- dirty-bits, last-written index for the set, and also the valids..
	constant dpmem_data_width : integer := 
		(DWORDS_PER_LINE*ASSOCIATIVITY) + LOG2_ASSOCIATIVITY + ASSOCIATIVITY;
	signal dpmem_write_data: std_logic_vector(dpmem_data_width-1 downto 0);
	signal dpmem_read_data: std_logic_vector(dpmem_data_width-1 downto 0);

	-- read will be from one port, write from the other.
	signal dpmem_read_enable, dpmem_write_enable: std_logic;
	signal dpmem_read_address : std_logic_vector(LOG2_NUMBER_OF_SETS-1 downto 0);
	signal dpmem_write_address : std_logic_vector(LOG2_NUMBER_OF_SETS-1 downto 0);

	signal is_two_cycle_operation, is_two_cycle_operation_reg: boolean;

	type FsmState is (INIT_STATE, IDLE_STATE, READ_AFTER_WRITE_STATE);
	signal fsm_state: FsmState;

	signal init_counter: unsigned (LOG2_NUMBER_OF_SETS-1 downto 0);

	signal latch_inputs: boolean;
    
	signal tag_mem_read_reg : std_logic_vector(0 downto 0);
    	signal tag_mem_write_reg : std_logic_vector(0 downto 0);
    	signal read_set_id_reg : std_logic_vector(LOG2_NUMBER_OF_SETS-1 downto 0);
    	signal write_set_id_reg : std_logic_vector(LOG2_NUMBER_OF_SETS-1  downto 0);

    	signal tags_have_been_modified_reg : std_logic_vector(0 downto 0);
    	signal lwi_has_been_modified_reg : std_logic_vector(0 downto 0);
    	signal valids_have_been_modified_reg : std_logic_vector(0 downto 0);
    	signal dirty_bits_have_been_modified_reg : std_logic_vector(0 downto 0);

    	signal tags_from_spmem, updated_set_tags_reg : std_logic_vector((PA_TAG_WIDTH*ASSOCIATIVITY)-1 downto 0);

    	signal lwi_from_dpmem, updated_set_lwi_reg : std_logic_vector(LOG2_ASSOCIATIVITY-1 downto 0);

    	signal valids_from_dpmem, updated_set_valids_reg : std_logic_vector(ASSOCIATIVITY-1 downto 0);

    	signal dirty_bits_from_dpmem, updated_set_dirty_dword_masks_reg : 
	     std_logic_vector((DWORDS_PER_LINE*ASSOCIATIVITY)-1 downto 0);

	signal tag_mem_response_pre_reg, tag_mem_response_reg: 
		std_logic_vector(tag_mem_response'length -1 downto 0);

	signal done_reg, is_nop: boolean;
	signal fin_ack_sig: std_logic;
	signal latch_outputs: boolean;
		

begin --  


	-- read and write are both specified on a single port memory..
	is_two_cycle_operation <= ((tag_mem_read(0) = '1') and 
					(tag_mem_write(0) = '1') and
					(tags_have_been_modified(0) = '1'));
	is_nop <= (tag_mem_read(0) = '0') and (tag_mem_write(0) = '0');

	process(clk, reset, latch_inputs)
	begin
		if(clk'event and (clk = '1')) then
			if(reset = '1') then
				is_two_cycle_operation_reg <= false;
			elsif (latch_inputs) then
				is_two_cycle_operation_reg <= is_two_cycle_operation;
				tag_mem_read_reg <= tag_mem_read;
    				tag_mem_write_reg <= tag_mem_write;
    				read_set_id_reg <= read_set_id;
    				tags_have_been_modified_reg <= tags_have_been_modified;
    				lwi_has_been_modified_reg <= lwi_has_been_modified;
    				valids_have_been_modified_reg <= valids_have_been_modified;
    				dirty_bits_have_been_modified_reg <= dirty_bits_have_been_modified;
    				write_set_id_reg <= write_set_id;
    				updated_set_tags_reg <= updated_set_tags;
    				updated_set_lwi_reg <= updated_set_lwi;
    				updated_set_valids_reg <= updated_set_valids;
    				updated_set_dirty_dword_masks_reg <= updated_set_dirty_dword_masks;
			end if;
		end if;
	end process;

	process(clk, reset, fsm_state, start_req, fin_req,
    			init_flag,
    			tag_mem_read,
    			tag_mem_write,
    			read_set_id,
    			write_set_id,
    			tags_have_been_modified,
    			lwi_has_been_modified,
    			valids_have_been_modified,
    			dirty_bits_have_been_modified,
			init_counter,
			is_two_cycle_operation,
			is_nop,
			is_two_cycle_operation_reg,
			tag_mem_read_reg,
    			tag_mem_write_reg,
    			read_set_id_reg,
    			write_set_id_reg,
    			updated_set_tags_reg,
    			updated_set_lwi_reg,
    			updated_set_valids_reg,
    			updated_set_dirty_dword_masks_reg
		)

		variable next_fsm_state_var: FsmState;

		variable spmem_address_var : std_logic_vector(LOG2_NUMBER_OF_SETS-1 downto 0);
		variable spmem_enable_var, spmem_write_bar_var: std_logic;
		variable spmem_write_data_var: std_logic_vector(spmem_data_width-1 downto 0);

		variable dpmem_read_address_var : std_logic_vector(LOG2_NUMBER_OF_SETS-1 downto 0);
		variable dpmem_write_address_var : std_logic_vector(LOG2_NUMBER_OF_SETS-1 downto 0);
		variable dpmem_read_enable_var, dpmem_write_enable_var: std_logic;
		variable dpmem_write_data_var: std_logic_vector(dpmem_data_width-1 downto 0);

		variable next_init_counter_var: unsigned (LOG2_NUMBER_OF_SETS-1 downto 0);

		variable start_ack_var, fin_ack_var: std_logic;
		variable latch_inputs_var : boolean;
		variable next_done_reg_var : boolean;
	begin
		next_fsm_state_var := fsm_state;

		spmem_address_var := (others => '0');
		spmem_write_data_var := (others => '0');
		spmem_enable_var := '0';
		spmem_write_bar_var := '1';

		dpmem_read_address_var := (others => '0');
		dpmem_write_address_var := (others => '0');
		dpmem_write_data_var := (others => '0');
		dpmem_read_enable_var := '0';
		dpmem_write_enable_var := '0';

		next_init_counter_var := init_counter;
		start_ack_var := '0';
		fin_ack_var := '0';

		latch_inputs_var := false;
		next_done_reg_var := done_reg;

		case fsm_state is 
			when INIT_STATE =>
				dpmem_write_enable_var := '1';
				dpmem_write_address_var := std_logic_vector(init_counter);

				spmem_enable_var := '1';
				spmem_write_bar_var := '0';
				spmem_address_var := std_logic_vector(init_counter);

				if(init_counter = (NUMBER_OF_SETS - 1)) then
					next_fsm_state_var := IDLE_STATE;
					next_init_counter_var := (others => '0');
				else
					next_init_counter_var := init_counter + 1;
				end if;
			when IDLE_STATE =>
				if(done_reg) then 
					fin_ack_var := '1';
					if(fin_req = '1') then
						next_done_reg_var := false;
					end if;
				end if; -- done_reg
				if (not next_done_reg_var)  then 
				   start_ack_var := '1';
				   if(start_req = '1') then
			            if(is_nop) then
					next_done_reg_var := true;
				    else
			
					latch_inputs_var := true;

					if(is_two_cycle_operation) then
						-- do the write on the single port mem.
						--
						spmem_enable_var := '1';
						spmem_write_bar_var := '0';
						spmem_write_data_var := updated_set_tags;
						spmem_address_var := write_set_id;

						next_fsm_state_var := READ_AFTER_WRITE_STATE;
						next_done_reg_var  := false;
					else
						next_done_reg_var  := true;
						spmem_enable_var := '1';
						if(tag_mem_read(0)  = '1') then
							spmem_address_var := read_set_id;
						elsif (tag_mem_write(0) = '1') then
							spmem_address_var := write_set_id;
							spmem_write_data_var := updated_set_tags;
							spmem_write_bar_var := '0';
						end if;
					end if; -- two cycle operation check...
				
					--
					-- dual port write/read always occurs..
					--
					dpmem_read_enable_var := '1';
					dpmem_read_address_var := read_set_id;
					if ((tag_mem_write(0) = '1') and
						((lwi_has_been_modified(0) = '1') or
							(dirty_bits_have_been_modified(0) = '1') or
							(valids_have_been_modified(0) = '1'))) then
						--
						-- Note: The DPMEM includes a write->read
						--       bypass path!!!
						dpmem_write_enable_var := '1';
						dpmem_write_address_var := write_set_id;
						dpmem_write_data_var := 
							(updated_set_dirty_dword_masks & 
									updated_set_lwi & updated_set_valids);
					end if; -- write
                                    end if; -- not nop
                                  end if; -- start_req
				end if; -- fin ack completed...
			when READ_AFTER_WRITE_STATE =>
				-- just do the read...
				spmem_enable_var   := '1';
				spmem_address_var  := read_set_id_reg;
				next_fsm_state_var := IDLE_STATE;	
				next_done_reg_var  := true;
		end case;

		start_ack <= start_ack_var;
		fin_ack_sig <= fin_ack_var;

		dpmem_read_enable  <= dpmem_read_enable_var;
		dpmem_write_enable <= dpmem_write_enable_var;
		dpmem_read_address <= dpmem_read_address_var;
		dpmem_write_address <= dpmem_write_address_var;
		dpmem_write_data <= dpmem_write_data_var;

		spmem_enable <= spmem_enable_var;
		spmem_write_bar <= spmem_write_bar_var;
		spmem_address <= spmem_address_var;
		spmem_write_data <= spmem_write_data_var;

		latch_inputs <= latch_inputs_var;	

		if (clk'event and (clk = '1')) then
			if(reset = '1') then
				fsm_state <= INIT_STATE;
				init_counter <= (others => '0');
				done_reg <= false;
			else
				fsm_state <= next_fsm_state_var;
				init_counter <= next_init_counter_var;
				done_reg <= next_done_reg_var;
			end if;
		end if;
	end process;

	fin_ack <= fin_ack_sig;
	latch_outputs <= (fin_req = '1') and done_reg;
		
	-- instantiate the spmem and dpmem..
	spmem_inst: 
		base_bank 
			generic map (name => "accessL2TagMemGeneric:SPMEM",
					g_addr_width => LOG2_NUMBER_OF_SETS,
					g_data_width => SPMEM_DATA_WIDTH)
			port map
				(datain => spmem_write_data,
					dataout => spmem_read_data,
					addrin => spmem_address,
					enable => spmem_enable,
					writebar => spmem_write_bar,
					clk => clk, reset => reset);

	dpmem_inst:
		register_file_1w_1r_port_with_bypass 
			generic map (name => "accessL2TagMemGeneric:DPMEM",
					g_addr_width => LOG2_NUMBER_OF_SETS,
					g_data_width => dpmem_data_width)
			port map
				(
					datain_0 => dpmem_write_data,
					addrin_0 => dpmem_write_address,
					enable_0 => dpmem_write_enable,
					dataout_1 => dpmem_read_data,
					addrin_1 => dpmem_read_address,
					enable_1 => dpmem_read_enable,
					clk => clk, reset => reset);

	tags_from_spmem <= spmem_read_data (spmem_read_data'length -1 downto 0);
	dirty_bits_from_dpmem <= 
		dpmem_read_data (dpmem_read_data'length-1 downto 
					(updated_set_lwi'length + updated_set_valids'length));
	lwi_from_dpmem <= 
		dpmem_read_data ((updated_set_lwi'length + updated_set_valids'length)-1 downto 
						updated_set_valids'length);
	valids_from_dpmem <= 
		dpmem_read_data(updated_set_valids'length-1 downto 0);
	
	
	tag_mem_response_pre_reg <= tags_from_spmem & lwi_from_dpmem & valids_from_dpmem & dirty_bits_from_dpmem;

	process(clk, reset)
	begin
		if(clk'event and (clk = '1')) then
			if(reset = '1') then 
				tag_mem_response_reg <= (others => '0');
			elsif(latch_outputs) then
				tag_mem_response_reg <= tag_mem_response_pre_reg;
			end if;
		end if;
	end process;
	tag_mem_response <= tag_mem_response_pre_reg when latch_outputs else tag_mem_response_reg;
end accessL2TagMemGeneric_arch;

library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.mem_component_pack.all;
use ahir.basecomponents.all;

library AjitCustom;
use AjitCustom.AjitGlobalConfigurationPackage.all;
use AjitCustom.AjitCustomComponents.all;
--
-- X1024X8 means  that this manages 1024 lines
-- and set associativity is 8.  Thus a total cache size of 
-- 64KB organized into 128 sets.
-- 
-- Thus, the PA tag width is 30-(log2 (1024/8)) = 30-7=23
--   
entity accessL2TagMemX1024X8_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    init_flag : in  std_logic_vector(0 downto 0);
    tag_mem_read : in  std_logic_vector(0 downto 0);
    tag_mem_write : in  std_logic_vector(0 downto 0);
    read_set_id : in  std_logic_vector(6 downto 0);
    write_set_id : in  std_logic_vector(6 downto 0);
    tags_have_been_modified : in  std_logic_vector(0 downto 0);
    lwi_has_been_modified : in  std_logic_vector(0 downto 0);
    valids_have_been_modified : in  std_logic_vector(0 downto 0);
    dirty_bits_have_been_modified : in  std_logic_vector(0 downto 0);
    updated_set_tags : in  std_logic_vector(183 downto 0);
    updated_set_lwi : in  std_logic_vector(2 downto 0);
    updated_set_valids : in  std_logic_vector(7 downto 0);
    updated_set_dirty_dword_masks : in  std_logic_vector(63 downto 0);
    tag_mem_response : out  std_logic_vector(258 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity accessL2TagMemX1024X8_Operator;
architecture accessL2TagMemX1024X8_Operator_arch of accessL2TagMemX1024X8_Operator is -- 
	signal start_req, start_ack, fin_req, fin_ack: std_logic;
begin --  
	p2lInst:
		Sample_Pulse_To_Level_Translate_Entity
			generic map ("accessL2TagMem_P2L")
			port map 
				( rL => sample_req,
					rR => start_req,
					aL => sample_ack,
					aR => start_ack,
					clk => clk, reset => reset);	
	l2pInst: 
		Level_To_Pulse_Translate_Entity
			generic map ("accessL2TagMem_L2P")
			port map (rL => fin_req,
					rR => update_req,
					aL => fin_ack,
					aR => update_ack,
					clk => clk, reset => reset);

	baseInst:
		accessL2TagMemGeneric
			generic map (LOG2_NUMBER_OF_LINES => 10,
						LOG2_ASSOCIATIVITY => 3,
						LOG2_DWORDS_PER_LINE => 3,
						PA_ADDRESS_WIDTH => 36)
			port map
				(
    					start_req => start_req,
    					start_ack => start_ack,
    					fin_req => fin_req,
    					fin_ack => fin_ack,
    					init_flag  => init_flag ,
    					tag_mem_read  => tag_mem_read ,
    					tag_mem_write  => tag_mem_write ,
    					read_set_id  => read_set_id ,
    					write_set_id  => write_set_id ,
    					tags_have_been_modified  => tags_have_been_modified ,
    					lwi_has_been_modified  => lwi_has_been_modified ,
    					valids_have_been_modified  => valids_have_been_modified ,
    					dirty_bits_have_been_modified  => dirty_bits_have_been_modified ,
    					updated_set_tags  => updated_set_tags ,
    					updated_set_lwi  => updated_set_lwi ,
    					updated_set_valids  => updated_set_valids ,
    					updated_set_dirty_dword_masks  => updated_set_dirty_dword_masks ,
    					tag_mem_response  => tag_mem_response ,
    					clk => clk, 
					reset => reset
				);

end accessL2TagMemX1024X8_Operator_arch;

library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.mem_component_pack.all;
use ahir.basecomponents.all;

library AjitCustom;
use AjitCustom.AjitGlobalConfigurationPackage.all;
use AjitCustom.AjitCustomComponents.all;
--
-- X2048X8 means  that this manages 2048 lines
-- and set associativity is 8.  Thus a total cache size of 
-- 128KB organized into 256 sets.
-- 
-- Thus, the PA tag width is 30-(log2 (2048/8)) = 30-8=22
--   
entity accessL2TagMemX2048X8_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    init_flag : in  std_logic_vector(0 downto 0);
    tag_mem_read : in  std_logic_vector(0 downto 0);
    tag_mem_write : in  std_logic_vector(0 downto 0);
    read_set_id : in  std_logic_vector(7 downto 0);
    write_set_id : in  std_logic_vector(7 downto 0);
    tags_have_been_modified : in  std_logic_vector(0 downto 0);
    lwi_has_been_modified : in  std_logic_vector(0 downto 0);
    valids_have_been_modified : in  std_logic_vector(0 downto 0);
    dirty_bits_have_been_modified : in  std_logic_vector(0 downto 0);
    updated_set_tags : in  std_logic_vector(175 downto 0);
    updated_set_lwi : in  std_logic_vector(2 downto 0);
    updated_set_valids : in  std_logic_vector(7 downto 0);
    updated_set_dirty_dword_masks : in  std_logic_vector(63 downto 0);
    tag_mem_response : out  std_logic_vector(250 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity accessL2TagMemX2048X8_Operator;
architecture accessL2TagMemX2048X8_Operator_arch of accessL2TagMemX2048X8_Operator is -- 
	signal start_req, start_ack, fin_req, fin_ack: std_logic;
begin --  
	p2lInst:
		Sample_Pulse_To_Level_Translate_Entity
			generic map ("accessL2TagMem_P2L")
			port map 
				( rL => sample_req,
					rR => start_req,
					aL => sample_ack,
					aR => start_ack,
					clk => clk, reset => reset);	
	l2pInst: 
		Level_To_Pulse_Translate_Entity
			generic map ("accessL2TagMem_L2P")
			port map (rL => fin_req,
					rR => update_req,
					aL => fin_ack,
					aR => update_ack,
					clk => clk, reset => reset);

	baseInst:
		accessL2TagMemGeneric
			generic map (LOG2_NUMBER_OF_LINES => 11,
						LOG2_ASSOCIATIVITY => 3,
						LOG2_DWORDS_PER_LINE => 3,
						PA_ADDRESS_WIDTH => 36)
			port map
				(
    					start_req => start_req,
    					start_ack => start_ack,
    					fin_req => fin_req,
    					fin_ack => fin_ack,
    					init_flag  => init_flag ,
    					tag_mem_read  => tag_mem_read ,
    					tag_mem_write  => tag_mem_write ,
    					read_set_id  => read_set_id ,
    					write_set_id  => write_set_id ,
    					tags_have_been_modified  => tags_have_been_modified ,
    					lwi_has_been_modified  => lwi_has_been_modified ,
    					valids_have_been_modified  => valids_have_been_modified ,
    					dirty_bits_have_been_modified  => dirty_bits_have_been_modified ,
    					updated_set_tags  => updated_set_tags ,
    					updated_set_lwi  => updated_set_lwi ,
    					updated_set_valids  => updated_set_valids ,
    					updated_set_dirty_dword_masks  => updated_set_dirty_dword_masks ,
    					tag_mem_response  => tag_mem_response ,
    					clk => clk, 
					reset => reset
				);

end accessL2TagMemX2048X8_Operator_arch;

library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library ahir;
use ahir.mem_component_pack.all;
use ahir.basecomponents.all;

library AjitCustom;
use AjitCustom.AjitGlobalConfigurationPackage.all;
use AjitCustom.AjitCustomComponents.all;
--
-- X4096X8 means  that this manages 4096 lines
-- and set associativity is 8.  Thus a total cache size of 
-- 256KB organized into 512 sets.
-- 
-- Thus, the PA tag width is 30-(log2 (4096/8)) = 30-9=21
--   
entity accessL2TagMemX4096X8_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    init_flag : in  std_logic_vector(0 downto 0);
    tag_mem_read : in  std_logic_vector(0 downto 0);
    tag_mem_write : in  std_logic_vector(0 downto 0);
    read_set_id : in  std_logic_vector(8 downto 0);
    write_set_id : in  std_logic_vector(8 downto 0);
    tags_have_been_modified : in  std_logic_vector(0 downto 0);
    lwi_has_been_modified : in  std_logic_vector(0 downto 0);
    valids_have_been_modified : in  std_logic_vector(0 downto 0);
    dirty_bits_have_been_modified : in  std_logic_vector(0 downto 0);
    updated_set_tags : in  std_logic_vector(167 downto 0);
    updated_set_lwi : in  std_logic_vector(2 downto 0);
    updated_set_valids : in  std_logic_vector(7 downto 0);
    updated_set_dirty_dword_masks : in  std_logic_vector(63 downto 0);
    tag_mem_response : out  std_logic_vector(242 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity accessL2TagMemX4096X8_Operator;
architecture accessL2TagMemX4096X8_Operator_arch of accessL2TagMemX4096X8_Operator is -- 
	signal start_req, start_ack, fin_req, fin_ack: std_logic;
begin --  
	p2lInst:
		Sample_Pulse_To_Level_Translate_Entity
			generic map ("accessL2TagMem_P2L")
			port map 
				( rL => sample_req,
					rR => start_req,
					aL => sample_ack,
					aR => start_ack,
					clk => clk, reset => reset);	
	l2pInst: 
		Level_To_Pulse_Translate_Entity
			generic map ("accessL2TagMem_L2P")
			port map (rL => fin_req,
					rR => update_req,
					aL => fin_ack,
					aR => update_ack,
					clk => clk, reset => reset);

	baseInst:
		accessL2TagMemGeneric
			generic map (LOG2_NUMBER_OF_LINES => 12,
						LOG2_ASSOCIATIVITY => 3,
						LOG2_DWORDS_PER_LINE => 3,
						PA_ADDRESS_WIDTH => 36)
			port map
				(
    					start_req => start_req,
    					start_ack => start_ack,
    					fin_req => fin_req,
    					fin_ack => fin_ack,
    					init_flag  => init_flag ,
    					tag_mem_read  => tag_mem_read ,
    					tag_mem_write  => tag_mem_write ,
    					read_set_id  => read_set_id ,
    					write_set_id  => write_set_id ,
    					tags_have_been_modified  => tags_have_been_modified ,
    					lwi_has_been_modified  => lwi_has_been_modified ,
    					valids_have_been_modified  => valids_have_been_modified ,
    					dirty_bits_have_been_modified  => dirty_bits_have_been_modified ,
    					updated_set_tags  => updated_set_tags ,
    					updated_set_lwi  => updated_set_lwi ,
    					updated_set_valids  => updated_set_valids ,
    					updated_set_dirty_dword_masks  => updated_set_dirty_dword_masks ,
    					tag_mem_response  => tag_mem_response ,
    					clk => clk, 
					reset => reset
				);

end accessL2TagMemX4096X8_Operator_arch;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;


entity rt_clock_counter is

	port (
			clk, reset: in std_logic;
			one_hz_rt_clock: in std_logic_vector(0 downto 0);
			count_value : out std_logic_vector(31 downto 0)
		);

end entity rt_clock_counter;


architecture Behave of rt_clock_counter is

	signal counter : integer;
	signal last_one_hz_rt_clock, one_hz_rt_clock_synch: std_logic_vector(0 downto 0);
	signal rt_rising, rt_falling: boolean;
	type FsmState is (IDLE, RT_HIGH, RT_LOW);
	signal fsm_state: FsmState;

begin
	process(clk, reset)
	begin
		if(clk'event and clk = '1') then
			one_hz_rt_clock_synch <= one_hz_rt_clock;
			last_one_hz_rt_clock  <= one_hz_rt_clock_synch;
		end if;
	end process;

	rt_rising  <= (one_hz_rt_clock_synch(0) = '1') and (last_one_hz_rt_clock(0) = '0');
	rt_falling <= (one_hz_rt_clock_synch(0) = '0') and (last_one_hz_rt_clock(0) = '1');

	-- counter
	process(clk, reset, fsm_state, counter, rt_rising, rt_falling)
		variable latch_counter_var: boolean;
		variable next_counter_var : integer;
		variable next_fsm_state_var : FsmState;
	begin
		latch_counter_var := false;
		next_counter_var  := counter;
		next_fsm_state_var := fsm_state;

		case fsm_state is 
			when IDLE => 
				if rt_rising then
					next_counter_var := 0;
					next_fsm_state_var := RT_HIGH;
				end if;
			when RT_HIGH =>
				next_counter_var := (counter + 1);
				if(rt_falling) then
					next_fsm_state_var := RT_LOW;
				end if;
			when RT_LOW =>
				if(rt_rising) then
					latch_counter_var := true;
					next_counter_var := 0;
					next_fsm_state_var := RT_HIGH;
				else
					next_counter_var := (counter + 1);
				end if;
		end case;

		if(clk'event and clk = '1') then
			if(reset = '1') then
				counter <= 0;
				count_value <= (others => '0');				
				fsm_state <= IDLE;
			else
				counter <= next_counter_var;
				fsm_state <= next_fsm_state_var;

				if(latch_counter_var) then
					count_value <= std_logic_vector(to_unsigned(counter, 32));
				end if;

			end if;
		end if;
	end process;

end Behave; 
-- VHDL global package produced by vc2vhdl from virtual circuit (vc) description 
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
package baud_control_calculator_global_package is -- 
  component baud_control_calculator is -- 
    port (-- 
      clk : in std_logic;
      reset : in std_logic;
      BAUD_CONTROL_WORD_SIG: out std_logic_vector(31 downto 0);
      BAUD_CONTROL_WORD_VALID: out std_logic_vector(0 downto 0);
      BAUD_RATE_SIG: in std_logic_vector(31 downto 0);
      CLK_FREQUENCY_SIG: in std_logic_vector(31 downto 0);
      CLOCK_FREQUENCY_VALID: in std_logic_vector(0 downto 0)); -- 
    -- 
  end component;
  -- 
end package baud_control_calculator_global_package;
-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library AjitCustom;
use AjitCustom.baud_control_calculator_global_package.all;
entity baudControlCalculatorDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    BAUD_RATE_SIG : in std_logic_vector(31 downto 0);
    CLK_FREQUENCY_SIG : in std_logic_vector(31 downto 0);
    CLOCK_FREQUENCY_VALID : in std_logic_vector(0 downto 0);
    BAUD_CONTROL_WORD_SIG_pipe_write_req : out  std_logic_vector(0 downto 0);
    BAUD_CONTROL_WORD_SIG_pipe_write_ack : in   std_logic_vector(0 downto 0);
    BAUD_CONTROL_WORD_SIG_pipe_write_data : out  std_logic_vector(31 downto 0);
    BAUD_CONTROL_WORD_VALID_pipe_write_req : out  std_logic_vector(0 downto 0);
    BAUD_CONTROL_WORD_VALID_pipe_write_ack : in   std_logic_vector(0 downto 0);
    BAUD_CONTROL_WORD_VALID_pipe_write_data : out  std_logic_vector(0 downto 0);
    my_gcd_call_reqs : out  std_logic_vector(0 downto 0);
    my_gcd_call_acks : in   std_logic_vector(0 downto 0);
    my_gcd_call_data : out  std_logic_vector(63 downto 0);
    my_gcd_call_tag  :  out  std_logic_vector(0 downto 0);
    my_gcd_return_reqs : out  std_logic_vector(0 downto 0);
    my_gcd_return_acks : in   std_logic_vector(0 downto 0);
    my_gcd_return_data : in   std_logic_vector(31 downto 0);
    my_gcd_return_tag :  in   std_logic_vector(0 downto 0);
    my_div_call_reqs : out  std_logic_vector(0 downto 0);
    my_div_call_acks : in   std_logic_vector(0 downto 0);
    my_div_call_data : out  std_logic_vector(63 downto 0);
    my_div_call_tag  :  out  std_logic_vector(1 downto 0);
    my_div_return_reqs : out  std_logic_vector(0 downto 0);
    my_div_return_acks : in   std_logic_vector(0 downto 0);
    my_div_return_data : in   std_logic_vector(31 downto 0);
    my_div_return_tag :  in   std_logic_vector(1 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity baudControlCalculatorDaemon;
architecture baudControlCalculatorDaemon_arch of baudControlCalculatorDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal baudControlCalculatorDaemon_CP_295_start: Boolean;
  signal baudControlCalculatorDaemon_CP_295_symbol: Boolean;
  -- volatile/operator module components. 
  component my_gcd is -- 
    generic (tag_length : integer); 
    port ( -- 
      A : in  std_logic_vector(31 downto 0);
      B : in  std_logic_vector(31 downto 0);
      GCD : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component my_div is -- 
    generic (tag_length : integer); 
    port ( -- 
      A : in  std_logic_vector(31 downto 0);
      B : in  std_logic_vector(31 downto 0);
      Q : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal WPIPE_BAUD_CONTROL_WORD_VALID_130_inst_req_0 : boolean;
  signal WPIPE_BAUD_CONTROL_WORD_VALID_130_inst_ack_0 : boolean;
  signal WPIPE_BAUD_CONTROL_WORD_VALID_130_inst_req_1 : boolean;
  signal WPIPE_BAUD_CONTROL_WORD_VALID_130_inst_ack_1 : boolean;
  signal W_clock_valid_135_inst_req_0 : boolean;
  signal W_clock_valid_135_inst_ack_0 : boolean;
  signal W_clock_valid_135_inst_req_1 : boolean;
  signal W_clock_valid_135_inst_ack_1 : boolean;
  signal if_stmt_138_branch_req_0 : boolean;
  signal if_stmt_138_branch_ack_1 : boolean;
  signal if_stmt_138_branch_ack_0 : boolean;
  signal CONCAT_u16_u32_150_inst_req_0 : boolean;
  signal CONCAT_u16_u32_150_inst_ack_0 : boolean;
  signal CONCAT_u16_u32_150_inst_req_1 : boolean;
  signal CONCAT_u16_u32_150_inst_ack_1 : boolean;
  signal CONCAT_u28_u32_159_inst_req_0 : boolean;
  signal CONCAT_u28_u32_159_inst_ack_0 : boolean;
  signal CONCAT_u28_u32_159_inst_req_1 : boolean;
  signal CONCAT_u28_u32_159_inst_ack_1 : boolean;
  signal call_stmt_164_call_req_0 : boolean;
  signal call_stmt_164_call_ack_0 : boolean;
  signal call_stmt_164_call_req_1 : boolean;
  signal call_stmt_164_call_ack_1 : boolean;
  signal call_stmt_168_call_req_0 : boolean;
  signal call_stmt_168_call_ack_0 : boolean;
  signal call_stmt_168_call_req_1 : boolean;
  signal call_stmt_168_call_ack_1 : boolean;
  signal call_stmt_172_call_req_0 : boolean;
  signal call_stmt_172_call_ack_0 : boolean;
  signal call_stmt_172_call_req_1 : boolean;
  signal call_stmt_172_call_ack_1 : boolean;
  signal SUB_u32_u32_176_inst_req_0 : boolean;
  signal SUB_u32_u32_176_inst_ack_0 : boolean;
  signal SUB_u32_u32_176_inst_req_1 : boolean;
  signal SUB_u32_u32_176_inst_ack_1 : boolean;
  signal CONCAT_u20_u32_188_inst_req_0 : boolean;
  signal CONCAT_u20_u32_188_inst_ack_0 : boolean;
  signal CONCAT_u20_u32_188_inst_req_1 : boolean;
  signal CONCAT_u20_u32_188_inst_ack_1 : boolean;
  signal WPIPE_BAUD_CONTROL_WORD_SIG_178_inst_req_0 : boolean;
  signal WPIPE_BAUD_CONTROL_WORD_SIG_178_inst_ack_0 : boolean;
  signal WPIPE_BAUD_CONTROL_WORD_SIG_178_inst_req_1 : boolean;
  signal WPIPE_BAUD_CONTROL_WORD_SIG_178_inst_ack_1 : boolean;
  signal WPIPE_BAUD_CONTROL_WORD_VALID_191_inst_req_0 : boolean;
  signal WPIPE_BAUD_CONTROL_WORD_VALID_191_inst_ack_0 : boolean;
  signal WPIPE_BAUD_CONTROL_WORD_VALID_191_inst_req_1 : boolean;
  signal WPIPE_BAUD_CONTROL_WORD_VALID_191_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "baudControlCalculatorDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  baudControlCalculatorDaemon_CP_295_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "baudControlCalculatorDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= baudControlCalculatorDaemon_CP_295_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= baudControlCalculatorDaemon_CP_295_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= baudControlCalculatorDaemon_CP_295_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  baudControlCalculatorDaemon_CP_295: Block -- control-path 
    signal baudControlCalculatorDaemon_CP_295_elements: BooleanArray(32 downto 0);
    -- 
  begin -- 
    baudControlCalculatorDaemon_CP_295_elements(0) <= baudControlCalculatorDaemon_CP_295_start;
    baudControlCalculatorDaemon_CP_295_symbol <= baudControlCalculatorDaemon_CP_295_elements(3);
    -- CP-element group 0:  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_132/$entry
      -- CP-element group 0: 	 assign_stmt_132/WPIPE_BAUD_CONTROL_WORD_VALID_130_sample_start_
      -- CP-element group 0: 	 assign_stmt_132/WPIPE_BAUD_CONTROL_WORD_VALID_130_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_132/WPIPE_BAUD_CONTROL_WORD_VALID_130_Sample/req
      -- 
    req_308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => baudControlCalculatorDaemon_CP_295_elements(0), ack => WPIPE_BAUD_CONTROL_WORD_VALID_130_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_132/WPIPE_BAUD_CONTROL_WORD_VALID_130_sample_completed_
      -- CP-element group 1: 	 assign_stmt_132/WPIPE_BAUD_CONTROL_WORD_VALID_130_update_start_
      -- CP-element group 1: 	 assign_stmt_132/WPIPE_BAUD_CONTROL_WORD_VALID_130_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_132/WPIPE_BAUD_CONTROL_WORD_VALID_130_Sample/ack
      -- CP-element group 1: 	 assign_stmt_132/WPIPE_BAUD_CONTROL_WORD_VALID_130_Update/$entry
      -- CP-element group 1: 	 assign_stmt_132/WPIPE_BAUD_CONTROL_WORD_VALID_130_Update/req
      -- 
    ack_309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_BAUD_CONTROL_WORD_VALID_130_inst_ack_0, ack => baudControlCalculatorDaemon_CP_295_elements(1)); -- 
    req_313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => baudControlCalculatorDaemon_CP_295_elements(1), ack => WPIPE_BAUD_CONTROL_WORD_VALID_130_inst_req_1); -- 
    -- CP-element group 2:  branch  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	31 
    -- CP-element group 2:  members (10) 
      -- CP-element group 2: 	 assign_stmt_132/$exit
      -- CP-element group 2: 	 assign_stmt_132/WPIPE_BAUD_CONTROL_WORD_VALID_130_update_completed_
      -- CP-element group 2: 	 assign_stmt_132/WPIPE_BAUD_CONTROL_WORD_VALID_130_Update/$exit
      -- CP-element group 2: 	 assign_stmt_132/WPIPE_BAUD_CONTROL_WORD_VALID_130_Update/ack
      -- CP-element group 2: 	 branch_block_stmt_133/$entry
      -- CP-element group 2: 	 branch_block_stmt_133/branch_block_stmt_133__entry__
      -- CP-element group 2: 	 branch_block_stmt_133/merge_stmt_134__entry__
      -- CP-element group 2: 	 branch_block_stmt_133/merge_stmt_134_dead_link/$entry
      -- CP-element group 2: 	 branch_block_stmt_133/merge_stmt_134__entry___PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_133/merge_stmt_134__entry___PhiReq/$exit
      -- 
    ack_314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_BAUD_CONTROL_WORD_VALID_130_inst_ack_1, ack => baudControlCalculatorDaemon_CP_295_elements(2)); -- 
    -- CP-element group 3:  transition  place  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 $exit
      -- CP-element group 3: 	 branch_block_stmt_133/$exit
      -- CP-element group 3: 	 branch_block_stmt_133/branch_block_stmt_133__exit__
      -- 
    baudControlCalculatorDaemon_CP_295_elements(3) <= false; 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	31 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_133/assign_stmt_137/assign_stmt_137_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_133/assign_stmt_137/assign_stmt_137_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_133/assign_stmt_137/assign_stmt_137_Sample/ack
      -- 
    ack_344_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_clock_valid_135_inst_ack_0, ack => baudControlCalculatorDaemon_CP_295_elements(4)); -- 
    -- CP-element group 5:  branch  transition  place  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	31 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5: 	7 
    -- CP-element group 5:  members (25) 
      -- CP-element group 5: 	 branch_block_stmt_133/assign_stmt_137__exit__
      -- CP-element group 5: 	 branch_block_stmt_133/if_stmt_138__entry__
      -- CP-element group 5: 	 branch_block_stmt_133/assign_stmt_137/$exit
      -- CP-element group 5: 	 branch_block_stmt_133/assign_stmt_137/assign_stmt_137_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_133/assign_stmt_137/assign_stmt_137_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_133/assign_stmt_137/assign_stmt_137_Update/ack
      -- CP-element group 5: 	 branch_block_stmt_133/if_stmt_138_dead_link/$entry
      -- CP-element group 5: 	 branch_block_stmt_133/if_stmt_138_eval_test/$entry
      -- CP-element group 5: 	 branch_block_stmt_133/if_stmt_138_eval_test/$exit
      -- CP-element group 5: 	 branch_block_stmt_133/if_stmt_138_eval_test/NOT_u1_u1_140/$entry
      -- CP-element group 5: 	 branch_block_stmt_133/if_stmt_138_eval_test/NOT_u1_u1_140/$exit
      -- CP-element group 5: 	 branch_block_stmt_133/if_stmt_138_eval_test/NOT_u1_u1_140/SplitProtocol/$entry
      -- CP-element group 5: 	 branch_block_stmt_133/if_stmt_138_eval_test/NOT_u1_u1_140/SplitProtocol/$exit
      -- CP-element group 5: 	 branch_block_stmt_133/if_stmt_138_eval_test/NOT_u1_u1_140/SplitProtocol/Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_133/if_stmt_138_eval_test/NOT_u1_u1_140/SplitProtocol/Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_133/if_stmt_138_eval_test/NOT_u1_u1_140/SplitProtocol/Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_133/if_stmt_138_eval_test/NOT_u1_u1_140/SplitProtocol/Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_133/if_stmt_138_eval_test/NOT_u1_u1_140/SplitProtocol/Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_133/if_stmt_138_eval_test/NOT_u1_u1_140/SplitProtocol/Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_133/if_stmt_138_eval_test/NOT_u1_u1_140/SplitProtocol/Update/cr
      -- CP-element group 5: 	 branch_block_stmt_133/if_stmt_138_eval_test/NOT_u1_u1_140/SplitProtocol/Update/ca
      -- CP-element group 5: 	 branch_block_stmt_133/if_stmt_138_eval_test/branch_req
      -- CP-element group 5: 	 branch_block_stmt_133/NOT_u1_u1_140_place
      -- CP-element group 5: 	 branch_block_stmt_133/if_stmt_138_if_link/$entry
      -- CP-element group 5: 	 branch_block_stmt_133/if_stmt_138_else_link/$entry
      -- 
    ack_349_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_clock_valid_135_inst_ack_1, ack => baudControlCalculatorDaemon_CP_295_elements(5)); -- 
    branch_req_373_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_373_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => baudControlCalculatorDaemon_CP_295_elements(5), ack => if_stmt_138_branch_req_0); -- 
    -- CP-element group 6:  transition  place  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	31 
    -- CP-element group 6:  members (5) 
      -- CP-element group 6: 	 branch_block_stmt_133/if_stmt_138_if_link/$exit
      -- CP-element group 6: 	 branch_block_stmt_133/if_stmt_138_if_link/if_choice_transition
      -- CP-element group 6: 	 branch_block_stmt_133/wait_on_clock
      -- CP-element group 6: 	 branch_block_stmt_133/wait_on_clock_PhiReq/$entry
      -- CP-element group 6: 	 branch_block_stmt_133/wait_on_clock_PhiReq/$exit
      -- 
    if_choice_transition_378_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_138_branch_ack_1, ack => baudControlCalculatorDaemon_CP_295_elements(6)); -- 
    -- CP-element group 7:  merge  branch  transition  place  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	5 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	32 
    -- CP-element group 7:  members (7) 
      -- CP-element group 7: 	 branch_block_stmt_133/if_stmt_138__exit__
      -- CP-element group 7: 	 branch_block_stmt_133/merge_stmt_143__entry__
      -- CP-element group 7: 	 branch_block_stmt_133/if_stmt_138_else_link/$exit
      -- CP-element group 7: 	 branch_block_stmt_133/if_stmt_138_else_link/else_choice_transition
      -- CP-element group 7: 	 branch_block_stmt_133/merge_stmt_143_dead_link/$entry
      -- CP-element group 7: 	 branch_block_stmt_133/merge_stmt_143__entry___PhiReq/$entry
      -- CP-element group 7: 	 branch_block_stmt_133/merge_stmt_143__entry___PhiReq/$exit
      -- 
    else_choice_transition_382_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_138_branch_ack_0, ack => baudControlCalculatorDaemon_CP_295_elements(7)); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	32 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u16_u32_150_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u16_u32_150_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u16_u32_150_Sample/ra
      -- 
    ra_395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u16_u32_150_inst_ack_0, ack => baudControlCalculatorDaemon_CP_295_elements(8)); -- 
    -- CP-element group 9:  fork  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	32 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	18 
    -- CP-element group 9: 	12 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u16_u32_150_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u16_u32_150_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u16_u32_150_Update/ca
      -- 
    ca_400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u16_u32_150_inst_ack_1, ack => baudControlCalculatorDaemon_CP_295_elements(9)); -- 
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	32 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u28_u32_159_sample_completed_
      -- CP-element group 10: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u28_u32_159_Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u28_u32_159_Sample/ra
      -- 
    ra_409_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u28_u32_159_inst_ack_0, ack => baudControlCalculatorDaemon_CP_295_elements(10)); -- 
    -- CP-element group 11:  fork  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	32 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u28_u32_159_update_completed_
      -- CP-element group 11: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u28_u32_159_Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u28_u32_159_Update/ca
      -- 
    ca_414_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u28_u32_159_inst_ack_1, ack => baudControlCalculatorDaemon_CP_295_elements(11)); -- 
    -- CP-element group 12:  join  transition  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_164_sample_start_
      -- CP-element group 12: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_164_Sample/$entry
      -- CP-element group 12: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_164_Sample/crr
      -- 
    crr_422_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_422_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => baudControlCalculatorDaemon_CP_295_elements(12), ack => call_stmt_164_call_req_0); -- 
    baudControlCalculatorDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 47) := "baudControlCalculatorDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= baudControlCalculatorDaemon_CP_295_elements(9) & baudControlCalculatorDaemon_CP_295_elements(11);
      gj_baudControlCalculatorDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => baudControlCalculatorDaemon_CP_295_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_164_sample_completed_
      -- CP-element group 13: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_164_Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_164_Sample/cra
      -- 
    cra_423_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_164_call_ack_0, ack => baudControlCalculatorDaemon_CP_295_elements(13)); -- 
    -- CP-element group 14:  fork  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	32 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_164_update_completed_
      -- CP-element group 14: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_164_Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_164_Update/cca
      -- 
    cca_428_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_164_call_ack_1, ack => baudControlCalculatorDaemon_CP_295_elements(14)); -- 
    -- CP-element group 15:  join  transition  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: 	11 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_168_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_168_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_168_Sample/crr
      -- 
    crr_436_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_436_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => baudControlCalculatorDaemon_CP_295_elements(15), ack => call_stmt_168_call_req_0); -- 
    baudControlCalculatorDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 47) := "baudControlCalculatorDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= baudControlCalculatorDaemon_CP_295_elements(14) & baudControlCalculatorDaemon_CP_295_elements(11);
      gj_baudControlCalculatorDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => baudControlCalculatorDaemon_CP_295_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_168_sample_completed_
      -- CP-element group 16: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_168_Sample/$exit
      -- CP-element group 16: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_168_Sample/cra
      -- 
    cra_437_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_168_call_ack_0, ack => baudControlCalculatorDaemon_CP_295_elements(16)); -- 
    -- CP-element group 17:  fork  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	32 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	24 
    -- CP-element group 17: 	21 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_168_update_completed_
      -- CP-element group 17: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_168_Update/$exit
      -- CP-element group 17: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_168_Update/cca
      -- 
    cca_442_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_168_call_ack_1, ack => baudControlCalculatorDaemon_CP_295_elements(17)); -- 
    -- CP-element group 18:  join  transition  output  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	9 
    -- CP-element group 18: 	14 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_172_sample_start_
      -- CP-element group 18: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_172_Sample/$entry
      -- CP-element group 18: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_172_Sample/crr
      -- 
    crr_450_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_450_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => baudControlCalculatorDaemon_CP_295_elements(18), ack => call_stmt_172_call_req_0); -- 
    baudControlCalculatorDaemon_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 47) := "baudControlCalculatorDaemon_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= baudControlCalculatorDaemon_CP_295_elements(9) & baudControlCalculatorDaemon_CP_295_elements(14);
      gj_baudControlCalculatorDaemon_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => baudControlCalculatorDaemon_CP_295_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_172_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_172_Sample/$exit
      -- CP-element group 19: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_172_Sample/cra
      -- 
    cra_451_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_172_call_ack_0, ack => baudControlCalculatorDaemon_CP_295_elements(19)); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	32 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_172_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_172_Update/$exit
      -- CP-element group 20: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_172_Update/cca
      -- 
    cca_456_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_172_call_ack_1, ack => baudControlCalculatorDaemon_CP_295_elements(20)); -- 
    -- CP-element group 21:  join  transition  output  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	17 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/SUB_u32_u32_176_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/SUB_u32_u32_176_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/SUB_u32_u32_176_Sample/rr
      -- 
    rr_464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => baudControlCalculatorDaemon_CP_295_elements(21), ack => SUB_u32_u32_176_inst_req_0); -- 
    baudControlCalculatorDaemon_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 47) := "baudControlCalculatorDaemon_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= baudControlCalculatorDaemon_CP_295_elements(17) & baudControlCalculatorDaemon_CP_295_elements(20);
      gj_baudControlCalculatorDaemon_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => baudControlCalculatorDaemon_CP_295_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/SUB_u32_u32_176_sample_completed_
      -- CP-element group 22: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/SUB_u32_u32_176_Sample/$exit
      -- CP-element group 22: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/SUB_u32_u32_176_Sample/ra
      -- 
    ra_465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_176_inst_ack_0, ack => baudControlCalculatorDaemon_CP_295_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	32 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/SUB_u32_u32_176_update_completed_
      -- CP-element group 23: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/SUB_u32_u32_176_Update/$exit
      -- CP-element group 23: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/SUB_u32_u32_176_Update/ca
      -- 
    ca_470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u32_u32_176_inst_ack_1, ack => baudControlCalculatorDaemon_CP_295_elements(23)); -- 
    -- CP-element group 24:  join  transition  output  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: 	17 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u20_u32_188_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u20_u32_188_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u20_u32_188_Sample/rr
      -- 
    rr_478_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_478_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => baudControlCalculatorDaemon_CP_295_elements(24), ack => CONCAT_u20_u32_188_inst_req_0); -- 
    baudControlCalculatorDaemon_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 47) := "baudControlCalculatorDaemon_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= baudControlCalculatorDaemon_CP_295_elements(23) & baudControlCalculatorDaemon_CP_295_elements(17);
      gj_baudControlCalculatorDaemon_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => baudControlCalculatorDaemon_CP_295_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u20_u32_188_sample_completed_
      -- CP-element group 25: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u20_u32_188_Sample/$exit
      -- CP-element group 25: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u20_u32_188_Sample/ra
      -- 
    ra_479_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u20_u32_188_inst_ack_0, ack => baudControlCalculatorDaemon_CP_295_elements(25)); -- 
    -- CP-element group 26:  transition  input  output  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	32 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (6) 
      -- CP-element group 26: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u20_u32_188_update_completed_
      -- CP-element group 26: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u20_u32_188_Update/$exit
      -- CP-element group 26: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u20_u32_188_Update/ca
      -- CP-element group 26: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/WPIPE_BAUD_CONTROL_WORD_SIG_178_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/WPIPE_BAUD_CONTROL_WORD_SIG_178_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/WPIPE_BAUD_CONTROL_WORD_SIG_178_Sample/req
      -- 
    ca_484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u20_u32_188_inst_ack_1, ack => baudControlCalculatorDaemon_CP_295_elements(26)); -- 
    req_492_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_492_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => baudControlCalculatorDaemon_CP_295_elements(26), ack => WPIPE_BAUD_CONTROL_WORD_SIG_178_inst_req_0); -- 
    -- CP-element group 27:  transition  input  output  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	28 
    -- CP-element group 27:  members (6) 
      -- CP-element group 27: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/WPIPE_BAUD_CONTROL_WORD_SIG_178_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/WPIPE_BAUD_CONTROL_WORD_SIG_178_update_start_
      -- CP-element group 27: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/WPIPE_BAUD_CONTROL_WORD_SIG_178_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/WPIPE_BAUD_CONTROL_WORD_SIG_178_Sample/ack
      -- CP-element group 27: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/WPIPE_BAUD_CONTROL_WORD_SIG_178_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/WPIPE_BAUD_CONTROL_WORD_SIG_178_Update/req
      -- 
    ack_493_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_BAUD_CONTROL_WORD_SIG_178_inst_ack_0, ack => baudControlCalculatorDaemon_CP_295_elements(27)); -- 
    req_497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => baudControlCalculatorDaemon_CP_295_elements(27), ack => WPIPE_BAUD_CONTROL_WORD_SIG_178_inst_req_1); -- 
    -- CP-element group 28:  transition  place  input  output  bypass 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	27 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28:  members (10) 
      -- CP-element group 28: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189__exit__
      -- CP-element group 28: 	 branch_block_stmt_133/assign_stmt_193__entry__
      -- CP-element group 28: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/$exit
      -- CP-element group 28: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/WPIPE_BAUD_CONTROL_WORD_SIG_178_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/WPIPE_BAUD_CONTROL_WORD_SIG_178_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/WPIPE_BAUD_CONTROL_WORD_SIG_178_Update/ack
      -- CP-element group 28: 	 branch_block_stmt_133/assign_stmt_193/$entry
      -- CP-element group 28: 	 branch_block_stmt_133/assign_stmt_193/WPIPE_BAUD_CONTROL_WORD_VALID_191_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_133/assign_stmt_193/WPIPE_BAUD_CONTROL_WORD_VALID_191_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_133/assign_stmt_193/WPIPE_BAUD_CONTROL_WORD_VALID_191_Sample/req
      -- 
    ack_498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_BAUD_CONTROL_WORD_SIG_178_inst_ack_1, ack => baudControlCalculatorDaemon_CP_295_elements(28)); -- 
    req_509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => baudControlCalculatorDaemon_CP_295_elements(28), ack => WPIPE_BAUD_CONTROL_WORD_VALID_191_inst_req_0); -- 
    -- CP-element group 29:  transition  input  output  bypass 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	30 
    -- CP-element group 29:  members (6) 
      -- CP-element group 29: 	 branch_block_stmt_133/assign_stmt_193/WPIPE_BAUD_CONTROL_WORD_VALID_191_sample_completed_
      -- CP-element group 29: 	 branch_block_stmt_133/assign_stmt_193/WPIPE_BAUD_CONTROL_WORD_VALID_191_update_start_
      -- CP-element group 29: 	 branch_block_stmt_133/assign_stmt_193/WPIPE_BAUD_CONTROL_WORD_VALID_191_Sample/$exit
      -- CP-element group 29: 	 branch_block_stmt_133/assign_stmt_193/WPIPE_BAUD_CONTROL_WORD_VALID_191_Sample/ack
      -- CP-element group 29: 	 branch_block_stmt_133/assign_stmt_193/WPIPE_BAUD_CONTROL_WORD_VALID_191_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_133/assign_stmt_193/WPIPE_BAUD_CONTROL_WORD_VALID_191_Update/req
      -- 
    ack_510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_BAUD_CONTROL_WORD_VALID_191_inst_ack_0, ack => baudControlCalculatorDaemon_CP_295_elements(29)); -- 
    req_514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => baudControlCalculatorDaemon_CP_295_elements(29), ack => WPIPE_BAUD_CONTROL_WORD_VALID_191_inst_req_1); -- 
    -- CP-element group 30:  transition  place  input  bypass 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	29 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (8) 
      -- CP-element group 30: 	 branch_block_stmt_133/assign_stmt_193__exit__
      -- CP-element group 30: 	 branch_block_stmt_133/loopback
      -- CP-element group 30: 	 branch_block_stmt_133/assign_stmt_193/$exit
      -- CP-element group 30: 	 branch_block_stmt_133/assign_stmt_193/WPIPE_BAUD_CONTROL_WORD_VALID_191_update_completed_
      -- CP-element group 30: 	 branch_block_stmt_133/assign_stmt_193/WPIPE_BAUD_CONTROL_WORD_VALID_191_Update/$exit
      -- CP-element group 30: 	 branch_block_stmt_133/assign_stmt_193/WPIPE_BAUD_CONTROL_WORD_VALID_191_Update/ack
      -- CP-element group 30: 	 branch_block_stmt_133/loopback_PhiReq/$entry
      -- CP-element group 30: 	 branch_block_stmt_133/loopback_PhiReq/$exit
      -- 
    ack_515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_BAUD_CONTROL_WORD_VALID_191_inst_ack_1, ack => baudControlCalculatorDaemon_CP_295_elements(30)); -- 
    -- CP-element group 31:  merge  fork  transition  place  output  bypass 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	6 
    -- CP-element group 31: 	2 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	5 
    -- CP-element group 31: 	4 
    -- CP-element group 31:  members (13) 
      -- CP-element group 31: 	 branch_block_stmt_133/merge_stmt_134__exit__
      -- CP-element group 31: 	 branch_block_stmt_133/assign_stmt_137__entry__
      -- CP-element group 31: 	 branch_block_stmt_133/assign_stmt_137/$entry
      -- CP-element group 31: 	 branch_block_stmt_133/assign_stmt_137/assign_stmt_137_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_133/assign_stmt_137/assign_stmt_137_update_start_
      -- CP-element group 31: 	 branch_block_stmt_133/assign_stmt_137/assign_stmt_137_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_133/assign_stmt_137/assign_stmt_137_Sample/req
      -- CP-element group 31: 	 branch_block_stmt_133/assign_stmt_137/assign_stmt_137_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_133/assign_stmt_137/assign_stmt_137_Update/req
      -- CP-element group 31: 	 branch_block_stmt_133/merge_stmt_134_PhiReqMerge
      -- CP-element group 31: 	 branch_block_stmt_133/merge_stmt_134_PhiAck/$entry
      -- CP-element group 31: 	 branch_block_stmt_133/merge_stmt_134_PhiAck/$exit
      -- CP-element group 31: 	 branch_block_stmt_133/merge_stmt_134_PhiAck/dummy
      -- 
    req_343_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_343_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => baudControlCalculatorDaemon_CP_295_elements(31), ack => W_clock_valid_135_inst_req_0); -- 
    req_348_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_348_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => baudControlCalculatorDaemon_CP_295_elements(31), ack => W_clock_valid_135_inst_req_1); -- 
    baudControlCalculatorDaemon_CP_295_elements(31) <= OrReduce(baudControlCalculatorDaemon_CP_295_elements(6) & baudControlCalculatorDaemon_CP_295_elements(2));
    -- CP-element group 32:  merge  fork  transition  place  output  bypass 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	7 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	23 
    -- CP-element group 32: 	10 
    -- CP-element group 32: 	17 
    -- CP-element group 32: 	9 
    -- CP-element group 32: 	8 
    -- CP-element group 32: 	14 
    -- CP-element group 32: 	11 
    -- CP-element group 32: 	20 
    -- CP-element group 32: 	26 
    -- CP-element group 32:  members (34) 
      -- CP-element group 32: 	 branch_block_stmt_133/merge_stmt_143__exit__
      -- CP-element group 32: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189__entry__
      -- CP-element group 32: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/$entry
      -- CP-element group 32: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u16_u32_150_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u16_u32_150_update_start_
      -- CP-element group 32: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u16_u32_150_Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u16_u32_150_Sample/rr
      -- CP-element group 32: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u16_u32_150_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u16_u32_150_Update/cr
      -- CP-element group 32: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u28_u32_159_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u28_u32_159_update_start_
      -- CP-element group 32: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u28_u32_159_Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u28_u32_159_Sample/rr
      -- CP-element group 32: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u28_u32_159_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u28_u32_159_Update/cr
      -- CP-element group 32: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_164_update_start_
      -- CP-element group 32: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_164_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_164_Update/ccr
      -- CP-element group 32: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_168_update_start_
      -- CP-element group 32: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_168_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_168_Update/ccr
      -- CP-element group 32: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_172_update_start_
      -- CP-element group 32: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_172_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/call_stmt_172_Update/ccr
      -- CP-element group 32: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/SUB_u32_u32_176_update_start_
      -- CP-element group 32: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/SUB_u32_u32_176_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/SUB_u32_u32_176_Update/cr
      -- CP-element group 32: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u20_u32_188_update_start_
      -- CP-element group 32: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u20_u32_188_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_133/assign_stmt_151_to_assign_stmt_189/CONCAT_u20_u32_188_Update/cr
      -- CP-element group 32: 	 branch_block_stmt_133/merge_stmt_143_PhiReqMerge
      -- CP-element group 32: 	 branch_block_stmt_133/merge_stmt_143_PhiAck/$entry
      -- CP-element group 32: 	 branch_block_stmt_133/merge_stmt_143_PhiAck/$exit
      -- CP-element group 32: 	 branch_block_stmt_133/merge_stmt_143_PhiAck/dummy
      -- 
    rr_394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => baudControlCalculatorDaemon_CP_295_elements(32), ack => CONCAT_u16_u32_150_inst_req_0); -- 
    cr_399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => baudControlCalculatorDaemon_CP_295_elements(32), ack => CONCAT_u16_u32_150_inst_req_1); -- 
    rr_408_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_408_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => baudControlCalculatorDaemon_CP_295_elements(32), ack => CONCAT_u28_u32_159_inst_req_0); -- 
    cr_413_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_413_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => baudControlCalculatorDaemon_CP_295_elements(32), ack => CONCAT_u28_u32_159_inst_req_1); -- 
    ccr_427_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_427_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => baudControlCalculatorDaemon_CP_295_elements(32), ack => call_stmt_164_call_req_1); -- 
    ccr_441_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_441_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => baudControlCalculatorDaemon_CP_295_elements(32), ack => call_stmt_168_call_req_1); -- 
    ccr_455_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_455_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => baudControlCalculatorDaemon_CP_295_elements(32), ack => call_stmt_172_call_req_1); -- 
    cr_469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => baudControlCalculatorDaemon_CP_295_elements(32), ack => SUB_u32_u32_176_inst_req_1); -- 
    cr_483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => baudControlCalculatorDaemon_CP_295_elements(32), ack => CONCAT_u20_u32_188_inst_req_1); -- 
    baudControlCalculatorDaemon_CP_295_elements(32) <= OrReduce(baudControlCalculatorDaemon_CP_295_elements(7) & baudControlCalculatorDaemon_CP_295_elements(30));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal BF_168 : std_logic_vector(31 downto 0);
    signal BL_177 : std_logic_vector(31 downto 0);
    signal BLx_172 : std_logic_vector(31 downto 0);
    signal BRx16_160 : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u20_183_wire : std_logic_vector(19 downto 0);
    signal CONCAT_u20_u32_188_wire : std_logic_vector(31 downto 0);
    signal GCD_164 : std_logic_vector(31 downto 0);
    signal NOT_u1_u1_140_wire : std_logic_vector(0 downto 0);
    signal RPIPE_BAUD_RATE_SIG_153_wire : std_logic_vector(31 downto 0);
    signal RPIPE_CLK_FREQUENCY_SIG_145_wire : std_logic_vector(31 downto 0);
    signal RPIPE_CLOCK_FREQUENCY_VALID_136_wire : std_logic_vector(0 downto 0);
    signal SS_151 : std_logic_vector(31 downto 0);
    signal clock_valid_137 : std_logic_vector(0 downto 0);
    signal konst_131_wire_constant : std_logic_vector(0 downto 0);
    signal konst_192_wire_constant : std_logic_vector(0 downto 0);
    signal slice_147_wire : std_logic_vector(15 downto 0);
    signal slice_155_wire : std_logic_vector(27 downto 0);
    signal slice_180_wire : std_logic_vector(15 downto 0);
    signal slice_187_wire : std_logic_vector(11 downto 0);
    signal type_cast_149_wire_constant : std_logic_vector(15 downto 0);
    signal type_cast_158_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_182_wire_constant : std_logic_vector(3 downto 0);
    -- 
  begin -- 
    konst_131_wire_constant <= "0";
    konst_192_wire_constant <= "1";
    type_cast_149_wire_constant <= "0000000000000000";
    type_cast_158_wire_constant <= "0000";
    type_cast_182_wire_constant <= "0000";
    -- flow-through slice operator slice_147_inst
    slice_147_wire <= RPIPE_CLK_FREQUENCY_SIG_145_wire(31 downto 16);
    -- flow-through slice operator slice_155_inst
    slice_155_wire <= RPIPE_BAUD_RATE_SIG_153_wire(27 downto 0);
    -- flow-through slice operator slice_180_inst
    slice_180_wire <= BL_177(15 downto 0);
    -- flow-through slice operator slice_187_inst
    slice_187_wire <= BF_168(11 downto 0);
    W_clock_valid_135_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_clock_valid_135_inst_req_0;
      W_clock_valid_135_inst_ack_0<= wack(0);
      rreq(0) <= W_clock_valid_135_inst_req_1;
      W_clock_valid_135_inst_ack_1<= rack(0);
      W_clock_valid_135_inst : InterlockBuffer generic map ( -- 
        name => "W_clock_valid_135_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => RPIPE_CLOCK_FREQUENCY_VALID_136_wire,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => clock_valid_137,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    if_stmt_138_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_140_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_138_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_138_branch_req_0,
          ack0 => if_stmt_138_branch_ack_0,
          ack1 => if_stmt_138_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- flow through binary operator CONCAT_u16_u20_183_inst
    process(slice_180_wire) -- 
      variable tmp_var : std_logic_vector(19 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_180_wire, type_cast_182_wire_constant, tmp_var);
      CONCAT_u16_u20_183_wire <= tmp_var; --
    end process;
    -- shared split operator group (1) : CONCAT_u16_u32_150_inst 
    ApConcat_group_1: Block -- 
      signal data_in: std_logic_vector(15 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= slice_147_wire;
      SS_151 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u16_u32_150_inst_req_0;
      CONCAT_u16_u32_150_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u16_u32_150_inst_req_1;
      CONCAT_u16_u32_150_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_1_gI: SplitGuardInterface generic map(name => "ApConcat_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0000000000000000",
          constant_width => 16,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- shared split operator group (2) : CONCAT_u20_u32_188_inst 
    ApConcat_group_2: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u16_u20_183_wire & slice_187_wire;
      CONCAT_u20_u32_188_wire <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u20_u32_188_inst_req_0;
      CONCAT_u20_u32_188_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u20_u32_188_inst_req_1;
      CONCAT_u20_u32_188_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_2_gI: SplitGuardInterface generic map(name => "ApConcat_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_2",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 20,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 12, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 2
    -- shared split operator group (3) : CONCAT_u28_u32_159_inst 
    ApConcat_group_3: Block -- 
      signal data_in: std_logic_vector(27 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= slice_155_wire;
      BRx16_160 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u28_u32_159_inst_req_0;
      CONCAT_u28_u32_159_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u28_u32_159_inst_req_1;
      CONCAT_u28_u32_159_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_3_gI: SplitGuardInterface generic map(name => "ApConcat_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 28,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0000",
          constant_width => 4,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- unary operator NOT_u1_u1_140_inst
    process(clock_valid_137) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", clock_valid_137, tmp_var);
      NOT_u1_u1_140_wire <= tmp_var; -- 
    end process;
    -- shared split operator group (5) : SUB_u32_u32_176_inst 
    ApIntSub_group_5: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= BLx_172 & BF_168;
      BL_177 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u32_u32_176_inst_req_0;
      SUB_u32_u32_176_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u32_u32_176_inst_req_1;
      SUB_u32_u32_176_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_5_gI: SplitGuardInterface generic map(name => "ApIntSub_group_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_5",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 32, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- read from input-signal BAUD_RATE_SIG
    RPIPE_BAUD_RATE_SIG_153_wire <= BAUD_RATE_SIG;
    -- read from input-signal CLK_FREQUENCY_SIG
    RPIPE_CLK_FREQUENCY_SIG_145_wire <= CLK_FREQUENCY_SIG;
    -- read from input-signal CLOCK_FREQUENCY_VALID
    RPIPE_CLOCK_FREQUENCY_VALID_136_wire <= CLOCK_FREQUENCY_VALID;
    -- shared outport operator group (0) : WPIPE_BAUD_CONTROL_WORD_SIG_178_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_BAUD_CONTROL_WORD_SIG_178_inst_req_0;
      WPIPE_BAUD_CONTROL_WORD_SIG_178_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_BAUD_CONTROL_WORD_SIG_178_inst_req_1;
      WPIPE_BAUD_CONTROL_WORD_SIG_178_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= CONCAT_u20_u32_188_wire;
      BAUD_CONTROL_WORD_SIG_write_0_gI: SplitGuardInterface generic map(name => "BAUD_CONTROL_WORD_SIG_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      BAUD_CONTROL_WORD_SIG_write_0: OutputPortRevised -- 
        generic map ( name => "BAUD_CONTROL_WORD_SIG", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => BAUD_CONTROL_WORD_SIG_pipe_write_req(0),
          oack => BAUD_CONTROL_WORD_SIG_pipe_write_ack(0),
          odata => BAUD_CONTROL_WORD_SIG_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_BAUD_CONTROL_WORD_VALID_130_inst WPIPE_BAUD_CONTROL_WORD_VALID_191_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal sample_req, sample_ack : BooleanArray( 1 downto 0);
      signal update_req, update_ack : BooleanArray( 1 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 1 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 0, 0 => 0);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      sample_req_unguarded(1) <= WPIPE_BAUD_CONTROL_WORD_VALID_130_inst_req_0;
      sample_req_unguarded(0) <= WPIPE_BAUD_CONTROL_WORD_VALID_191_inst_req_0;
      WPIPE_BAUD_CONTROL_WORD_VALID_130_inst_ack_0 <= sample_ack_unguarded(1);
      WPIPE_BAUD_CONTROL_WORD_VALID_191_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(1) <= WPIPE_BAUD_CONTROL_WORD_VALID_130_inst_req_1;
      update_req_unguarded(0) <= WPIPE_BAUD_CONTROL_WORD_VALID_191_inst_req_1;
      WPIPE_BAUD_CONTROL_WORD_VALID_130_inst_ack_1 <= update_ack_unguarded(1);
      WPIPE_BAUD_CONTROL_WORD_VALID_191_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      data_in <= konst_131_wire_constant & konst_192_wire_constant;
      BAUD_CONTROL_WORD_VALID_write_1_gI: SplitGuardInterface generic map(name => "BAUD_CONTROL_WORD_VALID_write_1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      BAUD_CONTROL_WORD_VALID_write_1: OutputPortRevised -- 
        generic map ( name => "BAUD_CONTROL_WORD_VALID", data_width => 1, num_reqs => 2, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => BAUD_CONTROL_WORD_VALID_pipe_write_req(0),
          oack => BAUD_CONTROL_WORD_VALID_pipe_write_ack(0),
          odata => BAUD_CONTROL_WORD_VALID_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_164_call 
    my_gcd_call_group_0: Block -- 
      signal data_in: std_logic_vector(63 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_164_call_req_0;
      call_stmt_164_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_164_call_req_1;
      call_stmt_164_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      my_gcd_call_group_0_gI: SplitGuardInterface generic map(name => "my_gcd_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= SS_151 & BRx16_160;
      GCD_164 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 64,
        owidth => 64,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => my_gcd_call_reqs(0),
          ackR => my_gcd_call_acks(0),
          dataR => my_gcd_call_data(63 downto 0),
          tagR => my_gcd_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => my_gcd_return_acks(0), -- cross-over
          ackL => my_gcd_return_reqs(0), -- cross-over
          dataL => my_gcd_return_data(31 downto 0),
          tagL => my_gcd_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_168_call call_stmt_172_call 
    my_div_call_group_1: Block -- 
      signal data_in: std_logic_vector(127 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_168_call_req_0;
      reqL_unguarded(0) <= call_stmt_172_call_req_0;
      call_stmt_168_call_ack_0 <= ackL_unguarded(1);
      call_stmt_172_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_168_call_req_1;
      reqR_unguarded(0) <= call_stmt_172_call_req_1;
      call_stmt_168_call_ack_1 <= ackR_unguarded(1);
      call_stmt_172_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      my_div_call_group_1_accessRegulator_0: access_regulator_base generic map (name => "my_div_call_group_1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      my_div_call_group_1_accessRegulator_1: access_regulator_base generic map (name => "my_div_call_group_1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      my_div_call_group_1_gI: SplitGuardInterface generic map(name => "my_div_call_group_1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= BRx16_160 & GCD_164 & SS_151 & GCD_164;
      BF_168 <= data_out(63 downto 32);
      BLx_172 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 128,
        owidth => 64,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => my_div_call_reqs(0),
          ackR => my_div_call_acks(0),
          dataR => my_div_call_data(63 downto 0),
          tagR => my_div_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => my_div_return_acks(0), -- cross-over
          ackL => my_div_return_reqs(0), -- cross-over
          dataL => my_div_return_data(31 downto 0),
          tagL => my_div_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end baudControlCalculatorDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library AjitCustom;
use AjitCustom.baud_control_calculator_global_package.all;
entity my_div is -- 
  generic (tag_length : integer); 
  port ( -- 
    A : in  std_logic_vector(31 downto 0);
    B : in  std_logic_vector(31 downto 0);
    Q : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity my_div;
architecture my_div_arch of my_div is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal A_buffer :  std_logic_vector(31 downto 0);
  signal A_update_enable: Boolean;
  signal B_buffer :  std_logic_vector(31 downto 0);
  signal B_update_enable: Boolean;
  -- output port buffer signals
  signal Q_buffer :  std_logic_vector(31 downto 0);
  signal Q_update_enable: Boolean;
  signal my_div_CP_159_start: Boolean;
  signal my_div_CP_159_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal phi_stmt_85_ack_0 : boolean;
  signal phi_stmt_89_ack_0 : boolean;
  signal W_Q_125_inst_req_0 : boolean;
  signal if_stmt_120_branch_req_0 : boolean;
  signal if_stmt_120_branch_ack_1 : boolean;
  signal if_stmt_120_branch_ack_0 : boolean;
  signal A_87_buf_req_0 : boolean;
  signal A_87_buf_ack_0 : boolean;
  signal A_87_buf_req_1 : boolean;
  signal A_87_buf_ack_1 : boolean;
  signal phi_stmt_85_req_0 : boolean;
  signal phi_stmt_89_req_0 : boolean;
  signal ntA_111_88_buf_req_0 : boolean;
  signal ntA_111_88_buf_ack_0 : boolean;
  signal ntA_111_88_buf_req_1 : boolean;
  signal ntA_111_88_buf_ack_1 : boolean;
  signal phi_stmt_85_req_1 : boolean;
  signal ntQ_119_93_buf_req_0 : boolean;
  signal ntQ_119_93_buf_ack_0 : boolean;
  signal ntQ_119_93_buf_req_1 : boolean;
  signal ntQ_119_93_buf_ack_1 : boolean;
  signal phi_stmt_89_req_1 : boolean;
  signal W_Q_125_inst_ack_0 : boolean;
  signal W_Q_125_inst_req_1 : boolean;
  signal W_Q_125_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "my_div_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 64) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= A;
  A_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(63 downto 32) <= B;
  B_buffer <= in_buffer_data_out(63 downto 32);
  in_buffer_data_in(tag_length + 63 downto 64) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 63 downto 64);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  my_div_CP_159_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "my_div_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= Q_buffer;
  Q <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= my_div_CP_159_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= my_div_CP_159_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= my_div_CP_159_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  my_div_CP_159: Block -- control-path 
    signal my_div_CP_159_elements: BooleanArray(22 downto 0);
    -- 
  begin -- 
    my_div_CP_159_elements(0) <= my_div_CP_159_start;
    my_div_CP_159_symbol <= my_div_CP_159_elements(22);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_83/$entry
      -- CP-element group 0: 	 branch_block_stmt_83/branch_block_stmt_83__entry__
      -- CP-element group 0: 	 branch_block_stmt_83/merge_stmt_84__entry__
      -- CP-element group 0: 	 branch_block_stmt_83/merge_stmt_84_dead_link/$entry
      -- 
    -- CP-element group 1:  merge  branch  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	20 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1: 	3 
    -- CP-element group 1:  members (13) 
      -- CP-element group 1: 	 branch_block_stmt_83/merge_stmt_84__exit__
      -- CP-element group 1: 	 branch_block_stmt_83/assign_stmt_103_to_assign_stmt_119__entry__
      -- CP-element group 1: 	 branch_block_stmt_83/assign_stmt_103_to_assign_stmt_119__exit__
      -- CP-element group 1: 	 branch_block_stmt_83/if_stmt_120__entry__
      -- CP-element group 1: 	 branch_block_stmt_83/assign_stmt_103_to_assign_stmt_119/$entry
      -- CP-element group 1: 	 branch_block_stmt_83/assign_stmt_103_to_assign_stmt_119/$exit
      -- CP-element group 1: 	 branch_block_stmt_83/if_stmt_120_dead_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_83/if_stmt_120_eval_test/$entry
      -- CP-element group 1: 	 branch_block_stmt_83/if_stmt_120_eval_test/$exit
      -- CP-element group 1: 	 branch_block_stmt_83/if_stmt_120_eval_test/branch_req
      -- CP-element group 1: 	 branch_block_stmt_83/R_continue_flag_121_place
      -- CP-element group 1: 	 branch_block_stmt_83/if_stmt_120_if_link/$entry
      -- CP-element group 1: 	 branch_block_stmt_83/if_stmt_120_else_link/$entry
      -- 
    branch_req_183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_div_CP_159_elements(1), ack => if_stmt_120_branch_req_0); -- 
    my_div_CP_159_elements(1) <= my_div_CP_159_elements(20);
    -- CP-element group 2:  fork  transition  place  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	10 
    -- CP-element group 2: 	14 
    -- CP-element group 2: 	13 
    -- CP-element group 2: 	11 
    -- CP-element group 2:  members (18) 
      -- CP-element group 2: 	 branch_block_stmt_83/if_stmt_120_if_link/$exit
      -- CP-element group 2: 	 branch_block_stmt_83/if_stmt_120_if_link/if_choice_transition
      -- CP-element group 2: 	 branch_block_stmt_83/loopback
      -- CP-element group 2: 	 branch_block_stmt_83/loopback_PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_83/loopback_PhiReq/phi_stmt_85/$entry
      -- CP-element group 2: 	 branch_block_stmt_83/loopback_PhiReq/phi_stmt_85/phi_stmt_85_sources/$entry
      -- CP-element group 2: 	 branch_block_stmt_83/loopback_PhiReq/phi_stmt_85/phi_stmt_85_sources/Interlock/$entry
      -- CP-element group 2: 	 branch_block_stmt_83/loopback_PhiReq/phi_stmt_85/phi_stmt_85_sources/Interlock/Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_83/loopback_PhiReq/phi_stmt_85/phi_stmt_85_sources/Interlock/Sample/req
      -- CP-element group 2: 	 branch_block_stmt_83/loopback_PhiReq/phi_stmt_85/phi_stmt_85_sources/Interlock/Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_83/loopback_PhiReq/phi_stmt_85/phi_stmt_85_sources/Interlock/Update/req
      -- CP-element group 2: 	 branch_block_stmt_83/loopback_PhiReq/phi_stmt_89/$entry
      -- CP-element group 2: 	 branch_block_stmt_83/loopback_PhiReq/phi_stmt_89/phi_stmt_89_sources/$entry
      -- CP-element group 2: 	 branch_block_stmt_83/loopback_PhiReq/phi_stmt_89/phi_stmt_89_sources/Interlock/$entry
      -- CP-element group 2: 	 branch_block_stmt_83/loopback_PhiReq/phi_stmt_89/phi_stmt_89_sources/Interlock/Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_83/loopback_PhiReq/phi_stmt_89/phi_stmt_89_sources/Interlock/Sample/req
      -- CP-element group 2: 	 branch_block_stmt_83/loopback_PhiReq/phi_stmt_89/phi_stmt_89_sources/Interlock/Update/$entry
      -- CP-element group 2: 	 branch_block_stmt_83/loopback_PhiReq/phi_stmt_89/phi_stmt_89_sources/Interlock/Update/req
      -- 
    if_choice_transition_188_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_120_branch_ack_1, ack => my_div_CP_159_elements(2)); -- 
    req_244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_div_CP_159_elements(2), ack => ntA_111_88_buf_req_0); -- 
    req_249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_div_CP_159_elements(2), ack => ntA_111_88_buf_req_1); -- 
    req_264_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_264_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_div_CP_159_elements(2), ack => ntQ_119_93_buf_req_0); -- 
    req_269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_div_CP_159_elements(2), ack => ntQ_119_93_buf_req_1); -- 
    -- CP-element group 3:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	1 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	22 
    -- CP-element group 3: 	21 
    -- CP-element group 3:  members (12) 
      -- CP-element group 3: 	 assign_stmt_127/$entry
      -- CP-element group 3: 	 assign_stmt_127/assign_stmt_127_sample_start_
      -- CP-element group 3: 	 assign_stmt_127/assign_stmt_127_update_start_
      -- CP-element group 3: 	 assign_stmt_127/assign_stmt_127_Sample/$entry
      -- CP-element group 3: 	 assign_stmt_127/assign_stmt_127_Sample/req
      -- CP-element group 3: 	 branch_block_stmt_83/$exit
      -- CP-element group 3: 	 branch_block_stmt_83/branch_block_stmt_83__exit__
      -- CP-element group 3: 	 branch_block_stmt_83/if_stmt_120__exit__
      -- CP-element group 3: 	 branch_block_stmt_83/if_stmt_120_else_link/$exit
      -- CP-element group 3: 	 branch_block_stmt_83/if_stmt_120_else_link/else_choice_transition
      -- CP-element group 3: 	 assign_stmt_127/assign_stmt_127_Update/$entry
      -- CP-element group 3: 	 assign_stmt_127/assign_stmt_127_Update/req
      -- 
    else_choice_transition_192_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_120_branch_ack_0, ack => my_div_CP_159_elements(3)); -- 
    req_288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_div_CP_159_elements(3), ack => W_Q_125_inst_req_0); -- 
    req_293_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_293_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_div_CP_159_elements(3), ack => W_Q_125_inst_req_1); -- 
    -- CP-element group 4:  fork  transition  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4: 	8 
    -- CP-element group 4: 	6 
    -- CP-element group 4:  members (10) 
      -- CP-element group 4: 	 branch_block_stmt_83/merge_stmt_84__entry___PhiReq/$entry
      -- CP-element group 4: 	 branch_block_stmt_83/merge_stmt_84__entry___PhiReq/phi_stmt_85/$entry
      -- CP-element group 4: 	 branch_block_stmt_83/merge_stmt_84__entry___PhiReq/phi_stmt_85/phi_stmt_85_sources/$entry
      -- CP-element group 4: 	 branch_block_stmt_83/merge_stmt_84__entry___PhiReq/phi_stmt_85/phi_stmt_85_sources/Interlock/$entry
      -- CP-element group 4: 	 branch_block_stmt_83/merge_stmt_84__entry___PhiReq/phi_stmt_85/phi_stmt_85_sources/Interlock/Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_83/merge_stmt_84__entry___PhiReq/phi_stmt_85/phi_stmt_85_sources/Interlock/Sample/req
      -- CP-element group 4: 	 branch_block_stmt_83/merge_stmt_84__entry___PhiReq/phi_stmt_85/phi_stmt_85_sources/Interlock/Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_83/merge_stmt_84__entry___PhiReq/phi_stmt_85/phi_stmt_85_sources/Interlock/Update/req
      -- CP-element group 4: 	 branch_block_stmt_83/merge_stmt_84__entry___PhiReq/phi_stmt_89/$entry
      -- CP-element group 4: 	 branch_block_stmt_83/merge_stmt_84__entry___PhiReq/phi_stmt_89/phi_stmt_89_sources/$entry
      -- 
    req_213_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_213_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_div_CP_159_elements(4), ack => A_87_buf_req_0); -- 
    req_218_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_218_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_div_CP_159_elements(4), ack => A_87_buf_req_1); -- 
    my_div_CP_159_elements(4) <= my_div_CP_159_elements(0);
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	7 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 branch_block_stmt_83/merge_stmt_84__entry___PhiReq/phi_stmt_85/phi_stmt_85_sources/Interlock/Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_83/merge_stmt_84__entry___PhiReq/phi_stmt_85/phi_stmt_85_sources/Interlock/Sample/ack
      -- 
    ack_214_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => A_87_buf_ack_0, ack => my_div_CP_159_elements(5)); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	4 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 branch_block_stmt_83/merge_stmt_84__entry___PhiReq/phi_stmt_85/phi_stmt_85_sources/Interlock/Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_83/merge_stmt_84__entry___PhiReq/phi_stmt_85/phi_stmt_85_sources/Interlock/Update/ack
      -- 
    ack_219_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => A_87_buf_ack_1, ack => my_div_CP_159_elements(6)); -- 
    -- CP-element group 7:  join  transition  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	5 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	9 
    -- CP-element group 7:  members (4) 
      -- CP-element group 7: 	 branch_block_stmt_83/merge_stmt_84__entry___PhiReq/phi_stmt_85/$exit
      -- CP-element group 7: 	 branch_block_stmt_83/merge_stmt_84__entry___PhiReq/phi_stmt_85/phi_stmt_85_sources/$exit
      -- CP-element group 7: 	 branch_block_stmt_83/merge_stmt_84__entry___PhiReq/phi_stmt_85/phi_stmt_85_sources/Interlock/$exit
      -- CP-element group 7: 	 branch_block_stmt_83/merge_stmt_84__entry___PhiReq/phi_stmt_85/phi_stmt_85_req
      -- 
    phi_stmt_85_req_220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_85_req_220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_div_CP_159_elements(7), ack => phi_stmt_85_req_0); -- 
    my_div_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "my_div_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= my_div_CP_159_elements(5) & my_div_CP_159_elements(6);
      gj_my_div_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => my_div_CP_159_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  transition  output  delay-element  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	4 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (4) 
      -- CP-element group 8: 	 branch_block_stmt_83/merge_stmt_84__entry___PhiReq/phi_stmt_89/$exit
      -- CP-element group 8: 	 branch_block_stmt_83/merge_stmt_84__entry___PhiReq/phi_stmt_89/phi_stmt_89_sources/$exit
      -- CP-element group 8: 	 branch_block_stmt_83/merge_stmt_84__entry___PhiReq/phi_stmt_89/phi_stmt_89_sources/type_cast_92_konst_delay_trans
      -- CP-element group 8: 	 branch_block_stmt_83/merge_stmt_84__entry___PhiReq/phi_stmt_89/phi_stmt_89_req
      -- 
    phi_stmt_89_req_228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_89_req_228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_div_CP_159_elements(8), ack => phi_stmt_89_req_0); -- 
    -- Element group my_div_CP_159_elements(8) is a control-delay.
    cp_element_8_delay: control_delay_element  generic map(name => " 8_delay", delay_value => 1)  port map(req => my_div_CP_159_elements(4), ack => my_div_CP_159_elements(8), clk => clk, reset =>reset);
    -- CP-element group 9:  join  transition  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: 	7 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	17 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_83/merge_stmt_84__entry___PhiReq/$exit
      -- 
    my_div_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "my_div_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= my_div_CP_159_elements(8) & my_div_CP_159_elements(7);
      gj_my_div_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => my_div_CP_159_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	2 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (2) 
      -- CP-element group 10: 	 branch_block_stmt_83/loopback_PhiReq/phi_stmt_85/phi_stmt_85_sources/Interlock/Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_83/loopback_PhiReq/phi_stmt_85/phi_stmt_85_sources/Interlock/Sample/ack
      -- 
    ack_245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ntA_111_88_buf_ack_0, ack => my_div_CP_159_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	2 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_83/loopback_PhiReq/phi_stmt_85/phi_stmt_85_sources/Interlock/Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_83/loopback_PhiReq/phi_stmt_85/phi_stmt_85_sources/Interlock/Update/ack
      -- 
    ack_250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ntA_111_88_buf_ack_1, ack => my_div_CP_159_elements(11)); -- 
    -- CP-element group 12:  join  transition  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	16 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 branch_block_stmt_83/loopback_PhiReq/phi_stmt_85/$exit
      -- CP-element group 12: 	 branch_block_stmt_83/loopback_PhiReq/phi_stmt_85/phi_stmt_85_sources/$exit
      -- CP-element group 12: 	 branch_block_stmt_83/loopback_PhiReq/phi_stmt_85/phi_stmt_85_sources/Interlock/$exit
      -- CP-element group 12: 	 branch_block_stmt_83/loopback_PhiReq/phi_stmt_85/phi_stmt_85_req
      -- 
    phi_stmt_85_req_251_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_85_req_251_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_div_CP_159_elements(12), ack => phi_stmt_85_req_1); -- 
    my_div_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "my_div_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= my_div_CP_159_elements(10) & my_div_CP_159_elements(11);
      gj_my_div_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => my_div_CP_159_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	15 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_83/loopback_PhiReq/phi_stmt_89/phi_stmt_89_sources/Interlock/Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_83/loopback_PhiReq/phi_stmt_89/phi_stmt_89_sources/Interlock/Sample/ack
      -- 
    ack_265_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ntQ_119_93_buf_ack_0, ack => my_div_CP_159_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	2 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_83/loopback_PhiReq/phi_stmt_89/phi_stmt_89_sources/Interlock/Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_83/loopback_PhiReq/phi_stmt_89/phi_stmt_89_sources/Interlock/Update/ack
      -- 
    ack_270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ntQ_119_93_buf_ack_1, ack => my_div_CP_159_elements(14)); -- 
    -- CP-element group 15:  join  transition  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: 	13 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (4) 
      -- CP-element group 15: 	 branch_block_stmt_83/loopback_PhiReq/phi_stmt_89/$exit
      -- CP-element group 15: 	 branch_block_stmt_83/loopback_PhiReq/phi_stmt_89/phi_stmt_89_sources/$exit
      -- CP-element group 15: 	 branch_block_stmt_83/loopback_PhiReq/phi_stmt_89/phi_stmt_89_sources/Interlock/$exit
      -- CP-element group 15: 	 branch_block_stmt_83/loopback_PhiReq/phi_stmt_89/phi_stmt_89_req
      -- 
    phi_stmt_89_req_271_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_89_req_271_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_div_CP_159_elements(15), ack => phi_stmt_89_req_1); -- 
    my_div_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "my_div_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= my_div_CP_159_elements(14) & my_div_CP_159_elements(13);
      gj_my_div_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => my_div_CP_159_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	12 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_83/loopback_PhiReq/$exit
      -- 
    my_div_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "my_div_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= my_div_CP_159_elements(12) & my_div_CP_159_elements(15);
      gj_my_div_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => my_div_CP_159_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  merge  fork  transition  place  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	16 
    -- CP-element group 17: 	9 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	19 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_83/merge_stmt_84_PhiReqMerge
      -- CP-element group 17: 	 branch_block_stmt_83/merge_stmt_84_PhiAck/$entry
      -- 
    my_div_CP_159_elements(17) <= OrReduce(my_div_CP_159_elements(16) & my_div_CP_159_elements(9));
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	20 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_83/merge_stmt_84_PhiAck/phi_stmt_85_ack
      -- 
    phi_stmt_85_ack_276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_85_ack_0, ack => my_div_CP_159_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_83/merge_stmt_84_PhiAck/phi_stmt_89_ack
      -- 
    phi_stmt_89_ack_277_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_89_ack_0, ack => my_div_CP_159_elements(19)); -- 
    -- CP-element group 20:  join  transition  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: 	18 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	1 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_83/merge_stmt_84_PhiAck/$exit
      -- 
    my_div_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "my_div_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= my_div_CP_159_elements(19) & my_div_CP_159_elements(18);
      gj_my_div_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => my_div_CP_159_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	3 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 assign_stmt_127/assign_stmt_127_sample_completed_
      -- CP-element group 21: 	 assign_stmt_127/assign_stmt_127_Sample/$exit
      -- CP-element group 21: 	 assign_stmt_127/assign_stmt_127_Sample/ack
      -- 
    ack_289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_Q_125_inst_ack_0, ack => my_div_CP_159_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	3 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (5) 
      -- CP-element group 22: 	 assign_stmt_127/$exit
      -- CP-element group 22: 	 assign_stmt_127/assign_stmt_127_update_completed_
      -- CP-element group 22: 	 $exit
      -- CP-element group 22: 	 assign_stmt_127/assign_stmt_127_Update/$exit
      -- CP-element group 22: 	 assign_stmt_127/assign_stmt_127_Update/ack
      -- 
    ack_294_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_Q_125_inst_ack_1, ack => my_div_CP_159_elements(22)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_116_wire : std_logic_vector(31 downto 0);
    signal A_87_buffered : std_logic_vector(31 downto 0);
    signal NEQ_u32_u1_98_wire : std_logic_vector(0 downto 0);
    signal SUB_u32_u32_108_wire : std_logic_vector(31 downto 0);
    signal UGE_u32_u1_101_wire : std_logic_vector(0 downto 0);
    signal continue_flag_103 : std_logic_vector(0 downto 0);
    signal konst_115_wire_constant : std_logic_vector(31 downto 0);
    signal konst_97_wire_constant : std_logic_vector(31 downto 0);
    signal ntA_111 : std_logic_vector(31 downto 0);
    signal ntA_111_88_buffered : std_logic_vector(31 downto 0);
    signal ntQ_119 : std_logic_vector(31 downto 0);
    signal ntQ_119_93_buffered : std_logic_vector(31 downto 0);
    signal tA_85 : std_logic_vector(31 downto 0);
    signal tQ_89 : std_logic_vector(31 downto 0);
    signal type_cast_92_wire_constant : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    konst_115_wire_constant <= "00000000000000000000000000000001";
    konst_97_wire_constant <= "00000000000000000000000000000000";
    type_cast_92_wire_constant <= "00000000000000000000000000000000";
    phi_stmt_85: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= A_87_buffered & ntA_111_88_buffered;
      req <= phi_stmt_85_req_0 & phi_stmt_85_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_85",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_85_ack_0,
          idata => idata,
          odata => tA_85,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_85
    phi_stmt_89: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_92_wire_constant & ntQ_119_93_buffered;
      req <= phi_stmt_89_req_0 & phi_stmt_89_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_89",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_89_ack_0,
          idata => idata,
          odata => tQ_89,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_89
    -- flow-through select operator MUX_110_inst
    ntA_111 <= SUB_u32_u32_108_wire when (continue_flag_103(0) /=  '0') else tA_85;
    -- flow-through select operator MUX_118_inst
    ntQ_119 <= ADD_u32_u32_116_wire when (continue_flag_103(0) /=  '0') else tQ_89;
    A_87_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= A_87_buf_req_0;
      A_87_buf_ack_0<= wack(0);
      rreq(0) <= A_87_buf_req_1;
      A_87_buf_ack_1<= rack(0);
      A_87_buf : InterlockBuffer generic map ( -- 
        name => "A_87_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => A_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => A_87_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_Q_125_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_Q_125_inst_req_0;
      W_Q_125_inst_ack_0<= wack(0);
      rreq(0) <= W_Q_125_inst_req_1;
      W_Q_125_inst_ack_1<= rack(0);
      W_Q_125_inst : InterlockBuffer generic map ( -- 
        name => "W_Q_125_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false ,
        in_phi =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tQ_89,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => Q_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    ntA_111_88_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= ntA_111_88_buf_req_0;
      ntA_111_88_buf_ack_0<= wack(0);
      rreq(0) <= ntA_111_88_buf_req_1;
      ntA_111_88_buf_ack_1<= rack(0);
      ntA_111_88_buf : InterlockBuffer generic map ( -- 
        name => "ntA_111_88_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ntA_111,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ntA_111_88_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    ntQ_119_93_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= ntQ_119_93_buf_req_0;
      ntQ_119_93_buf_ack_0<= wack(0);
      rreq(0) <= ntQ_119_93_buf_req_1;
      ntQ_119_93_buf_ack_1<= rack(0);
      ntQ_119_93_buf : InterlockBuffer generic map ( -- 
        name => "ntQ_119_93_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ntQ_119,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ntQ_119_93_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    if_stmt_120_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= continue_flag_103;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_120_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_120_branch_req_0,
          ack0 => if_stmt_120_branch_ack_0,
          ack1 => if_stmt_120_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- flow through binary operator ADD_u32_u32_116_inst
    ADD_u32_u32_116_wire <= std_logic_vector(unsigned(tQ_89) + unsigned(konst_115_wire_constant));
    -- flow through binary operator AND_u1_u1_102_inst
    continue_flag_103 <= (NEQ_u32_u1_98_wire and UGE_u32_u1_101_wire);
    -- flow through binary operator NEQ_u32_u1_98_inst
    process(tA_85) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(tA_85, konst_97_wire_constant, tmp_var);
      NEQ_u32_u1_98_wire <= tmp_var; --
    end process;
    -- flow through binary operator SUB_u32_u32_108_inst
    SUB_u32_u32_108_wire <= std_logic_vector(unsigned(tA_85) - unsigned(B_buffer));
    -- flow through binary operator UGE_u32_u1_101_inst
    process(tA_85, B_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUge_proc(tA_85, B_buffer, tmp_var);
      UGE_u32_u1_101_wire <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end my_div_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library AjitCustom;
use AjitCustom.baud_control_calculator_global_package.all;
entity my_gcd is -- 
  generic (tag_length : integer); 
  port ( -- 
    A : in  std_logic_vector(31 downto 0);
    B : in  std_logic_vector(31 downto 0);
    GCD : out  std_logic_vector(31 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity my_gcd;
architecture my_gcd_arch of my_gcd is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal A_buffer :  std_logic_vector(31 downto 0);
  signal A_update_enable: Boolean;
  signal B_buffer :  std_logic_vector(31 downto 0);
  signal B_update_enable: Boolean;
  -- output port buffer signals
  signal GCD_buffer :  std_logic_vector(31 downto 0);
  signal GCD_update_enable: Boolean;
  signal my_gcd_CP_0_start: Boolean;
  signal my_gcd_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal AND_u1_u1_33_inst_req_0 : boolean;
  signal MUX_51_inst_req_0 : boolean;
  signal MUX_51_inst_ack_0 : boolean;
  signal MUX_51_inst_req_1 : boolean;
  signal MUX_51_inst_ack_1 : boolean;
  signal AND_u1_u1_33_inst_ack_0 : boolean;
  signal AND_u1_u1_33_inst_req_1 : boolean;
  signal AND_u1_u1_33_inst_ack_1 : boolean;
  signal ntA_62_16_buf_req_0 : boolean;
  signal ntA_62_16_buf_ack_0 : boolean;
  signal if_stmt_73_branch_req_0 : boolean;
  signal if_stmt_73_branch_ack_1 : boolean;
  signal if_stmt_73_branch_ack_0 : boolean;
  signal A_15_buf_req_0 : boolean;
  signal A_15_buf_ack_0 : boolean;
  signal A_15_buf_req_1 : boolean;
  signal A_15_buf_ack_1 : boolean;
  signal phi_stmt_13_req_0 : boolean;
  signal B_19_buf_req_0 : boolean;
  signal B_19_buf_ack_0 : boolean;
  signal B_19_buf_req_1 : boolean;
  signal B_19_buf_ack_1 : boolean;
  signal phi_stmt_17_req_0 : boolean;
  signal ntA_62_16_buf_req_1 : boolean;
  signal ntA_62_16_buf_ack_1 : boolean;
  signal phi_stmt_13_req_1 : boolean;
  signal ntB_72_20_buf_req_0 : boolean;
  signal ntB_72_20_buf_ack_0 : boolean;
  signal ntB_72_20_buf_req_1 : boolean;
  signal ntB_72_20_buf_ack_1 : boolean;
  signal phi_stmt_17_req_1 : boolean;
  signal phi_stmt_13_ack_0 : boolean;
  signal phi_stmt_17_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "my_gcd_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 64) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= A;
  A_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(63 downto 32) <= B;
  B_buffer <= in_buffer_data_out(63 downto 32);
  in_buffer_data_in(tag_length + 63 downto 64) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 63 downto 64);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  my_gcd_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "my_gcd_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= GCD_buffer;
  GCD <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= my_gcd_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= my_gcd_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= my_gcd_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  my_gcd_CP_0: Block -- control-path 
    signal my_gcd_CP_0_elements: BooleanArray(27 downto 0);
    -- 
  begin -- 
    my_gcd_CP_0_elements(0) <= my_gcd_CP_0_start;
    my_gcd_CP_0_symbol <= my_gcd_CP_0_elements(8);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	9 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_11/$entry
      -- CP-element group 0: 	 branch_block_stmt_11/branch_block_stmt_11__entry__
      -- CP-element group 0: 	 branch_block_stmt_11/merge_stmt_12__entry__
      -- CP-element group 0: 	 branch_block_stmt_11/merge_stmt_12_dead_link/$entry
      -- 
    -- CP-element group 1:  merge  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	27 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1: 	3 
    -- CP-element group 1: 	4 
    -- CP-element group 1: 	5 
    -- CP-element group 1:  members (15) 
      -- CP-element group 1: 	 branch_block_stmt_11/assign_stmt_34_to_assign_stmt_72/AND_u1_u1_33_update_start_
      -- CP-element group 1: 	 branch_block_stmt_11/assign_stmt_34_to_assign_stmt_72/AND_u1_u1_33_sample_start_
      -- CP-element group 1: 	 branch_block_stmt_11/assign_stmt_34_to_assign_stmt_72/AND_u1_u1_33_Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_11/assign_stmt_34_to_assign_stmt_72/AND_u1_u1_33_Sample/rr
      -- CP-element group 1: 	 branch_block_stmt_11/merge_stmt_12__exit__
      -- CP-element group 1: 	 branch_block_stmt_11/assign_stmt_34_to_assign_stmt_72__entry__
      -- CP-element group 1: 	 branch_block_stmt_11/assign_stmt_34_to_assign_stmt_72/$entry
      -- CP-element group 1: 	 branch_block_stmt_11/assign_stmt_34_to_assign_stmt_72/MUX_51_sample_start_
      -- CP-element group 1: 	 branch_block_stmt_11/assign_stmt_34_to_assign_stmt_72/MUX_51_update_start_
      -- CP-element group 1: 	 branch_block_stmt_11/assign_stmt_34_to_assign_stmt_72/MUX_51_start/$entry
      -- CP-element group 1: 	 branch_block_stmt_11/assign_stmt_34_to_assign_stmt_72/MUX_51_start/req
      -- CP-element group 1: 	 branch_block_stmt_11/assign_stmt_34_to_assign_stmt_72/MUX_51_complete/$entry
      -- CP-element group 1: 	 branch_block_stmt_11/assign_stmt_34_to_assign_stmt_72/MUX_51_complete/req
      -- CP-element group 1: 	 branch_block_stmt_11/assign_stmt_34_to_assign_stmt_72/AND_u1_u1_33_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_11/assign_stmt_34_to_assign_stmt_72/AND_u1_u1_33_Update/cr
      -- 
    rr_24_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_24_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_gcd_CP_0_elements(1), ack => AND_u1_u1_33_inst_req_0); -- 
    req_38_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_38_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_gcd_CP_0_elements(1), ack => MUX_51_inst_req_0); -- 
    req_43_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_43_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_gcd_CP_0_elements(1), ack => MUX_51_inst_req_1); -- 
    cr_29_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_29_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_gcd_CP_0_elements(1), ack => AND_u1_u1_33_inst_req_1); -- 
    my_gcd_CP_0_elements(1) <= my_gcd_CP_0_elements(27);
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 branch_block_stmt_11/assign_stmt_34_to_assign_stmt_72/AND_u1_u1_33_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_11/assign_stmt_34_to_assign_stmt_72/AND_u1_u1_33_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_11/assign_stmt_34_to_assign_stmt_72/AND_u1_u1_33_Sample/ra
      -- 
    ra_25_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_33_inst_ack_0, ack => my_gcd_CP_0_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	1 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	6 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_11/assign_stmt_34_to_assign_stmt_72/AND_u1_u1_33_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_11/assign_stmt_34_to_assign_stmt_72/AND_u1_u1_33_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_11/assign_stmt_34_to_assign_stmt_72/AND_u1_u1_33_Update/ca
      -- 
    ca_30_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_33_inst_ack_1, ack => my_gcd_CP_0_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	1 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_11/assign_stmt_34_to_assign_stmt_72/MUX_51_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_11/assign_stmt_34_to_assign_stmt_72/MUX_51_start/$exit
      -- CP-element group 4: 	 branch_block_stmt_11/assign_stmt_34_to_assign_stmt_72/MUX_51_start/ack
      -- 
    ack_39_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_51_inst_ack_0, ack => my_gcd_CP_0_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	1 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_11/assign_stmt_34_to_assign_stmt_72/MUX_51_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_11/assign_stmt_34_to_assign_stmt_72/MUX_51_complete/$exit
      -- CP-element group 5: 	 branch_block_stmt_11/assign_stmt_34_to_assign_stmt_72/MUX_51_complete/ack
      -- 
    ack_44_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_51_inst_ack_1, ack => my_gcd_CP_0_elements(5)); -- 
    -- CP-element group 6:  branch  join  transition  place  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	3 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	8 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (10) 
      -- CP-element group 6: 	 branch_block_stmt_11/assign_stmt_34_to_assign_stmt_72__exit__
      -- CP-element group 6: 	 branch_block_stmt_11/if_stmt_73__entry__
      -- CP-element group 6: 	 branch_block_stmt_11/assign_stmt_34_to_assign_stmt_72/$exit
      -- CP-element group 6: 	 branch_block_stmt_11/if_stmt_73_dead_link/$entry
      -- CP-element group 6: 	 branch_block_stmt_11/if_stmt_73_eval_test/$entry
      -- CP-element group 6: 	 branch_block_stmt_11/if_stmt_73_eval_test/$exit
      -- CP-element group 6: 	 branch_block_stmt_11/if_stmt_73_eval_test/branch_req
      -- CP-element group 6: 	 branch_block_stmt_11/R_continue_flag_74_place
      -- CP-element group 6: 	 branch_block_stmt_11/if_stmt_73_if_link/$entry
      -- CP-element group 6: 	 branch_block_stmt_11/if_stmt_73_else_link/$entry
      -- 
    branch_req_52_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_52_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_gcd_CP_0_elements(6), ack => if_stmt_73_branch_req_0); -- 
    my_gcd_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 25) := "my_gcd_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= my_gcd_CP_0_elements(3) & my_gcd_CP_0_elements(5);
      gj_my_gcd_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => my_gcd_CP_0_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  fork  transition  place  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	20 
    -- CP-element group 7: 	18 
    -- CP-element group 7: 	17 
    -- CP-element group 7: 	21 
    -- CP-element group 7:  members (18) 
      -- CP-element group 7: 	 branch_block_stmt_11/loopback_PhiReq/phi_stmt_13/phi_stmt_13_sources/Interlock/Sample/req
      -- CP-element group 7: 	 branch_block_stmt_11/loopback_PhiReq/phi_stmt_13/phi_stmt_13_sources/Interlock/Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_11/if_stmt_73_if_link/$exit
      -- CP-element group 7: 	 branch_block_stmt_11/if_stmt_73_if_link/if_choice_transition
      -- CP-element group 7: 	 branch_block_stmt_11/loopback
      -- CP-element group 7: 	 branch_block_stmt_11/loopback_PhiReq/$entry
      -- CP-element group 7: 	 branch_block_stmt_11/loopback_PhiReq/phi_stmt_13/$entry
      -- CP-element group 7: 	 branch_block_stmt_11/loopback_PhiReq/phi_stmt_13/phi_stmt_13_sources/$entry
      -- CP-element group 7: 	 branch_block_stmt_11/loopback_PhiReq/phi_stmt_13/phi_stmt_13_sources/Interlock/$entry
      -- CP-element group 7: 	 branch_block_stmt_11/loopback_PhiReq/phi_stmt_13/phi_stmt_13_sources/Interlock/Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_11/loopback_PhiReq/phi_stmt_13/phi_stmt_13_sources/Interlock/Update/req
      -- CP-element group 7: 	 branch_block_stmt_11/loopback_PhiReq/phi_stmt_17/$entry
      -- CP-element group 7: 	 branch_block_stmt_11/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/$entry
      -- CP-element group 7: 	 branch_block_stmt_11/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/$entry
      -- CP-element group 7: 	 branch_block_stmt_11/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_11/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Sample/req
      -- CP-element group 7: 	 branch_block_stmt_11/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_11/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Update/req
      -- 
    if_choice_transition_57_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_73_branch_ack_1, ack => my_gcd_CP_0_elements(7)); -- 
    req_125_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_125_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_gcd_CP_0_elements(7), ack => ntA_62_16_buf_req_0); -- 
    req_130_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_130_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_gcd_CP_0_elements(7), ack => ntA_62_16_buf_req_1); -- 
    req_145_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_145_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_gcd_CP_0_elements(7), ack => ntB_72_20_buf_req_0); -- 
    req_150_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_150_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_gcd_CP_0_elements(7), ack => ntB_72_20_buf_req_1); -- 
    -- CP-element group 8:  merge  transition  place  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	6 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 $exit
      -- CP-element group 8: 	 branch_block_stmt_11/$exit
      -- CP-element group 8: 	 branch_block_stmt_11/branch_block_stmt_11__exit__
      -- CP-element group 8: 	 branch_block_stmt_11/if_stmt_73__exit__
      -- CP-element group 8: 	 branch_block_stmt_11/if_stmt_73_else_link/$exit
      -- CP-element group 8: 	 branch_block_stmt_11/if_stmt_73_else_link/else_choice_transition
      -- 
    else_choice_transition_61_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_73_branch_ack_0, ack => my_gcd_CP_0_elements(8)); -- 
    -- CP-element group 9:  fork  transition  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	0 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	10 
    -- CP-element group 9: 	14 
    -- CP-element group 9: 	13 
    -- CP-element group 9:  members (15) 
      -- CP-element group 9: 	 branch_block_stmt_11/merge_stmt_12__entry___PhiReq/$entry
      -- CP-element group 9: 	 branch_block_stmt_11/merge_stmt_12__entry___PhiReq/phi_stmt_13/$entry
      -- CP-element group 9: 	 branch_block_stmt_11/merge_stmt_12__entry___PhiReq/phi_stmt_13/phi_stmt_13_sources/$entry
      -- CP-element group 9: 	 branch_block_stmt_11/merge_stmt_12__entry___PhiReq/phi_stmt_13/phi_stmt_13_sources/Interlock/$entry
      -- CP-element group 9: 	 branch_block_stmt_11/merge_stmt_12__entry___PhiReq/phi_stmt_13/phi_stmt_13_sources/Interlock/Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_11/merge_stmt_12__entry___PhiReq/phi_stmt_13/phi_stmt_13_sources/Interlock/Sample/req
      -- CP-element group 9: 	 branch_block_stmt_11/merge_stmt_12__entry___PhiReq/phi_stmt_13/phi_stmt_13_sources/Interlock/Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_11/merge_stmt_12__entry___PhiReq/phi_stmt_13/phi_stmt_13_sources/Interlock/Update/req
      -- CP-element group 9: 	 branch_block_stmt_11/merge_stmt_12__entry___PhiReq/phi_stmt_17/$entry
      -- CP-element group 9: 	 branch_block_stmt_11/merge_stmt_12__entry___PhiReq/phi_stmt_17/phi_stmt_17_sources/$entry
      -- CP-element group 9: 	 branch_block_stmt_11/merge_stmt_12__entry___PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/$entry
      -- CP-element group 9: 	 branch_block_stmt_11/merge_stmt_12__entry___PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_11/merge_stmt_12__entry___PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Sample/req
      -- CP-element group 9: 	 branch_block_stmt_11/merge_stmt_12__entry___PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_11/merge_stmt_12__entry___PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Update/req
      -- 
    req_102_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_102_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_gcd_CP_0_elements(9), ack => B_19_buf_req_0); -- 
    req_107_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_107_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_gcd_CP_0_elements(9), ack => B_19_buf_req_1); -- 
    req_82_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_82_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_gcd_CP_0_elements(9), ack => A_15_buf_req_0); -- 
    req_87_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_87_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_gcd_CP_0_elements(9), ack => A_15_buf_req_1); -- 
    my_gcd_CP_0_elements(9) <= my_gcd_CP_0_elements(0);
    -- CP-element group 10:  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (2) 
      -- CP-element group 10: 	 branch_block_stmt_11/merge_stmt_12__entry___PhiReq/phi_stmt_13/phi_stmt_13_sources/Interlock/Sample/$exit
      -- CP-element group 10: 	 branch_block_stmt_11/merge_stmt_12__entry___PhiReq/phi_stmt_13/phi_stmt_13_sources/Interlock/Sample/ack
      -- 
    ack_83_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => A_15_buf_ack_0, ack => my_gcd_CP_0_elements(10)); -- 
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_11/merge_stmt_12__entry___PhiReq/phi_stmt_13/phi_stmt_13_sources/Interlock/Update/$exit
      -- CP-element group 11: 	 branch_block_stmt_11/merge_stmt_12__entry___PhiReq/phi_stmt_13/phi_stmt_13_sources/Interlock/Update/ack
      -- 
    ack_88_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => A_15_buf_ack_1, ack => my_gcd_CP_0_elements(11)); -- 
    -- CP-element group 12:  join  transition  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	16 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 branch_block_stmt_11/merge_stmt_12__entry___PhiReq/phi_stmt_13/$exit
      -- CP-element group 12: 	 branch_block_stmt_11/merge_stmt_12__entry___PhiReq/phi_stmt_13/phi_stmt_13_sources/$exit
      -- CP-element group 12: 	 branch_block_stmt_11/merge_stmt_12__entry___PhiReq/phi_stmt_13/phi_stmt_13_sources/Interlock/$exit
      -- CP-element group 12: 	 branch_block_stmt_11/merge_stmt_12__entry___PhiReq/phi_stmt_13/phi_stmt_13_req
      -- 
    phi_stmt_13_req_89_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_13_req_89_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_gcd_CP_0_elements(12), ack => phi_stmt_13_req_0); -- 
    my_gcd_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "my_gcd_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= my_gcd_CP_0_elements(11) & my_gcd_CP_0_elements(10);
      gj_my_gcd_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => my_gcd_CP_0_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	15 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_11/merge_stmt_12__entry___PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Sample/$exit
      -- CP-element group 13: 	 branch_block_stmt_11/merge_stmt_12__entry___PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Sample/ack
      -- 
    ack_103_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => B_19_buf_ack_0, ack => my_gcd_CP_0_elements(13)); -- 
    -- CP-element group 14:  transition  input  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	9 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_11/merge_stmt_12__entry___PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_11/merge_stmt_12__entry___PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Update/ack
      -- 
    ack_108_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => B_19_buf_ack_1, ack => my_gcd_CP_0_elements(14)); -- 
    -- CP-element group 15:  join  transition  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: 	13 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (4) 
      -- CP-element group 15: 	 branch_block_stmt_11/merge_stmt_12__entry___PhiReq/phi_stmt_17/$exit
      -- CP-element group 15: 	 branch_block_stmt_11/merge_stmt_12__entry___PhiReq/phi_stmt_17/phi_stmt_17_sources/$exit
      -- CP-element group 15: 	 branch_block_stmt_11/merge_stmt_12__entry___PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/$exit
      -- CP-element group 15: 	 branch_block_stmt_11/merge_stmt_12__entry___PhiReq/phi_stmt_17/phi_stmt_17_req
      -- 
    phi_stmt_17_req_109_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_17_req_109_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_gcd_CP_0_elements(15), ack => phi_stmt_17_req_0); -- 
    my_gcd_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "my_gcd_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= my_gcd_CP_0_elements(14) & my_gcd_CP_0_elements(13);
      gj_my_gcd_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => my_gcd_CP_0_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	12 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	24 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_11/merge_stmt_12__entry___PhiReq/$exit
      -- 
    my_gcd_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "my_gcd_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= my_gcd_CP_0_elements(12) & my_gcd_CP_0_elements(15);
      gj_my_gcd_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => my_gcd_CP_0_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  transition  input  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	7 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	19 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_11/loopback_PhiReq/phi_stmt_13/phi_stmt_13_sources/Interlock/Sample/ack
      -- CP-element group 17: 	 branch_block_stmt_11/loopback_PhiReq/phi_stmt_13/phi_stmt_13_sources/Interlock/Sample/$exit
      -- 
    ack_126_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 17_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ntA_62_16_buf_ack_0, ack => my_gcd_CP_0_elements(17)); -- 
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	7 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	19 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_11/loopback_PhiReq/phi_stmt_13/phi_stmt_13_sources/Interlock/Update/$exit
      -- CP-element group 18: 	 branch_block_stmt_11/loopback_PhiReq/phi_stmt_13/phi_stmt_13_sources/Interlock/Update/ack
      -- 
    ack_131_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ntA_62_16_buf_ack_1, ack => my_gcd_CP_0_elements(18)); -- 
    -- CP-element group 19:  join  transition  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	18 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	23 
    -- CP-element group 19:  members (4) 
      -- CP-element group 19: 	 branch_block_stmt_11/loopback_PhiReq/phi_stmt_13/$exit
      -- CP-element group 19: 	 branch_block_stmt_11/loopback_PhiReq/phi_stmt_13/phi_stmt_13_sources/$exit
      -- CP-element group 19: 	 branch_block_stmt_11/loopback_PhiReq/phi_stmt_13/phi_stmt_13_sources/Interlock/$exit
      -- CP-element group 19: 	 branch_block_stmt_11/loopback_PhiReq/phi_stmt_13/phi_stmt_13_req
      -- 
    phi_stmt_13_req_132_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_13_req_132_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_gcd_CP_0_elements(19), ack => phi_stmt_13_req_1); -- 
    my_gcd_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "my_gcd_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= my_gcd_CP_0_elements(18) & my_gcd_CP_0_elements(17);
      gj_my_gcd_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => my_gcd_CP_0_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	7 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	22 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_11/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Sample/$exit
      -- CP-element group 20: 	 branch_block_stmt_11/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Sample/ack
      -- 
    ack_146_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ntB_72_20_buf_ack_0, ack => my_gcd_CP_0_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	7 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_11/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Update/$exit
      -- CP-element group 21: 	 branch_block_stmt_11/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/Update/ack
      -- 
    ack_151_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ntB_72_20_buf_ack_1, ack => my_gcd_CP_0_elements(21)); -- 
    -- CP-element group 22:  join  transition  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	20 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	23 
    -- CP-element group 22:  members (4) 
      -- CP-element group 22: 	 branch_block_stmt_11/loopback_PhiReq/phi_stmt_17/$exit
      -- CP-element group 22: 	 branch_block_stmt_11/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/$exit
      -- CP-element group 22: 	 branch_block_stmt_11/loopback_PhiReq/phi_stmt_17/phi_stmt_17_sources/Interlock/$exit
      -- CP-element group 22: 	 branch_block_stmt_11/loopback_PhiReq/phi_stmt_17/phi_stmt_17_req
      -- 
    phi_stmt_17_req_152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_17_req_152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => my_gcd_CP_0_elements(22), ack => phi_stmt_17_req_1); -- 
    my_gcd_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "my_gcd_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= my_gcd_CP_0_elements(20) & my_gcd_CP_0_elements(21);
      gj_my_gcd_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => my_gcd_CP_0_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	19 
    -- CP-element group 23: 	22 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_11/loopback_PhiReq/$exit
      -- 
    my_gcd_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "my_gcd_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= my_gcd_CP_0_elements(19) & my_gcd_CP_0_elements(22);
      gj_my_gcd_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => my_gcd_CP_0_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  merge  fork  transition  place  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	16 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_11/merge_stmt_12_PhiReqMerge
      -- CP-element group 24: 	 branch_block_stmt_11/merge_stmt_12_PhiAck/$entry
      -- 
    my_gcd_CP_0_elements(24) <= OrReduce(my_gcd_CP_0_elements(16) & my_gcd_CP_0_elements(23));
    -- CP-element group 25:  transition  input  bypass 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_11/merge_stmt_12_PhiAck/phi_stmt_13_ack
      -- 
    phi_stmt_13_ack_157_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_13_ack_0, ack => my_gcd_CP_0_elements(25)); -- 
    -- CP-element group 26:  transition  input  bypass 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	27 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_11/merge_stmt_12_PhiAck/phi_stmt_17_ack
      -- 
    phi_stmt_17_ack_158_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_17_ack_0, ack => my_gcd_CP_0_elements(26)); -- 
    -- CP-element group 27:  join  transition  bypass 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: 	26 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	1 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_11/merge_stmt_12_PhiAck/$exit
      -- 
    my_gcd_cp_element_group_27: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 26) := "my_gcd_cp_element_group_27"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= my_gcd_CP_0_elements(25) & my_gcd_CP_0_elements(26);
      gj_my_gcd_cp_element_group_27 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => my_gcd_CP_0_elements(27), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_29_wire : std_logic_vector(0 downto 0);
    signal A_15_buffered : std_logic_vector(31 downto 0);
    signal B_19_buffered : std_logic_vector(31 downto 0);
    signal EQ_u32_u1_38_wire : std_logic_vector(0 downto 0);
    signal EQ_u32_u1_42_wire : std_logic_vector(0 downto 0);
    signal EQ_u32_u1_45_wire : std_logic_vector(0 downto 0);
    signal MUX_50_wire : std_logic_vector(31 downto 0);
    signal NEQ_u32_u1_32_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_46_wire : std_logic_vector(0 downto 0);
    signal SUB_u32_u32_59_wire : std_logic_vector(31 downto 0);
    signal SUB_u32_u32_69_wire : std_logic_vector(31 downto 0);
    signal UGT_u32_u1_25_wire : std_logic_vector(0 downto 0);
    signal UGT_u32_u1_28_wire : std_logic_vector(0 downto 0);
    signal UGT_u32_u1_56_wire : std_logic_vector(0 downto 0);
    signal UGT_u32_u1_66_wire : std_logic_vector(0 downto 0);
    signal continue_flag_34 : std_logic_vector(0 downto 0);
    signal konst_24_wire_constant : std_logic_vector(31 downto 0);
    signal konst_27_wire_constant : std_logic_vector(31 downto 0);
    signal konst_41_wire_constant : std_logic_vector(31 downto 0);
    signal konst_44_wire_constant : std_logic_vector(31 downto 0);
    signal konst_47_wire_constant : std_logic_vector(31 downto 0);
    signal ntA_62 : std_logic_vector(31 downto 0);
    signal ntA_62_16_buffered : std_logic_vector(31 downto 0);
    signal ntB_72 : std_logic_vector(31 downto 0);
    signal ntB_72_20_buffered : std_logic_vector(31 downto 0);
    signal tA_13 : std_logic_vector(31 downto 0);
    signal tB_17 : std_logic_vector(31 downto 0);
    signal type_cast_49_wire_constant : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    konst_24_wire_constant <= "00000000000000000000000000000001";
    konst_27_wire_constant <= "00000000000000000000000000000001";
    konst_41_wire_constant <= "00000000000000000000000000000001";
    konst_44_wire_constant <= "00000000000000000000000000000001";
    konst_47_wire_constant <= "00000000000000000000000000000001";
    type_cast_49_wire_constant <= "00000000000000000000000000000000";
    phi_stmt_13: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= A_15_buffered & ntA_62_16_buffered;
      req <= phi_stmt_13_req_0 & phi_stmt_13_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_13",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_13_ack_0,
          idata => idata,
          odata => tA_13,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_13
    phi_stmt_17: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= B_19_buffered & ntB_72_20_buffered;
      req <= phi_stmt_17_req_0 & phi_stmt_17_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_17",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_17_ack_0,
          idata => idata,
          odata => tB_17,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_17
    -- flow-through select operator MUX_50_inst
    MUX_50_wire <= konst_47_wire_constant when (OR_u1_u1_46_wire(0) /=  '0') else type_cast_49_wire_constant;
    MUX_51_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_51_inst_req_0;
      MUX_51_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_51_inst_req_1;
      MUX_51_inst_ack_1<= update_ack(0);
      MUX_51_inst: SelectSplitProtocol generic map(name => "MUX_51_inst", data_width => 32, buffering => 1, flow_through => false, full_rate => false) -- 
        port map( x => tA_13, y => MUX_50_wire, sel => EQ_u32_u1_38_wire, z => GCD_buffer, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through select operator MUX_61_inst
    ntA_62 <= SUB_u32_u32_59_wire when (UGT_u32_u1_56_wire(0) /=  '0') else tA_13;
    -- flow-through select operator MUX_71_inst
    ntB_72 <= SUB_u32_u32_69_wire when (UGT_u32_u1_66_wire(0) /=  '0') else tB_17;
    A_15_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= A_15_buf_req_0;
      A_15_buf_ack_0<= wack(0);
      rreq(0) <= A_15_buf_req_1;
      A_15_buf_ack_1<= rack(0);
      A_15_buf : InterlockBuffer generic map ( -- 
        name => "A_15_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => A_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => A_15_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    B_19_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= B_19_buf_req_0;
      B_19_buf_ack_0<= wack(0);
      rreq(0) <= B_19_buf_req_1;
      B_19_buf_ack_1<= rack(0);
      B_19_buf : InterlockBuffer generic map ( -- 
        name => "B_19_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => B_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => B_19_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    ntA_62_16_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= ntA_62_16_buf_req_0;
      ntA_62_16_buf_ack_0<= wack(0);
      rreq(0) <= ntA_62_16_buf_req_1;
      ntA_62_16_buf_ack_1<= rack(0);
      ntA_62_16_buf : InterlockBuffer generic map ( -- 
        name => "ntA_62_16_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ntA_62,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ntA_62_16_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    ntB_72_20_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= ntB_72_20_buf_req_0;
      ntB_72_20_buf_ack_0<= wack(0);
      rreq(0) <= ntB_72_20_buf_req_1;
      ntB_72_20_buf_ack_1<= rack(0);
      ntB_72_20_buf : InterlockBuffer generic map ( -- 
        name => "ntB_72_20_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false ,
        in_phi =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ntB_72,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ntB_72_20_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    if_stmt_73_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= continue_flag_34;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_73_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_73_branch_req_0,
          ack0 => if_stmt_73_branch_ack_0,
          ack1 => if_stmt_73_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- flow through binary operator AND_u1_u1_29_inst
    AND_u1_u1_29_wire <= (UGT_u32_u1_25_wire and UGT_u32_u1_28_wire);
    -- shared split operator group (1) : AND_u1_u1_33_inst 
    ApIntAnd_group_1: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= AND_u1_u1_29_wire & NEQ_u32_u1_32_wire;
      continue_flag_34 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u1_u1_33_inst_req_0;
      AND_u1_u1_33_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u1_u1_33_inst_req_1;
      AND_u1_u1_33_inst_ack_1 <= ackR_unguarded(0);
      ApIntAnd_group_1_gI: SplitGuardInterface generic map(name => "ApIntAnd_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_1",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 1, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 1
    -- flow through binary operator EQ_u32_u1_38_inst
    process(tA_13, tB_17) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(tA_13, tB_17, tmp_var);
      EQ_u32_u1_38_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u32_u1_42_inst
    process(tA_13) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(tA_13, konst_41_wire_constant, tmp_var);
      EQ_u32_u1_42_wire <= tmp_var; --
    end process;
    -- flow through binary operator EQ_u32_u1_45_inst
    process(tB_17) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(tB_17, konst_44_wire_constant, tmp_var);
      EQ_u32_u1_45_wire <= tmp_var; --
    end process;
    -- flow through binary operator NEQ_u32_u1_32_inst
    process(tA_13, tB_17) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(tA_13, tB_17, tmp_var);
      NEQ_u32_u1_32_wire <= tmp_var; --
    end process;
    -- flow through binary operator OR_u1_u1_46_inst
    OR_u1_u1_46_wire <= (EQ_u32_u1_42_wire or EQ_u32_u1_45_wire);
    -- flow through binary operator SUB_u32_u32_59_inst
    SUB_u32_u32_59_wire <= std_logic_vector(unsigned(tA_13) - unsigned(tB_17));
    -- flow through binary operator SUB_u32_u32_69_inst
    SUB_u32_u32_69_wire <= std_logic_vector(unsigned(tB_17) - unsigned(tA_13));
    -- flow through binary operator UGT_u32_u1_25_inst
    process(tA_13) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tA_13, konst_24_wire_constant, tmp_var);
      UGT_u32_u1_25_wire <= tmp_var; --
    end process;
    -- flow through binary operator UGT_u32_u1_28_inst
    process(tB_17) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tB_17, konst_27_wire_constant, tmp_var);
      UGT_u32_u1_28_wire <= tmp_var; --
    end process;
    -- flow through binary operator UGT_u32_u1_56_inst
    process(tA_13, tB_17) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tA_13, tB_17, tmp_var);
      UGT_u32_u1_56_wire <= tmp_var; --
    end process;
    -- flow through binary operator UGT_u32_u1_66_inst
    process(tB_17, tA_13) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(tB_17, tA_13, tmp_var);
      UGT_u32_u1_66_wire <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end my_gcd_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library AjitCustom;
use AjitCustom.baud_control_calculator_global_package.all;
entity baud_control_calculator is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    BAUD_CONTROL_WORD_SIG: out std_logic_vector(31 downto 0);
    BAUD_CONTROL_WORD_VALID: out std_logic_vector(0 downto 0);
    BAUD_RATE_SIG: in std_logic_vector(31 downto 0);
    CLK_FREQUENCY_SIG: in std_logic_vector(31 downto 0);
    CLOCK_FREQUENCY_VALID: in std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture baud_control_calculator_arch  of baud_control_calculator is -- system-architecture 
  -- declarations related to module baudControlCalculatorDaemon
  component baudControlCalculatorDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      BAUD_RATE_SIG : in std_logic_vector(31 downto 0);
      CLK_FREQUENCY_SIG : in std_logic_vector(31 downto 0);
      CLOCK_FREQUENCY_VALID : in std_logic_vector(0 downto 0);
      BAUD_CONTROL_WORD_SIG_pipe_write_req : out  std_logic_vector(0 downto 0);
      BAUD_CONTROL_WORD_SIG_pipe_write_ack : in   std_logic_vector(0 downto 0);
      BAUD_CONTROL_WORD_SIG_pipe_write_data : out  std_logic_vector(31 downto 0);
      BAUD_CONTROL_WORD_VALID_pipe_write_req : out  std_logic_vector(0 downto 0);
      BAUD_CONTROL_WORD_VALID_pipe_write_ack : in   std_logic_vector(0 downto 0);
      BAUD_CONTROL_WORD_VALID_pipe_write_data : out  std_logic_vector(0 downto 0);
      my_gcd_call_reqs : out  std_logic_vector(0 downto 0);
      my_gcd_call_acks : in   std_logic_vector(0 downto 0);
      my_gcd_call_data : out  std_logic_vector(63 downto 0);
      my_gcd_call_tag  :  out  std_logic_vector(0 downto 0);
      my_gcd_return_reqs : out  std_logic_vector(0 downto 0);
      my_gcd_return_acks : in   std_logic_vector(0 downto 0);
      my_gcd_return_data : in   std_logic_vector(31 downto 0);
      my_gcd_return_tag :  in   std_logic_vector(0 downto 0);
      my_div_call_reqs : out  std_logic_vector(0 downto 0);
      my_div_call_acks : in   std_logic_vector(0 downto 0);
      my_div_call_data : out  std_logic_vector(63 downto 0);
      my_div_call_tag  :  out  std_logic_vector(1 downto 0);
      my_div_return_reqs : out  std_logic_vector(0 downto 0);
      my_div_return_acks : in   std_logic_vector(0 downto 0);
      my_div_return_data : in   std_logic_vector(31 downto 0);
      my_div_return_tag :  in   std_logic_vector(1 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module baudControlCalculatorDaemon
  signal baudControlCalculatorDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal baudControlCalculatorDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal baudControlCalculatorDaemon_start_req : std_logic;
  signal baudControlCalculatorDaemon_start_ack : std_logic;
  signal baudControlCalculatorDaemon_fin_req   : std_logic;
  signal baudControlCalculatorDaemon_fin_ack : std_logic;
  -- declarations related to module my_div
  component my_div is -- 
    generic (tag_length : integer); 
    port ( -- 
      A : in  std_logic_vector(31 downto 0);
      B : in  std_logic_vector(31 downto 0);
      Q : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module my_div
  signal my_div_A :  std_logic_vector(31 downto 0);
  signal my_div_B :  std_logic_vector(31 downto 0);
  signal my_div_Q :  std_logic_vector(31 downto 0);
  signal my_div_in_args    : std_logic_vector(63 downto 0);
  signal my_div_out_args   : std_logic_vector(31 downto 0);
  signal my_div_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal my_div_tag_out   : std_logic_vector(2 downto 0);
  signal my_div_start_req : std_logic;
  signal my_div_start_ack : std_logic;
  signal my_div_fin_req   : std_logic;
  signal my_div_fin_ack : std_logic;
  -- caller side aggregated signals for module my_div
  signal my_div_call_reqs: std_logic_vector(0 downto 0);
  signal my_div_call_acks: std_logic_vector(0 downto 0);
  signal my_div_return_reqs: std_logic_vector(0 downto 0);
  signal my_div_return_acks: std_logic_vector(0 downto 0);
  signal my_div_call_data: std_logic_vector(63 downto 0);
  signal my_div_call_tag: std_logic_vector(1 downto 0);
  signal my_div_return_data: std_logic_vector(31 downto 0);
  signal my_div_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module my_gcd
  component my_gcd is -- 
    generic (tag_length : integer); 
    port ( -- 
      A : in  std_logic_vector(31 downto 0);
      B : in  std_logic_vector(31 downto 0);
      GCD : out  std_logic_vector(31 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module my_gcd
  signal my_gcd_A :  std_logic_vector(31 downto 0);
  signal my_gcd_B :  std_logic_vector(31 downto 0);
  signal my_gcd_GCD :  std_logic_vector(31 downto 0);
  signal my_gcd_in_args    : std_logic_vector(63 downto 0);
  signal my_gcd_out_args   : std_logic_vector(31 downto 0);
  signal my_gcd_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal my_gcd_tag_out   : std_logic_vector(1 downto 0);
  signal my_gcd_start_req : std_logic;
  signal my_gcd_start_ack : std_logic;
  signal my_gcd_fin_req   : std_logic;
  signal my_gcd_fin_ack : std_logic;
  -- caller side aggregated signals for module my_gcd
  signal my_gcd_call_reqs: std_logic_vector(0 downto 0);
  signal my_gcd_call_acks: std_logic_vector(0 downto 0);
  signal my_gcd_return_reqs: std_logic_vector(0 downto 0);
  signal my_gcd_return_acks: std_logic_vector(0 downto 0);
  signal my_gcd_call_data: std_logic_vector(63 downto 0);
  signal my_gcd_call_tag: std_logic_vector(0 downto 0);
  signal my_gcd_return_data: std_logic_vector(31 downto 0);
  signal my_gcd_return_tag: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe BAUD_CONTROL_WORD_SIG
  signal BAUD_CONTROL_WORD_SIG_pipe_write_data: std_logic_vector(31 downto 0);
  signal BAUD_CONTROL_WORD_SIG_pipe_write_req: std_logic_vector(0 downto 0);
  signal BAUD_CONTROL_WORD_SIG_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe BAUD_CONTROL_WORD_VALID
  signal BAUD_CONTROL_WORD_VALID_pipe_write_data: std_logic_vector(0 downto 0);
  signal BAUD_CONTROL_WORD_VALID_pipe_write_req: std_logic_vector(0 downto 0);
  signal BAUD_CONTROL_WORD_VALID_pipe_write_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module baudControlCalculatorDaemon
  baudControlCalculatorDaemon_instance:baudControlCalculatorDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => baudControlCalculatorDaemon_start_req,
      start_ack => baudControlCalculatorDaemon_start_ack,
      fin_req => baudControlCalculatorDaemon_fin_req,
      fin_ack => baudControlCalculatorDaemon_fin_ack,
      clk => clk,
      reset => reset,
      BAUD_RATE_SIG => BAUD_RATE_SIG,
      CLK_FREQUENCY_SIG => CLK_FREQUENCY_SIG,
      CLOCK_FREQUENCY_VALID => CLOCK_FREQUENCY_VALID,
      BAUD_CONTROL_WORD_SIG_pipe_write_req => BAUD_CONTROL_WORD_SIG_pipe_write_req(0 downto 0),
      BAUD_CONTROL_WORD_SIG_pipe_write_ack => BAUD_CONTROL_WORD_SIG_pipe_write_ack(0 downto 0),
      BAUD_CONTROL_WORD_SIG_pipe_write_data => BAUD_CONTROL_WORD_SIG_pipe_write_data(31 downto 0),
      BAUD_CONTROL_WORD_VALID_pipe_write_req => BAUD_CONTROL_WORD_VALID_pipe_write_req(0 downto 0),
      BAUD_CONTROL_WORD_VALID_pipe_write_ack => BAUD_CONTROL_WORD_VALID_pipe_write_ack(0 downto 0),
      BAUD_CONTROL_WORD_VALID_pipe_write_data => BAUD_CONTROL_WORD_VALID_pipe_write_data(0 downto 0),
      my_gcd_call_reqs => my_gcd_call_reqs(0 downto 0),
      my_gcd_call_acks => my_gcd_call_acks(0 downto 0),
      my_gcd_call_data => my_gcd_call_data(63 downto 0),
      my_gcd_call_tag => my_gcd_call_tag(0 downto 0),
      my_gcd_return_reqs => my_gcd_return_reqs(0 downto 0),
      my_gcd_return_acks => my_gcd_return_acks(0 downto 0),
      my_gcd_return_data => my_gcd_return_data(31 downto 0),
      my_gcd_return_tag => my_gcd_return_tag(0 downto 0),
      my_div_call_reqs => my_div_call_reqs(0 downto 0),
      my_div_call_acks => my_div_call_acks(0 downto 0),
      my_div_call_data => my_div_call_data(63 downto 0),
      my_div_call_tag => my_div_call_tag(1 downto 0),
      my_div_return_reqs => my_div_return_reqs(0 downto 0),
      my_div_return_acks => my_div_return_acks(0 downto 0),
      my_div_return_data => my_div_return_data(31 downto 0),
      my_div_return_tag => my_div_return_tag(1 downto 0),
      tag_in => baudControlCalculatorDaemon_tag_in,
      tag_out => baudControlCalculatorDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  baudControlCalculatorDaemon_tag_in <= (others => '0');
  baudControlCalculatorDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => baudControlCalculatorDaemon_start_req, start_ack => baudControlCalculatorDaemon_start_ack,  fin_req => baudControlCalculatorDaemon_fin_req,  fin_ack => baudControlCalculatorDaemon_fin_ack);
  -- module my_div
  my_div_A <= my_div_in_args(63 downto 32);
  my_div_B <= my_div_in_args(31 downto 0);
  my_div_out_args <= my_div_Q ;
  -- call arbiter for module my_div
  my_div_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 64,
      return_data_width => 32,
      callee_tag_length => 1,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => my_div_call_reqs,
      call_acks => my_div_call_acks,
      return_reqs => my_div_return_reqs,
      return_acks => my_div_return_acks,
      call_data  => my_div_call_data,
      call_tag  => my_div_call_tag,
      return_tag  => my_div_return_tag,
      call_mtag => my_div_tag_in,
      return_mtag => my_div_tag_out,
      return_data =>my_div_return_data,
      call_mreq => my_div_start_req,
      call_mack => my_div_start_ack,
      return_mreq => my_div_fin_req,
      return_mack => my_div_fin_ack,
      call_mdata => my_div_in_args,
      return_mdata => my_div_out_args,
      clk => clk, 
      reset => reset --
    ); --
  my_div_instance:my_div-- 
    generic map(tag_length => 3)
    port map(-- 
      A => my_div_A,
      B => my_div_B,
      Q => my_div_Q,
      start_req => my_div_start_req,
      start_ack => my_div_start_ack,
      fin_req => my_div_fin_req,
      fin_ack => my_div_fin_ack,
      clk => clk,
      reset => reset,
      tag_in => my_div_tag_in,
      tag_out => my_div_tag_out-- 
    ); -- 
  -- module my_gcd
  my_gcd_A <= my_gcd_in_args(63 downto 32);
  my_gcd_B <= my_gcd_in_args(31 downto 0);
  my_gcd_out_args <= my_gcd_GCD ;
  -- call arbiter for module my_gcd
  my_gcd_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 64,
      return_data_width => 32,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => my_gcd_call_reqs,
      call_acks => my_gcd_call_acks,
      return_reqs => my_gcd_return_reqs,
      return_acks => my_gcd_return_acks,
      call_data  => my_gcd_call_data,
      call_tag  => my_gcd_call_tag,
      return_tag  => my_gcd_return_tag,
      call_mtag => my_gcd_tag_in,
      return_mtag => my_gcd_tag_out,
      return_data =>my_gcd_return_data,
      call_mreq => my_gcd_start_req,
      call_mack => my_gcd_start_ack,
      return_mreq => my_gcd_fin_req,
      return_mack => my_gcd_fin_ack,
      call_mdata => my_gcd_in_args,
      return_mdata => my_gcd_out_args,
      clk => clk, 
      reset => reset --
    ); --
  my_gcd_instance:my_gcd-- 
    generic map(tag_length => 2)
    port map(-- 
      A => my_gcd_A,
      B => my_gcd_B,
      GCD => my_gcd_GCD,
      start_req => my_gcd_start_req,
      start_ack => my_gcd_start_ack,
      fin_req => my_gcd_fin_req,
      fin_ack => my_gcd_fin_ack,
      clk => clk,
      reset => reset,
      tag_in => my_gcd_tag_in,
      tag_out => my_gcd_tag_out-- 
    ); -- 
  BAUD_CONTROL_WORD_SIG_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe BAUD_CONTROL_WORD_SIG",
      volatile_flag => false,
      num_writes => 1,
      data_width => 32 --
    ) 
    port map( -- 
      read_data => BAUD_CONTROL_WORD_SIG,
      write_req => BAUD_CONTROL_WORD_SIG_pipe_write_req,
      write_ack => BAUD_CONTROL_WORD_SIG_pipe_write_ack,
      write_data => BAUD_CONTROL_WORD_SIG_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  BAUD_CONTROL_WORD_VALID_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe BAUD_CONTROL_WORD_VALID",
      volatile_flag => false,
      num_writes => 1,
      data_width => 1 --
    ) 
    port map( -- 
      read_data => BAUD_CONTROL_WORD_VALID,
      write_req => BAUD_CONTROL_WORD_VALID_pipe_write_req,
      write_ack => BAUD_CONTROL_WORD_VALID_pipe_write_ack,
      write_data => BAUD_CONTROL_WORD_VALID_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- input signal-pipe BAUD_RATE_SIG accessed directly. 
  -- input signal-pipe CLK_FREQUENCY_SIG accessed directly. 
  -- input signal-pipe CLOCK_FREQUENCY_VALID accessed directly. 
  -- gated clock generators 
  -- 
end baud_control_calculator_arch;
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

library AjitCustom;
use AjitCustom.AjitCustomComponents.all;

library simpleUartLib;
use simpleUartLib.uartPackage.all;

entity configurable_self_tuning_uart is
	port (clk, reset: in std_logic; 
		rt_1Hz: in std_logic_vector(0 downto 0); 

		BAUD_RATE: in std_logic_vector(31 downto 0);
		UART_RX: in std_logic_vector(0 downto 0); 
		UART_TX: out std_logic_vector(0 downto 0);

		TX_to_CONSOLE_pipe_write_data: in std_logic_vector(7 downto 0);
		TX_to_CONSOLE_pipe_write_req:  in std_logic_vector(0 downto 0);
		TX_to_CONSOLE_pipe_write_ack:  out std_logic_vector(0 downto 0);

		CONSOLE_to_RX_pipe_read_data : out std_logic_vector(7 downto 0);
		CONSOLE_to_RX_pipe_read_req :  in std_logic_vector(0 downto 0);
		CONSOLE_to_RX_pipe_read_ack :  out std_logic_vector(0 downto 0));
end entity configurable_self_tuning_uart;


architecture Struct of configurable_self_tuning_uart is

	signal baud_control_word: std_logic_vector(31 downto 0);
	signal baud_control_word_valid: std_logic;
	signal clock_frequency_valid: std_logic;
        signal clock_frequency  : std_logic_vector(31 downto 0);
    				
	signal counter : integer;
	signal reset_uart: std_logic;

	constant Z32: std_logic_vector(31 downto 0) := (others => '0');
	signal soft_reset: std_logic;
begin

	--------------------------------------------------------------
	-- soft reset
	--------------------------------------------------------------
	process(clk, reset)
	begin
		if(clk'event and clk = '1') then
			if(reset_uart = '1') then
				counter <= 0;
				soft_reset <= '1';
			else 
				if(counter = 255) then
					soft_reset <= '0';
					counter <= 0;
				else
					counter <= counter + 1;
				end if;
			end if;
		end if;
	end process;

	-------------------------------------------------------
	-- estimate the clock frequency
	-------------------------------------------------------
	rt_ctr_inst: rt_clock_counter
		port map (clk => clk, 
				reset => reset,
				one_hz_rt_clock => rt_1Hz,
				count_value => clock_frequency);	
	clock_frequency_valid <= '1' when (clock_frequency /= Z32) else '0';
	reset_uart <= '1' when ((reset = '1') or  (baud_control_word_valid = '0')) else '0';

	-------------------------------------------------------
	-- calculate the baud control word.
	-------------------------------------------------------
	bcc_inst: baud_control_calculator
		port map (clk => clk, reset => reset,
				BAUD_CONTROL_WORD_SIG => baud_control_word,
				BAUD_CONTROL_WORD_VALID(0) => baud_control_word_valid,
				BAUD_RATE_SIG => BAUD_RATE,
				CLK_FREQUENCY_SIG => clock_frequency,
				CLOCK_FREQUENCY_VALID(0) => clock_frequency_valid);

	-------------------------------------------------------
	-- The UART!
	-------------------------------------------------------
	uart_inst: uartTopPortConfigurable
		port map (
				reset => reset_uart,
				clk => clk,
				soft_reset => soft_reset,
				serIn     => UART_RX(0),	
				serOut    => UART_TX(0),	
				baudFreq  =>  baud_control_word(11 downto 0),
				baudLimit => baud_control_word(31 downto 16),
	 			uart_rx_pipe_read_data => CONSOLE_to_RX_pipe_read_data,
	 			uart_rx_pipe_read_req => CONSOLE_to_RX_pipe_read_req,
	 			uart_rx_pipe_read_ack => CONSOLE_to_RX_pipe_read_ack,
	 			uart_tx_pipe_write_data => TX_to_CONSOLE_pipe_write_data,
	 			uart_tx_pipe_write_req => TX_to_CONSOLE_pipe_write_req,
	 			uart_tx_pipe_write_ack => TX_to_CONSOLE_pipe_write_ack
		);
end Struct;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
use AjitCustom.AjitCoreConfigurationPackage.all;

entity access_instruction_buffer_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    clear_flag : in  std_logic_vector(0 downto 0);
    insert_flag : in  std_logic_vector(0 downto 0);
    insert_addr : in  std_logic_vector(28 downto 0);
    insert_acc  : in  std_logic_vector(2 downto 0);
    insert_ipair : in  std_logic_vector(63 downto 0);
    lookup_flag : in  std_logic_vector(0 downto 0);
    lookup_addr : in  std_logic_vector(28 downto 0);
    lookup_match : out  std_logic_vector(0 downto 0);
    lookup_acc  : out  std_logic_vector(2 downto 0);
    lookup_ipair : out  std_logic_vector(63 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity access_instruction_buffer_Operator;
architecture access_instruction_buffer_Operator_arch of access_instruction_buffer_Operator is -- 
	signal lookup_tag, insert_tag: std_logic_vector(28 downto 0);
	signal lookup_data, insert_data: std_logic_vector(66 downto 0);
begin --  
	insert_tag  <= insert_addr (28 downto 0);
	insert_data <= insert_acc & insert_ipair;
	
	lookup_tag <= lookup_addr (28 downto 0);
	basemem:genericDirectMappedAssociativeMemory
			generic map(
					tag_width => insert_tag'length,
					data_width => insert_data'length,
					log2_number_of_entries => INSTRUCTION_BUFFER_LOG_MEMORY_SIZE
				    )
			port map(
					sample_req => sample_req,
					sample_ack => sample_ack,
					update_req => update_req,
					update_ack => update_ack,
					init_flag => clear_flag,
					insert_flag => insert_flag,
					insert_data => insert_data,
					insert_tag =>  insert_tag,
					lookup_flag => lookup_flag,
					lookup_tag => lookup_tag,
					lookup_match => lookup_match,
					lookup_data => lookup_data,
					clk => clk, reset => reset);
	
	lookup_acc <= lookup_data (66 downto 64);
	lookup_ipair <= lookup_data (63 downto 0);

end access_instruction_buffer_Operator_arch;
-- Optimized version of instruction buffer.
-- The instruction buffer is used in the icache path of the
-- dual threaded CPU's in order to reduce blocking on the
-- icache (for example a tight spin-loop can be absorbed into
-- the instruction buffer thus reducing the pressure on the shared
-- icache)
--
-- Author: Madhav Desai, January 25, 2023.
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.basecomponents.all;
use ahir.Utilities.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
use AjitCustom.AjitCoreConfigurationPackage.all;
use AjitCustom.UsefulFunctions.all;

entity instruction_buffer_optimized is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    icache_to_instruction_buffer_response_pipe_write_data: in std_logic_vector(89 downto 0);
    icache_to_instruction_buffer_response_pipe_write_req : in std_logic_vector(0 downto 0);
    icache_to_instruction_buffer_response_pipe_write_ack : out std_logic_vector(0 downto 0);
    instruction_buffer_to_cpu_response_pipe_read_data: out std_logic_vector(89 downto 0);
    instruction_buffer_to_cpu_response_pipe_read_req : in std_logic_vector(0 downto 0);
    instruction_buffer_to_cpu_response_pipe_read_ack : out std_logic_vector(0 downto 0);
    noblock_cpu_to_instruction_buffer_request_pipe_write_data: in std_logic_vector(40 downto 0);
    noblock_cpu_to_instruction_buffer_request_pipe_write_req : in std_logic_vector(0 downto 0);
    noblock_cpu_to_instruction_buffer_request_pipe_write_ack : out std_logic_vector(0 downto 0);
    noblock_instruction_buffer_to_icache_request_pipe_read_data: out std_logic_vector(40 downto 0);
    noblock_instruction_buffer_to_icache_request_pipe_read_req : in std_logic_vector(0 downto 0);
    noblock_instruction_buffer_to_icache_request_pipe_read_ack : out std_logic_vector(0 downto 0);
    core_id: std_logic_Vector(3 downto 0);
    cpu_id: std_logic_vector(3 downto 0)); -- 
  -- 
end entity; 

architecture instruction_buffer_arch  of instruction_buffer_optimized is -- system-architecture 

  	constant ASI_SUPERVISOR_INSTRUCTION : std_logic_vector(3 downto 0) := "1001";
  	constant ASI_USER_INSTRUCTION : std_logic_vector(3 downto 0) := "1000";


	signal cpu_has_request, cpu_ready_for_response: boolean;
	signal icache_ready_for_request, icache_has_response, icache_response_is_awaited: boolean;

	signal pending_queue_has_room, pending_queue_has_data: boolean;
	signal pending_queue_push_data, pending_queue_pop_data: std_logic_vector(93 downto 0);
	signal pending_queue_push_req, pending_queue_push_ack,
			pending_queue_pop_req, pending_queue_pop_ack: std_logic;

	signal ipair_from_lookup_data, ipair_from_pending_queue, 
		ipair_from_icache_response, ipair_to_cpu : std_logic_vector(63 downto 0);
	signal acc_from_lookup_data, acc_from_icache_response: std_logic_vector(2 downto 0);
	signal cacheable_from_icache_response: std_logic_vector(0 downto 0);

	signal cpu_request_is_flush, is_cacheable_non_mae_icache_response: boolean;

	signal cpu_request_valid, cpu_request_valid_d: std_logic;
	signal cpu_request_asi_4_d: std_logic_vector(3 downto 0);
	signal cpu_request_addr, cpu_request_addr_d: std_logic_vector(31 downto 0);

	signal lookup_flag, insert_flag, init_flag, lookup_match:  std_logic_vector(0 downto 0);
	signal lookup_addr, insert_addr: std_logic_vector(28 downto 0);
	signal lookup_data, lookup_data_reg, lookup_data_qualified, insert_data: std_logic_vector(66 downto 0);

	signal access_permissions_ok: std_logic;
	signal send_to_icache, send_to_cpu: boolean;
	signal forward_pending_to_cpu: boolean;
	signal accept_cpu_request, accept_icache_response: boolean;
	signal privileges_ok: boolean;

	constant PENDING_QUEUE_DEPTH: integer := 4;

	
	signal is_S, is_U, is_ifetch, is_read: std_logic;
	signal is_tlb_hit, is_tlb_hit_reg, is_tlb_hit_qualified: boolean;
	signal fsr_from_icache_response, fsr_to_cpu: std_logic_vector(17 downto 0);
	signal mae_8_from_icache_response, mae_8_from_lookup,  mae_8_to_cpu: std_logic_vector(7 downto 0);

	signal cpu_request_started: boolean;

	signal tlb_sample_req, tlb_sample_ack, tlb_update_req, tlb_update_ack: boolean;
    
	signal icache_response_data: std_logic_vector(89 downto 0);
	signal icache_response_ready, icache_response_accept: boolean;
    
	signal cpu_response_data: std_logic_vector(89 downto 0);
    	signal cpu_response_ready, cpu_hit_response_ready, cpu_miss_response_ready : boolean;

    	signal cpu_request_data, cpu_request_data_reg: std_logic_vector(40 downto 0);
    	signal cpu_request_ready, cpu_request_accept: boolean;

   	signal icache_request_data: std_logic_vector(40 downto 0);
    	signal icache_request_ready: boolean;

	signal exec_tlb_lookup, exec_tlb_insert, exec_tlb_clear: boolean;


	type FsmState is (IDLE, RUNNING, STALLED);
	signal fsm_state: FsmState;

	signal save_lookup_results: boolean;

begin -- 
	-----------------------------------------------------------------------
	-- handles.
	-----------------------------------------------------------------------

	-- icache response to instruction buffer.
	icache_response_data <= icache_to_instruction_buffer_response_pipe_write_data;
	icache_response_ready <= icache_to_instruction_buffer_response_pipe_write_req(0) = '1';
	icache_to_instruction_buffer_response_pipe_write_ack(0) <= '1' when icache_response_accept else '0';

	-- instruction buffer response to cpu.
    	instruction_buffer_to_cpu_response_pipe_read_data <= cpu_response_data;
    	cpu_ready_for_response <= instruction_buffer_to_cpu_response_pipe_read_req(0) = '1';
    	instruction_buffer_to_cpu_response_pipe_read_ack(0) <= '1' when cpu_response_ready else '0';

	-- request data from the cpu.
    	cpu_request_data <= noblock_cpu_to_instruction_buffer_request_pipe_write_data;
    	cpu_request_ready <= noblock_cpu_to_instruction_buffer_request_pipe_write_req(0) = '1' and
    				noblock_cpu_to_instruction_buffer_request_pipe_write_data(40) = '1';
	noblock_cpu_to_instruction_buffer_request_pipe_write_ack(0) <= '1' when cpu_request_accept else '0';
	
	-- instruction buffer request to icache.
    	noblock_instruction_buffer_to_icache_request_pipe_read_data <= icache_request_data;
    	icache_ready_for_request <= (noblock_instruction_buffer_to_icache_request_pipe_read_req(0) = '1');
    	noblock_instruction_buffer_to_icache_request_pipe_read_ack(0) <= '1' when icache_request_ready else '0';

	-- is the cpu request a flush?
    	cpu_request_is_flush <= (cpu_request_data(39) = '1');


	-- delayed version of cpu request updated whenever cpu request is accepted.
	process(clk, cpu_request_data, cpu_request_started)
	begin
		if(clk'event and (clk = '1')) then
			if(cpu_request_started) then
				cpu_request_data_reg <= cpu_request_data;
			end if;
		end if;
	end process;


	cpu_request_started <= cpu_request_ready and cpu_request_accept;

	--------------------------------------------------------------------------------
	-- FSM to determine when a cpu request can be accepted.
	--------------------------------------------------------------------------------
	process(clk, reset, fsm_state, 
			cpu_request_ready, 
			icache_ready_for_request,
			pending_queue_has_room)
		variable next_fsm_state_var: FsmState;
		variable cpu_request_accept_var: boolean;
		variable exec_tlb_lookup_var: boolean;
		variable save_lookup_results_var: boolean;
		variable icache_request_ready_var : boolean;
		variable pending_queue_push_req_var: std_logic;
		variable stall_var: boolean;
	begin
		next_fsm_state_var := fsm_state;
		cpu_request_accept_var := false;
		exec_tlb_lookup_var := false;
		save_lookup_results_var := false;
		icache_request_ready_var := false;
		pending_queue_push_req_var := '0';
		stall_var := false;
	

		case fsm_state is 
			when IDLE =>
				cpu_request_accept_var := true;
				if(cpu_request_ready) then 
					exec_tlb_lookup_var := true;
					next_fsm_state_var := RUNNING;
				end if;
			when RUNNING =>
				-- pending queue must have room... and if needed,
				-- icache must be ready to accept request..
				stall_var := (not pending_queue_has_room) or
							((not is_tlb_hit) and (not icache_ready_for_request));
							
				icache_request_ready_var := (not is_tlb_hit) and pending_queue_has_room;

				if(stall_var) then
					save_lookup_results_var := true;
					next_fsm_state_var := STALLED;
				else
					pending_queue_push_req_var := '1';
					cpu_request_accept_var := true;

					if(cpu_request_ready) then 
						exec_tlb_lookup_var := true;
					else
						next_fsm_state_var := IDLE;
					end if;
				end if;
			when STALLED =>
				stall_var := (not pending_queue_has_room) or
							((not is_tlb_hit_reg) and (not icache_ready_for_request));
				icache_request_ready_var := (not is_tlb_hit_reg) and pending_queue_has_room;

				if(not stall_var) then
					next_fsm_state_var := IDLE;
					pending_queue_push_req_var := '1';
				end if;
		end case;

		exec_tlb_lookup <= exec_tlb_lookup_var;
		save_lookup_results <= save_lookup_results_var;
		cpu_request_accept <= cpu_request_accept_var;
		icache_request_ready <= icache_request_ready_var;
		pending_queue_push_req <= pending_queue_push_req_var;

		if(clk'event and (clk = '1')) then
			if(reset = '1') then
				fsm_state <= IDLE;
			else
				fsm_state <= next_fsm_state_var;
			end if;
		end if;
	end process;

	--------------------------------------------------------------------------------
	-- TLB... 
	--------------------------------------------------------------------------------
	exec_tlb_clear <= cpu_request_is_flush and cpu_request_started;
	exec_tlb_insert <= 
		(icache_response_ready and icache_response_accept and is_cacheable_non_mae_icache_response);
	insert_flag(0) <= '1' when exec_tlb_insert else '0';


	process(clk, reset, is_tlb_hit, lookup_data, save_lookup_results)
	begin
		if(clk'event and (clk = '1')) then
			if(reset ='1') then
				is_tlb_hit_reg <= is_tlb_hit;
				lookup_data_reg  <= (others => '0');
			else
				if(save_lookup_results) then
					is_tlb_hit_reg <= is_tlb_hit;
					lookup_data_reg <= lookup_data;
				end if;
			end if;
		end if;
	end process;

	-- lookup if cpu request started and cpu request is not a flush.
	lookup_flag(0) <= '1' when exec_tlb_lookup else '0';
	lookup_addr <= cpu_request_data(31 downto 3);


	-- clear all when it is a flush.
	init_flag(0) <= '1' when exec_tlb_clear else '0';

	-- trigger the tlb.
	tlb_sample_req <= (exec_tlb_lookup or exec_tlb_insert or exec_tlb_clear);
	tlb_update_req <= tlb_sample_req;
	
	tlb_inst:
		genericDirectMappedAssociativeMemory
			generic map (data_width => 67, tag_width => 29,
						log2_number_of_entries => INSTRUCTION_BUFFER_LOG_MEMORY_SIZE)
			port map (
					sample_req => tlb_sample_req,
					sample_ack => tlb_sample_ack,
					update_req => tlb_update_req,
					update_ack => tlb_update_ack,
					init_flag => init_flag,
					insert_flag => insert_flag,
					insert_tag => insert_addr,
					insert_data => insert_data,
					lookup_flag => lookup_flag,
					lookup_tag => lookup_addr, 
					lookup_match => lookup_match,
					lookup_data => lookup_data,
					clk => clk, reset => reset
				);
					

	lookup_data_qualified  <= lookup_data  when (fsm_state = RUNNING) else lookup_data_reg;
	is_tlb_hit_qualified   <= is_tlb_hit   when (fsm_state = RUNNING) else is_tlb_hit_reg;


	acc_from_lookup_data <= lookup_data_qualified(66 downto 64);
	ipair_from_lookup_data <= lookup_data_qualified(63 downto 0);

	-- the cpu request asi (delayed!).
	cpu_request_asi_4_d <= cpu_request_data_reg(35 downto 32);

	is_S <= '1' when (cpu_request_asi_4_d = ASI_SUPERVISOR_INSTRUCTION) else '0';
	is_U <= '1' when (cpu_request_asi_4_d = ASI_USER_INSTRUCTION) else '0';

	is_ifetch <= '1';
	is_read   <= '0';

	access_permissions_ok <= accessPermissionsOk(is_S, is_ifetch, is_read, acc_from_lookup_data); 

	is_tlb_hit <= (lookup_match(0) = '1') and (access_permissions_ok = '1');
	icache_request_data <= cpu_request_data_reg;

	--------------------------------------------------------------------------------
	-- Pending queue
	--      is-hit lookup-ipair addr
	--         1       64        29
	--------------------------------------------------------------------------------
	pq: QueueWithBypass
		generic map (name => "pending_queue", data_width => 94, queue_depth => PENDING_QUEUE_DEPTH)
		port map (
			data_in => pending_queue_push_data,
			push_req => pending_queue_push_req,
			push_ack => pending_queue_push_ack,
			data_out => pending_queue_pop_data,
			pop_req => pending_queue_pop_req,
			pop_ack => pending_queue_pop_ack,
			clk => clk, reset => reset
		);

	pending_queue_push_data(93)  <=  '1' when is_tlb_hit_qualified else '0';
	pending_queue_push_data(92 downto 0)  <=  (cpu_request_data_reg(31 downto 3) & ipair_from_lookup_data);

	pending_queue_has_room <= (pending_queue_push_ack = '1');
	pending_queue_has_data <= (pending_queue_pop_ack  = '1');

	pending_queue_pop_req  <= '1' when 
				(pending_queue_has_data and cpu_ready_for_response and 
						((not icache_response_is_awaited) or icache_response_ready))  else '0';

	
	--------------------------------------------------------------------------------
	-- reverse path logic.
	--------------------------------------------------------------------------------
	icache_response_accept <=  pending_queue_has_data and cpu_ready_for_response and icache_response_is_awaited;
	cpu_response_ready <= (pending_queue_has_data and 
						((not icache_response_is_awaited) or icache_response_ready));

	process(clk, reset)
		variable a32: std_logic_vector(31 downto 0);
	begin

		if(clk'event and clk = '1') then
			if((reset = '0') and cpu_response_ready and cpu_ready_for_response) then
				a32(2 downto 0) := (others => '0');
				a32(31 downto 3) := insert_addr;
				assert false report "IBUFFER " & Convert_SLV_To_Hex_String (core_id) & " " 
						& Convert_SLV_To_Hex_String(cpu_id) & " " 
						& Convert_SLV_To_Hex_String(a32) & " "
						& Convert_SLV_to_Hex_String(ipair_to_cpu) & " " 
						& Convert_To_String(is_tlb_hit_qualified)
					severity note;
			end if;
		end if;
	end process;

	-- insert information..
	-- 18     1          3   2        1  1     64
	-- fsr   cacheable  acc unused   err mae   ipair
	acc_from_icache_response <= icache_response_data (70 downto 68);
	ipair_from_icache_response <= icache_response_data (63 downto 0);
	fsr_from_icache_response <= icache_response_data (89 downto 72);
	mae_8_from_icache_response <= icache_response_data (71 downto 64);

	-- insert addr indicated by pending queue.
	insert_addr <= pending_queue_pop_data((64 + 29 - 1)  downto 64);

	-- acc ipair from the icache response..
	insert_data <= acc_from_icache_response & ipair_from_icache_response;

	icache_response_is_awaited <= pending_queue_has_data and (pending_queue_pop_data(93) = '0');
	ipair_from_pending_queue <= pending_queue_pop_data (63 downto 0);

	-- icache response must be cacheable, without mae.
	is_cacheable_non_mae_icache_response <= 
		(icache_response_data (71) = '1') and
			(icache_response_data (65) = '0') and
			(icache_response_data (64) = '0');
			

	-- Response is either from icache or from pending queue..

	-- fsr? non-zero only from icache.
	fsr_to_cpu <= fsr_from_icache_response when  icache_response_is_awaited else (others => '0');

	-- mae? from icache or indicate ibuf hit and cache hit from lookup.
	mae_8_from_lookup <= "00001100";
	mae_8_to_cpu <= mae_8_from_icache_response when icache_response_is_awaited else mae_8_from_lookup;

	-- ipair? from icache or from pending queue.
	ipair_to_cpu <= ipair_from_icache_response when icache_response_is_awaited else ipair_from_pending_queue;

    	cpu_response_data <= fsr_to_cpu & mae_8_to_cpu & ipair_to_cpu;
			
	
end instruction_buffer_arch;

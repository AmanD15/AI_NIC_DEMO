-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.nic_system_global_package.all;
entity AccessRegister is -- 
  generic (tag_length : integer); 
  port ( -- 
    rwbar : in  std_logic_vector(0 downto 0);
    bmask : in  std_logic_vector(3 downto 0);
    register_index : in  std_logic_vector(5 downto 0);
    wdata : in  std_logic_vector(31 downto 0);
    rdata : out  std_logic_vector(31 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity AccessRegister;
architecture AccessRegister_arch of AccessRegister is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 43)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rwbar_buffer :  std_logic_vector(0 downto 0);
  signal rwbar_update_enable: Boolean;
  signal bmask_buffer :  std_logic_vector(3 downto 0);
  signal bmask_update_enable: Boolean;
  signal register_index_buffer :  std_logic_vector(5 downto 0);
  signal register_index_update_enable: Boolean;
  signal wdata_buffer :  std_logic_vector(31 downto 0);
  signal wdata_update_enable: Boolean;
  -- output port buffer signals
  signal rdata_buffer :  std_logic_vector(31 downto 0);
  signal rdata_update_enable: Boolean;
  signal AccessRegister_CP_0_start: Boolean;
  signal AccessRegister_CP_0_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_203_inst_req_0 : boolean;
  signal WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_203_inst_ack_0 : boolean;
  signal WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_203_inst_req_1 : boolean;
  signal WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_203_inst_ack_1 : boolean;
  signal RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_208_inst_req_0 : boolean;
  signal RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_208_inst_ack_0 : boolean;
  signal RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_208_inst_req_1 : boolean;
  signal RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_208_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "AccessRegister_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 43) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= rwbar;
  rwbar_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(4 downto 1) <= bmask;
  bmask_buffer <= in_buffer_data_out(4 downto 1);
  in_buffer_data_in(10 downto 5) <= register_index;
  register_index_buffer <= in_buffer_data_out(10 downto 5);
  in_buffer_data_in(42 downto 11) <= wdata;
  wdata_buffer <= in_buffer_data_out(42 downto 11);
  in_buffer_data_in(tag_length + 42 downto 43) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 42 downto 43);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  AccessRegister_CP_0_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "AccessRegister_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= rdata_buffer;
  rdata <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= AccessRegister_CP_0_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= AccessRegister_CP_0_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= AccessRegister_CP_0_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  AccessRegister_CP_0: Block -- control-path 
    signal AccessRegister_CP_0_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    AccessRegister_CP_0_elements(0) <= AccessRegister_CP_0_start;
    AccessRegister_CP_0_symbol <= AccessRegister_CP_0_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_197_to_assign_stmt_215/$entry
      -- CP-element group 0: 	 assign_stmt_197_to_assign_stmt_215/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_203_sample_start_
      -- CP-element group 0: 	 assign_stmt_197_to_assign_stmt_215/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_203_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_197_to_assign_stmt_215/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_203_Sample/req
      -- CP-element group 0: 	 assign_stmt_197_to_assign_stmt_215/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_208_sample_start_
      -- CP-element group 0: 	 assign_stmt_197_to_assign_stmt_215/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_208_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_197_to_assign_stmt_215/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_208_Sample/rr
      -- 
    req_13_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_13_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AccessRegister_CP_0_elements(0), ack => WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_203_inst_req_0); -- 
    rr_27_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_27_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AccessRegister_CP_0_elements(0), ack => RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_208_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_197_to_assign_stmt_215/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_203_sample_completed_
      -- CP-element group 1: 	 assign_stmt_197_to_assign_stmt_215/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_203_update_start_
      -- CP-element group 1: 	 assign_stmt_197_to_assign_stmt_215/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_203_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_197_to_assign_stmt_215/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_203_Sample/ack
      -- CP-element group 1: 	 assign_stmt_197_to_assign_stmt_215/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_203_Update/$entry
      -- CP-element group 1: 	 assign_stmt_197_to_assign_stmt_215/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_203_Update/req
      -- 
    ack_14_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_203_inst_ack_0, ack => AccessRegister_CP_0_elements(1)); -- 
    req_18_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_18_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AccessRegister_CP_0_elements(1), ack => WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_203_inst_req_1); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_197_to_assign_stmt_215/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_203_update_completed_
      -- CP-element group 2: 	 assign_stmt_197_to_assign_stmt_215/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_203_Update/$exit
      -- CP-element group 2: 	 assign_stmt_197_to_assign_stmt_215/WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_203_Update/ack
      -- 
    ack_19_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_203_inst_ack_1, ack => AccessRegister_CP_0_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 assign_stmt_197_to_assign_stmt_215/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_208_sample_completed_
      -- CP-element group 3: 	 assign_stmt_197_to_assign_stmt_215/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_208_update_start_
      -- CP-element group 3: 	 assign_stmt_197_to_assign_stmt_215/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_208_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_197_to_assign_stmt_215/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_208_Sample/ra
      -- CP-element group 3: 	 assign_stmt_197_to_assign_stmt_215/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_208_Update/$entry
      -- CP-element group 3: 	 assign_stmt_197_to_assign_stmt_215/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_208_Update/cr
      -- 
    ra_28_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_208_inst_ack_0, ack => AccessRegister_CP_0_elements(3)); -- 
    cr_32_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_32_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AccessRegister_CP_0_elements(3), ack => RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_208_inst_req_1); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 assign_stmt_197_to_assign_stmt_215/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_208_update_completed_
      -- CP-element group 4: 	 assign_stmt_197_to_assign_stmt_215/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_208_Update/$exit
      -- CP-element group 4: 	 assign_stmt_197_to_assign_stmt_215/RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_208_Update/ca
      -- 
    ca_33_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_208_inst_ack_1, ack => AccessRegister_CP_0_elements(4)); -- 
    -- CP-element group 5:  join  transition  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 $exit
      -- CP-element group 5: 	 assign_stmt_197_to_assign_stmt_215/$exit
      -- 
    AccessRegister_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "AccessRegister_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= AccessRegister_CP_0_elements(2) & AccessRegister_CP_0_elements(4);
      gj_AccessRegister_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => AccessRegister_CP_0_elements(5), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u1_u5_192_wire : std_logic_vector(4 downto 0);
    signal CONCAT_u6_u38_195_wire : std_logic_vector(37 downto 0);
    signal request_197 : std_logic_vector(42 downto 0);
    signal response_209 : std_logic_vector(32 downto 0);
    -- 
  begin -- 
    -- flow-through slice operator slice_214_inst
    rdata_buffer <= response_209(31 downto 0);
    -- binary operator CONCAT_u1_u5_192_inst
    process(rwbar_buffer, bmask_buffer) -- 
      variable tmp_var : std_logic_vector(4 downto 0); -- 
    begin -- 
      ApConcat_proc(rwbar_buffer, bmask_buffer, tmp_var);
      CONCAT_u1_u5_192_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u5_u43_196_inst
    process(CONCAT_u1_u5_192_wire, CONCAT_u6_u38_195_wire) -- 
      variable tmp_var : std_logic_vector(42 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u5_192_wire, CONCAT_u6_u38_195_wire, tmp_var);
      request_197 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u6_u38_195_inst
    process(register_index_buffer, wdata_buffer) -- 
      variable tmp_var : std_logic_vector(37 downto 0); -- 
    begin -- 
      ApConcat_proc(register_index_buffer, wdata_buffer, tmp_var);
      CONCAT_u6_u38_195_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_208_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(32 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_208_inst_req_0;
      RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_208_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_208_inst_req_1;
      RPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_208_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      response_209 <= data_out(32 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_read_0_gI: SplitGuardInterface generic map(name => "NIC_RESPONSE_REGISTER_ACCESS_PIPE_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_read_0: InputPortRevised -- 
        generic map ( name => "NIC_RESPONSE_REGISTER_ACCESS_PIPE_read_0", data_width => 33,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req(0),
          oack => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack(0),
          odata => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data(32 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_203_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(42 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_203_inst_req_0;
      WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_203_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_203_inst_req_1;
      WPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_203_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= request_197;
      NIC_REQUEST_REGISTER_ACCESS_PIPE_write_0_gI: SplitGuardInterface generic map(name => "NIC_REQUEST_REGISTER_ACCESS_PIPE_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      NIC_REQUEST_REGISTER_ACCESS_PIPE_write_0: OutputPortRevised -- 
        generic map ( name => "NIC_REQUEST_REGISTER_ACCESS_PIPE", data_width => 43, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req(0),
          oack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack(0),
          odata => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data(42 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end AccessRegister_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.nic_system_global_package.all;
entity NicRegisterAccessDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(5 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(5 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(2 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(42 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(32 downto 0);
    MAC_ENABLE_pipe_write_req : out  std_logic_vector(0 downto 0);
    MAC_ENABLE_pipe_write_ack : in   std_logic_vector(0 downto 0);
    MAC_ENABLE_pipe_write_data : out  std_logic_vector(0 downto 0);
    UpdateRegister_call_reqs : out  std_logic_vector(0 downto 0);
    UpdateRegister_call_acks : in   std_logic_vector(0 downto 0);
    UpdateRegister_call_data : out  std_logic_vector(73 downto 0);
    UpdateRegister_call_tag  :  out  std_logic_vector(0 downto 0);
    UpdateRegister_return_reqs : out  std_logic_vector(0 downto 0);
    UpdateRegister_return_acks : in   std_logic_vector(0 downto 0);
    UpdateRegister_return_data : in   std_logic_vector(31 downto 0);
    UpdateRegister_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity NicRegisterAccessDaemon;
architecture NicRegisterAccessDaemon_arch of NicRegisterAccessDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal NicRegisterAccessDaemon_CP_516_start: Boolean;
  signal NicRegisterAccessDaemon_CP_516_symbol: Boolean;
  -- volatile/operator module components. 
  component UpdateRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      bmask : in  std_logic_vector(3 downto 0);
      rval : in  std_logic_vector(31 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      index : in  std_logic_vector(5 downto 0);
      wval : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(5 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal MUX_428_inst_ack_1 : boolean;
  signal phi_stmt_405_ack_0 : boolean;
  signal phi_stmt_405_req_1 : boolean;
  signal nI_421_410_buf_ack_1 : boolean;
  signal nI_421_410_buf_req_1 : boolean;
  signal nI_421_410_buf_ack_0 : boolean;
  signal nI_421_410_buf_req_0 : boolean;
  signal phi_stmt_405_req_0 : boolean;
  signal MUX_428_inst_req_1 : boolean;
  signal if_stmt_430_branch_ack_0 : boolean;
  signal if_stmt_430_branch_ack_1 : boolean;
  signal if_stmt_430_branch_req_0 : boolean;
  signal RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_442_inst_ack_1 : boolean;
  signal RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_442_inst_ack_0 : boolean;
  signal MUX_428_inst_ack_0 : boolean;
  signal RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_442_inst_req_1 : boolean;
  signal MUX_428_inst_req_0 : boolean;
  signal WPIPE_MAC_ENABLE_422_inst_ack_0 : boolean;
  signal WPIPE_MAC_ENABLE_422_inst_req_0 : boolean;
  signal array_obj_ref_413_store_0_ack_1 : boolean;
  signal array_obj_ref_413_store_0_req_1 : boolean;
  signal RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_442_inst_req_0 : boolean;
  signal do_while_stmt_439_branch_req_0 : boolean;
  signal WPIPE_MAC_ENABLE_422_inst_ack_1 : boolean;
  signal array_obj_ref_413_store_0_ack_0 : boolean;
  signal WPIPE_MAC_ENABLE_422_inst_req_1 : boolean;
  signal array_obj_ref_413_store_0_req_0 : boolean;
  signal array_obj_ref_463_load_0_req_0 : boolean;
  signal array_obj_ref_463_load_0_ack_0 : boolean;
  signal array_obj_ref_463_load_0_req_1 : boolean;
  signal array_obj_ref_463_load_0_ack_1 : boolean;
  signal W_rwbar_468_delayed_5_0_468_inst_req_0 : boolean;
  signal W_rwbar_468_delayed_5_0_468_inst_ack_0 : boolean;
  signal W_rwbar_468_delayed_5_0_468_inst_req_1 : boolean;
  signal W_rwbar_468_delayed_5_0_468_inst_ack_1 : boolean;
  signal W_bmask_469_delayed_5_0_471_inst_req_0 : boolean;
  signal W_bmask_469_delayed_5_0_471_inst_ack_0 : boolean;
  signal W_bmask_469_delayed_5_0_471_inst_req_1 : boolean;
  signal W_bmask_469_delayed_5_0_471_inst_ack_1 : boolean;
  signal W_wdata_471_delayed_5_0_474_inst_req_0 : boolean;
  signal W_wdata_471_delayed_5_0_474_inst_ack_0 : boolean;
  signal W_wdata_471_delayed_5_0_474_inst_req_1 : boolean;
  signal W_wdata_471_delayed_5_0_474_inst_ack_1 : boolean;
  signal W_index_472_delayed_5_0_477_inst_req_0 : boolean;
  signal W_index_472_delayed_5_0_477_inst_ack_0 : boolean;
  signal W_index_472_delayed_5_0_477_inst_req_1 : boolean;
  signal W_index_472_delayed_5_0_477_inst_ack_1 : boolean;
  signal call_stmt_486_call_req_0 : boolean;
  signal call_stmt_486_call_ack_0 : boolean;
  signal call_stmt_486_call_req_1 : boolean;
  signal call_stmt_486_call_ack_1 : boolean;
  signal W_rwbar_476_delayed_5_0_487_inst_req_0 : boolean;
  signal W_rwbar_476_delayed_5_0_487_inst_ack_0 : boolean;
  signal W_rwbar_476_delayed_5_0_487_inst_req_1 : boolean;
  signal W_rwbar_476_delayed_5_0_487_inst_ack_1 : boolean;
  signal WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_503_inst_req_0 : boolean;
  signal WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_503_inst_ack_0 : boolean;
  signal WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_503_inst_req_1 : boolean;
  signal WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_503_inst_ack_1 : boolean;
  signal do_while_stmt_439_branch_ack_0 : boolean;
  signal do_while_stmt_439_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "NicRegisterAccessDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  NicRegisterAccessDaemon_CP_516_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "NicRegisterAccessDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= NicRegisterAccessDaemon_CP_516_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= NicRegisterAccessDaemon_CP_516_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= NicRegisterAccessDaemon_CP_516_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  NicRegisterAccessDaemon_CP_516: Block -- control-path 
    signal NicRegisterAccessDaemon_CP_516_elements: BooleanArray(65 downto 0);
    -- 
  begin -- 
    NicRegisterAccessDaemon_CP_516_elements(0) <= NicRegisterAccessDaemon_CP_516_start;
    NicRegisterAccessDaemon_CP_516_symbol <= NicRegisterAccessDaemon_CP_516_elements(16);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	10 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 branch_block_stmt_403/merge_stmt_404__entry___PhiReq/phi_stmt_405/phi_stmt_405_sources/$entry
      -- CP-element group 0: 	 branch_block_stmt_403/merge_stmt_404__entry___PhiReq/phi_stmt_405/$entry
      -- CP-element group 0: 	 branch_block_stmt_403/merge_stmt_404__entry___PhiReq/$entry
      -- CP-element group 0: 	 branch_block_stmt_403/merge_stmt_404_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_403/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_403/merge_stmt_404__entry__
      -- CP-element group 0: 	 branch_block_stmt_403/branch_block_stmt_403__entry__
      -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	15 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (5) 
      -- CP-element group 1: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_Sample/word_access_start/word_0/$exit
      -- CP-element group 1: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_Sample/word_access_start/$exit
      -- CP-element group 1: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_Sample/$exit
      -- CP-element group 1: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_Sample/word_access_start/word_0/ra
      -- 
    ra_583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_413_store_0_ack_0, ack => NicRegisterAccessDaemon_CP_516_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	15 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	7 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_Update/word_access_complete/word_0/ca
      -- CP-element group 2: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_Update/word_access_complete/word_0/$exit
      -- CP-element group 2: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_Update/word_access_complete/$exit
      -- CP-element group 2: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_Update/$exit
      -- 
    ca_594_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_413_store_0_ack_1, ack => NicRegisterAccessDaemon_CP_516_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	15 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/MUX_428_start/ack
      -- CP-element group 3: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/MUX_428_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/MUX_428_start/$exit
      -- 
    ack_603_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_428_inst_ack_0, ack => NicRegisterAccessDaemon_CP_516_elements(3)); -- 
    -- CP-element group 4:  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	15 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4:  members (6) 
      -- CP-element group 4: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/MUX_428_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/MUX_428_complete/ack
      -- CP-element group 4: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/MUX_428_complete/$exit
      -- CP-element group 4: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/WPIPE_MAC_ENABLE_422_Sample/req
      -- CP-element group 4: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/WPIPE_MAC_ENABLE_422_Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/WPIPE_MAC_ENABLE_422_sample_start_
      -- 
    ack_608_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_428_inst_ack_1, ack => NicRegisterAccessDaemon_CP_516_elements(4)); -- 
    req_616_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_616_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_516_elements(4), ack => WPIPE_MAC_ENABLE_422_inst_req_0); -- 
    -- CP-element group 5:  transition  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5:  members (6) 
      -- CP-element group 5: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/WPIPE_MAC_ENABLE_422_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/WPIPE_MAC_ENABLE_422_Sample/ack
      -- CP-element group 5: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/WPIPE_MAC_ENABLE_422_Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/WPIPE_MAC_ENABLE_422_update_start_
      -- CP-element group 5: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/WPIPE_MAC_ENABLE_422_sample_completed_
      -- CP-element group 5: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/WPIPE_MAC_ENABLE_422_Update/req
      -- 
    ack_617_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_MAC_ENABLE_422_inst_ack_0, ack => NicRegisterAccessDaemon_CP_516_elements(5)); -- 
    req_621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_516_elements(5), ack => WPIPE_MAC_ENABLE_422_inst_req_1); -- 
    -- CP-element group 6:  transition  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/WPIPE_MAC_ENABLE_422_Update/$exit
      -- CP-element group 6: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/WPIPE_MAC_ENABLE_422_update_completed_
      -- CP-element group 6: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/WPIPE_MAC_ENABLE_422_Update/ack
      -- 
    ack_622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_MAC_ENABLE_422_inst_ack_1, ack => NicRegisterAccessDaemon_CP_516_elements(6)); -- 
    -- CP-element group 7:  branch  join  transition  place  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7: 	9 
    -- CP-element group 7:  members (24) 
      -- CP-element group 7: 	 branch_block_stmt_403/if_stmt_430_eval_test/ULT_u7_u1_433/SplitProtocol/Sample/rr
      -- CP-element group 7: 	 branch_block_stmt_403/if_stmt_430_eval_test/ULT_u7_u1_433/SplitProtocol/Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_403/if_stmt_430_eval_test/ULT_u7_u1_433/ULT_u7_u1_433_inputs/$exit
      -- CP-element group 7: 	 branch_block_stmt_403/if_stmt_430_else_link/$entry
      -- CP-element group 7: 	 branch_block_stmt_403/if_stmt_430_if_link/$entry
      -- CP-element group 7: 	 branch_block_stmt_403/ULT_u7_u1_433_place
      -- CP-element group 7: 	 branch_block_stmt_403/if_stmt_430_eval_test/branch_req
      -- CP-element group 7: 	 branch_block_stmt_403/if_stmt_430_eval_test/ULT_u7_u1_433/SplitProtocol/Update/ca
      -- CP-element group 7: 	 branch_block_stmt_403/if_stmt_430_eval_test/ULT_u7_u1_433/ULT_u7_u1_433_inputs/$entry
      -- CP-element group 7: 	 branch_block_stmt_403/if_stmt_430_eval_test/ULT_u7_u1_433/SplitProtocol/Update/cr
      -- CP-element group 7: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429__exit__
      -- CP-element group 7: 	 branch_block_stmt_403/if_stmt_430_eval_test/ULT_u7_u1_433/SplitProtocol/$exit
      -- CP-element group 7: 	 branch_block_stmt_403/if_stmt_430_dead_link/$entry
      -- CP-element group 7: 	 branch_block_stmt_403/if_stmt_430_eval_test/ULT_u7_u1_433/$entry
      -- CP-element group 7: 	 branch_block_stmt_403/if_stmt_430_eval_test/ULT_u7_u1_433/SplitProtocol/Update/$entry
      -- CP-element group 7: 	 branch_block_stmt_403/if_stmt_430_eval_test/ULT_u7_u1_433/SplitProtocol/Update/$exit
      -- CP-element group 7: 	 branch_block_stmt_403/if_stmt_430_eval_test/ULT_u7_u1_433/SplitProtocol/Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_403/if_stmt_430_eval_test/$exit
      -- CP-element group 7: 	 branch_block_stmt_403/if_stmt_430_eval_test/$entry
      -- CP-element group 7: 	 branch_block_stmt_403/if_stmt_430_eval_test/ULT_u7_u1_433/SplitProtocol/Sample/ra
      -- CP-element group 7: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/$exit
      -- CP-element group 7: 	 branch_block_stmt_403/if_stmt_430__entry__
      -- CP-element group 7: 	 branch_block_stmt_403/if_stmt_430_eval_test/ULT_u7_u1_433/$exit
      -- CP-element group 7: 	 branch_block_stmt_403/if_stmt_430_eval_test/ULT_u7_u1_433/SplitProtocol/$entry
      -- 
    branch_req_649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_516_elements(7), ack => if_stmt_430_branch_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 42) := "NicRegisterAccessDaemon_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_516_elements(2) & NicRegisterAccessDaemon_CP_516_elements(6);
      gj_NicRegisterAccessDaemon_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_516_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  fork  transition  place  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	11 
    -- CP-element group 8: 	12 
    -- CP-element group 8:  members (11) 
      -- CP-element group 8: 	 branch_block_stmt_403/loopback_PhiReq/phi_stmt_405/$entry
      -- CP-element group 8: 	 branch_block_stmt_403/loopback_PhiReq/phi_stmt_405/phi_stmt_405_sources/Interlock/Update/req
      -- CP-element group 8: 	 branch_block_stmt_403/loopback_PhiReq/phi_stmt_405/phi_stmt_405_sources/Interlock/Update/$entry
      -- CP-element group 8: 	 branch_block_stmt_403/loopback_PhiReq/phi_stmt_405/phi_stmt_405_sources/Interlock/Sample/req
      -- CP-element group 8: 	 branch_block_stmt_403/loopback_PhiReq/phi_stmt_405/phi_stmt_405_sources/Interlock/Sample/$entry
      -- CP-element group 8: 	 branch_block_stmt_403/loopback_PhiReq/phi_stmt_405/phi_stmt_405_sources/Interlock/$entry
      -- CP-element group 8: 	 branch_block_stmt_403/loopback_PhiReq/phi_stmt_405/phi_stmt_405_sources/$entry
      -- CP-element group 8: 	 branch_block_stmt_403/loopback_PhiReq/$entry
      -- CP-element group 8: 	 branch_block_stmt_403/loopback
      -- CP-element group 8: 	 branch_block_stmt_403/if_stmt_430_if_link/if_choice_transition
      -- CP-element group 8: 	 branch_block_stmt_403/if_stmt_430_if_link/$exit
      -- 
    if_choice_transition_654_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_430_branch_ack_1, ack => NicRegisterAccessDaemon_CP_516_elements(8)); -- 
    req_695_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_695_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_516_elements(8), ack => nI_421_410_buf_req_1); -- 
    req_690_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_690_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_516_elements(8), ack => nI_421_410_buf_req_0); -- 
    -- CP-element group 9:  merge  transition  place  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	7 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	17 
    -- CP-element group 9:  members (8) 
      -- CP-element group 9: 	 branch_block_stmt_438/$entry
      -- CP-element group 9: 	 branch_block_stmt_438/do_while_stmt_439__entry__
      -- CP-element group 9: 	 branch_block_stmt_438/branch_block_stmt_438__entry__
      -- CP-element group 9: 	 branch_block_stmt_403/if_stmt_430_else_link/else_choice_transition
      -- CP-element group 9: 	 branch_block_stmt_403/if_stmt_430_else_link/$exit
      -- CP-element group 9: 	 branch_block_stmt_403/$exit
      -- CP-element group 9: 	 branch_block_stmt_403/if_stmt_430__exit__
      -- CP-element group 9: 	 branch_block_stmt_403/branch_block_stmt_403__exit__
      -- 
    else_choice_transition_658_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_430_branch_ack_0, ack => NicRegisterAccessDaemon_CP_516_elements(9)); -- 
    -- CP-element group 10:  transition  output  delay-element  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	0 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	14 
    -- CP-element group 10:  members (5) 
      -- CP-element group 10: 	 branch_block_stmt_403/merge_stmt_404__entry___PhiReq/phi_stmt_405/phi_stmt_405_req
      -- CP-element group 10: 	 branch_block_stmt_403/merge_stmt_404__entry___PhiReq/phi_stmt_405/phi_stmt_405_sources/type_cast_409_konst_delay_trans
      -- CP-element group 10: 	 branch_block_stmt_403/merge_stmt_404__entry___PhiReq/phi_stmt_405/phi_stmt_405_sources/$exit
      -- CP-element group 10: 	 branch_block_stmt_403/merge_stmt_404__entry___PhiReq/phi_stmt_405/$exit
      -- CP-element group 10: 	 branch_block_stmt_403/merge_stmt_404__entry___PhiReq/$exit
      -- 
    phi_stmt_405_req_674_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_405_req_674_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_516_elements(10), ack => phi_stmt_405_req_0); -- 
    -- Element group NicRegisterAccessDaemon_CP_516_elements(10) is a control-delay.
    cp_element_10_delay: control_delay_element  generic map(name => " 10_delay", delay_value => 1)  port map(req => NicRegisterAccessDaemon_CP_516_elements(0), ack => NicRegisterAccessDaemon_CP_516_elements(10), clk => clk, reset =>reset);
    -- CP-element group 11:  transition  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	8 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_403/loopback_PhiReq/phi_stmt_405/phi_stmt_405_sources/Interlock/Sample/ack
      -- CP-element group 11: 	 branch_block_stmt_403/loopback_PhiReq/phi_stmt_405/phi_stmt_405_sources/Interlock/Sample/$exit
      -- 
    ack_691_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nI_421_410_buf_ack_0, ack => NicRegisterAccessDaemon_CP_516_elements(11)); -- 
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	8 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (2) 
      -- CP-element group 12: 	 branch_block_stmt_403/loopback_PhiReq/phi_stmt_405/phi_stmt_405_sources/Interlock/Update/ack
      -- CP-element group 12: 	 branch_block_stmt_403/loopback_PhiReq/phi_stmt_405/phi_stmt_405_sources/Interlock/Update/$exit
      -- 
    ack_696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nI_421_410_buf_ack_1, ack => NicRegisterAccessDaemon_CP_516_elements(12)); -- 
    -- CP-element group 13:  join  transition  output  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 branch_block_stmt_403/loopback_PhiReq/phi_stmt_405/$exit
      -- CP-element group 13: 	 branch_block_stmt_403/loopback_PhiReq/phi_stmt_405/phi_stmt_405_req
      -- CP-element group 13: 	 branch_block_stmt_403/loopback_PhiReq/phi_stmt_405/phi_stmt_405_sources/Interlock/$exit
      -- CP-element group 13: 	 branch_block_stmt_403/loopback_PhiReq/phi_stmt_405/phi_stmt_405_sources/$exit
      -- CP-element group 13: 	 branch_block_stmt_403/loopback_PhiReq/$exit
      -- 
    phi_stmt_405_req_697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_405_req_697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_516_elements(13), ack => phi_stmt_405_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_516_elements(11) & NicRegisterAccessDaemon_CP_516_elements(12);
      gj_NicRegisterAccessDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_516_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  merge  transition  place  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_403/merge_stmt_404_PhiAck/$entry
      -- CP-element group 14: 	 branch_block_stmt_403/merge_stmt_404_PhiReqMerge
      -- 
    NicRegisterAccessDaemon_CP_516_elements(14) <= OrReduce(NicRegisterAccessDaemon_CP_516_elements(10) & NicRegisterAccessDaemon_CP_516_elements(13));
    -- CP-element group 15:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: 	3 
    -- CP-element group 15: 	4 
    -- CP-element group 15: 	1 
    -- CP-element group 15:  members (51) 
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/MUX_428_update_start_
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_final_index_sum_regn/$exit
      -- CP-element group 15: 	 branch_block_stmt_403/merge_stmt_404_PhiAck/phi_stmt_405_ack
      -- CP-element group 15: 	 branch_block_stmt_403/merge_stmt_404_PhiAck/$exit
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/MUX_428_complete/req
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/MUX_428_complete/$entry
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_word_addrgen/root_register_ack
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_final_index_sum_regn/$entry
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_root_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_index_scaled_0
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_word_address_calculated
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_index_scale_0/scale_rename_ack
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_index_scale_0/scale_rename_req
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_update_start_
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_Sample/word_access_start/word_0/$entry
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_Sample/word_access_start/$entry
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/MUX_428_start/req
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_Sample/array_obj_ref_413_Split/split_ack
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_Sample/array_obj_ref_413_Split/split_req
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_Sample/array_obj_ref_413_Split/$exit
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_Sample/array_obj_ref_413_Split/$entry
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_index_scale_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_Sample/$entry
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/$entry
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/MUX_428_sample_start_
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_index_scale_0/$entry
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_word_addrgen/root_register_req
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_index_resized_0
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_word_addrgen/$exit
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_word_addrgen/$entry
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_base_plus_offset/sum_rename_ack
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429__entry__
      -- CP-element group 15: 	 branch_block_stmt_403/merge_stmt_404__exit__
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_base_plus_offset/sum_rename_req
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_Update/word_access_complete/word_0/cr
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_base_plus_offset/$exit
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/MUX_428_start/$entry
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_base_plus_offset/$entry
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_index_resize_0/index_resize_ack
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_offset_calculated
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_Update/word_access_complete/word_0/$entry
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_index_resize_0/index_resize_req
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_Update/word_access_complete/$entry
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_index_resize_0/$exit
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_index_resize_0/$entry
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_index_computed_0
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_final_index_sum_regn/ack
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_Sample/word_access_start/word_0/rr
      -- CP-element group 15: 	 branch_block_stmt_403/assign_stmt_416_to_assign_stmt_429/array_obj_ref_413_final_index_sum_regn/req
      -- 
    phi_stmt_405_ack_702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_405_ack_0, ack => NicRegisterAccessDaemon_CP_516_elements(15)); -- 
    req_607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_516_elements(15), ack => MUX_428_inst_req_1); -- 
    req_602_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_602_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_516_elements(15), ack => MUX_428_inst_req_0); -- 
    cr_593_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_593_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_516_elements(15), ack => array_obj_ref_413_store_0_req_1); -- 
    rr_582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_516_elements(15), ack => array_obj_ref_413_store_0_req_0); -- 
    -- CP-element group 16:  transition  place  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	65 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (4) 
      -- CP-element group 16: 	 branch_block_stmt_438/$exit
      -- CP-element group 16: 	 branch_block_stmt_438/do_while_stmt_439__exit__
      -- CP-element group 16: 	 branch_block_stmt_438/branch_block_stmt_438__exit__
      -- CP-element group 16: 	 $exit
      -- 
    NicRegisterAccessDaemon_CP_516_elements(16) <= NicRegisterAccessDaemon_CP_516_elements(65);
    -- CP-element group 17:  transition  place  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	9 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	23 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439__entry__
      -- CP-element group 17: 	 branch_block_stmt_438/do_while_stmt_439/$entry
      -- 
    NicRegisterAccessDaemon_CP_516_elements(17) <= NicRegisterAccessDaemon_CP_516_elements(9);
    -- CP-element group 18:  merge  place  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	65 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439__exit__
      -- 
    -- Element group NicRegisterAccessDaemon_CP_516_elements(18) is bound as output of CP function.
    -- CP-element group 19:  merge  place  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	22 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_438/do_while_stmt_439/loop_back
      -- 
    -- Element group NicRegisterAccessDaemon_CP_516_elements(19) is bound as output of CP function.
    -- CP-element group 20:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	60 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	63 
    -- CP-element group 20: 	64 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_438/do_while_stmt_439/condition_done
      -- CP-element group 20: 	 branch_block_stmt_438/do_while_stmt_439/loop_exit/$entry
      -- CP-element group 20: 	 branch_block_stmt_438/do_while_stmt_439/loop_taken/$entry
      -- 
    NicRegisterAccessDaemon_CP_516_elements(20) <= NicRegisterAccessDaemon_CP_516_elements(60);
    -- CP-element group 21:  branch  place  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	62 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_438/do_while_stmt_439/loop_body_done
      -- 
    NicRegisterAccessDaemon_CP_516_elements(21) <= NicRegisterAccessDaemon_CP_516_elements(62);
    -- CP-element group 22:  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/back_edge_to_loop_body
      -- 
    NicRegisterAccessDaemon_CP_516_elements(22) <= NicRegisterAccessDaemon_CP_516_elements(19);
    -- CP-element group 23:  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	17 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/first_time_through_loop_body
      -- 
    NicRegisterAccessDaemon_CP_516_elements(23) <= NicRegisterAccessDaemon_CP_516_elements(17);
    -- CP-element group 24:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	25 
    -- CP-element group 24: 	60 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/$entry
      -- CP-element group 24: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/loop_body_start
      -- 
    -- Element group NicRegisterAccessDaemon_CP_516_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	24 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	28 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_442_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_442_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_442_Sample/rr
      -- 
    rr_733_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_733_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_516_elements(25), ack => RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_442_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_516_elements(24) & NicRegisterAccessDaemon_CP_516_elements(28);
      gj_NicRegisterAccessDaemon_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_516_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	27 
    -- CP-element group 26: marked-predecessors 
    -- CP-element group 26: 	31 
    -- CP-element group 26: 	35 
    -- CP-element group 26: 	39 
    -- CP-element group 26: 	43 
    -- CP-element group 26: 	47 
    -- CP-element group 26: 	55 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_442_update_start_
      -- CP-element group 26: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_442_Update/cr
      -- CP-element group 26: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_442_Update/$entry
      -- 
    cr_738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_516_elements(26), ack => RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_442_inst_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_516_elements(27) & NicRegisterAccessDaemon_CP_516_elements(31) & NicRegisterAccessDaemon_CP_516_elements(35) & NicRegisterAccessDaemon_CP_516_elements(39) & NicRegisterAccessDaemon_CP_516_elements(43) & NicRegisterAccessDaemon_CP_516_elements(47) & NicRegisterAccessDaemon_CP_516_elements(55);
      gj_NicRegisterAccessDaemon_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_516_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	26 
    -- CP-element group 27:  members (3) 
      -- CP-element group 27: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_442_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_442_Sample/ra
      -- CP-element group 27: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_442_Sample/$exit
      -- 
    ra_734_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_442_inst_ack_0, ack => NicRegisterAccessDaemon_CP_516_elements(27)); -- 
    -- CP-element group 28:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	29 
    -- CP-element group 28: 	33 
    -- CP-element group 28: 	37 
    -- CP-element group 28: 	41 
    -- CP-element group 28: 	45 
    -- CP-element group 28: 	53 
    -- CP-element group 28: marked-successors 
    -- CP-element group 28: 	25 
    -- CP-element group 28:  members (29) 
      -- CP-element group 28: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_final_index_sum_regn/ack
      -- CP-element group 28: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_index_resize_0/$entry
      -- CP-element group 28: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_index_resize_0/$exit
      -- CP-element group 28: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_442_Update/ca
      -- CP-element group 28: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_index_scale_0/scale_rename_req
      -- CP-element group 28: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_index_scale_0/$entry
      -- CP-element group 28: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_index_scale_0/$exit
      -- CP-element group 28: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_index_scale_0/scale_rename_ack
      -- CP-element group 28: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_base_plus_offset/sum_rename_req
      -- CP-element group 28: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_base_plus_offset/sum_rename_ack
      -- CP-element group 28: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_word_addrgen/$entry
      -- CP-element group 28: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_word_addrgen/$exit
      -- CP-element group 28: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_word_addrgen/root_register_req
      -- CP-element group 28: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_index_resize_0/index_resize_ack
      -- CP-element group 28: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_root_address_calculated
      -- CP-element group 28: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_offset_calculated
      -- CP-element group 28: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_442_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_base_plus_offset/$entry
      -- CP-element group 28: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_base_plus_offset/$exit
      -- CP-element group 28: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_index_scaled_0
      -- CP-element group 28: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_442_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_final_index_sum_regn/$entry
      -- CP-element group 28: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_index_resized_0
      -- CP-element group 28: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_index_resize_0/index_resize_req
      -- CP-element group 28: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_index_computed_0
      -- CP-element group 28: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_final_index_sum_regn/$exit
      -- CP-element group 28: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_final_index_sum_regn/req
      -- CP-element group 28: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_word_address_calculated
      -- CP-element group 28: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_word_addrgen/root_register_ack
      -- 
    ca_739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_442_inst_ack_1, ack => NicRegisterAccessDaemon_CP_516_elements(28)); -- 
    -- CP-element group 29:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	28 
    -- CP-element group 29: marked-predecessors 
    -- CP-element group 29: 	31 
    -- CP-element group 29: 	52 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (5) 
      -- CP-element group 29: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_sample_start_
      -- CP-element group 29: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_Sample/$entry
      -- CP-element group 29: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_Sample/word_access_start/$entry
      -- CP-element group 29: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_Sample/word_access_start/word_0/$entry
      -- CP-element group 29: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_Sample/word_access_start/word_0/rr
      -- 
    rr_785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_516_elements(29), ack => array_obj_ref_463_load_0_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_516_elements(28) & NicRegisterAccessDaemon_CP_516_elements(31) & NicRegisterAccessDaemon_CP_516_elements(52);
      gj_NicRegisterAccessDaemon_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_516_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	32 
    -- CP-element group 30: 	51 
    -- CP-element group 30: 	58 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (5) 
      -- CP-element group 30: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_update_start_
      -- CP-element group 30: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_Update/$entry
      -- CP-element group 30: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_Update/word_access_complete/$entry
      -- CP-element group 30: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_Update/word_access_complete/word_0/$entry
      -- CP-element group 30: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_Update/word_access_complete/word_0/cr
      -- 
    cr_796_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_796_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_516_elements(30), ack => array_obj_ref_463_load_0_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_516_elements(32) & NicRegisterAccessDaemon_CP_516_elements(51) & NicRegisterAccessDaemon_CP_516_elements(58);
      gj_NicRegisterAccessDaemon_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_516_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	61 
    -- CP-element group 31: marked-successors 
    -- CP-element group 31: 	26 
    -- CP-element group 31: 	29 
    -- CP-element group 31:  members (5) 
      -- CP-element group 31: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_sample_completed_
      -- CP-element group 31: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_Sample/$exit
      -- CP-element group 31: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_Sample/word_access_start/$exit
      -- CP-element group 31: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_Sample/word_access_start/word_0/$exit
      -- CP-element group 31: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_Sample/word_access_start/word_0/ra
      -- 
    ra_786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_463_load_0_ack_0, ack => NicRegisterAccessDaemon_CP_516_elements(31)); -- 
    -- CP-element group 32:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	49 
    -- CP-element group 32: 	57 
    -- CP-element group 32: marked-successors 
    -- CP-element group 32: 	30 
    -- CP-element group 32:  members (9) 
      -- CP-element group 32: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_update_completed_
      -- CP-element group 32: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_Update/$exit
      -- CP-element group 32: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_Update/word_access_complete/$exit
      -- CP-element group 32: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_Update/word_access_complete/word_0/$exit
      -- CP-element group 32: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_Update/word_access_complete/word_0/ca
      -- CP-element group 32: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_Update/array_obj_ref_463_Merge/$entry
      -- CP-element group 32: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_Update/array_obj_ref_463_Merge/$exit
      -- CP-element group 32: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_Update/array_obj_ref_463_Merge/merge_req
      -- CP-element group 32: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_Update/array_obj_ref_463_Merge/merge_ack
      -- 
    ca_797_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_463_load_0_ack_1, ack => NicRegisterAccessDaemon_CP_516_elements(32)); -- 
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	28 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	35 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_470_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_470_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_470_Sample/req
      -- 
    req_810_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_810_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_516_elements(33), ack => W_rwbar_468_delayed_5_0_468_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_516_elements(28) & NicRegisterAccessDaemon_CP_516_elements(35);
      gj_NicRegisterAccessDaemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_516_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	36 
    -- CP-element group 34: 	51 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_470_update_start_
      -- CP-element group 34: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_470_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_470_Update/req
      -- 
    req_815_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_815_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_516_elements(34), ack => W_rwbar_468_delayed_5_0_468_inst_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_516_elements(36) & NicRegisterAccessDaemon_CP_516_elements(51);
      gj_NicRegisterAccessDaemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_516_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: marked-successors 
    -- CP-element group 35: 	26 
    -- CP-element group 35: 	33 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_470_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_470_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_470_Sample/ack
      -- 
    ack_811_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_468_delayed_5_0_468_inst_ack_0, ack => NicRegisterAccessDaemon_CP_516_elements(35)); -- 
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	49 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	34 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_470_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_470_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_470_Update/ack
      -- 
    ack_816_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_468_delayed_5_0_468_inst_ack_1, ack => NicRegisterAccessDaemon_CP_516_elements(36)); -- 
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	28 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_473_sample_start_
      -- CP-element group 37: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_473_Sample/$entry
      -- CP-element group 37: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_473_Sample/req
      -- 
    req_824_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_824_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_516_elements(37), ack => W_bmask_469_delayed_5_0_471_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_516_elements(28) & NicRegisterAccessDaemon_CP_516_elements(39);
      gj_NicRegisterAccessDaemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_516_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	40 
    -- CP-element group 38: 	51 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_473_update_start_
      -- CP-element group 38: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_473_Update/$entry
      -- CP-element group 38: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_473_Update/req
      -- 
    req_829_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_829_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_516_elements(38), ack => W_bmask_469_delayed_5_0_471_inst_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_516_elements(40) & NicRegisterAccessDaemon_CP_516_elements(51);
      gj_NicRegisterAccessDaemon_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_516_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	26 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_473_sample_completed_
      -- CP-element group 39: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_473_Sample/$exit
      -- CP-element group 39: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_473_Sample/ack
      -- 
    ack_825_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bmask_469_delayed_5_0_471_inst_ack_0, ack => NicRegisterAccessDaemon_CP_516_elements(39)); -- 
    -- CP-element group 40:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	49 
    -- CP-element group 40: marked-successors 
    -- CP-element group 40: 	38 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_473_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_473_Update/$exit
      -- CP-element group 40: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_473_Update/ack
      -- 
    ack_830_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bmask_469_delayed_5_0_471_inst_ack_1, ack => NicRegisterAccessDaemon_CP_516_elements(40)); -- 
    -- CP-element group 41:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	28 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	43 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	43 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_476_sample_start_
      -- CP-element group 41: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_476_Sample/$entry
      -- CP-element group 41: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_476_Sample/req
      -- 
    req_838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_516_elements(41), ack => W_wdata_471_delayed_5_0_474_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_516_elements(28) & NicRegisterAccessDaemon_CP_516_elements(43);
      gj_NicRegisterAccessDaemon_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_516_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	44 
    -- CP-element group 42: 	51 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	44 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_476_update_start_
      -- CP-element group 42: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_476_Update/$entry
      -- CP-element group 42: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_476_Update/req
      -- 
    req_843_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_843_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_516_elements(42), ack => W_wdata_471_delayed_5_0_474_inst_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_516_elements(44) & NicRegisterAccessDaemon_CP_516_elements(51);
      gj_NicRegisterAccessDaemon_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_516_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43: marked-successors 
    -- CP-element group 43: 	26 
    -- CP-element group 43: 	41 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_476_sample_completed_
      -- CP-element group 43: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_476_Sample/$exit
      -- CP-element group 43: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_476_Sample/ack
      -- 
    ack_839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_wdata_471_delayed_5_0_474_inst_ack_0, ack => NicRegisterAccessDaemon_CP_516_elements(43)); -- 
    -- CP-element group 44:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	49 
    -- CP-element group 44: marked-successors 
    -- CP-element group 44: 	42 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_476_update_completed_
      -- CP-element group 44: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_476_Update/$exit
      -- CP-element group 44: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_476_Update/ack
      -- 
    ack_844_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_wdata_471_delayed_5_0_474_inst_ack_1, ack => NicRegisterAccessDaemon_CP_516_elements(44)); -- 
    -- CP-element group 45:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	28 
    -- CP-element group 45: marked-predecessors 
    -- CP-element group 45: 	47 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	47 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_479_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_479_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_479_Sample/req
      -- 
    req_852_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_852_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_516_elements(45), ack => W_index_472_delayed_5_0_477_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_516_elements(28) & NicRegisterAccessDaemon_CP_516_elements(47);
      gj_NicRegisterAccessDaemon_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_516_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: marked-predecessors 
    -- CP-element group 46: 	48 
    -- CP-element group 46: 	51 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_479_update_start_
      -- CP-element group 46: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_479_Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_479_Update/req
      -- 
    req_857_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_857_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_516_elements(46), ack => W_index_472_delayed_5_0_477_inst_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_516_elements(48) & NicRegisterAccessDaemon_CP_516_elements(51);
      gj_NicRegisterAccessDaemon_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_516_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	45 
    -- CP-element group 47: successors 
    -- CP-element group 47: marked-successors 
    -- CP-element group 47: 	26 
    -- CP-element group 47: 	45 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_479_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_479_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_479_Sample/ack
      -- 
    ack_853_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_index_472_delayed_5_0_477_inst_ack_0, ack => NicRegisterAccessDaemon_CP_516_elements(47)); -- 
    -- CP-element group 48:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	49 
    -- CP-element group 48: marked-successors 
    -- CP-element group 48: 	46 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_479_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_479_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_479_Update/ack
      -- 
    ack_858_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_index_472_delayed_5_0_477_inst_ack_1, ack => NicRegisterAccessDaemon_CP_516_elements(48)); -- 
    -- CP-element group 49:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	32 
    -- CP-element group 49: 	36 
    -- CP-element group 49: 	40 
    -- CP-element group 49: 	44 
    -- CP-element group 49: 	48 
    -- CP-element group 49: 	61 
    -- CP-element group 49: marked-predecessors 
    -- CP-element group 49: 	51 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/call_stmt_486_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/call_stmt_486_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/call_stmt_486_Sample/crr
      -- 
    crr_866_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_866_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_516_elements(49), ack => call_stmt_486_call_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 31,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_516_elements(32) & NicRegisterAccessDaemon_CP_516_elements(36) & NicRegisterAccessDaemon_CP_516_elements(40) & NicRegisterAccessDaemon_CP_516_elements(44) & NicRegisterAccessDaemon_CP_516_elements(48) & NicRegisterAccessDaemon_CP_516_elements(61) & NicRegisterAccessDaemon_CP_516_elements(51);
      gj_NicRegisterAccessDaemon_cp_element_group_49 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_516_elements(49), clk => clk, reset => reset); --
    end block;
    -- CP-element group 50:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: marked-predecessors 
    -- CP-element group 50: 	52 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/call_stmt_486_update_start_
      -- CP-element group 50: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/call_stmt_486_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/call_stmt_486_Update/ccr
      -- 
    ccr_871_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_871_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_516_elements(50), ack => call_stmt_486_call_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= NicRegisterAccessDaemon_CP_516_elements(52);
      gj_NicRegisterAccessDaemon_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_516_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: marked-successors 
    -- CP-element group 51: 	30 
    -- CP-element group 51: 	34 
    -- CP-element group 51: 	38 
    -- CP-element group 51: 	42 
    -- CP-element group 51: 	46 
    -- CP-element group 51: 	49 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/call_stmt_486_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/call_stmt_486_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/call_stmt_486_Sample/cra
      -- 
    cra_867_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_486_call_ack_0, ack => NicRegisterAccessDaemon_CP_516_elements(51)); -- 
    -- CP-element group 52:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	62 
    -- CP-element group 52: marked-successors 
    -- CP-element group 52: 	29 
    -- CP-element group 52: 	50 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/call_stmt_486_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/call_stmt_486_Update/$exit
      -- CP-element group 52: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/call_stmt_486_Update/cca
      -- CP-element group 52: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/ring_reenable_memory_space_2
      -- 
    cca_872_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_486_call_ack_1, ack => NicRegisterAccessDaemon_CP_516_elements(52)); -- 
    -- CP-element group 53:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	28 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	55 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_489_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_489_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_489_Sample/req
      -- 
    req_880_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_880_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_516_elements(53), ack => W_rwbar_476_delayed_5_0_487_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_516_elements(28) & NicRegisterAccessDaemon_CP_516_elements(55);
      gj_NicRegisterAccessDaemon_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_516_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	56 
    -- CP-element group 54: 	58 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_489_update_start_
      -- CP-element group 54: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_489_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_489_Update/req
      -- 
    req_885_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_885_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_516_elements(54), ack => W_rwbar_476_delayed_5_0_487_inst_req_1); -- 
    NicRegisterAccessDaemon_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_516_elements(56) & NicRegisterAccessDaemon_CP_516_elements(58);
      gj_NicRegisterAccessDaemon_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_516_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: marked-successors 
    -- CP-element group 55: 	26 
    -- CP-element group 55: 	53 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_489_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_489_Sample/$exit
      -- CP-element group 55: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_489_Sample/ack
      -- 
    ack_881_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_476_delayed_5_0_487_inst_ack_0, ack => NicRegisterAccessDaemon_CP_516_elements(55)); -- 
    -- CP-element group 56:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	57 
    -- CP-element group 56: marked-successors 
    -- CP-element group 56: 	54 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_489_update_completed_
      -- CP-element group 56: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_489_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/assign_stmt_489_Update/ack
      -- 
    ack_886_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_476_delayed_5_0_487_inst_ack_1, ack => NicRegisterAccessDaemon_CP_516_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	32 
    -- CP-element group 57: 	56 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	59 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_503_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_503_Sample/$entry
      -- CP-element group 57: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_503_Sample/req
      -- 
    req_894_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_894_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_516_elements(57), ack => WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_503_inst_req_0); -- 
    NicRegisterAccessDaemon_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_516_elements(32) & NicRegisterAccessDaemon_CP_516_elements(56) & NicRegisterAccessDaemon_CP_516_elements(59);
      gj_NicRegisterAccessDaemon_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_516_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	59 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	30 
    -- CP-element group 58: 	54 
    -- CP-element group 58:  members (6) 
      -- CP-element group 58: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_503_sample_completed_
      -- CP-element group 58: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_503_update_start_
      -- CP-element group 58: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_503_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_503_Sample/ack
      -- CP-element group 58: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_503_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_503_Update/req
      -- 
    ack_895_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_503_inst_ack_0, ack => NicRegisterAccessDaemon_CP_516_elements(58)); -- 
    req_899_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_899_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_516_elements(58), ack => WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_503_inst_req_1); -- 
    -- CP-element group 59:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	58 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	62 
    -- CP-element group 59: marked-successors 
    -- CP-element group 59: 	57 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_503_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_503_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_503_Update/ack
      -- 
    ack_900_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_503_inst_ack_1, ack => NicRegisterAccessDaemon_CP_516_elements(59)); -- 
    -- CP-element group 60:  transition  output  delay-element  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	24 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	20 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/condition_evaluated
      -- CP-element group 60: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/loop_body_delay_to_condition_start
      -- 
    condition_evaluated_724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NicRegisterAccessDaemon_CP_516_elements(60), ack => do_while_stmt_439_branch_req_0); -- 
    -- Element group NicRegisterAccessDaemon_CP_516_elements(60) is a control-delay.
    cp_element_60_delay: control_delay_element  generic map(name => " 60_delay", delay_value => 1)  port map(req => NicRegisterAccessDaemon_CP_516_elements(24), ack => NicRegisterAccessDaemon_CP_516_elements(60), clk => clk, reset =>reset);
    -- CP-element group 61:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	31 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	49 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/array_obj_ref_463_call_stmt_486_delay
      -- 
    -- Element group NicRegisterAccessDaemon_CP_516_elements(61) is a control-delay.
    cp_element_61_delay: control_delay_element  generic map(name => " 61_delay", delay_value => 1)  port map(req => NicRegisterAccessDaemon_CP_516_elements(31), ack => NicRegisterAccessDaemon_CP_516_elements(61), clk => clk, reset =>reset);
    -- CP-element group 62:  join  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	52 
    -- CP-element group 62: 	59 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	21 
    -- CP-element group 62:  members (1) 
      -- CP-element group 62: 	 branch_block_stmt_438/do_while_stmt_439/do_while_stmt_439_loop_body/$exit
      -- 
    NicRegisterAccessDaemon_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 43) := "NicRegisterAccessDaemon_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= NicRegisterAccessDaemon_CP_516_elements(52) & NicRegisterAccessDaemon_CP_516_elements(59);
      gj_NicRegisterAccessDaemon_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => NicRegisterAccessDaemon_CP_516_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	20 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_438/do_while_stmt_439/loop_exit/$exit
      -- CP-element group 63: 	 branch_block_stmt_438/do_while_stmt_439/loop_exit/ack
      -- 
    ack_907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_439_branch_ack_0, ack => NicRegisterAccessDaemon_CP_516_elements(63)); -- 
    -- CP-element group 64:  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	20 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_438/do_while_stmt_439/loop_taken/$exit
      -- CP-element group 64: 	 branch_block_stmt_438/do_while_stmt_439/loop_taken/ack
      -- 
    ack_911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_439_branch_ack_1, ack => NicRegisterAccessDaemon_CP_516_elements(64)); -- 
    -- CP-element group 65:  transition  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	18 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	16 
    -- CP-element group 65:  members (1) 
      -- CP-element group 65: 	 branch_block_stmt_438/do_while_stmt_439/$exit
      -- 
    NicRegisterAccessDaemon_CP_516_elements(65) <= NicRegisterAccessDaemon_CP_516_elements(18);
    NicRegisterAccessDaemon_do_while_stmt_439_terminator_912: loop_terminator -- 
      generic map (name => " NicRegisterAccessDaemon_do_while_stmt_439_terminator_912", max_iterations_in_flight =>31) 
      port map(loop_body_exit => NicRegisterAccessDaemon_CP_516_elements(21),loop_continue => NicRegisterAccessDaemon_CP_516_elements(64),loop_terminate => NicRegisterAccessDaemon_CP_516_elements(63),loop_back => NicRegisterAccessDaemon_CP_516_elements(19),loop_exit => NicRegisterAccessDaemon_CP_516_elements(18),clk => clk, reset => reset); -- 
    entry_tmerge_725_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= NicRegisterAccessDaemon_CP_516_elements(22);
        preds(1)  <= NicRegisterAccessDaemon_CP_516_elements(23);
        entry_tmerge_725 : transition_merge -- 
          generic map(name => " entry_tmerge_725")
          port map (preds => preds, symbol_out => NicRegisterAccessDaemon_CP_516_elements(24));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal EQ_u7_u1_425_wire : std_logic_vector(0 downto 0);
    signal I_405 : std_logic_vector(6 downto 0);
    signal MUX_428_wire : std_logic_vector(0 downto 0);
    signal R_I_412_resized : std_logic_vector(5 downto 0);
    signal R_I_412_scaled : std_logic_vector(5 downto 0);
    signal R_index_462_resized : std_logic_vector(5 downto 0);
    signal R_index_462_scaled : std_logic_vector(5 downto 0);
    signal ULT_u7_u1_433_wire : std_logic_vector(0 downto 0);
    signal array_obj_ref_413_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_413_final_offset : std_logic_vector(5 downto 0);
    signal array_obj_ref_413_offset_scale_factor_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_413_resized_base_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_413_root_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_413_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_413_word_offset_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_463_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_463_final_offset : std_logic_vector(5 downto 0);
    signal array_obj_ref_463_offset_scale_factor_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_463_resized_base_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_463_root_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_463_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_463_word_offset_0 : std_logic_vector(5 downto 0);
    signal bmask_452 : std_logic_vector(3 downto 0);
    signal bmask_469_delayed_5_0_473 : std_logic_vector(3 downto 0);
    signal index_456 : std_logic_vector(5 downto 0);
    signal index_472_delayed_5_0_479 : std_logic_vector(5 downto 0);
    signal konst_419_wire_constant : std_logic_vector(6 downto 0);
    signal konst_424_wire_constant : std_logic_vector(6 downto 0);
    signal konst_426_wire_constant : std_logic_vector(0 downto 0);
    signal konst_427_wire_constant : std_logic_vector(0 downto 0);
    signal konst_432_wire_constant : std_logic_vector(6 downto 0);
    signal konst_507_wire_constant : std_logic_vector(0 downto 0);
    signal nI_421 : std_logic_vector(6 downto 0);
    signal nI_421_410_buffered : std_logic_vector(6 downto 0);
    signal rdata_496 : std_logic_vector(31 downto 0);
    signal req_443 : std_logic_vector(42 downto 0);
    signal resp_502 : std_logic_vector(32 downto 0);
    signal rval_464 : std_logic_vector(31 downto 0);
    signal rwbar_448 : std_logic_vector(0 downto 0);
    signal rwbar_468_delayed_5_0_470 : std_logic_vector(0 downto 0);
    signal rwbar_476_delayed_5_0_489 : std_logic_vector(0 downto 0);
    signal type_cast_409_wire_constant : std_logic_vector(6 downto 0);
    signal type_cast_415_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_494_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_499_wire_constant : std_logic_vector(0 downto 0);
    signal wdata_460 : std_logic_vector(31 downto 0);
    signal wdata_471_delayed_5_0_476 : std_logic_vector(31 downto 0);
    signal wval_486 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_413_offset_scale_factor_0 <= "000001";
    array_obj_ref_413_resized_base_address <= "000000";
    array_obj_ref_413_word_offset_0 <= "000000";
    array_obj_ref_463_offset_scale_factor_0 <= "000001";
    array_obj_ref_463_resized_base_address <= "000000";
    array_obj_ref_463_word_offset_0 <= "000000";
    konst_419_wire_constant <= "0000001";
    konst_424_wire_constant <= "0111111";
    konst_426_wire_constant <= "1";
    konst_427_wire_constant <= "0";
    konst_432_wire_constant <= "0111111";
    konst_507_wire_constant <= "1";
    type_cast_409_wire_constant <= "0000000";
    type_cast_415_wire_constant <= "00000000000000000000000000000000";
    type_cast_494_wire_constant <= "00000000000000000000000000000000";
    type_cast_499_wire_constant <= "0";
    phi_stmt_405: Block -- phi operator 
      signal idata: std_logic_vector(13 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_409_wire_constant & nI_421_410_buffered;
      req <= phi_stmt_405_req_0 & phi_stmt_405_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_405",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 7) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_405_ack_0,
          idata => idata,
          odata => I_405,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_405
    MUX_428_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_428_inst_req_0;
      MUX_428_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_428_inst_req_1;
      MUX_428_inst_ack_1<= update_ack(0);
      MUX_428_inst: SelectSplitProtocol generic map(name => "MUX_428_inst", data_width => 1, buffering => 1, flow_through => false, full_rate => false) -- 
        port map( x => konst_426_wire_constant, y => konst_427_wire_constant, sel => EQ_u7_u1_425_wire, z => MUX_428_wire, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through select operator MUX_495_inst
    rdata_496 <= rval_464 when (rwbar_476_delayed_5_0_489(0) /=  '0') else type_cast_494_wire_constant;
    -- flow-through slice operator slice_447_inst
    rwbar_448 <= req_443(42 downto 42);
    -- flow-through slice operator slice_451_inst
    bmask_452 <= req_443(41 downto 38);
    -- flow-through slice operator slice_455_inst
    index_456 <= req_443(37 downto 32);
    -- flow-through slice operator slice_459_inst
    wdata_460 <= req_443(31 downto 0);
    W_bmask_469_delayed_5_0_471_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_bmask_469_delayed_5_0_471_inst_req_0;
      W_bmask_469_delayed_5_0_471_inst_ack_0<= wack(0);
      rreq(0) <= W_bmask_469_delayed_5_0_471_inst_req_1;
      W_bmask_469_delayed_5_0_471_inst_ack_1<= rack(0);
      W_bmask_469_delayed_5_0_471_inst : InterlockBuffer generic map ( -- 
        name => "W_bmask_469_delayed_5_0_471_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 4,
        out_data_width => 4,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => bmask_452,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => bmask_469_delayed_5_0_473,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_index_472_delayed_5_0_477_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_index_472_delayed_5_0_477_inst_req_0;
      W_index_472_delayed_5_0_477_inst_ack_0<= wack(0);
      rreq(0) <= W_index_472_delayed_5_0_477_inst_req_1;
      W_index_472_delayed_5_0_477_inst_ack_1<= rack(0);
      W_index_472_delayed_5_0_477_inst : InterlockBuffer generic map ( -- 
        name => "W_index_472_delayed_5_0_477_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 6,
        out_data_width => 6,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => index_456,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => index_472_delayed_5_0_479,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rwbar_468_delayed_5_0_468_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rwbar_468_delayed_5_0_468_inst_req_0;
      W_rwbar_468_delayed_5_0_468_inst_ack_0<= wack(0);
      rreq(0) <= W_rwbar_468_delayed_5_0_468_inst_req_1;
      W_rwbar_468_delayed_5_0_468_inst_ack_1<= rack(0);
      W_rwbar_468_delayed_5_0_468_inst : InterlockBuffer generic map ( -- 
        name => "W_rwbar_468_delayed_5_0_468_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rwbar_448,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rwbar_468_delayed_5_0_470,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rwbar_476_delayed_5_0_487_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rwbar_476_delayed_5_0_487_inst_req_0;
      W_rwbar_476_delayed_5_0_487_inst_ack_0<= wack(0);
      rreq(0) <= W_rwbar_476_delayed_5_0_487_inst_req_1;
      W_rwbar_476_delayed_5_0_487_inst_ack_1<= rack(0);
      W_rwbar_476_delayed_5_0_487_inst : InterlockBuffer generic map ( -- 
        name => "W_rwbar_476_delayed_5_0_487_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rwbar_448,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rwbar_476_delayed_5_0_489,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_wdata_471_delayed_5_0_474_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_wdata_471_delayed_5_0_474_inst_req_0;
      W_wdata_471_delayed_5_0_474_inst_ack_0<= wack(0);
      rreq(0) <= W_wdata_471_delayed_5_0_474_inst_req_1;
      W_wdata_471_delayed_5_0_474_inst_ack_1<= rack(0);
      W_wdata_471_delayed_5_0_474_inst : InterlockBuffer generic map ( -- 
        name => "W_wdata_471_delayed_5_0_474_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => wdata_460,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => wdata_471_delayed_5_0_476,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nI_421_410_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nI_421_410_buf_req_0;
      nI_421_410_buf_ack_0<= wack(0);
      rreq(0) <= nI_421_410_buf_req_1;
      nI_421_410_buf_ack_1<= rack(0);
      nI_421_410_buf : InterlockBuffer generic map ( -- 
        name => "nI_421_410_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 7,
        out_data_width => 7,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nI_421,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nI_421_410_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_413_addr_0
    process(array_obj_ref_413_root_address) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_413_root_address;
      ov(5 downto 0) := iv;
      array_obj_ref_413_word_address_0 <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_413_gather_scatter
    process(type_cast_415_wire_constant) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := type_cast_415_wire_constant;
      ov(31 downto 0) := iv;
      array_obj_ref_413_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_413_index_0_rename
    process(R_I_412_resized) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_I_412_resized;
      ov(5 downto 0) := iv;
      R_I_412_scaled <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_413_index_0_resize
    process(I_405) --
      variable iv : std_logic_vector(6 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := I_405;
      ov := iv(5 downto 0);
      R_I_412_resized <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_413_index_offset
    process(R_I_412_scaled) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_I_412_scaled;
      ov(5 downto 0) := iv;
      array_obj_ref_413_final_offset <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_413_root_address_inst
    process(array_obj_ref_413_final_offset) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_413_final_offset;
      ov(5 downto 0) := iv;
      array_obj_ref_413_root_address <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_463_addr_0
    process(array_obj_ref_463_root_address) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_463_root_address;
      ov(5 downto 0) := iv;
      array_obj_ref_463_word_address_0 <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_463_gather_scatter
    process(array_obj_ref_463_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_463_data_0;
      ov(31 downto 0) := iv;
      rval_464 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_463_index_0_rename
    process(R_index_462_resized) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_462_resized;
      ov(5 downto 0) := iv;
      R_index_462_scaled <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_463_index_0_resize
    process(index_456) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := index_456;
      ov(5 downto 0) := iv;
      R_index_462_resized <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_463_index_offset
    process(R_index_462_scaled) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_462_scaled;
      ov(5 downto 0) := iv;
      array_obj_ref_463_final_offset <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_463_root_address_inst
    process(array_obj_ref_463_final_offset) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_463_final_offset;
      ov(5 downto 0) := iv;
      array_obj_ref_463_root_address <= ov(5 downto 0);
      --
    end process;
    do_while_stmt_439_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_507_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_439_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_439_branch_req_0,
          ack0 => do_while_stmt_439_branch_ack_0,
          ack1 => do_while_stmt_439_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_430_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULT_u7_u1_433_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_430_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_430_branch_req_0,
          ack0 => if_stmt_430_branch_ack_0,
          ack1 => if_stmt_430_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u7_u7_420_inst
    process(I_405) -- 
      variable tmp_var : std_logic_vector(6 downto 0); -- 
    begin -- 
      ApIntAdd_proc(I_405, konst_419_wire_constant, tmp_var);
      nI_421 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u33_501_inst
    process(type_cast_499_wire_constant, rdata_496) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_499_wire_constant, rdata_496, tmp_var);
      resp_502 <= tmp_var; --
    end process;
    -- binary operator EQ_u7_u1_425_inst
    process(I_405) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(I_405, konst_424_wire_constant, tmp_var);
      EQ_u7_u1_425_wire <= tmp_var; --
    end process;
    -- binary operator ULT_u7_u1_433_inst
    process(I_405) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(I_405, konst_432_wire_constant, tmp_var);
      ULT_u7_u1_433_wire <= tmp_var; --
    end process;
    -- shared load operator group (0) : array_obj_ref_463_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 5);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_463_load_0_req_0;
      array_obj_ref_463_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_463_load_0_req_1;
      array_obj_ref_463_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_463_word_address_0;
      array_obj_ref_463_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 6,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(5 downto 0),
          mtag => memory_space_2_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 1,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared store operator group (0) : array_obj_ref_413_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(5 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_413_store_0_req_0;
      array_obj_ref_413_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_413_store_0_req_1;
      array_obj_ref_413_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_413_word_address_0;
      data_in <= array_obj_ref_413_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 6,
        data_width => 32,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(5 downto 0),
          mdata => memory_space_2_sr_data(31 downto 0),
          mtag => memory_space_2_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- shared inport operator group (0) : RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_442_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(42 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_442_inst_req_0;
      RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_442_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_442_inst_req_1;
      RPIPE_NIC_REQUEST_REGISTER_ACCESS_PIPE_442_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      req_443 <= data_out(42 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_read_0_gI: SplitGuardInterface generic map(name => "NIC_REQUEST_REGISTER_ACCESS_PIPE_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      NIC_REQUEST_REGISTER_ACCESS_PIPE_read_0: InputPortRevised -- 
        generic map ( name => "NIC_REQUEST_REGISTER_ACCESS_PIPE_read_0", data_width => 43,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req(0),
          oack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack(0),
          odata => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data(42 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_MAC_ENABLE_422_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_MAC_ENABLE_422_inst_req_0;
      WPIPE_MAC_ENABLE_422_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_MAC_ENABLE_422_inst_req_1;
      WPIPE_MAC_ENABLE_422_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= MUX_428_wire;
      MAC_ENABLE_write_0_gI: SplitGuardInterface generic map(name => "MAC_ENABLE_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      MAC_ENABLE_write_0: OutputPortRevised -- 
        generic map ( name => "MAC_ENABLE", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => MAC_ENABLE_pipe_write_req(0),
          oack => MAC_ENABLE_pipe_write_ack(0),
          odata => MAC_ENABLE_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_503_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_503_inst_req_0;
      WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_503_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_503_inst_req_1;
      WPIPE_NIC_RESPONSE_REGISTER_ACCESS_PIPE_503_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= resp_502;
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_write_1_gI: SplitGuardInterface generic map(name => "NIC_RESPONSE_REGISTER_ACCESS_PIPE_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_write_1: OutputPortRevised -- 
        generic map ( name => "NIC_RESPONSE_REGISTER_ACCESS_PIPE", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req(0),
          oack => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack(0),
          odata => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_486_call 
    UpdateRegister_call_group_0: Block -- 
      signal data_in: std_logic_vector(73 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_486_call_req_0;
      call_stmt_486_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_486_call_req_1;
      call_stmt_486_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not rwbar_468_delayed_5_0_470(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      UpdateRegister_call_group_0_gI: SplitGuardInterface generic map(name => "UpdateRegister_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= bmask_469_delayed_5_0_473 & rval_464 & wdata_471_delayed_5_0_476 & index_472_delayed_5_0_479;
      wval_486 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 74,
        owidth => 74,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => UpdateRegister_call_reqs(0),
          ackR => UpdateRegister_call_acks(0),
          dataR => UpdateRegister_call_data(73 downto 0),
          tagR => UpdateRegister_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => UpdateRegister_return_acks(0), -- cross-over
          ackL => UpdateRegister_return_reqs(0), -- cross-over
          dataL => UpdateRegister_return_data(31 downto 0),
          tagL => UpdateRegister_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end NicRegisterAccessDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.nic_system_global_package.all;
entity ReceiveEngineDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    CONTROL_REGISTER : in std_logic_vector(31 downto 0);
    FREE_Q : in std_logic_vector(35 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(5 downto 0);
    AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_call_data : out  std_logic_vector(42 downto 0);
    AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
    AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_return_data : in   std_logic_vector(31 downto 0);
    AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
    popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
    popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
    popFromQueue_call_data : out  std_logic_vector(36 downto 0);
    popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
    popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
    popFromQueue_return_data : in   std_logic_vector(32 downto 0);
    popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
    pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
    pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
    loadBuffer_call_reqs : out  std_logic_vector(0 downto 0);
    loadBuffer_call_acks : in   std_logic_vector(0 downto 0);
    loadBuffer_call_data : out  std_logic_vector(35 downto 0);
    loadBuffer_call_tag  :  out  std_logic_vector(0 downto 0);
    loadBuffer_return_reqs : out  std_logic_vector(0 downto 0);
    loadBuffer_return_acks : in   std_logic_vector(0 downto 0);
    loadBuffer_return_data : in   std_logic_vector(0 downto 0);
    loadBuffer_return_tag :  in   std_logic_vector(0 downto 0);
    populateRxQueue_call_reqs : out  std_logic_vector(0 downto 0);
    populateRxQueue_call_acks : in   std_logic_vector(0 downto 0);
    populateRxQueue_call_data : out  std_logic_vector(35 downto 0);
    populateRxQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    populateRxQueue_return_reqs : out  std_logic_vector(0 downto 0);
    populateRxQueue_return_acks : in   std_logic_vector(0 downto 0);
    populateRxQueue_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity ReceiveEngineDaemon;
architecture ReceiveEngineDaemon_arch of ReceiveEngineDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal ReceiveEngineDaemon_CP_2495_start: Boolean;
  signal ReceiveEngineDaemon_CP_2495_symbol: Boolean;
  -- volatile/operator module components. 
  component AccessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      register_index : in  std_logic_vector(5 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component popFromQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_r_data : out  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_call_acks : in   std_logic_vector(0 downto 0);
      releaseLock_call_data : out  std_logic_vector(35 downto 0);
      releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_return_acks : in   std_logic_vector(0 downto 0);
      releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_call_acks : in   std_logic_vector(0 downto 0);
      acquireLock_call_data : out  std_logic_vector(35 downto 0);
      acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_return_acks : in   std_logic_vector(0 downto 0);
      acquireLock_return_data : in   std_logic_vector(0 downto 0);
      acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      updateTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_data : out  std_logic_vector(67 downto 0);
      updateTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_call_data : out  std_logic_vector(67 downto 0);
      getQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_return_data : in   std_logic_vector(31 downto 0);
      getQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_call_data : out  std_logic_vector(35 downto 0);
      getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
      getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_call_data : out  std_logic_vector(35 downto 0);
      getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_return_data : in   std_logic_vector(31 downto 0);
      getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component pushIntoQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_call_acks : in   std_logic_vector(0 downto 0);
      releaseLock_call_data : out  std_logic_vector(35 downto 0);
      releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_return_acks : in   std_logic_vector(0 downto 0);
      releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_call_acks : in   std_logic_vector(0 downto 0);
      acquireLock_call_data : out  std_logic_vector(35 downto 0);
      acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_return_acks : in   std_logic_vector(0 downto 0);
      acquireLock_return_data : in   std_logic_vector(0 downto 0);
      acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      updateTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_data : out  std_logic_vector(67 downto 0);
      updateTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_call_data : out  std_logic_vector(35 downto 0);
      getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
      getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_call_data : out  std_logic_vector(35 downto 0);
      getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_return_data : in   std_logic_vector(31 downto 0);
      getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_call_data : out  std_logic_vector(99 downto 0);
      setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component loadBuffer is -- 
    generic (tag_length : integer); 
    port ( -- 
      rx_buffer_pointer : in  std_logic_vector(35 downto 0);
      bad_packet_identifier : out  std_logic_vector(0 downto 0);
      writePayloadToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writePayloadToMem_call_acks : in   std_logic_vector(0 downto 0);
      writePayloadToMem_call_data : out  std_logic_vector(71 downto 0);
      writePayloadToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writePayloadToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writePayloadToMem_return_acks : in   std_logic_vector(0 downto 0);
      writePayloadToMem_return_data : in   std_logic_vector(19 downto 0);
      writePayloadToMem_return_tag :  in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_acks : in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_data : out  std_logic_vector(35 downto 0);
      writeEthernetHeaderToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_acks : in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_data : in   std_logic_vector(35 downto 0);
      writeEthernetHeaderToMem_return_tag :  in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_acks : in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_data : out  std_logic_vector(54 downto 0);
      writeControlInformationToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_acks : in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component populateRxQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      rx_buffer_pointer : in  std_logic_vector(35 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX : in std_logic_vector(5 downto 0);
      NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(5 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
      pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal NOT_u1_u1_1789_inst_req_1 : boolean;
  signal NOT_u1_u1_1779_inst_req_0 : boolean;
  signal NOT_u1_u1_1779_inst_ack_0 : boolean;
  signal phi_stmt_1735_req_0 : boolean;
  signal npkt_cnt_1828_1737_buf_ack_0 : boolean;
  signal NOT_u1_u1_1789_inst_ack_1 : boolean;
  signal call_stmt_1759_call_req_0 : boolean;
  signal NOT_u1_u1_1789_inst_req_0 : boolean;
  signal NOT_u1_u1_1789_inst_ack_0 : boolean;
  signal W_pkt_cnt_1778_delayed_13_0_1801_inst_ack_1 : boolean;
  signal W_pkt_cnt_1778_delayed_13_0_1801_inst_req_0 : boolean;
  signal phi_stmt_1735_req_1 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1719_inst_req_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1719_inst_ack_0 : boolean;
  signal phi_stmt_1735_ack_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1719_inst_req_1 : boolean;
  signal W_pkt_cnt_1778_delayed_13_0_1801_inst_ack_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1719_inst_ack_1 : boolean;
  signal do_while_stmt_1733_branch_req_0 : boolean;
  signal npkt_cnt_1828_1737_buf_req_0 : boolean;
  signal NOT_u1_u1_1779_inst_req_1 : boolean;
  signal call_stmt_1747_call_ack_1 : boolean;
  signal call_stmt_1747_call_req_1 : boolean;
  signal call_stmt_1747_call_ack_0 : boolean;
  signal call_stmt_1747_call_req_0 : boolean;
  signal call_stmt_1776_call_ack_1 : boolean;
  signal call_stmt_1776_call_req_1 : boolean;
  signal if_stmt_1725_branch_ack_0 : boolean;
  signal call_stmt_1759_call_ack_1 : boolean;
  signal call_stmt_1776_call_ack_0 : boolean;
  signal NOT_u1_u1_1779_inst_ack_1 : boolean;
  signal call_stmt_1813_call_ack_0 : boolean;
  signal W_pkt_cnt_1778_delayed_13_0_1801_inst_req_1 : boolean;
  signal if_stmt_1725_branch_ack_1 : boolean;
  signal call_stmt_1813_call_req_0 : boolean;
  signal call_stmt_1813_call_req_1 : boolean;
  signal call_stmt_1813_call_ack_1 : boolean;
  signal call_stmt_1776_call_req_0 : boolean;
  signal if_stmt_1725_branch_req_0 : boolean;
  signal call_stmt_1759_call_req_1 : boolean;
  signal call_stmt_1759_call_ack_0 : boolean;
  signal npkt_cnt_1828_1737_buf_ack_1 : boolean;
  signal npkt_cnt_1828_1737_buf_req_1 : boolean;
  signal W_pkt_cnt_1787_delayed_13_0_1814_inst_req_0 : boolean;
  signal W_pkt_cnt_1787_delayed_13_0_1814_inst_ack_0 : boolean;
  signal W_pkt_cnt_1787_delayed_13_0_1814_inst_req_1 : boolean;
  signal W_pkt_cnt_1787_delayed_13_0_1814_inst_ack_1 : boolean;
  signal ADD_u32_u32_1821_inst_req_0 : boolean;
  signal ADD_u32_u32_1821_inst_ack_0 : boolean;
  signal ADD_u32_u32_1821_inst_req_1 : boolean;
  signal ADD_u32_u32_1821_inst_ack_1 : boolean;
  signal W_rx_buffer_pointer_36_1795_delayed_10_0_1833_inst_req_0 : boolean;
  signal W_rx_buffer_pointer_36_1795_delayed_10_0_1833_inst_ack_0 : boolean;
  signal W_rx_buffer_pointer_36_1795_delayed_10_0_1833_inst_req_1 : boolean;
  signal W_rx_buffer_pointer_36_1795_delayed_10_0_1833_inst_ack_1 : boolean;
  signal call_stmt_1838_call_req_0 : boolean;
  signal call_stmt_1838_call_ack_0 : boolean;
  signal call_stmt_1838_call_req_1 : boolean;
  signal call_stmt_1838_call_ack_1 : boolean;
  signal W_rx_buffer_pointer_36_1803_delayed_10_0_1841_inst_req_0 : boolean;
  signal W_rx_buffer_pointer_36_1803_delayed_10_0_1841_inst_ack_0 : boolean;
  signal W_rx_buffer_pointer_36_1803_delayed_10_0_1841_inst_req_1 : boolean;
  signal W_rx_buffer_pointer_36_1803_delayed_10_0_1841_inst_ack_1 : boolean;
  signal call_stmt_1851_call_req_0 : boolean;
  signal call_stmt_1851_call_ack_0 : boolean;
  signal call_stmt_1851_call_req_1 : boolean;
  signal call_stmt_1851_call_ack_1 : boolean;
  signal do_while_stmt_1733_branch_ack_0 : boolean;
  signal do_while_stmt_1733_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "ReceiveEngineDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  ReceiveEngineDaemon_CP_2495_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "ReceiveEngineDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= ReceiveEngineDaemon_CP_2495_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= ReceiveEngineDaemon_CP_2495_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= ReceiveEngineDaemon_CP_2495_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  ReceiveEngineDaemon_CP_2495: Block -- control-path 
    signal ReceiveEngineDaemon_CP_2495_elements: BooleanArray(91 downto 0);
    -- 
  begin -- 
    ReceiveEngineDaemon_CP_2495_elements(0) <= ReceiveEngineDaemon_CP_2495_start;
    ReceiveEngineDaemon_CP_2495_symbol <= ReceiveEngineDaemon_CP_2495_elements(3);
    -- CP-element group 0:  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 assign_stmt_1721/$entry
      -- CP-element group 0: 	 assign_stmt_1721/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1719_sample_start_
      -- CP-element group 0: 	 assign_stmt_1721/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1719_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_1721/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1719_Sample/req
      -- CP-element group 0: 	 $entry
      -- 
    req_2508_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2508_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2495_elements(0), ack => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1719_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_1721/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1719_update_start_
      -- CP-element group 1: 	 assign_stmt_1721/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1719_sample_completed_
      -- CP-element group 1: 	 assign_stmt_1721/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1719_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_1721/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1719_Sample/ack
      -- CP-element group 1: 	 assign_stmt_1721/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1719_Update/$entry
      -- CP-element group 1: 	 assign_stmt_1721/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1719_Update/req
      -- 
    ack_2509_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1719_inst_ack_0, ack => ReceiveEngineDaemon_CP_2495_elements(1)); -- 
    req_2513_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2513_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2495_elements(1), ack => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1719_inst_req_1); -- 
    -- CP-element group 2:  branch  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	91 
    -- CP-element group 2:  members (10) 
      -- CP-element group 2: 	 assign_stmt_1721/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1719_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_1722/merge_stmt_1724__entry__
      -- CP-element group 2: 	 assign_stmt_1721/$exit
      -- CP-element group 2: 	 assign_stmt_1721/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1719_Update/$exit
      -- CP-element group 2: 	 assign_stmt_1721/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1719_Update/ack
      -- CP-element group 2: 	 branch_block_stmt_1722/branch_block_stmt_1722__entry__
      -- CP-element group 2: 	 branch_block_stmt_1722/$entry
      -- CP-element group 2: 	 branch_block_stmt_1722/merge_stmt_1724_dead_link/$entry
      -- CP-element group 2: 	 branch_block_stmt_1722/merge_stmt_1724__entry___PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_1722/merge_stmt_1724__entry___PhiReq/$exit
      -- 
    ack_2514_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1719_inst_ack_1, ack => ReceiveEngineDaemon_CP_2495_elements(2)); -- 
    -- CP-element group 3:  transition  place  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 $exit
      -- CP-element group 3: 	 branch_block_stmt_1722/branch_block_stmt_1722__exit__
      -- CP-element group 3: 	 branch_block_stmt_1722/$exit
      -- 
    ReceiveEngineDaemon_CP_2495_elements(3) <= false; 
    -- CP-element group 4:  transition  place  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	90 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	91 
    -- CP-element group 4:  members (4) 
      -- CP-element group 4: 	 branch_block_stmt_1722/do_while_stmt_1733__exit__
      -- CP-element group 4: 	 branch_block_stmt_1722/disable_loopback
      -- CP-element group 4: 	 branch_block_stmt_1722/disable_loopback_PhiReq/$entry
      -- CP-element group 4: 	 branch_block_stmt_1722/disable_loopback_PhiReq/$exit
      -- 
    ReceiveEngineDaemon_CP_2495_elements(4) <= ReceiveEngineDaemon_CP_2495_elements(90);
    -- CP-element group 5:  transition  place  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	91 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	91 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_1722/not_enabled_yet_loopback
      -- CP-element group 5: 	 branch_block_stmt_1722/if_stmt_1725_if_link/if_choice_transition
      -- CP-element group 5: 	 branch_block_stmt_1722/if_stmt_1725_if_link/$exit
      -- CP-element group 5: 	 branch_block_stmt_1722/not_enabled_yet_loopback_PhiReq/$entry
      -- CP-element group 5: 	 branch_block_stmt_1722/not_enabled_yet_loopback_PhiReq/$exit
      -- 
    if_choice_transition_2587_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1725_branch_ack_1, ack => ReceiveEngineDaemon_CP_2495_elements(5)); -- 
    -- CP-element group 6:  merge  transition  place  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	91 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (4) 
      -- CP-element group 6: 	 branch_block_stmt_1722/do_while_stmt_1733__entry__
      -- CP-element group 6: 	 branch_block_stmt_1722/if_stmt_1725__exit__
      -- CP-element group 6: 	 branch_block_stmt_1722/if_stmt_1725_else_link/else_choice_transition
      -- CP-element group 6: 	 branch_block_stmt_1722/if_stmt_1725_else_link/$exit
      -- 
    else_choice_transition_2591_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1725_branch_ack_0, ack => ReceiveEngineDaemon_CP_2495_elements(6)); -- 
    -- CP-element group 7:  transition  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	13 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733__entry__
      -- CP-element group 7: 	 branch_block_stmt_1722/do_while_stmt_1733/$entry
      -- 
    ReceiveEngineDaemon_CP_2495_elements(7) <= ReceiveEngineDaemon_CP_2495_elements(6);
    -- CP-element group 8:  merge  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	90 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733__exit__
      -- 
    -- Element group ReceiveEngineDaemon_CP_2495_elements(8) is bound as output of CP function.
    -- CP-element group 9:  merge  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_1722/do_while_stmt_1733/loop_back
      -- 
    -- Element group ReceiveEngineDaemon_CP_2495_elements(9) is bound as output of CP function.
    -- CP-element group 10:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	88 
    -- CP-element group 10: 	89 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_1722/do_while_stmt_1733/condition_done
      -- CP-element group 10: 	 branch_block_stmt_1722/do_while_stmt_1733/loop_exit/$entry
      -- CP-element group 10: 	 branch_block_stmt_1722/do_while_stmt_1733/loop_taken/$entry
      -- 
    ReceiveEngineDaemon_CP_2495_elements(10) <= ReceiveEngineDaemon_CP_2495_elements(15);
    -- CP-element group 11:  branch  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	87 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_1722/do_while_stmt_1733/loop_body_done
      -- 
    ReceiveEngineDaemon_CP_2495_elements(11) <= ReceiveEngineDaemon_CP_2495_elements(87);
    -- CP-element group 12:  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	21 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/back_edge_to_loop_body
      -- 
    ReceiveEngineDaemon_CP_2495_elements(12) <= ReceiveEngineDaemon_CP_2495_elements(9);
    -- CP-element group 13:  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	7 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	23 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/first_time_through_loop_body
      -- 
    ReceiveEngineDaemon_CP_2495_elements(13) <= ReceiveEngineDaemon_CP_2495_elements(7);
    -- CP-element group 14:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	86 
    -- CP-element group 14: 	17 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	34 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/loop_body_start
      -- CP-element group 14: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/$entry
      -- 
    -- Element group ReceiveEngineDaemon_CP_2495_elements(14) is bound as output of CP function.
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	86 
    -- CP-element group 15: 	20 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/condition_evaluated
      -- 
    condition_evaluated_2607_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2607_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2495_elements(15), ack => do_while_stmt_1733_branch_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2495_elements(86) & ReceiveEngineDaemon_CP_2495_elements(20);
      gj_ReceiveEngineDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2495_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	17 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	20 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/aggregated_phi_sample_req
      -- CP-element group 16: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/phi_stmt_1735_sample_start__ps
      -- 
    ReceiveEngineDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2495_elements(17) & ReceiveEngineDaemon_CP_2495_elements(20);
      gj_ReceiveEngineDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2495_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	69 
    -- CP-element group 17: 	49 
    -- CP-element group 17: 	45 
    -- CP-element group 17: 	65 
    -- CP-element group 17: 	19 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	16 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/phi_stmt_1735_sample_start_
      -- 
    ReceiveEngineDaemon_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 31,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2495_elements(14) & ReceiveEngineDaemon_CP_2495_elements(69) & ReceiveEngineDaemon_CP_2495_elements(49) & ReceiveEngineDaemon_CP_2495_elements(45) & ReceiveEngineDaemon_CP_2495_elements(65) & ReceiveEngineDaemon_CP_2495_elements(19);
      gj_ReceiveEngineDaemon_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2495_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	68 
    -- CP-element group 18: 	56 
    -- CP-element group 18: 	64 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/aggregated_phi_update_req
      -- CP-element group 18: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/phi_stmt_1735_update_start_
      -- CP-element group 18: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/phi_stmt_1735_update_start__ps
      -- 
    ReceiveEngineDaemon_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2495_elements(14) & ReceiveEngineDaemon_CP_2495_elements(68) & ReceiveEngineDaemon_CP_2495_elements(56) & ReceiveEngineDaemon_CP_2495_elements(64);
      gj_ReceiveEngineDaemon_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2495_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	67 
    -- CP-element group 19: 	47 
    -- CP-element group 19: 	63 
    -- CP-element group 19: 	43 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	17 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/aggregated_phi_sample_ack
      -- CP-element group 19: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/phi_stmt_1735_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/phi_stmt_1735_sample_completed__ps
      -- 
    -- Element group ReceiveEngineDaemon_CP_2495_elements(19) is bound as output of CP function.
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	66 
    -- CP-element group 20: 	54 
    -- CP-element group 20: 	62 
    -- CP-element group 20: 	15 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	16 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/aggregated_phi_update_ack
      -- CP-element group 20: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/phi_stmt_1735_update_completed__ps
      -- CP-element group 20: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/phi_stmt_1735_update_completed_
      -- 
    -- Element group ReceiveEngineDaemon_CP_2495_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	12 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/phi_stmt_1735_loopback_trigger
      -- 
    ReceiveEngineDaemon_CP_2495_elements(21) <= ReceiveEngineDaemon_CP_2495_elements(12);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/phi_stmt_1735_loopback_sample_req
      -- CP-element group 22: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/phi_stmt_1735_loopback_sample_req_ps
      -- 
    phi_stmt_1735_loopback_sample_req_2622_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1735_loopback_sample_req_2622_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2495_elements(22), ack => phi_stmt_1735_req_0); -- 
    -- Element group ReceiveEngineDaemon_CP_2495_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	13 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/phi_stmt_1735_entry_trigger
      -- 
    ReceiveEngineDaemon_CP_2495_elements(23) <= ReceiveEngineDaemon_CP_2495_elements(13);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/phi_stmt_1735_entry_sample_req_ps
      -- CP-element group 24: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/phi_stmt_1735_entry_sample_req
      -- 
    phi_stmt_1735_entry_sample_req_2625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1735_entry_sample_req_2625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2495_elements(24), ack => phi_stmt_1735_req_1); -- 
    -- Element group ReceiveEngineDaemon_CP_2495_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/phi_stmt_1735_phi_mux_ack
      -- CP-element group 25: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/phi_stmt_1735_phi_mux_ack_ps
      -- 
    phi_stmt_1735_phi_mux_ack_2628_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1735_ack_0, ack => ReceiveEngineDaemon_CP_2495_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/R_npkt_cnt_1737_sample_start__ps
      -- CP-element group 26: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/R_npkt_cnt_1737_Sample/req
      -- CP-element group 26: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/R_npkt_cnt_1737_Sample/$entry
      -- CP-element group 26: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/R_npkt_cnt_1737_sample_start_
      -- 
    req_2641_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2641_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2495_elements(26), ack => npkt_cnt_1828_1737_buf_req_0); -- 
    -- Element group ReceiveEngineDaemon_CP_2495_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/R_npkt_cnt_1737_Update/$entry
      -- CP-element group 27: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/R_npkt_cnt_1737_update_start_
      -- CP-element group 27: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/R_npkt_cnt_1737_update_start__ps
      -- CP-element group 27: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/R_npkt_cnt_1737_Update/req
      -- 
    req_2646_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2646_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2495_elements(27), ack => npkt_cnt_1828_1737_buf_req_1); -- 
    -- Element group ReceiveEngineDaemon_CP_2495_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/R_npkt_cnt_1737_Sample/ack
      -- CP-element group 28: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/R_npkt_cnt_1737_Sample/$exit
      -- CP-element group 28: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/R_npkt_cnt_1737_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/R_npkt_cnt_1737_sample_completed__ps
      -- 
    ack_2642_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => npkt_cnt_1828_1737_buf_ack_0, ack => ReceiveEngineDaemon_CP_2495_elements(28)); -- 
    -- CP-element group 29:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (4) 
      -- CP-element group 29: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/R_npkt_cnt_1737_Update/$exit
      -- CP-element group 29: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/R_npkt_cnt_1737_update_completed_
      -- CP-element group 29: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/R_npkt_cnt_1737_update_completed__ps
      -- CP-element group 29: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/R_npkt_cnt_1737_Update/ack
      -- 
    ack_2647_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 29_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => npkt_cnt_1828_1737_buf_ack_1, ack => ReceiveEngineDaemon_CP_2495_elements(29)); -- 
    -- CP-element group 30:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/type_cast_1739_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/type_cast_1739_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/type_cast_1739_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/type_cast_1739_sample_start__ps
      -- 
    -- Element group ReceiveEngineDaemon_CP_2495_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/type_cast_1739_update_start_
      -- CP-element group 31: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/type_cast_1739_update_start__ps
      -- 
    -- Element group ReceiveEngineDaemon_CP_2495_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	33 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/type_cast_1739_update_completed__ps
      -- 
    ReceiveEngineDaemon_CP_2495_elements(32) <= ReceiveEngineDaemon_CP_2495_elements(33);
    -- CP-element group 33:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	32 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/type_cast_1739_update_completed_
      -- 
    -- Element group ReceiveEngineDaemon_CP_2495_elements(33) is a control-delay.
    cp_element_33_delay: control_delay_element  generic map(name => " 33_delay", delay_value => 1)  port map(req => ReceiveEngineDaemon_CP_2495_elements(31), ack => ReceiveEngineDaemon_CP_2495_elements(33), clk => clk, reset =>reset);
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	14 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	85 
    -- CP-element group 34: 	36 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1747_Sample/crr
      -- CP-element group 34: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1747_Sample/$entry
      -- CP-element group 34: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1747_sample_start_
      -- 
    crr_2664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2495_elements(34), ack => call_stmt_1747_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2495_elements(14) & ReceiveEngineDaemon_CP_2495_elements(85) & ReceiveEngineDaemon_CP_2495_elements(36);
      gj_ReceiveEngineDaemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2495_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	72 
    -- CP-element group 35: 	80 
    -- CP-element group 35: 	85 
    -- CP-element group 35: 	52 
    -- CP-element group 35: 	48 
    -- CP-element group 35: 	40 
    -- CP-element group 35: 	44 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1747_Update/ccr
      -- CP-element group 35: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1747_Update/$entry
      -- CP-element group 35: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1747_update_start_
      -- 
    ccr_2669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2495_elements(35), ack => call_stmt_1747_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2495_elements(72) & ReceiveEngineDaemon_CP_2495_elements(80) & ReceiveEngineDaemon_CP_2495_elements(85) & ReceiveEngineDaemon_CP_2495_elements(52) & ReceiveEngineDaemon_CP_2495_elements(48) & ReceiveEngineDaemon_CP_2495_elements(40) & ReceiveEngineDaemon_CP_2495_elements(44);
      gj_ReceiveEngineDaemon_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2495_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	34 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1747_Sample/cra
      -- CP-element group 36: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1747_Sample/$exit
      -- CP-element group 36: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1747_sample_completed_
      -- 
    cra_2665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1747_call_ack_0, ack => ReceiveEngineDaemon_CP_2495_elements(36)); -- 
    -- CP-element group 37:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	70 
    -- CP-element group 37: 	78 
    -- CP-element group 37: 	50 
    -- CP-element group 37: 	46 
    -- CP-element group 37: 	38 
    -- CP-element group 37: 	42 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1747_Update/cca
      -- CP-element group 37: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1747_Update/$exit
      -- CP-element group 37: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1747_update_completed_
      -- 
    cca_2670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1747_call_ack_1, ack => ReceiveEngineDaemon_CP_2495_elements(37)); -- 
    -- CP-element group 38:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	37 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	77 
    -- CP-element group 38: 	40 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1759_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1759_Sample/crr
      -- CP-element group 38: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1759_sample_start_
      -- 
    crr_2678_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2678_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2495_elements(38), ack => call_stmt_1759_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2495_elements(37) & ReceiveEngineDaemon_CP_2495_elements(77) & ReceiveEngineDaemon_CP_2495_elements(40);
      gj_ReceiveEngineDaemon_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2495_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	77 
    -- CP-element group 39: 	41 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1759_update_start_
      -- CP-element group 39: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1759_Update/ccr
      -- CP-element group 39: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1759_Update/$entry
      -- 
    ccr_2683_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2683_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2495_elements(39), ack => call_stmt_1759_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2495_elements(77) & ReceiveEngineDaemon_CP_2495_elements(41);
      gj_ReceiveEngineDaemon_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2495_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40: marked-successors 
    -- CP-element group 40: 	35 
    -- CP-element group 40: 	38 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1759_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1759_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1759_Sample/cra
      -- 
    cra_2679_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1759_call_ack_0, ack => ReceiveEngineDaemon_CP_2495_elements(40)); -- 
    -- CP-element group 41:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	58 
    -- CP-element group 41: marked-successors 
    -- CP-element group 41: 	39 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1759_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1759_Update/cca
      -- CP-element group 41: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1759_Update/$exit
      -- 
    cca_2684_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1759_call_ack_1, ack => ReceiveEngineDaemon_CP_2495_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	37 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	44 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	44 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1776_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1776_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1776_Sample/crr
      -- 
    crr_2692_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2692_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2495_elements(42), ack => call_stmt_1776_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2495_elements(37) & ReceiveEngineDaemon_CP_2495_elements(44);
      gj_ReceiveEngineDaemon_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2495_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	19 
    -- CP-element group 43: marked-predecessors 
    -- CP-element group 43: 	76 
    -- CP-element group 43: 	84 
    -- CP-element group 43: 	60 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	45 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1776_update_start_
      -- CP-element group 43: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1776_Update/ccr
      -- CP-element group 43: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1776_Update/$entry
      -- 
    ccr_2697_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2697_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2495_elements(43), ack => call_stmt_1776_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2495_elements(19) & ReceiveEngineDaemon_CP_2495_elements(76) & ReceiveEngineDaemon_CP_2495_elements(84) & ReceiveEngineDaemon_CP_2495_elements(60);
      gj_ReceiveEngineDaemon_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2495_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: successors 
    -- CP-element group 44: marked-successors 
    -- CP-element group 44: 	35 
    -- CP-element group 44: 	42 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1776_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1776_Sample/cra
      -- CP-element group 44: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1776_Sample/$exit
      -- 
    cra_2693_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1776_call_ack_0, ack => ReceiveEngineDaemon_CP_2495_elements(44)); -- 
    -- CP-element group 45:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	43 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	74 
    -- CP-element group 45: 	82 
    -- CP-element group 45: 	58 
    -- CP-element group 45: marked-successors 
    -- CP-element group 45: 	17 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1776_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1776_Update/cca
      -- CP-element group 45: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1776_Update/$exit
      -- 
    cca_2698_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1776_call_ack_1, ack => ReceiveEngineDaemon_CP_2495_elements(45)); -- 
    -- CP-element group 46:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	37 
    -- CP-element group 46: marked-predecessors 
    -- CP-element group 46: 	48 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/NOT_u1_u1_1779_Sample/rr
      -- CP-element group 46: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/NOT_u1_u1_1779_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/NOT_u1_u1_1779_sample_start_
      -- 
    rr_2706_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2706_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2495_elements(46), ack => NOT_u1_u1_1779_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2495_elements(37) & ReceiveEngineDaemon_CP_2495_elements(48);
      gj_ReceiveEngineDaemon_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2495_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	19 
    -- CP-element group 47: marked-predecessors 
    -- CP-element group 47: 	76 
    -- CP-element group 47: 	60 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/NOT_u1_u1_1779_update_start_
      -- CP-element group 47: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/NOT_u1_u1_1779_Update/cr
      -- CP-element group 47: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/NOT_u1_u1_1779_Update/$entry
      -- 
    cr_2711_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2711_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2495_elements(47), ack => NOT_u1_u1_1779_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2495_elements(19) & ReceiveEngineDaemon_CP_2495_elements(76) & ReceiveEngineDaemon_CP_2495_elements(60);
      gj_ReceiveEngineDaemon_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2495_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: marked-successors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: 	35 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/NOT_u1_u1_1779_Sample/ra
      -- CP-element group 48: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/NOT_u1_u1_1779_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/NOT_u1_u1_1779_sample_completed_
      -- 
    ra_2707_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1779_inst_ack_0, ack => ReceiveEngineDaemon_CP_2495_elements(48)); -- 
    -- CP-element group 49:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	74 
    -- CP-element group 49: 	58 
    -- CP-element group 49: marked-successors 
    -- CP-element group 49: 	17 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/NOT_u1_u1_1779_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/NOT_u1_u1_1779_Update/ca
      -- CP-element group 49: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/NOT_u1_u1_1779_update_completed_
      -- 
    ca_2712_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1779_inst_ack_1, ack => ReceiveEngineDaemon_CP_2495_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	37 
    -- CP-element group 50: marked-predecessors 
    -- CP-element group 50: 	52 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/NOT_u1_u1_1789_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/NOT_u1_u1_1789_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/NOT_u1_u1_1789_Sample/$entry
      -- 
    rr_2720_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2720_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2495_elements(50), ack => NOT_u1_u1_1789_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2495_elements(37) & ReceiveEngineDaemon_CP_2495_elements(52);
      gj_ReceiveEngineDaemon_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2495_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	84 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/NOT_u1_u1_1789_Update/cr
      -- CP-element group 51: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/NOT_u1_u1_1789_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/NOT_u1_u1_1789_update_start_
      -- 
    cr_2725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2495_elements(51), ack => NOT_u1_u1_1789_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_2495_elements(84);
      gj_ReceiveEngineDaemon_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2495_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: marked-successors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: 	35 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/NOT_u1_u1_1789_Sample/ra
      -- CP-element group 52: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/NOT_u1_u1_1789_sample_completed_
      -- CP-element group 52: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/NOT_u1_u1_1789_Sample/$exit
      -- 
    ra_2721_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1789_inst_ack_0, ack => ReceiveEngineDaemon_CP_2495_elements(52)); -- 
    -- CP-element group 53:  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	82 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/NOT_u1_u1_1789_Update/ca
      -- CP-element group 53: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/NOT_u1_u1_1789_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/NOT_u1_u1_1789_Update/$exit
      -- 
    ca_2726_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1789_inst_ack_1, ack => ReceiveEngineDaemon_CP_2495_elements(53)); -- 
    -- CP-element group 54:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	20 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	56 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1803_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1803_Sample/req
      -- CP-element group 54: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1803_sample_start_
      -- 
    req_2734_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2734_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2495_elements(54), ack => W_pkt_cnt_1778_delayed_13_0_1801_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2495_elements(20) & ReceiveEngineDaemon_CP_2495_elements(56);
      gj_ReceiveEngineDaemon_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2495_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: marked-predecessors 
    -- CP-element group 55: 	60 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1803_update_start_
      -- CP-element group 55: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1803_Update/req
      -- CP-element group 55: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1803_Update/$entry
      -- 
    req_2739_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2739_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2495_elements(55), ack => W_pkt_cnt_1778_delayed_13_0_1801_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_2495_elements(60);
      gj_ReceiveEngineDaemon_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2495_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: marked-successors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: 	18 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1803_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1803_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1803_Sample/ack
      -- 
    ack_2735_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_pkt_cnt_1778_delayed_13_0_1801_inst_ack_0, ack => ReceiveEngineDaemon_CP_2495_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1803_Update/ack
      -- CP-element group 57: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1803_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1803_Update/$exit
      -- 
    ack_2740_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_pkt_cnt_1778_delayed_13_0_1801_inst_ack_1, ack => ReceiveEngineDaemon_CP_2495_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: 	49 
    -- CP-element group 58: 	45 
    -- CP-element group 58: 	41 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	60 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1813_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1813_Sample/crr
      -- CP-element group 58: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1813_sample_start_
      -- 
    crr_2748_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2748_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2495_elements(58), ack => call_stmt_1813_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 31,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2495_elements(57) & ReceiveEngineDaemon_CP_2495_elements(49) & ReceiveEngineDaemon_CP_2495_elements(45) & ReceiveEngineDaemon_CP_2495_elements(41) & ReceiveEngineDaemon_CP_2495_elements(60);
      gj_ReceiveEngineDaemon_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2495_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1813_Update/ccr
      -- CP-element group 59: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1813_update_start_
      -- CP-element group 59: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1813_Update/$entry
      -- 
    ccr_2753_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2753_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2495_elements(59), ack => call_stmt_1813_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_2495_elements(61);
      gj_ReceiveEngineDaemon_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2495_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	55 
    -- CP-element group 60: 	58 
    -- CP-element group 60: 	47 
    -- CP-element group 60: 	43 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1813_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1813_Sample/cra
      -- CP-element group 60: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1813_Sample/$exit
      -- 
    cra_2749_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1813_call_ack_0, ack => ReceiveEngineDaemon_CP_2495_elements(60)); -- 
    -- CP-element group 61:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	74 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	59 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1813_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1813_Update/cca
      -- CP-element group 61: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1813_Update/$exit
      -- 
    cca_2754_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1813_call_ack_1, ack => ReceiveEngineDaemon_CP_2495_elements(61)); -- 
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	20 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	64 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1816_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1816_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1816_Sample/req
      -- 
    req_2762_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2762_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2495_elements(62), ack => W_pkt_cnt_1787_delayed_13_0_1814_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2495_elements(20) & ReceiveEngineDaemon_CP_2495_elements(64);
      gj_ReceiveEngineDaemon_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2495_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	19 
    -- CP-element group 63: marked-predecessors 
    -- CP-element group 63: 	65 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1816_update_start_
      -- CP-element group 63: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1816_Update/$entry
      -- CP-element group 63: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1816_Update/req
      -- 
    req_2767_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2767_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2495_elements(63), ack => W_pkt_cnt_1787_delayed_13_0_1814_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2495_elements(19) & ReceiveEngineDaemon_CP_2495_elements(65);
      gj_ReceiveEngineDaemon_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2495_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: 	18 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1816_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1816_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1816_Sample/ack
      -- 
    ack_2763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_pkt_cnt_1787_delayed_13_0_1814_inst_ack_0, ack => ReceiveEngineDaemon_CP_2495_elements(64)); -- 
    -- CP-element group 65:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	87 
    -- CP-element group 65: marked-successors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: 	17 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1816_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1816_Update/$exit
      -- CP-element group 65: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1816_Update/ack
      -- 
    ack_2768_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_pkt_cnt_1787_delayed_13_0_1814_inst_ack_1, ack => ReceiveEngineDaemon_CP_2495_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	20 
    -- CP-element group 66: marked-predecessors 
    -- CP-element group 66: 	68 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/ADD_u32_u32_1821_sample_start_
      -- CP-element group 66: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/ADD_u32_u32_1821_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/ADD_u32_u32_1821_Sample/rr
      -- 
    rr_2776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2495_elements(66), ack => ADD_u32_u32_1821_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2495_elements(20) & ReceiveEngineDaemon_CP_2495_elements(68);
      gj_ReceiveEngineDaemon_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2495_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	19 
    -- CP-element group 67: marked-predecessors 
    -- CP-element group 67: 	69 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/ADD_u32_u32_1821_update_start_
      -- CP-element group 67: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/ADD_u32_u32_1821_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/ADD_u32_u32_1821_Update/cr
      -- 
    cr_2781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2495_elements(67), ack => ADD_u32_u32_1821_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2495_elements(19) & ReceiveEngineDaemon_CP_2495_elements(69);
      gj_ReceiveEngineDaemon_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2495_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: marked-successors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: 	18 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/ADD_u32_u32_1821_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/ADD_u32_u32_1821_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/ADD_u32_u32_1821_Sample/ra
      -- 
    ra_2777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_1821_inst_ack_0, ack => ReceiveEngineDaemon_CP_2495_elements(68)); -- 
    -- CP-element group 69:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	87 
    -- CP-element group 69: marked-successors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: 	17 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/ADD_u32_u32_1821_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/ADD_u32_u32_1821_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/ADD_u32_u32_1821_Update/ca
      -- 
    ca_2782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_1821_inst_ack_1, ack => ReceiveEngineDaemon_CP_2495_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	37 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	72 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1835_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1835_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1835_Sample/req
      -- 
    req_2790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2495_elements(70), ack => W_rx_buffer_pointer_36_1795_delayed_10_0_1833_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2495_elements(37) & ReceiveEngineDaemon_CP_2495_elements(72);
      gj_ReceiveEngineDaemon_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2495_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	76 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1835_update_start_
      -- CP-element group 71: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1835_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1835_Update/req
      -- 
    req_2795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2495_elements(71), ack => W_rx_buffer_pointer_36_1795_delayed_10_0_1833_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_2495_elements(76);
      gj_ReceiveEngineDaemon_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2495_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: marked-successors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: 	35 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1835_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1835_Sample/$exit
      -- CP-element group 72: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1835_Sample/ack
      -- 
    ack_2791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_36_1795_delayed_10_0_1833_inst_ack_0, ack => ReceiveEngineDaemon_CP_2495_elements(72)); -- 
    -- CP-element group 73:  transition  input  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	74 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1835_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1835_Update/$exit
      -- CP-element group 73: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1835_Update/ack
      -- 
    ack_2796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_36_1795_delayed_10_0_1833_inst_ack_1, ack => ReceiveEngineDaemon_CP_2495_elements(73)); -- 
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	73 
    -- CP-element group 74: 	61 
    -- CP-element group 74: 	49 
    -- CP-element group 74: 	45 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	76 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1838_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1838_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1838_Sample/crr
      -- 
    crr_2804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2495_elements(74), ack => call_stmt_1838_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 31,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2495_elements(73) & ReceiveEngineDaemon_CP_2495_elements(61) & ReceiveEngineDaemon_CP_2495_elements(49) & ReceiveEngineDaemon_CP_2495_elements(45) & ReceiveEngineDaemon_CP_2495_elements(76);
      gj_ReceiveEngineDaemon_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2495_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: marked-predecessors 
    -- CP-element group 75: 	77 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1838_update_start_
      -- CP-element group 75: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1838_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1838_Update/ccr
      -- 
    ccr_2809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2495_elements(75), ack => call_stmt_1838_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_2495_elements(77);
      gj_ReceiveEngineDaemon_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2495_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: marked-successors 
    -- CP-element group 76: 	71 
    -- CP-element group 76: 	74 
    -- CP-element group 76: 	47 
    -- CP-element group 76: 	43 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1838_sample_completed_
      -- CP-element group 76: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1838_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1838_Sample/cra
      -- 
    cra_2805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1838_call_ack_0, ack => ReceiveEngineDaemon_CP_2495_elements(76)); -- 
    -- CP-element group 77:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	82 
    -- CP-element group 77: marked-successors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: 	38 
    -- CP-element group 77: 	39 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1838_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1838_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1838_Update/cca
      -- 
    cca_2810_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1838_call_ack_1, ack => ReceiveEngineDaemon_CP_2495_elements(77)); -- 
    -- CP-element group 78:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	37 
    -- CP-element group 78: marked-predecessors 
    -- CP-element group 78: 	80 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	80 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1843_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1843_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1843_Sample/req
      -- 
    req_2818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2495_elements(78), ack => W_rx_buffer_pointer_36_1803_delayed_10_0_1841_inst_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2495_elements(37) & ReceiveEngineDaemon_CP_2495_elements(80);
      gj_ReceiveEngineDaemon_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2495_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: marked-predecessors 
    -- CP-element group 79: 	84 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	81 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1843_update_start_
      -- CP-element group 79: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1843_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1843_Update/req
      -- 
    req_2823_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2823_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2495_elements(79), ack => W_rx_buffer_pointer_36_1803_delayed_10_0_1841_inst_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_79: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_79"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_2495_elements(84);
      gj_ReceiveEngineDaemon_cp_element_group_79 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2495_elements(79), clk => clk, reset => reset); --
    end block;
    -- CP-element group 80:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: successors 
    -- CP-element group 80: marked-successors 
    -- CP-element group 80: 	78 
    -- CP-element group 80: 	35 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1843_sample_completed_
      -- CP-element group 80: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1843_Sample/$exit
      -- CP-element group 80: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1843_Sample/ack
      -- 
    ack_2819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_36_1803_delayed_10_0_1841_inst_ack_0, ack => ReceiveEngineDaemon_CP_2495_elements(80)); -- 
    -- CP-element group 81:  transition  input  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	79 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1843_update_completed_
      -- CP-element group 81: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1843_Update/$exit
      -- CP-element group 81: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/assign_stmt_1843_Update/ack
      -- 
    ack_2824_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_36_1803_delayed_10_0_1841_inst_ack_1, ack => ReceiveEngineDaemon_CP_2495_elements(81)); -- 
    -- CP-element group 82:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	77 
    -- CP-element group 82: 	81 
    -- CP-element group 82: 	53 
    -- CP-element group 82: 	45 
    -- CP-element group 82: marked-predecessors 
    -- CP-element group 82: 	84 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	84 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1851_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1851_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1851_Sample/crr
      -- 
    crr_2832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2495_elements(82), ack => call_stmt_1851_call_req_0); -- 
    ReceiveEngineDaemon_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 31,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2495_elements(77) & ReceiveEngineDaemon_CP_2495_elements(81) & ReceiveEngineDaemon_CP_2495_elements(53) & ReceiveEngineDaemon_CP_2495_elements(45) & ReceiveEngineDaemon_CP_2495_elements(84);
      gj_ReceiveEngineDaemon_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2495_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: marked-predecessors 
    -- CP-element group 83: 	85 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1851_update_start_
      -- CP-element group 83: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1851_Update/$entry
      -- CP-element group 83: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1851_Update/ccr
      -- 
    ccr_2837_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2837_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2495_elements(83), ack => call_stmt_1851_call_req_1); -- 
    ReceiveEngineDaemon_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= ReceiveEngineDaemon_CP_2495_elements(85);
      gj_ReceiveEngineDaemon_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2495_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	82 
    -- CP-element group 84: successors 
    -- CP-element group 84: marked-successors 
    -- CP-element group 84: 	79 
    -- CP-element group 84: 	82 
    -- CP-element group 84: 	51 
    -- CP-element group 84: 	43 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1851_sample_completed_
      -- CP-element group 84: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1851_Sample/$exit
      -- CP-element group 84: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1851_Sample/cra
      -- 
    cra_2833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1851_call_ack_0, ack => ReceiveEngineDaemon_CP_2495_elements(84)); -- 
    -- CP-element group 85:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85: marked-successors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: 	34 
    -- CP-element group 85: 	35 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1851_update_completed_
      -- CP-element group 85: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1851_Update/$exit
      -- CP-element group 85: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/call_stmt_1851_Update/cca
      -- 
    cca_2838_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1851_call_ack_1, ack => ReceiveEngineDaemon_CP_2495_elements(85)); -- 
    -- CP-element group 86:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	14 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	15 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group ReceiveEngineDaemon_CP_2495_elements(86) is a control-delay.
    cp_element_86_delay: control_delay_element  generic map(name => " 86_delay", delay_value => 1)  port map(req => ReceiveEngineDaemon_CP_2495_elements(14), ack => ReceiveEngineDaemon_CP_2495_elements(86), clk => clk, reset =>reset);
    -- CP-element group 87:  join  transition  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	69 
    -- CP-element group 87: 	85 
    -- CP-element group 87: 	65 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	11 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_1722/do_while_stmt_1733/do_while_stmt_1733_loop_body/$exit
      -- 
    ReceiveEngineDaemon_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 31,2 => 31);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 39) := "ReceiveEngineDaemon_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= ReceiveEngineDaemon_CP_2495_elements(69) & ReceiveEngineDaemon_CP_2495_elements(85) & ReceiveEngineDaemon_CP_2495_elements(65);
      gj_ReceiveEngineDaemon_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => ReceiveEngineDaemon_CP_2495_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  transition  input  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	10 
    -- CP-element group 88: successors 
    -- CP-element group 88:  members (2) 
      -- CP-element group 88: 	 branch_block_stmt_1722/do_while_stmt_1733/loop_exit/$exit
      -- CP-element group 88: 	 branch_block_stmt_1722/do_while_stmt_1733/loop_exit/ack
      -- 
    ack_2843_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 88_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1733_branch_ack_0, ack => ReceiveEngineDaemon_CP_2495_elements(88)); -- 
    -- CP-element group 89:  transition  input  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	10 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (2) 
      -- CP-element group 89: 	 branch_block_stmt_1722/do_while_stmt_1733/loop_taken/$exit
      -- CP-element group 89: 	 branch_block_stmt_1722/do_while_stmt_1733/loop_taken/ack
      -- 
    ack_2847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1733_branch_ack_1, ack => ReceiveEngineDaemon_CP_2495_elements(89)); -- 
    -- CP-element group 90:  transition  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	8 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	4 
    -- CP-element group 90:  members (1) 
      -- CP-element group 90: 	 branch_block_stmt_1722/do_while_stmt_1733/$exit
      -- 
    ReceiveEngineDaemon_CP_2495_elements(90) <= ReceiveEngineDaemon_CP_2495_elements(8);
    -- CP-element group 91:  merge  branch  transition  place  output  bypass 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	2 
    -- CP-element group 91: 	4 
    -- CP-element group 91: 	5 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	5 
    -- CP-element group 91: 	6 
    -- CP-element group 91:  members (49) 
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725__entry__
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/SplitProtocol/$exit
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/BITSEL_u32_u1_1728/$entry
      -- CP-element group 91: 	 branch_block_stmt_1722/NOT_u1_u1_1729_place
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/SplitProtocol/Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/SplitProtocol/Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_1722/merge_stmt_1724__exit__
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/SplitProtocol/Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/BITSEL_u32_u1_1728/$exit
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/BITSEL_u32_u1_1728/BITSEL_u32_u1_1728_inputs/$entry
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/SplitProtocol/Sample/ra
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/SplitProtocol/Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/SplitProtocol/$entry
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/BITSEL_u32_u1_1728/SplitProtocol/Update/ca
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/BITSEL_u32_u1_1728/SplitProtocol/Update/cr
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/$exit
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/BITSEL_u32_u1_1728/SplitProtocol/Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/BITSEL_u32_u1_1728/SplitProtocol/Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/BITSEL_u32_u1_1728/SplitProtocol/Sample/ra
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/BITSEL_u32_u1_1728/SplitProtocol/Sample/rr
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/BITSEL_u32_u1_1728/SplitProtocol/Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/BITSEL_u32_u1_1728/SplitProtocol/Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/BITSEL_u32_u1_1728/SplitProtocol/$exit
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_else_link/$entry
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/BITSEL_u32_u1_1728/SplitProtocol/$entry
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/BITSEL_u32_u1_1728/BITSEL_u32_u1_1728_inputs/RPIPE_CONTROL_REGISTER_1726/Update/ack
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/$entry
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_if_link/$entry
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/BITSEL_u32_u1_1728/BITSEL_u32_u1_1728_inputs/RPIPE_CONTROL_REGISTER_1726/Update/req
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/BITSEL_u32_u1_1728/BITSEL_u32_u1_1728_inputs/RPIPE_CONTROL_REGISTER_1726/Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/branch_req
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/BITSEL_u32_u1_1728/BITSEL_u32_u1_1728_inputs/RPIPE_CONTROL_REGISTER_1726/Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/BITSEL_u32_u1_1728/BITSEL_u32_u1_1728_inputs/RPIPE_CONTROL_REGISTER_1726/Sample/ack
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/SplitProtocol/Update/ca
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/SplitProtocol/Update/cr
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/$exit
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/BITSEL_u32_u1_1728/BITSEL_u32_u1_1728_inputs/RPIPE_CONTROL_REGISTER_1726/Sample/req
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/BITSEL_u32_u1_1728/BITSEL_u32_u1_1728_inputs/RPIPE_CONTROL_REGISTER_1726/Sample/$exit
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/$entry
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/BITSEL_u32_u1_1728/BITSEL_u32_u1_1728_inputs/RPIPE_CONTROL_REGISTER_1726/Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/BITSEL_u32_u1_1728/BITSEL_u32_u1_1728_inputs/RPIPE_CONTROL_REGISTER_1726/$exit
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_dead_link/$entry
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/SplitProtocol/Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/BITSEL_u32_u1_1728/BITSEL_u32_u1_1728_inputs/RPIPE_CONTROL_REGISTER_1726/$entry
      -- CP-element group 91: 	 branch_block_stmt_1722/if_stmt_1725_eval_test/NOT_u1_u1_1729/BITSEL_u32_u1_1728/BITSEL_u32_u1_1728_inputs/$exit
      -- CP-element group 91: 	 branch_block_stmt_1722/merge_stmt_1724_PhiReqMerge
      -- CP-element group 91: 	 branch_block_stmt_1722/merge_stmt_1724_PhiAck/$entry
      -- CP-element group 91: 	 branch_block_stmt_1722/merge_stmt_1724_PhiAck/$exit
      -- CP-element group 91: 	 branch_block_stmt_1722/merge_stmt_1724_PhiAck/dummy
      -- 
    branch_req_2582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ReceiveEngineDaemon_CP_2495_elements(91), ack => if_stmt_1725_branch_req_0); -- 
    ReceiveEngineDaemon_CP_2495_elements(91) <= OrReduce(ReceiveEngineDaemon_CP_2495_elements(2) & ReceiveEngineDaemon_CP_2495_elements(4) & ReceiveEngineDaemon_CP_2495_elements(5));
    ReceiveEngineDaemon_do_while_stmt_1733_terminator_2848: loop_terminator -- 
      generic map (name => " ReceiveEngineDaemon_do_while_stmt_1733_terminator_2848", max_iterations_in_flight =>31) 
      port map(loop_body_exit => ReceiveEngineDaemon_CP_2495_elements(11),loop_continue => ReceiveEngineDaemon_CP_2495_elements(89),loop_terminate => ReceiveEngineDaemon_CP_2495_elements(88),loop_back => ReceiveEngineDaemon_CP_2495_elements(9),loop_exit => ReceiveEngineDaemon_CP_2495_elements(8),clk => clk, reset => reset); -- 
    phi_stmt_1735_phi_seq_2656_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= ReceiveEngineDaemon_CP_2495_elements(21);
      ReceiveEngineDaemon_CP_2495_elements(26)<= src_sample_reqs(0);
      src_sample_acks(0)  <= ReceiveEngineDaemon_CP_2495_elements(28);
      ReceiveEngineDaemon_CP_2495_elements(27)<= src_update_reqs(0);
      src_update_acks(0)  <= ReceiveEngineDaemon_CP_2495_elements(29);
      ReceiveEngineDaemon_CP_2495_elements(22) <= phi_mux_reqs(0);
      triggers(1)  <= ReceiveEngineDaemon_CP_2495_elements(23);
      ReceiveEngineDaemon_CP_2495_elements(30)<= src_sample_reqs(1);
      src_sample_acks(1)  <= ReceiveEngineDaemon_CP_2495_elements(30);
      ReceiveEngineDaemon_CP_2495_elements(31)<= src_update_reqs(1);
      src_update_acks(1)  <= ReceiveEngineDaemon_CP_2495_elements(32);
      ReceiveEngineDaemon_CP_2495_elements(24) <= phi_mux_reqs(1);
      phi_stmt_1735_phi_seq_2656 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_1735_phi_seq_2656") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => ReceiveEngineDaemon_CP_2495_elements(16), 
          phi_sample_ack => ReceiveEngineDaemon_CP_2495_elements(19), 
          phi_update_req => ReceiveEngineDaemon_CP_2495_elements(18), 
          phi_update_ack => ReceiveEngineDaemon_CP_2495_elements(20), 
          phi_mux_ack => ReceiveEngineDaemon_CP_2495_elements(25), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_2608_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= ReceiveEngineDaemon_CP_2495_elements(12);
        preds(1)  <= ReceiveEngineDaemon_CP_2495_elements(13);
        entry_tmerge_2608 : transition_merge -- 
          generic map(name => " entry_tmerge_2608")
          port map (preds => preds, symbol_out => ReceiveEngineDaemon_CP_2495_elements(14));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_1786_1786_delayed_13_0_1822 : std_logic_vector(31 downto 0);
    signal BITSEL_u32_u1_1728_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_1856_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1729_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1755_1755_delayed_10_0_1780 : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1762_1762_delayed_10_0_1790 : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1784_wire : std_logic_vector(0 downto 0);
    signal NOT_u4_u4_1755_wire_constant : std_logic_vector(3 downto 0);
    signal NOT_u4_u4_1809_wire_constant : std_logic_vector(3 downto 0);
    signal RPIPE_CONTROL_REGISTER_1726_wire : std_logic_vector(31 downto 0);
    signal RPIPE_CONTROL_REGISTER_1854_wire : std_logic_vector(31 downto 0);
    signal RPIPE_FREE_Q_1744_wire : std_logic_vector(35 downto 0);
    signal RPIPE_FREE_Q_1847_wire : std_logic_vector(35 downto 0);
    signal bad_packet_identifier_1776 : std_logic_vector(0 downto 0);
    signal cond_1800 : std_logic_vector(0 downto 0);
    signal free_flag_1795 : std_logic_vector(0 downto 0);
    signal ignore_resp0_1759 : std_logic_vector(31 downto 0);
    signal ignore_resp1_1813 : std_logic_vector(31 downto 0);
    signal konst_1720_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1727_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1756_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1798_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1810_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1855_wire_constant : std_logic_vector(31 downto 0);
    signal npkt_cnt_1828 : std_logic_vector(31 downto 0);
    signal npkt_cnt_1828_1737_buffered : std_logic_vector(31 downto 0);
    signal ok_flag_1786 : std_logic_vector(0 downto 0);
    signal pkt_cnt_1735 : std_logic_vector(31 downto 0);
    signal pkt_cnt_1778_delayed_13_0_1803 : std_logic_vector(31 downto 0);
    signal pkt_cnt_1787_delayed_13_0_1816 : std_logic_vector(31 downto 0);
    signal push_status_1851 : std_logic_vector(0 downto 0);
    signal rx_buffer_pointer_32_1747 : std_logic_vector(31 downto 0);
    signal rx_buffer_pointer_36_1765 : std_logic_vector(35 downto 0);
    signal rx_buffer_pointer_36_1795_delayed_10_0_1835 : std_logic_vector(35 downto 0);
    signal rx_buffer_pointer_36_1803_delayed_10_0_1843 : std_logic_vector(35 downto 0);
    signal slice_1849_wire : std_logic_vector(31 downto 0);
    signal status_1747 : std_logic_vector(0 downto 0);
    signal type_cast_1739_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1743_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1752_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1762_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_1806_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1820_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1846_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    NOT_u4_u4_1755_wire_constant <= "1111";
    NOT_u4_u4_1809_wire_constant <= "1111";
    konst_1720_wire_constant <= "000000";
    konst_1727_wire_constant <= "00000000000000000000000000000000";
    konst_1756_wire_constant <= "011000";
    konst_1798_wire_constant <= "1";
    konst_1810_wire_constant <= "011001";
    konst_1855_wire_constant <= "00000000000000000000000000000000";
    type_cast_1739_wire_constant <= "00000000000000000000000000000000";
    type_cast_1743_wire_constant <= "1";
    type_cast_1752_wire_constant <= "0";
    type_cast_1762_wire_constant <= "0000";
    type_cast_1806_wire_constant <= "0";
    type_cast_1820_wire_constant <= "00000000000000000000000000000001";
    type_cast_1846_wire_constant <= "1";
    phi_stmt_1735: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= npkt_cnt_1828_1737_buffered & type_cast_1739_wire_constant;
      req <= phi_stmt_1735_req_0 & phi_stmt_1735_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1735",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1735_ack_0,
          idata => idata,
          odata => pkt_cnt_1735,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1735
    -- flow-through select operator MUX_1827_inst
    npkt_cnt_1828 <= ADD_u32_u32_1786_1786_delayed_13_0_1822 when (ok_flag_1786(0) /=  '0') else pkt_cnt_1787_delayed_13_0_1816;
    -- flow-through slice operator slice_1849_inst
    slice_1849_wire <= rx_buffer_pointer_36_1803_delayed_10_0_1843(31 downto 0);
    W_pkt_cnt_1778_delayed_13_0_1801_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_pkt_cnt_1778_delayed_13_0_1801_inst_req_0;
      W_pkt_cnt_1778_delayed_13_0_1801_inst_ack_0<= wack(0);
      rreq(0) <= W_pkt_cnt_1778_delayed_13_0_1801_inst_req_1;
      W_pkt_cnt_1778_delayed_13_0_1801_inst_ack_1<= rack(0);
      W_pkt_cnt_1778_delayed_13_0_1801_inst : InterlockBuffer generic map ( -- 
        name => "W_pkt_cnt_1778_delayed_13_0_1801_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => pkt_cnt_1735,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pkt_cnt_1778_delayed_13_0_1803,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_pkt_cnt_1787_delayed_13_0_1814_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_pkt_cnt_1787_delayed_13_0_1814_inst_req_0;
      W_pkt_cnt_1787_delayed_13_0_1814_inst_ack_0<= wack(0);
      rreq(0) <= W_pkt_cnt_1787_delayed_13_0_1814_inst_req_1;
      W_pkt_cnt_1787_delayed_13_0_1814_inst_ack_1<= rack(0);
      W_pkt_cnt_1787_delayed_13_0_1814_inst : InterlockBuffer generic map ( -- 
        name => "W_pkt_cnt_1787_delayed_13_0_1814_inst",
        buffer_size => 13,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => pkt_cnt_1735,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pkt_cnt_1787_delayed_13_0_1816,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rx_buffer_pointer_36_1795_delayed_10_0_1833_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rx_buffer_pointer_36_1795_delayed_10_0_1833_inst_req_0;
      W_rx_buffer_pointer_36_1795_delayed_10_0_1833_inst_ack_0<= wack(0);
      rreq(0) <= W_rx_buffer_pointer_36_1795_delayed_10_0_1833_inst_req_1;
      W_rx_buffer_pointer_36_1795_delayed_10_0_1833_inst_ack_1<= rack(0);
      W_rx_buffer_pointer_36_1795_delayed_10_0_1833_inst : InterlockBuffer generic map ( -- 
        name => "W_rx_buffer_pointer_36_1795_delayed_10_0_1833_inst",
        buffer_size => 10,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rx_buffer_pointer_36_1765,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rx_buffer_pointer_36_1795_delayed_10_0_1835,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rx_buffer_pointer_36_1803_delayed_10_0_1841_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rx_buffer_pointer_36_1803_delayed_10_0_1841_inst_req_0;
      W_rx_buffer_pointer_36_1803_delayed_10_0_1841_inst_ack_0<= wack(0);
      rreq(0) <= W_rx_buffer_pointer_36_1803_delayed_10_0_1841_inst_req_1;
      W_rx_buffer_pointer_36_1803_delayed_10_0_1841_inst_ack_1<= rack(0);
      W_rx_buffer_pointer_36_1803_delayed_10_0_1841_inst : InterlockBuffer generic map ( -- 
        name => "W_rx_buffer_pointer_36_1803_delayed_10_0_1841_inst",
        buffer_size => 10,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rx_buffer_pointer_36_1765,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rx_buffer_pointer_36_1803_delayed_10_0_1843,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    npkt_cnt_1828_1737_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= npkt_cnt_1828_1737_buf_req_0;
      npkt_cnt_1828_1737_buf_ack_0<= wack(0);
      rreq(0) <= npkt_cnt_1828_1737_buf_req_1;
      npkt_cnt_1828_1737_buf_ack_1<= rack(0);
      npkt_cnt_1828_1737_buf : InterlockBuffer generic map ( -- 
        name => "npkt_cnt_1828_1737_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => npkt_cnt_1828,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => npkt_cnt_1828_1737_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_1733_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= BITSEL_u32_u1_1856_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1733_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1733_branch_req_0,
          ack0 => do_while_stmt_1733_branch_ack_0,
          ack1 => do_while_stmt_1733_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1725_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_1729_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1725_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1725_branch_req_0,
          ack0 => if_stmt_1725_branch_ack_0,
          ack1 => if_stmt_1725_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u32_u32_1821_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 13);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= pkt_cnt_1735;
      ADD_u32_u32_1786_1786_delayed_13_0_1822 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_1821_inst_req_0;
      ADD_u32_u32_1821_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_1821_inst_req_1;
      ADD_u32_u32_1821_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 13,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- binary operator AND_u1_u1_1785_inst
    process(NOT_u1_u1_1755_1755_delayed_10_0_1780, NOT_u1_u1_1784_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_1755_1755_delayed_10_0_1780, NOT_u1_u1_1784_wire, tmp_var);
      ok_flag_1786 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1794_inst
    process(NOT_u1_u1_1762_1762_delayed_10_0_1790, bad_packet_identifier_1776) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_1762_1762_delayed_10_0_1790, bad_packet_identifier_1776, tmp_var);
      free_flag_1795 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_1728_inst
    process(RPIPE_CONTROL_REGISTER_1726_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_CONTROL_REGISTER_1726_wire, konst_1727_wire_constant, tmp_var);
      BITSEL_u32_u1_1728_wire <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_1856_inst
    process(RPIPE_CONTROL_REGISTER_1854_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_CONTROL_REGISTER_1854_wire, konst_1855_wire_constant, tmp_var);
      BITSEL_u32_u1_1856_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u4_u36_1764_inst
    process(type_cast_1762_wire_constant, rx_buffer_pointer_32_1747) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1762_wire_constant, rx_buffer_pointer_32_1747, tmp_var);
      rx_buffer_pointer_36_1765 <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_1799_inst
    process(ok_flag_1786) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(ok_flag_1786, konst_1798_wire_constant, tmp_var);
      cond_1800 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1729_inst
    process(BITSEL_u32_u1_1728_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", BITSEL_u32_u1_1728_wire, tmp_var);
      NOT_u1_u1_1729_wire <= tmp_var; -- 
    end process;
    -- shared split operator group (8) : NOT_u1_u1_1779_inst 
    ApIntNot_group_8: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 10);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= status_1747;
      NOT_u1_u1_1755_1755_delayed_10_0_1780 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NOT_u1_u1_1779_inst_req_0;
      NOT_u1_u1_1779_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NOT_u1_u1_1779_inst_req_1;
      NOT_u1_u1_1779_inst_ack_1 <= ackR_unguarded(0);
      ApIntNot_group_8_gI: SplitGuardInterface generic map(name => "ApIntNot_group_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNot",
          name => "ApIntNot_group_8",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 10,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 8
    -- unary operator NOT_u1_u1_1784_inst
    process(bad_packet_identifier_1776) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", bad_packet_identifier_1776, tmp_var);
      NOT_u1_u1_1784_wire <= tmp_var; -- 
    end process;
    -- shared split operator group (10) : NOT_u1_u1_1789_inst 
    ApIntNot_group_10: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 10);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= status_1747;
      NOT_u1_u1_1762_1762_delayed_10_0_1790 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NOT_u1_u1_1789_inst_req_0;
      NOT_u1_u1_1789_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NOT_u1_u1_1789_inst_req_1;
      NOT_u1_u1_1789_inst_ack_1 <= ackR_unguarded(0);
      ApIntNot_group_10_gI: SplitGuardInterface generic map(name => "ApIntNot_group_10_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNot",
          name => "ApIntNot_group_10",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 10,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 10
    -- read from input-signal CONTROL_REGISTER
    RPIPE_CONTROL_REGISTER_1726_wire <= CONTROL_REGISTER;
    -- read from input-signal CONTROL_REGISTER
    RPIPE_CONTROL_REGISTER_1854_wire <= CONTROL_REGISTER;
    -- read from input-signal FREE_Q
    RPIPE_FREE_Q_1744_wire <= FREE_Q;
    RPIPE_FREE_Q_1847_wire <= FREE_Q;
    -- shared outport operator group (0) : WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1719_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1719_inst_req_0;
      WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1719_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1719_inst_req_1;
      WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1719_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= konst_1720_wire_constant;
      LAST_WRITTEN_RX_QUEUE_INDEX_write_0_gI: SplitGuardInterface generic map(name => "LAST_WRITTEN_RX_QUEUE_INDEX_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      LAST_WRITTEN_RX_QUEUE_INDEX_write_0: OutputPortRevised -- 
        generic map ( name => "LAST_WRITTEN_RX_QUEUE_INDEX", data_width => 6, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req(0),
          oack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack(0),
          odata => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data(5 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_1747_call 
    popFromQueue_call_group_0: Block -- 
      signal data_in: std_logic_vector(36 downto 0);
      signal data_out: std_logic_vector(32 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1747_call_req_0;
      call_stmt_1747_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1747_call_req_1;
      call_stmt_1747_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      popFromQueue_call_group_0_gI: SplitGuardInterface generic map(name => "popFromQueue_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1743_wire_constant & RPIPE_FREE_Q_1744_wire;
      rx_buffer_pointer_32_1747 <= data_out(32 downto 1);
      status_1747 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 37,
        owidth => 37,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => popFromQueue_call_reqs(0),
          ackR => popFromQueue_call_acks(0),
          dataR => popFromQueue_call_data(36 downto 0),
          tagR => popFromQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 33,
          owidth => 33,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => popFromQueue_return_acks(0), -- cross-over
          ackL => popFromQueue_return_reqs(0), -- cross-over
          dataL => popFromQueue_return_data(32 downto 0),
          tagL => popFromQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1759_call call_stmt_1813_call 
    AccessRegister_call_group_1: Block -- 
      signal data_in: std_logic_vector(85 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => true, 1 => true);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 4, 1 => 4);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1759_call_req_0;
      reqL_unguarded(0) <= call_stmt_1813_call_req_0;
      call_stmt_1759_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1813_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1759_call_req_1;
      reqR_unguarded(0) <= call_stmt_1813_call_req_1;
      call_stmt_1759_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1813_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= ok_flag_1786(0);
      guard_vector(1)  <=  not status_1747(0);
      AccessRegister_call_group_1_accessRegulator_0: access_regulator_base generic map (name => "AccessRegister_call_group_1_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      AccessRegister_call_group_1_accessRegulator_1: access_regulator_base generic map (name => "AccessRegister_call_group_1_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      AccessRegister_call_group_1_gI: SplitGuardInterface generic map(name => "AccessRegister_call_group_1_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1752_wire_constant & NOT_u4_u4_1755_wire_constant & konst_1756_wire_constant & rx_buffer_pointer_32_1747 & type_cast_1806_wire_constant & NOT_u4_u4_1809_wire_constant & konst_1810_wire_constant & pkt_cnt_1778_delayed_13_0_1803;
      ignore_resp0_1759 <= data_out(63 downto 32);
      ignore_resp1_1813 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 86,
        owidth => 43,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 2,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => AccessRegister_call_reqs(0),
          ackR => AccessRegister_call_acks(0),
          dataR => AccessRegister_call_data(42 downto 0),
          tagR => AccessRegister_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => AccessRegister_return_acks(0), -- cross-over
          ackL => AccessRegister_return_reqs(0), -- cross-over
          dataL => AccessRegister_return_data(31 downto 0),
          tagL => AccessRegister_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1776_call 
    loadBuffer_call_group_2: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 10);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1776_call_req_0;
      call_stmt_1776_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1776_call_req_1;
      call_stmt_1776_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not status_1747(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      loadBuffer_call_group_2_gI: SplitGuardInterface generic map(name => "loadBuffer_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_buffer_pointer_36_1765;
      bad_packet_identifier_1776 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => loadBuffer_call_reqs(0),
          ackR => loadBuffer_call_acks(0),
          dataR => loadBuffer_call_data(35 downto 0),
          tagR => loadBuffer_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => loadBuffer_return_acks(0), -- cross-over
          ackL => loadBuffer_return_reqs(0), -- cross-over
          dataL => loadBuffer_return_data(0 downto 0),
          tagL => loadBuffer_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_1838_call 
    populateRxQueue_call_group_3: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1838_call_req_0;
      call_stmt_1838_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1838_call_req_1;
      call_stmt_1838_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= ok_flag_1786(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      populateRxQueue_call_group_3_gI: SplitGuardInterface generic map(name => "populateRxQueue_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_buffer_pointer_36_1795_delayed_10_0_1835;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => populateRxQueue_call_reqs(0),
          ackR => populateRxQueue_call_acks(0),
          dataR => populateRxQueue_call_data(35 downto 0),
          tagR => populateRxQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => populateRxQueue_return_acks(0), -- cross-over
          ackL => populateRxQueue_return_reqs(0), -- cross-over
          tagL => populateRxQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- shared call operator group (4) : call_stmt_1851_call 
    pushIntoQueue_call_group_4: Block -- 
      signal data_in: std_logic_vector(68 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1851_call_req_0;
      call_stmt_1851_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1851_call_req_1;
      call_stmt_1851_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= free_flag_1795(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      pushIntoQueue_call_group_4_gI: SplitGuardInterface generic map(name => "pushIntoQueue_call_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1846_wire_constant & RPIPE_FREE_Q_1847_wire & slice_1849_wire;
      push_status_1851 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 69,
        owidth => 69,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => pushIntoQueue_call_reqs(0),
          ackR => pushIntoQueue_call_acks(0),
          dataR => pushIntoQueue_call_data(68 downto 0),
          tagR => pushIntoQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => pushIntoQueue_return_acks(0), -- cross-over
          ackL => pushIntoQueue_return_reqs(0), -- cross-over
          dataL => pushIntoQueue_return_data(0 downto 0),
          tagL => pushIntoQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 4
    -- 
  end Block; -- data_path
  -- 
end ReceiveEngineDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.nic_system_global_package.all;
entity SoftwareRegisterAccessDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lr_addr : out  std_logic_vector(5 downto 0);
    memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
    memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
    AFB_NIC_REQUEST_pipe_read_req : out  std_logic_vector(0 downto 0);
    AFB_NIC_REQUEST_pipe_read_ack : in   std_logic_vector(0 downto 0);
    AFB_NIC_REQUEST_pipe_read_data : in   std_logic_vector(73 downto 0);
    MAC_ENABLE : in std_logic_vector(0 downto 0);
    AFB_NIC_RESPONSE_pipe_write_req : out  std_logic_vector(0 downto 0);
    AFB_NIC_RESPONSE_pipe_write_ack : in   std_logic_vector(0 downto 0);
    AFB_NIC_RESPONSE_pipe_write_data : out  std_logic_vector(32 downto 0);
    CONTROL_REGISTER_pipe_write_req : out  std_logic_vector(0 downto 0);
    CONTROL_REGISTER_pipe_write_ack : in   std_logic_vector(0 downto 0);
    CONTROL_REGISTER_pipe_write_data : out  std_logic_vector(31 downto 0);
    FREE_Q_pipe_write_req : out  std_logic_vector(0 downto 0);
    FREE_Q_pipe_write_ack : in   std_logic_vector(0 downto 0);
    FREE_Q_pipe_write_data : out  std_logic_vector(35 downto 0);
    NUMBER_OF_SERVERS_pipe_write_req : out  std_logic_vector(0 downto 0);
    NUMBER_OF_SERVERS_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NUMBER_OF_SERVERS_pipe_write_data : out  std_logic_vector(31 downto 0);
    enable_mac_pipe_write_req : out  std_logic_vector(0 downto 0);
    enable_mac_pipe_write_ack : in   std_logic_vector(0 downto 0);
    enable_mac_pipe_write_data : out  std_logic_vector(0 downto 0);
    UpdateRegister_call_reqs : out  std_logic_vector(0 downto 0);
    UpdateRegister_call_acks : in   std_logic_vector(0 downto 0);
    UpdateRegister_call_data : out  std_logic_vector(73 downto 0);
    UpdateRegister_call_tag  :  out  std_logic_vector(0 downto 0);
    UpdateRegister_return_reqs : out  std_logic_vector(0 downto 0);
    UpdateRegister_return_acks : in   std_logic_vector(0 downto 0);
    UpdateRegister_return_data : in   std_logic_vector(31 downto 0);
    UpdateRegister_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity SoftwareRegisterAccessDaemon;
architecture SoftwareRegisterAccessDaemon_arch of SoftwareRegisterAccessDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal SoftwareRegisterAccessDaemon_CP_2867_start: Boolean;
  signal SoftwareRegisterAccessDaemon_CP_2867_symbol: Boolean;
  -- volatile/operator module components. 
  component UpdateRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      bmask : in  std_logic_vector(3 downto 0);
      rval : in  std_logic_vector(31 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      index : in  std_logic_vector(5 downto 0);
      wval : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(5 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal array_obj_ref_1899_load_0_ack_1 : boolean;
  signal phi_stmt_1874_ack_0 : boolean;
  signal WPIPE_CONTROL_REGISTER_1928_inst_ack_1 : boolean;
  signal phi_stmt_1880_req_1 : boolean;
  signal phi_stmt_1890_ack_0 : boolean;
  signal phi_stmt_1890_req_0 : boolean;
  signal array_obj_ref_1930_load_0_ack_0 : boolean;
  signal WPIPE_CONTROL_REGISTER_1928_inst_ack_0 : boolean;
  signal phi_stmt_1880_req_0 : boolean;
  signal array_obj_ref_1899_load_0_req_1 : boolean;
  signal phi_stmt_1874_req_1 : boolean;
  signal check_free_q_2003_1889_buf_req_0 : boolean;
  signal W_update_control_register_pipe_1887_delayed_5_0_1932_inst_req_0 : boolean;
  signal WPIPE_CONTROL_REGISTER_1928_inst_req_1 : boolean;
  signal check_num_server_2012_1894_buf_ack_1 : boolean;
  signal check_num_server_2012_1894_buf_req_1 : boolean;
  signal phi_stmt_1890_req_1 : boolean;
  signal check_num_server_2012_1894_buf_ack_0 : boolean;
  signal check_num_server_2012_1894_buf_req_0 : boolean;
  signal check_control_regsiter_1994_1882_buf_ack_1 : boolean;
  signal array_obj_ref_1930_load_0_req_0 : boolean;
  signal array_obj_ref_1930_load_0_ack_1 : boolean;
  signal check_control_regsiter_1994_1882_buf_req_1 : boolean;
  signal check_control_regsiter_1994_1882_buf_ack_0 : boolean;
  signal phi_stmt_1885_ack_0 : boolean;
  signal array_obj_ref_1930_load_0_req_1 : boolean;
  signal check_control_regsiter_1994_1882_buf_req_0 : boolean;
  signal phi_stmt_1885_req_0 : boolean;
  signal check_free_q_2003_1889_buf_ack_1 : boolean;
  signal check_free_q_2003_1889_buf_req_1 : boolean;
  signal do_while_stmt_1872_branch_req_0 : boolean;
  signal phi_stmt_1885_req_1 : boolean;
  signal WPIPE_CONTROL_REGISTER_1928_inst_req_0 : boolean;
  signal array_obj_ref_1899_load_0_ack_0 : boolean;
  signal array_obj_ref_1899_load_0_req_0 : boolean;
  signal phi_stmt_1880_ack_0 : boolean;
  signal check_free_q_2003_1889_buf_ack_0 : boolean;
  signal W_update_control_register_pipe_1887_delayed_5_0_1932_inst_ack_0 : boolean;
  signal phi_stmt_1874_req_0 : boolean;
  signal if_stmt_1866_branch_req_0 : boolean;
  signal if_stmt_1866_branch_ack_1 : boolean;
  signal if_stmt_1866_branch_ack_0 : boolean;
  signal W_update_control_register_pipe_1887_delayed_5_0_1932_inst_req_1 : boolean;
  signal W_update_control_register_pipe_1887_delayed_5_0_1932_inst_ack_1 : boolean;
  signal array_obj_ref_1938_load_0_req_0 : boolean;
  signal array_obj_ref_1938_load_0_ack_0 : boolean;
  signal array_obj_ref_1938_load_0_req_1 : boolean;
  signal array_obj_ref_1938_load_0_ack_1 : boolean;
  signal EQ_u32_u1_1941_inst_req_0 : boolean;
  signal EQ_u32_u1_1941_inst_ack_0 : boolean;
  signal EQ_u32_u1_1941_inst_req_1 : boolean;
  signal EQ_u32_u1_1941_inst_ack_1 : boolean;
  signal WPIPE_enable_mac_1936_inst_req_0 : boolean;
  signal WPIPE_enable_mac_1936_inst_ack_0 : boolean;
  signal WPIPE_enable_mac_1936_inst_req_1 : boolean;
  signal WPIPE_enable_mac_1936_inst_ack_1 : boolean;
  signal array_obj_ref_1946_load_0_req_0 : boolean;
  signal array_obj_ref_1946_load_0_ack_0 : boolean;
  signal array_obj_ref_1946_load_0_req_1 : boolean;
  signal array_obj_ref_1946_load_0_ack_1 : boolean;
  signal W_update_free_q_pipe_1900_delayed_5_0_1948_inst_req_0 : boolean;
  signal W_update_free_q_pipe_1900_delayed_5_0_1948_inst_ack_0 : boolean;
  signal W_update_free_q_pipe_1900_delayed_5_0_1948_inst_req_1 : boolean;
  signal W_update_free_q_pipe_1900_delayed_5_0_1948_inst_ack_1 : boolean;
  signal type_cast_1954_inst_req_0 : boolean;
  signal type_cast_1954_inst_ack_0 : boolean;
  signal type_cast_1954_inst_req_1 : boolean;
  signal type_cast_1954_inst_ack_1 : boolean;
  signal WPIPE_FREE_Q_1952_inst_req_0 : boolean;
  signal WPIPE_FREE_Q_1952_inst_ack_0 : boolean;
  signal WPIPE_FREE_Q_1952_inst_req_1 : boolean;
  signal WPIPE_FREE_Q_1952_inst_ack_1 : boolean;
  signal array_obj_ref_1959_load_0_req_0 : boolean;
  signal array_obj_ref_1959_load_0_ack_0 : boolean;
  signal array_obj_ref_1959_load_0_req_1 : boolean;
  signal array_obj_ref_1959_load_0_ack_1 : boolean;
  signal WPIPE_NUMBER_OF_SERVERS_1957_inst_req_0 : boolean;
  signal WPIPE_NUMBER_OF_SERVERS_1957_inst_ack_0 : boolean;
  signal WPIPE_NUMBER_OF_SERVERS_1957_inst_req_1 : boolean;
  signal WPIPE_NUMBER_OF_SERVERS_1957_inst_ack_1 : boolean;
  signal RPIPE_AFB_NIC_REQUEST_1962_inst_req_0 : boolean;
  signal RPIPE_AFB_NIC_REQUEST_1962_inst_ack_0 : boolean;
  signal RPIPE_AFB_NIC_REQUEST_1962_inst_req_1 : boolean;
  signal RPIPE_AFB_NIC_REQUEST_1962_inst_ack_1 : boolean;
  signal array_obj_ref_2015_load_0_req_0 : boolean;
  signal array_obj_ref_2015_load_0_ack_0 : boolean;
  signal array_obj_ref_2015_load_0_req_1 : boolean;
  signal array_obj_ref_2015_load_0_ack_1 : boolean;
  signal W_rwbar_1966_delayed_5_0_2017_inst_req_0 : boolean;
  signal W_rwbar_1966_delayed_5_0_2017_inst_ack_0 : boolean;
  signal W_rwbar_1966_delayed_5_0_2017_inst_req_1 : boolean;
  signal W_rwbar_1966_delayed_5_0_2017_inst_ack_1 : boolean;
  signal W_bmask_1967_delayed_5_0_2020_inst_req_0 : boolean;
  signal W_bmask_1967_delayed_5_0_2020_inst_ack_0 : boolean;
  signal W_bmask_1967_delayed_5_0_2020_inst_req_1 : boolean;
  signal W_bmask_1967_delayed_5_0_2020_inst_ack_1 : boolean;
  signal W_wdata_1969_delayed_5_0_2023_inst_req_0 : boolean;
  signal W_wdata_1969_delayed_5_0_2023_inst_ack_0 : boolean;
  signal W_wdata_1969_delayed_5_0_2023_inst_req_1 : boolean;
  signal W_wdata_1969_delayed_5_0_2023_inst_ack_1 : boolean;
  signal W_index_1970_delayed_5_0_2026_inst_req_0 : boolean;
  signal W_index_1970_delayed_5_0_2026_inst_ack_0 : boolean;
  signal W_index_1970_delayed_5_0_2026_inst_req_1 : boolean;
  signal W_index_1970_delayed_5_0_2026_inst_ack_1 : boolean;
  signal call_stmt_2035_call_req_0 : boolean;
  signal call_stmt_2035_call_ack_0 : boolean;
  signal call_stmt_2035_call_req_1 : boolean;
  signal call_stmt_2035_call_ack_1 : boolean;
  signal W_rwbar_1974_delayed_5_0_2036_inst_req_0 : boolean;
  signal W_rwbar_1974_delayed_5_0_2036_inst_ack_0 : boolean;
  signal W_rwbar_1974_delayed_5_0_2036_inst_req_1 : boolean;
  signal W_rwbar_1974_delayed_5_0_2036_inst_ack_1 : boolean;
  signal WPIPE_AFB_NIC_RESPONSE_2052_inst_req_0 : boolean;
  signal WPIPE_AFB_NIC_RESPONSE_2052_inst_ack_0 : boolean;
  signal WPIPE_AFB_NIC_RESPONSE_2052_inst_req_1 : boolean;
  signal WPIPE_AFB_NIC_RESPONSE_2052_inst_ack_1 : boolean;
  signal do_while_stmt_1872_branch_ack_0 : boolean;
  signal do_while_stmt_1872_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "SoftwareRegisterAccessDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  SoftwareRegisterAccessDaemon_CP_2867_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "SoftwareRegisterAccessDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= SoftwareRegisterAccessDaemon_CP_2867_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= SoftwareRegisterAccessDaemon_CP_2867_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= SoftwareRegisterAccessDaemon_CP_2867_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  SoftwareRegisterAccessDaemon_CP_2867: Block -- control-path 
    signal SoftwareRegisterAccessDaemon_CP_2867_elements: BooleanArray(185 downto 0);
    -- 
  begin -- 
    SoftwareRegisterAccessDaemon_CP_2867_elements(0) <= SoftwareRegisterAccessDaemon_CP_2867_start;
    SoftwareRegisterAccessDaemon_CP_2867_symbol <= SoftwareRegisterAccessDaemon_CP_2867_elements(1);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	185 
    -- CP-element group 0:  members (7) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1862/$entry
      -- CP-element group 0: 	 branch_block_stmt_1862/branch_block_stmt_1862__entry__
      -- CP-element group 0: 	 branch_block_stmt_1862/merge_stmt_1863__entry__
      -- CP-element group 0: 	 branch_block_stmt_1862/merge_stmt_1863_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_1862/merge_stmt_1863__entry___PhiReq/$entry
      -- CP-element group 0: 	 branch_block_stmt_1862/merge_stmt_1863__entry___PhiReq/$exit
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	184 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1862/$exit
      -- CP-element group 1: 	 branch_block_stmt_1862/branch_block_stmt_1862__exit__
      -- CP-element group 1: 	 branch_block_stmt_1862/do_while_stmt_1872__exit__
      -- 
    SoftwareRegisterAccessDaemon_CP_2867_elements(1) <= SoftwareRegisterAccessDaemon_CP_2867_elements(184);
    -- CP-element group 2:  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	185 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	185 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 branch_block_stmt_1862/if_stmt_1866_if_link/$exit
      -- CP-element group 2: 	 branch_block_stmt_1862/if_stmt_1866_if_link/if_choice_transition
      -- CP-element group 2: 	 branch_block_stmt_1862/not_mac_enable_loopback
      -- CP-element group 2: 	 branch_block_stmt_1862/not_mac_enable_loopback_PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_1862/not_mac_enable_loopback_PhiReq/$exit
      -- 
    if_choice_transition_2925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1866_branch_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(2)); -- 
    -- CP-element group 3:  merge  transition  place  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	185 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (4) 
      -- CP-element group 3: 	 branch_block_stmt_1862/if_stmt_1866__exit__
      -- CP-element group 3: 	 branch_block_stmt_1862/do_while_stmt_1872__entry__
      -- CP-element group 3: 	 branch_block_stmt_1862/if_stmt_1866_else_link/$exit
      -- CP-element group 3: 	 branch_block_stmt_1862/if_stmt_1866_else_link/else_choice_transition
      -- 
    else_choice_transition_2929_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1866_branch_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(3)); -- 
    -- CP-element group 4:  transition  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	10 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 branch_block_stmt_1862/do_while_stmt_1872/$entry
      -- CP-element group 4: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872__entry__
      -- 
    SoftwareRegisterAccessDaemon_CP_2867_elements(4) <= SoftwareRegisterAccessDaemon_CP_2867_elements(3);
    -- CP-element group 5:  merge  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	184 
    -- CP-element group 5:  members (1) 
      -- CP-element group 5: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872__exit__
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(5) is bound as output of CP function.
    -- CP-element group 6:  merge  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1862/do_while_stmt_1872/loop_back
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(6) is bound as output of CP function.
    -- CP-element group 7:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	12 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	182 
    -- CP-element group 7: 	183 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_1862/do_while_stmt_1872/condition_done
      -- CP-element group 7: 	 branch_block_stmt_1862/do_while_stmt_1872/loop_exit/$entry
      -- CP-element group 7: 	 branch_block_stmt_1862/do_while_stmt_1872/loop_taken/$entry
      -- 
    SoftwareRegisterAccessDaemon_CP_2867_elements(7) <= SoftwareRegisterAccessDaemon_CP_2867_elements(12);
    -- CP-element group 8:  branch  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	181 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1862/do_while_stmt_1872/loop_body_done
      -- 
    SoftwareRegisterAccessDaemon_CP_2867_elements(8) <= SoftwareRegisterAccessDaemon_CP_2867_elements(181);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	21 
    -- CP-element group 9: 	40 
    -- CP-element group 9: 	59 
    -- CP-element group 9: 	78 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/back_edge_to_loop_body
      -- 
    SoftwareRegisterAccessDaemon_CP_2867_elements(9) <= SoftwareRegisterAccessDaemon_CP_2867_elements(6);
    -- CP-element group 10:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	4 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	23 
    -- CP-element group 10: 	42 
    -- CP-element group 10: 	61 
    -- CP-element group 10: 	80 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/first_time_through_loop_body
      -- 
    SoftwareRegisterAccessDaemon_CP_2867_elements(10) <= SoftwareRegisterAccessDaemon_CP_2867_elements(4);
    -- CP-element group 11:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	95 
    -- CP-element group 11: 	17 
    -- CP-element group 11: 	18 
    -- CP-element group 11: 	117 
    -- CP-element group 11: 	132 
    -- CP-element group 11: 	174 
    -- CP-element group 11: 	139 
    -- CP-element group 11: 	91 
    -- CP-element group 11: 	108 
    -- CP-element group 11: 	34 
    -- CP-element group 11: 	35 
    -- CP-element group 11: 	53 
    -- CP-element group 11: 	54 
    -- CP-element group 11: 	72 
    -- CP-element group 11: 	73 
    -- CP-element group 11:  members (12) 
      -- CP-element group 11: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1899_word_address_calculated
      -- CP-element group 11: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1899_root_address_calculated
      -- CP-element group 11: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1930_word_address_calculated
      -- CP-element group 11: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1930_root_address_calculated
      -- CP-element group 11: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/$entry
      -- CP-element group 11: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/loop_body_start
      -- CP-element group 11: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1938_word_address_calculated
      -- CP-element group 11: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1938_root_address_calculated
      -- CP-element group 11: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1946_word_address_calculated
      -- CP-element group 11: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1946_root_address_calculated
      -- CP-element group 11: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1959_word_address_calculated
      -- CP-element group 11: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1959_root_address_calculated
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(11) is bound as output of CP function.
    -- CP-element group 12:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	16 
    -- CP-element group 12: 	174 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	7 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/condition_evaluated
      -- 
    condition_evaluated_2945_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2945_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(12), ack => do_while_stmt_1872_branch_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(16) & SoftwareRegisterAccessDaemon_CP_2867_elements(174);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	17 
    -- CP-element group 13: 	34 
    -- CP-element group 13: 	53 
    -- CP-element group 13: 	72 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	36 
    -- CP-element group 13: 	55 
    -- CP-element group 13: 	74 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1874_sample_start__ps
      -- CP-element group 13: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/aggregated_phi_sample_req
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 31,1 => 31,2 => 31,3 => 31,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(17) & SoftwareRegisterAccessDaemon_CP_2867_elements(34) & SoftwareRegisterAccessDaemon_CP_2867_elements(53) & SoftwareRegisterAccessDaemon_CP_2867_elements(72) & SoftwareRegisterAccessDaemon_CP_2867_elements(16);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	19 
    -- CP-element group 14: 	37 
    -- CP-element group 14: 	56 
    -- CP-element group 14: 	75 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	140 
    -- CP-element group 14: 	181 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	17 
    -- CP-element group 14: 	34 
    -- CP-element group 14: 	53 
    -- CP-element group 14: 	72 
    -- CP-element group 14:  members (5) 
      -- CP-element group 14: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1885_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1880_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1874_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1890_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/aggregated_phi_sample_ack
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 31,2 => 31,3 => 31);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(19) & SoftwareRegisterAccessDaemon_CP_2867_elements(37) & SoftwareRegisterAccessDaemon_CP_2867_elements(56) & SoftwareRegisterAccessDaemon_CP_2867_elements(75);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	18 
    -- CP-element group 15: 	35 
    -- CP-element group 15: 	54 
    -- CP-element group 15: 	73 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	38 
    -- CP-element group 15: 	57 
    -- CP-element group 15: 	76 
    -- CP-element group 15:  members (2) 
      -- CP-element group 15: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1874_update_start__ps
      -- CP-element group 15: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/aggregated_phi_update_req
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 31,2 => 31,3 => 31);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(18) & SoftwareRegisterAccessDaemon_CP_2867_elements(35) & SoftwareRegisterAccessDaemon_CP_2867_elements(54) & SoftwareRegisterAccessDaemon_CP_2867_elements(73);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	20 
    -- CP-element group 16: 	39 
    -- CP-element group 16: 	58 
    -- CP-element group 16: 	77 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	12 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/aggregated_phi_update_ack
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 31,2 => 31,3 => 31);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(20) & SoftwareRegisterAccessDaemon_CP_2867_elements(39) & SoftwareRegisterAccessDaemon_CP_2867_elements(58) & SoftwareRegisterAccessDaemon_CP_2867_elements(77);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	13 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1874_sample_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(11) & SoftwareRegisterAccessDaemon_CP_2867_elements(14);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	11 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	97 
    -- CP-element group 18: 	119 
    -- CP-element group 18: 	134 
    -- CP-element group 18: 	137 
    -- CP-element group 18: 	123 
    -- CP-element group 18: 	104 
    -- CP-element group 18: 	100 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	15 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1874_update_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 31,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(11) & SoftwareRegisterAccessDaemon_CP_2867_elements(97) & SoftwareRegisterAccessDaemon_CP_2867_elements(119) & SoftwareRegisterAccessDaemon_CP_2867_elements(134) & SoftwareRegisterAccessDaemon_CP_2867_elements(137) & SoftwareRegisterAccessDaemon_CP_2867_elements(123) & SoftwareRegisterAccessDaemon_CP_2867_elements(104) & SoftwareRegisterAccessDaemon_CP_2867_elements(100);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	14 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1874_sample_completed__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(19) is bound as output of CP function.
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	95 
    -- CP-element group 20: 	16 
    -- CP-element group 20: 	117 
    -- CP-element group 20: 	136 
    -- CP-element group 20: 	132 
    -- CP-element group 20: 	121 
    -- CP-element group 20: 	102 
    -- CP-element group 20: 	99 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1874_update_completed__ps
      -- CP-element group 20: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1874_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	9 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1874_loopback_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_2867_elements(21) <= SoftwareRegisterAccessDaemon_CP_2867_elements(9);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1874_loopback_sample_req
      -- CP-element group 22: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1874_loopback_sample_req_ps
      -- 
    phi_stmt_1874_loopback_sample_req_2960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1874_loopback_sample_req_2960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(22), ack => phi_stmt_1874_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	10 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1874_entry_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_2867_elements(23) <= SoftwareRegisterAccessDaemon_CP_2867_elements(10);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1874_entry_sample_req_ps
      -- CP-element group 24: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1874_entry_sample_req
      -- 
    phi_stmt_1874_entry_sample_req_2963_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1874_entry_sample_req_2963_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(24), ack => phi_stmt_1874_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1874_phi_mux_ack
      -- CP-element group 25: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1874_phi_mux_ack_ps
      -- 
    phi_stmt_1874_phi_mux_ack_2966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1874_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1877_sample_start__ps
      -- CP-element group 26: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1877_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1877_sample_start_
      -- CP-element group 26: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1877_sample_completed__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1877_update_start_
      -- CP-element group 27: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1877_update_start__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	29 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1877_update_completed__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_2867_elements(28) <= SoftwareRegisterAccessDaemon_CP_2867_elements(29);
    -- CP-element group 29:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	28 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1877_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(29) is a control-delay.
    cp_element_29_delay: control_delay_element  generic map(name => " 29_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2867_elements(27), ack => SoftwareRegisterAccessDaemon_CP_2867_elements(29), clk => clk, reset =>reset);
    -- CP-element group 30:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1879_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1879_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1879_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1879_sample_start__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1879_update_start_
      -- CP-element group 31: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1879_update_start__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	33 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1879_update_completed__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_2867_elements(32) <= SoftwareRegisterAccessDaemon_CP_2867_elements(33);
    -- CP-element group 33:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	32 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1879_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(33) is a control-delay.
    cp_element_33_delay: control_delay_element  generic map(name => " 33_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2867_elements(31), ack => SoftwareRegisterAccessDaemon_CP_2867_elements(33), clk => clk, reset =>reset);
    -- CP-element group 34:  join  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	11 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	14 
    -- CP-element group 34: 	142 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	13 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1880_sample_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(11) & SoftwareRegisterAccessDaemon_CP_2867_elements(14) & SoftwareRegisterAccessDaemon_CP_2867_elements(142);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	11 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	97 
    -- CP-element group 35: 	104 
    -- CP-element group 35: 	100 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	15 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1880_update_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(11) & SoftwareRegisterAccessDaemon_CP_2867_elements(97) & SoftwareRegisterAccessDaemon_CP_2867_elements(104) & SoftwareRegisterAccessDaemon_CP_2867_elements(100);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	13 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1880_sample_start__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_2867_elements(36) <= SoftwareRegisterAccessDaemon_CP_2867_elements(13);
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	14 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1880_sample_completed__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(37) is bound as output of CP function.
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	15 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1880_update_start__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_2867_elements(38) <= SoftwareRegisterAccessDaemon_CP_2867_elements(15);
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	95 
    -- CP-element group 39: 	16 
    -- CP-element group 39: 	102 
    -- CP-element group 39: 	99 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1880_update_completed__ps
      -- CP-element group 39: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1880_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	9 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1880_loopback_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_2867_elements(40) <= SoftwareRegisterAccessDaemon_CP_2867_elements(9);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1880_loopback_sample_req
      -- CP-element group 41: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1880_loopback_sample_req_ps
      -- 
    phi_stmt_1880_loopback_sample_req_2994_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1880_loopback_sample_req_2994_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(41), ack => phi_stmt_1880_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	10 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1880_entry_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_2867_elements(42) <= SoftwareRegisterAccessDaemon_CP_2867_elements(10);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1880_entry_sample_req
      -- CP-element group 43: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1880_entry_sample_req_ps
      -- 
    phi_stmt_1880_entry_sample_req_2997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1880_entry_sample_req_2997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(43), ack => phi_stmt_1880_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1880_phi_mux_ack_ps
      -- CP-element group 44: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1880_phi_mux_ack
      -- 
    phi_stmt_1880_phi_mux_ack_3000_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1880_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(44)); -- 
    -- CP-element group 45:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	47 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_control_regsiter_1882_Sample/req
      -- CP-element group 45: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_control_regsiter_1882_Sample/$entry
      -- CP-element group 45: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_control_regsiter_1882_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_control_regsiter_1882_sample_start__ps
      -- 
    req_3013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(45), ack => check_control_regsiter_1994_1882_buf_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (4) 
      -- CP-element group 46: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_control_regsiter_1882_Update/req
      -- CP-element group 46: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_control_regsiter_1882_Update/$entry
      -- CP-element group 46: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_control_regsiter_1882_update_start_
      -- CP-element group 46: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_control_regsiter_1882_update_start__ps
      -- 
    req_3018_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3018_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(46), ack => check_control_regsiter_1994_1882_buf_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	45 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (4) 
      -- CP-element group 47: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_control_regsiter_1882_Sample/ack
      -- CP-element group 47: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_control_regsiter_1882_Sample/$exit
      -- CP-element group 47: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_control_regsiter_1882_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_control_regsiter_1882_sample_completed__ps
      -- 
    ack_3014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_control_regsiter_1994_1882_buf_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(47)); -- 
    -- CP-element group 48:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (4) 
      -- CP-element group 48: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_control_regsiter_1882_Update/ack
      -- CP-element group 48: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_control_regsiter_1882_Update/$exit
      -- CP-element group 48: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_control_regsiter_1882_update_completed_
      -- CP-element group 48: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_control_regsiter_1882_update_completed__ps
      -- 
    ack_3019_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_control_regsiter_1994_1882_buf_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(48)); -- 
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1884_sample_completed_
      -- CP-element group 49: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1884_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1884_sample_completed__ps
      -- CP-element group 49: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1884_sample_start__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (2) 
      -- CP-element group 50: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1884_update_start_
      -- CP-element group 50: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1884_update_start__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	52 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1884_update_completed__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_2867_elements(51) <= SoftwareRegisterAccessDaemon_CP_2867_elements(52);
    -- CP-element group 52:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	51 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1884_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(52) is a control-delay.
    cp_element_52_delay: control_delay_element  generic map(name => " 52_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2867_elements(50), ack => SoftwareRegisterAccessDaemon_CP_2867_elements(52), clk => clk, reset =>reset);
    -- CP-element group 53:  join  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	11 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	14 
    -- CP-element group 53: 	142 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	13 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1885_sample_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(11) & SoftwareRegisterAccessDaemon_CP_2867_elements(14) & SoftwareRegisterAccessDaemon_CP_2867_elements(142);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	11 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	119 
    -- CP-element group 54: 	123 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	15 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1885_update_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(11) & SoftwareRegisterAccessDaemon_CP_2867_elements(119) & SoftwareRegisterAccessDaemon_CP_2867_elements(123);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	13 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1885_sample_start__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_2867_elements(55) <= SoftwareRegisterAccessDaemon_CP_2867_elements(13);
    -- CP-element group 56:  join  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	14 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1885_sample_completed__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(56) is bound as output of CP function.
    -- CP-element group 57:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	15 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1885_update_start__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_2867_elements(57) <= SoftwareRegisterAccessDaemon_CP_2867_elements(15);
    -- CP-element group 58:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	16 
    -- CP-element group 58: 	117 
    -- CP-element group 58: 	121 
    -- CP-element group 58:  members (2) 
      -- CP-element group 58: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1885_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1885_update_completed__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(58) is bound as output of CP function.
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	9 
    -- CP-element group 59: successors 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1885_loopback_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_2867_elements(59) <= SoftwareRegisterAccessDaemon_CP_2867_elements(9);
    -- CP-element group 60:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (2) 
      -- CP-element group 60: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1885_loopback_sample_req_ps
      -- CP-element group 60: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1885_loopback_sample_req
      -- 
    phi_stmt_1885_loopback_sample_req_3038_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1885_loopback_sample_req_3038_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(60), ack => phi_stmt_1885_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(60) is bound as output of CP function.
    -- CP-element group 61:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	10 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1885_entry_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_2867_elements(61) <= SoftwareRegisterAccessDaemon_CP_2867_elements(10);
    -- CP-element group 62:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1885_entry_sample_req_ps
      -- CP-element group 62: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1885_entry_sample_req
      -- 
    phi_stmt_1885_entry_sample_req_3041_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1885_entry_sample_req_3041_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(62), ack => phi_stmt_1885_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(62) is bound as output of CP function.
    -- CP-element group 63:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1885_phi_mux_ack_ps
      -- CP-element group 63: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1885_phi_mux_ack
      -- 
    phi_stmt_1885_phi_mux_ack_3044_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1885_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(63)); -- 
    -- CP-element group 64:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (4) 
      -- CP-element group 64: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1888_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1888_sample_start_
      -- CP-element group 64: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1888_sample_completed__ps
      -- CP-element group 64: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1888_sample_start__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(64) is bound as output of CP function.
    -- CP-element group 65:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1888_update_start_
      -- CP-element group 65: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1888_update_start__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(65) is bound as output of CP function.
    -- CP-element group 66:  join  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (1) 
      -- CP-element group 66: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1888_update_completed__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_2867_elements(66) <= SoftwareRegisterAccessDaemon_CP_2867_elements(67);
    -- CP-element group 67:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	66 
    -- CP-element group 67:  members (1) 
      -- CP-element group 67: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1888_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(67) is a control-delay.
    cp_element_67_delay: control_delay_element  generic map(name => " 67_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2867_elements(65), ack => SoftwareRegisterAccessDaemon_CP_2867_elements(67), clk => clk, reset =>reset);
    -- CP-element group 68:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_free_q_1889_sample_start_
      -- CP-element group 68: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_free_q_1889_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_free_q_1889_sample_start__ps
      -- CP-element group 68: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_free_q_1889_Sample/req
      -- 
    req_3065_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3065_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(68), ack => check_free_q_2003_1889_buf_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(68) is bound as output of CP function.
    -- CP-element group 69:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_free_q_1889_update_start__ps
      -- CP-element group 69: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_free_q_1889_update_start_
      -- CP-element group 69: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_free_q_1889_Update/req
      -- CP-element group 69: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_free_q_1889_Update/$entry
      -- 
    req_3070_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3070_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(69), ack => check_free_q_2003_1889_buf_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(69) is bound as output of CP function.
    -- CP-element group 70:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70:  members (4) 
      -- CP-element group 70: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_free_q_1889_sample_completed_
      -- CP-element group 70: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_free_q_1889_sample_completed__ps
      -- CP-element group 70: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_free_q_1889_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_free_q_1889_Sample/ack
      -- 
    ack_3066_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_free_q_2003_1889_buf_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(70)); -- 
    -- CP-element group 71:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (4) 
      -- CP-element group 71: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_free_q_1889_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_free_q_1889_update_completed__ps
      -- CP-element group 71: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_free_q_1889_Update/ack
      -- CP-element group 71: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_free_q_1889_Update/$exit
      -- 
    ack_3071_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_free_q_2003_1889_buf_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(71)); -- 
    -- CP-element group 72:  join  transition  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	11 
    -- CP-element group 72: marked-predecessors 
    -- CP-element group 72: 	14 
    -- CP-element group 72: 	142 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	13 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1890_sample_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(11) & SoftwareRegisterAccessDaemon_CP_2867_elements(14) & SoftwareRegisterAccessDaemon_CP_2867_elements(142);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  join  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	11 
    -- CP-element group 73: marked-predecessors 
    -- CP-element group 73: 	134 
    -- CP-element group 73: 	137 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	15 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1890_update_start_
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(11) & SoftwareRegisterAccessDaemon_CP_2867_elements(134) & SoftwareRegisterAccessDaemon_CP_2867_elements(137);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	13 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1890_sample_start__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_2867_elements(74) <= SoftwareRegisterAccessDaemon_CP_2867_elements(13);
    -- CP-element group 75:  join  transition  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	14 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1890_sample_completed__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(75) is bound as output of CP function.
    -- CP-element group 76:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	15 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1890_update_start__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_2867_elements(76) <= SoftwareRegisterAccessDaemon_CP_2867_elements(15);
    -- CP-element group 77:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	16 
    -- CP-element group 77: 	136 
    -- CP-element group 77: 	132 
    -- CP-element group 77:  members (2) 
      -- CP-element group 77: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1890_update_completed__ps
      -- CP-element group 77: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1890_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(77) is bound as output of CP function.
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	9 
    -- CP-element group 78: successors 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1890_loopback_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_2867_elements(78) <= SoftwareRegisterAccessDaemon_CP_2867_elements(9);
    -- CP-element group 79:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1890_loopback_sample_req_ps
      -- CP-element group 79: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1890_loopback_sample_req
      -- 
    phi_stmt_1890_loopback_sample_req_3082_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1890_loopback_sample_req_3082_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(79), ack => phi_stmt_1890_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(79) is bound as output of CP function.
    -- CP-element group 80:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	10 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (1) 
      -- CP-element group 80: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1890_entry_trigger
      -- 
    SoftwareRegisterAccessDaemon_CP_2867_elements(80) <= SoftwareRegisterAccessDaemon_CP_2867_elements(10);
    -- CP-element group 81:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (2) 
      -- CP-element group 81: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1890_entry_sample_req_ps
      -- CP-element group 81: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1890_entry_sample_req
      -- 
    phi_stmt_1890_entry_sample_req_3085_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1890_entry_sample_req_3085_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(81), ack => phi_stmt_1890_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(81) is bound as output of CP function.
    -- CP-element group 82:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1890_phi_mux_ack
      -- CP-element group 82: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/phi_stmt_1890_phi_mux_ack_ps
      -- 
    phi_stmt_1890_phi_mux_ack_3088_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1890_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(82)); -- 
    -- CP-element group 83:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (4) 
      -- CP-element group 83: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1893_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1893_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1893_sample_completed__ps
      -- CP-element group 83: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1893_sample_start__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(83) is bound as output of CP function.
    -- CP-element group 84:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1893_update_start_
      -- CP-element group 84: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1893_update_start__ps
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(84) is bound as output of CP function.
    -- CP-element group 85:  join  transition  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	86 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1893_update_completed__ps
      -- 
    SoftwareRegisterAccessDaemon_CP_2867_elements(85) <= SoftwareRegisterAccessDaemon_CP_2867_elements(86);
    -- CP-element group 86:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	85 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1893_update_completed_
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(86) is a control-delay.
    cp_element_86_delay: control_delay_element  generic map(name => " 86_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2867_elements(84), ack => SoftwareRegisterAccessDaemon_CP_2867_elements(86), clk => clk, reset =>reset);
    -- CP-element group 87:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (4) 
      -- CP-element group 87: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_num_server_1894_sample_start__ps
      -- CP-element group 87: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_num_server_1894_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_num_server_1894_Sample/req
      -- CP-element group 87: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_num_server_1894_Sample/$entry
      -- 
    req_3109_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3109_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(87), ack => check_num_server_2012_1894_buf_req_0); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(87) is bound as output of CP function.
    -- CP-element group 88:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (4) 
      -- CP-element group 88: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_num_server_1894_update_start__ps
      -- CP-element group 88: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_num_server_1894_update_start_
      -- CP-element group 88: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_num_server_1894_Update/req
      -- CP-element group 88: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_num_server_1894_Update/$entry
      -- 
    req_3114_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3114_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(88), ack => check_num_server_2012_1894_buf_req_1); -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(88) is bound as output of CP function.
    -- CP-element group 89:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: successors 
    -- CP-element group 89:  members (4) 
      -- CP-element group 89: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_num_server_1894_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_num_server_1894_sample_completed__ps
      -- CP-element group 89: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_num_server_1894_Sample/ack
      -- CP-element group 89: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_num_server_1894_Sample/$exit
      -- 
    ack_3110_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_num_server_2012_1894_buf_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(89)); -- 
    -- CP-element group 90:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90:  members (4) 
      -- CP-element group 90: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_num_server_1894_update_completed__ps
      -- CP-element group 90: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_num_server_1894_Update/ack
      -- CP-element group 90: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_num_server_1894_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/R_check_num_server_1894_update_completed_
      -- 
    ack_3115_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => check_num_server_2012_1894_buf_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(90)); -- 
    -- CP-element group 91:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	11 
    -- CP-element group 91: marked-predecessors 
    -- CP-element group 91: 	93 
    -- CP-element group 91: 	166 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (5) 
      -- CP-element group 91: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1899_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1899_Sample/word_access_start/$entry
      -- CP-element group 91: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1899_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1899_Sample/word_access_start/word_0/rr
      -- CP-element group 91: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1899_Sample/word_access_start/word_0/$entry
      -- 
    rr_3133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(91), ack => array_obj_ref_1899_load_0_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(11) & SoftwareRegisterAccessDaemon_CP_2867_elements(93) & SoftwareRegisterAccessDaemon_CP_2867_elements(166);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: marked-predecessors 
    -- CP-element group 92: 	94 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (5) 
      -- CP-element group 92: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1899_Update/word_access_complete/word_0/$entry
      -- CP-element group 92: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1899_Update/word_access_complete/$entry
      -- CP-element group 92: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1899_update_start_
      -- CP-element group 92: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1899_Update/word_access_complete/word_0/cr
      -- CP-element group 92: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1899_Update/$entry
      -- 
    cr_3144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(92), ack => array_obj_ref_1899_load_0_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2867_elements(94);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	175 
    -- CP-element group 93: marked-successors 
    -- CP-element group 93: 	91 
    -- CP-element group 93:  members (5) 
      -- CP-element group 93: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1899_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1899_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1899_Sample/word_access_start/word_0/ra
      -- CP-element group 93: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1899_Sample/word_access_start/word_0/$exit
      -- CP-element group 93: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1899_Sample/word_access_start/$exit
      -- 
    ra_3134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1899_load_0_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(93)); -- 
    -- CP-element group 94:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	181 
    -- CP-element group 94: marked-successors 
    -- CP-element group 94: 	92 
    -- CP-element group 94:  members (9) 
      -- CP-element group 94: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1899_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1899_Update/word_access_complete/word_0/ca
      -- CP-element group 94: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1899_Update/word_access_complete/word_0/$exit
      -- CP-element group 94: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1899_Update/array_obj_ref_1899_Merge/$entry
      -- CP-element group 94: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1899_Update/array_obj_ref_1899_Merge/merge_req
      -- CP-element group 94: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1899_Update/word_access_complete/$exit
      -- CP-element group 94: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1899_Update/array_obj_ref_1899_Merge/merge_ack
      -- CP-element group 94: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1899_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1899_Update/array_obj_ref_1899_Merge/$exit
      -- 
    ca_3145_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1899_load_0_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(94)); -- 
    -- CP-element group 95:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	11 
    -- CP-element group 95: 	20 
    -- CP-element group 95: 	39 
    -- CP-element group 95: marked-predecessors 
    -- CP-element group 95: 	97 
    -- CP-element group 95: 	166 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (5) 
      -- CP-element group 95: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1930_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1930_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1930_Sample/word_access_start/$entry
      -- CP-element group 95: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1930_Sample/word_access_start/word_0/rr
      -- CP-element group 95: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1930_Sample/word_access_start/word_0/$entry
      -- 
    rr_3167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(95), ack => array_obj_ref_1930_load_0_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 31,1 => 31,2 => 31,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(11) & SoftwareRegisterAccessDaemon_CP_2867_elements(20) & SoftwareRegisterAccessDaemon_CP_2867_elements(39) & SoftwareRegisterAccessDaemon_CP_2867_elements(97) & SoftwareRegisterAccessDaemon_CP_2867_elements(166);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: marked-predecessors 
    -- CP-element group 96: 	100 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	98 
    -- CP-element group 96:  members (5) 
      -- CP-element group 96: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1930_update_start_
      -- CP-element group 96: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1930_Update/$entry
      -- CP-element group 96: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1930_Update/word_access_complete/$entry
      -- CP-element group 96: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1930_Update/word_access_complete/word_0/cr
      -- CP-element group 96: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1930_Update/word_access_complete/word_0/$entry
      -- 
    cr_3178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(96), ack => array_obj_ref_1930_load_0_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2867_elements(100);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	176 
    -- CP-element group 97: marked-successors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: 	18 
    -- CP-element group 97: 	35 
    -- CP-element group 97:  members (5) 
      -- CP-element group 97: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1930_sample_completed_
      -- CP-element group 97: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1930_Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1930_Sample/word_access_start/$exit
      -- CP-element group 97: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1930_Sample/word_access_start/word_0/ra
      -- CP-element group 97: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1930_Sample/word_access_start/word_0/$exit
      -- 
    ra_3168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1930_load_0_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(97)); -- 
    -- CP-element group 98:  transition  input  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	96 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	99 
    -- CP-element group 98:  members (9) 
      -- CP-element group 98: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1930_update_completed_
      -- CP-element group 98: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1930_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1930_Update/array_obj_ref_1930_Merge/merge_ack
      -- CP-element group 98: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1930_Update/array_obj_ref_1930_Merge/merge_req
      -- CP-element group 98: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1930_Update/array_obj_ref_1930_Merge/$exit
      -- CP-element group 98: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1930_Update/array_obj_ref_1930_Merge/$entry
      -- CP-element group 98: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1930_Update/word_access_complete/word_0/ca
      -- CP-element group 98: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1930_Update/word_access_complete/word_0/$exit
      -- CP-element group 98: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1930_Update/word_access_complete/$exit
      -- 
    ca_3179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1930_load_0_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(98)); -- 
    -- CP-element group 99:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	20 
    -- CP-element group 99: 	98 
    -- CP-element group 99: 	39 
    -- CP-element group 99: marked-predecessors 
    -- CP-element group 99: 	101 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	100 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_CONTROL_REGISTER_1928_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_CONTROL_REGISTER_1928_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_CONTROL_REGISTER_1928_Sample/req
      -- 
    req_3192_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3192_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(99), ack => WPIPE_CONTROL_REGISTER_1928_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_99: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 1,2 => 31,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 48) := "SoftwareRegisterAccessDaemon_cp_element_group_99"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(20) & SoftwareRegisterAccessDaemon_CP_2867_elements(98) & SoftwareRegisterAccessDaemon_CP_2867_elements(39) & SoftwareRegisterAccessDaemon_CP_2867_elements(101);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_99 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(99), clk => clk, reset => reset); --
    end block;
    -- CP-element group 100:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	99 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	101 
    -- CP-element group 100: marked-successors 
    -- CP-element group 100: 	96 
    -- CP-element group 100: 	18 
    -- CP-element group 100: 	35 
    -- CP-element group 100:  members (6) 
      -- CP-element group 100: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_CONTROL_REGISTER_1928_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_CONTROL_REGISTER_1928_update_start_
      -- CP-element group 100: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_CONTROL_REGISTER_1928_Sample/$exit
      -- CP-element group 100: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_CONTROL_REGISTER_1928_Sample/ack
      -- CP-element group 100: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_CONTROL_REGISTER_1928_Update/req
      -- CP-element group 100: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_CONTROL_REGISTER_1928_sample_completed_
      -- 
    ack_3193_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 100_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_CONTROL_REGISTER_1928_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(100)); -- 
    req_3197_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3197_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(100), ack => WPIPE_CONTROL_REGISTER_1928_inst_req_1); -- 
    -- CP-element group 101:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	100 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	181 
    -- CP-element group 101: marked-successors 
    -- CP-element group 101: 	99 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_CONTROL_REGISTER_1928_Update/ack
      -- CP-element group 101: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_CONTROL_REGISTER_1928_update_completed_
      -- CP-element group 101: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_CONTROL_REGISTER_1928_Update/$exit
      -- 
    ack_3198_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_CONTROL_REGISTER_1928_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(101)); -- 
    -- CP-element group 102:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	20 
    -- CP-element group 102: 	39 
    -- CP-element group 102: marked-predecessors 
    -- CP-element group 102: 	104 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	104 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_1934_sample_start_
      -- CP-element group 102: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_1934_Sample/$entry
      -- CP-element group 102: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_1934_Sample/req
      -- 
    req_3206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(102), ack => W_update_control_register_pipe_1887_delayed_5_0_1932_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_102: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 31,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_102"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(20) & SoftwareRegisterAccessDaemon_CP_2867_elements(39) & SoftwareRegisterAccessDaemon_CP_2867_elements(104);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_102 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(102), clk => clk, reset => reset); --
    end block;
    -- CP-element group 103:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: marked-predecessors 
    -- CP-element group 103: 	115 
    -- CP-element group 103: 	110 
    -- CP-element group 103: 	112 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	105 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_1934_update_start_
      -- CP-element group 103: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_1934_Update/$entry
      -- CP-element group 103: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_1934_Update/req
      -- 
    req_3211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(103), ack => W_update_control_register_pipe_1887_delayed_5_0_1932_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_103: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_103"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(115) & SoftwareRegisterAccessDaemon_CP_2867_elements(110) & SoftwareRegisterAccessDaemon_CP_2867_elements(112);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_103 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(103), clk => clk, reset => reset); --
    end block;
    -- CP-element group 104:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	102 
    -- CP-element group 104: successors 
    -- CP-element group 104: marked-successors 
    -- CP-element group 104: 	18 
    -- CP-element group 104: 	102 
    -- CP-element group 104: 	35 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_1934_sample_completed_
      -- CP-element group 104: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_1934_Sample/$exit
      -- CP-element group 104: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_1934_Sample/ack
      -- 
    ack_3207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_update_control_register_pipe_1887_delayed_5_0_1932_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(104)); -- 
    -- CP-element group 105:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	103 
    -- CP-element group 105: successors 
    -- CP-element group 105: 	106 
    -- CP-element group 105: 	108 
    -- CP-element group 105: 	114 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_1934_update_completed_
      -- CP-element group 105: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_1934_Update/$exit
      -- CP-element group 105: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_1934_Update/ack
      -- 
    ack_3212_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_update_control_register_pipe_1887_delayed_5_0_1932_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(105)); -- 
    -- CP-element group 106:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	105 
    -- CP-element group 106: 	111 
    -- CP-element group 106: marked-predecessors 
    -- CP-element group 106: 	112 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	112 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/EQ_u32_u1_1941_sample_start_
      -- CP-element group 106: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/EQ_u32_u1_1941_Sample/$entry
      -- CP-element group 106: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/EQ_u32_u1_1941_Sample/rr
      -- 
    rr_3254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(106), ack => EQ_u32_u1_1941_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_106: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_106"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(105) & SoftwareRegisterAccessDaemon_CP_2867_elements(111) & SoftwareRegisterAccessDaemon_CP_2867_elements(112);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_106 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(106), clk => clk, reset => reset); --
    end block;
    -- CP-element group 107:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: marked-predecessors 
    -- CP-element group 107: 	115 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	113 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/EQ_u32_u1_1941_update_start_
      -- CP-element group 107: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/EQ_u32_u1_1941_Update/$entry
      -- CP-element group 107: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/EQ_u32_u1_1941_Update/cr
      -- 
    cr_3259_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3259_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(107), ack => EQ_u32_u1_1941_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2867_elements(115);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	11 
    -- CP-element group 108: 	105 
    -- CP-element group 108: marked-predecessors 
    -- CP-element group 108: 	166 
    -- CP-element group 108: 	110 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (5) 
      -- CP-element group 108: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1938_sample_start_
      -- CP-element group 108: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1938_Sample/$entry
      -- CP-element group 108: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1938_Sample/word_access_start/$entry
      -- CP-element group 108: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1938_Sample/word_access_start/word_0/$entry
      -- CP-element group 108: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1938_Sample/word_access_start/word_0/rr
      -- 
    rr_3233_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3233_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(108), ack => array_obj_ref_1938_load_0_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 1,3 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(11) & SoftwareRegisterAccessDaemon_CP_2867_elements(105) & SoftwareRegisterAccessDaemon_CP_2867_elements(166) & SoftwareRegisterAccessDaemon_CP_2867_elements(110);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: marked-predecessors 
    -- CP-element group 109: 	112 
    -- CP-element group 109: successors 
    -- CP-element group 109: 	111 
    -- CP-element group 109:  members (5) 
      -- CP-element group 109: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1938_update_start_
      -- CP-element group 109: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1938_Update/$entry
      -- CP-element group 109: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1938_Update/word_access_complete/$entry
      -- CP-element group 109: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1938_Update/word_access_complete/word_0/$entry
      -- CP-element group 109: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1938_Update/word_access_complete/word_0/cr
      -- 
    cr_3244_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3244_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(109), ack => array_obj_ref_1938_load_0_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_109: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_109"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2867_elements(112);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_109 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(109), clk => clk, reset => reset); --
    end block;
    -- CP-element group 110:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	177 
    -- CP-element group 110: marked-successors 
    -- CP-element group 110: 	103 
    -- CP-element group 110: 	108 
    -- CP-element group 110:  members (5) 
      -- CP-element group 110: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1938_sample_completed_
      -- CP-element group 110: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1938_Sample/$exit
      -- CP-element group 110: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1938_Sample/word_access_start/$exit
      -- CP-element group 110: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1938_Sample/word_access_start/word_0/$exit
      -- CP-element group 110: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1938_Sample/word_access_start/word_0/ra
      -- 
    ra_3234_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1938_load_0_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(110)); -- 
    -- CP-element group 111:  transition  input  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	109 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	106 
    -- CP-element group 111:  members (9) 
      -- CP-element group 111: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1938_update_completed_
      -- CP-element group 111: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1938_Update/$exit
      -- CP-element group 111: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1938_Update/word_access_complete/$exit
      -- CP-element group 111: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1938_Update/word_access_complete/word_0/$exit
      -- CP-element group 111: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1938_Update/word_access_complete/word_0/ca
      -- CP-element group 111: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1938_Update/array_obj_ref_1938_Merge/$entry
      -- CP-element group 111: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1938_Update/array_obj_ref_1938_Merge/$exit
      -- CP-element group 111: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1938_Update/array_obj_ref_1938_Merge/merge_req
      -- CP-element group 111: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1938_Update/array_obj_ref_1938_Merge/merge_ack
      -- 
    ca_3245_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 111_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1938_load_0_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(111)); -- 
    -- CP-element group 112:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	106 
    -- CP-element group 112: successors 
    -- CP-element group 112: marked-successors 
    -- CP-element group 112: 	103 
    -- CP-element group 112: 	106 
    -- CP-element group 112: 	109 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/EQ_u32_u1_1941_sample_completed_
      -- CP-element group 112: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/EQ_u32_u1_1941_Sample/$exit
      -- CP-element group 112: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/EQ_u32_u1_1941_Sample/ra
      -- 
    ra_3255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 112_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_1941_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(112)); -- 
    -- CP-element group 113:  transition  input  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	107 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/EQ_u32_u1_1941_update_completed_
      -- CP-element group 113: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/EQ_u32_u1_1941_Update/$exit
      -- CP-element group 113: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/EQ_u32_u1_1941_Update/ca
      -- 
    ca_3260_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u32_u1_1941_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(113)); -- 
    -- CP-element group 114:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	105 
    -- CP-element group 114: 	113 
    -- CP-element group 114: marked-predecessors 
    -- CP-element group 114: 	116 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_enable_mac_1936_sample_start_
      -- CP-element group 114: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_enable_mac_1936_Sample/$entry
      -- CP-element group 114: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_enable_mac_1936_Sample/req
      -- 
    req_3268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(114), ack => WPIPE_enable_mac_1936_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_114: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_114"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(105) & SoftwareRegisterAccessDaemon_CP_2867_elements(113) & SoftwareRegisterAccessDaemon_CP_2867_elements(116);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_114 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(114), clk => clk, reset => reset); --
    end block;
    -- CP-element group 115:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	116 
    -- CP-element group 115: marked-successors 
    -- CP-element group 115: 	103 
    -- CP-element group 115: 	107 
    -- CP-element group 115:  members (6) 
      -- CP-element group 115: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_enable_mac_1936_sample_completed_
      -- CP-element group 115: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_enable_mac_1936_update_start_
      -- CP-element group 115: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_enable_mac_1936_Sample/$exit
      -- CP-element group 115: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_enable_mac_1936_Sample/ack
      -- CP-element group 115: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_enable_mac_1936_Update/$entry
      -- CP-element group 115: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_enable_mac_1936_Update/req
      -- 
    ack_3269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_enable_mac_1936_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(115)); -- 
    req_3273_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3273_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(115), ack => WPIPE_enable_mac_1936_inst_req_1); -- 
    -- CP-element group 116:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	115 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	181 
    -- CP-element group 116: marked-successors 
    -- CP-element group 116: 	114 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_enable_mac_1936_update_completed_
      -- CP-element group 116: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_enable_mac_1936_Update/$exit
      -- CP-element group 116: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_enable_mac_1936_Update/ack
      -- 
    ack_3274_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 116_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_enable_mac_1936_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(116)); -- 
    -- CP-element group 117:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	11 
    -- CP-element group 117: 	20 
    -- CP-element group 117: 	58 
    -- CP-element group 117: marked-predecessors 
    -- CP-element group 117: 	119 
    -- CP-element group 117: 	166 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	119 
    -- CP-element group 117:  members (5) 
      -- CP-element group 117: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1946_sample_start_
      -- CP-element group 117: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1946_Sample/$entry
      -- CP-element group 117: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1946_Sample/word_access_start/$entry
      -- CP-element group 117: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1946_Sample/word_access_start/word_0/$entry
      -- CP-element group 117: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1946_Sample/word_access_start/word_0/rr
      -- 
    rr_3291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(117), ack => array_obj_ref_1946_load_0_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 31,1 => 31,2 => 31,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(11) & SoftwareRegisterAccessDaemon_CP_2867_elements(20) & SoftwareRegisterAccessDaemon_CP_2867_elements(58) & SoftwareRegisterAccessDaemon_CP_2867_elements(119) & SoftwareRegisterAccessDaemon_CP_2867_elements(166);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: marked-predecessors 
    -- CP-element group 118: 	127 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	120 
    -- CP-element group 118:  members (5) 
      -- CP-element group 118: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1946_update_start_
      -- CP-element group 118: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1946_Update/$entry
      -- CP-element group 118: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1946_Update/word_access_complete/$entry
      -- CP-element group 118: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1946_Update/word_access_complete/word_0/$entry
      -- CP-element group 118: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1946_Update/word_access_complete/word_0/cr
      -- 
    cr_3302_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3302_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(118), ack => array_obj_ref_1946_load_0_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_118: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_118"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2867_elements(127);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_118 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(118), clk => clk, reset => reset); --
    end block;
    -- CP-element group 119:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	117 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	178 
    -- CP-element group 119: marked-successors 
    -- CP-element group 119: 	18 
    -- CP-element group 119: 	117 
    -- CP-element group 119: 	54 
    -- CP-element group 119:  members (5) 
      -- CP-element group 119: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1946_sample_completed_
      -- CP-element group 119: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1946_Sample/$exit
      -- CP-element group 119: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1946_Sample/word_access_start/$exit
      -- CP-element group 119: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1946_Sample/word_access_start/word_0/$exit
      -- CP-element group 119: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1946_Sample/word_access_start/word_0/ra
      -- 
    ra_3292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1946_load_0_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(119)); -- 
    -- CP-element group 120:  transition  input  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	118 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	125 
    -- CP-element group 120:  members (9) 
      -- CP-element group 120: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1946_update_completed_
      -- CP-element group 120: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1946_Update/$exit
      -- CP-element group 120: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1946_Update/word_access_complete/$exit
      -- CP-element group 120: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1946_Update/word_access_complete/word_0/$exit
      -- CP-element group 120: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1946_Update/word_access_complete/word_0/ca
      -- CP-element group 120: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1946_Update/array_obj_ref_1946_Merge/$entry
      -- CP-element group 120: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1946_Update/array_obj_ref_1946_Merge/$exit
      -- CP-element group 120: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1946_Update/array_obj_ref_1946_Merge/merge_req
      -- CP-element group 120: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1946_Update/array_obj_ref_1946_Merge/merge_ack
      -- 
    ca_3303_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 120_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1946_load_0_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(120)); -- 
    -- CP-element group 121:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	20 
    -- CP-element group 121: 	58 
    -- CP-element group 121: marked-predecessors 
    -- CP-element group 121: 	123 
    -- CP-element group 121: successors 
    -- CP-element group 121: 	123 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_1950_sample_start_
      -- CP-element group 121: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_1950_Sample/$entry
      -- CP-element group 121: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_1950_Sample/req
      -- 
    req_3316_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3316_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(121), ack => W_update_free_q_pipe_1900_delayed_5_0_1948_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_121: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 31,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_121"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(20) & SoftwareRegisterAccessDaemon_CP_2867_elements(58) & SoftwareRegisterAccessDaemon_CP_2867_elements(123);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_121 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(121), clk => clk, reset => reset); --
    end block;
    -- CP-element group 122:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: marked-predecessors 
    -- CP-element group 122: 	127 
    -- CP-element group 122: 	130 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	124 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_1950_update_start_
      -- CP-element group 122: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_1950_Update/$entry
      -- CP-element group 122: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_1950_Update/req
      -- 
    req_3321_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3321_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(122), ack => W_update_free_q_pipe_1900_delayed_5_0_1948_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_122: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_122"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(127) & SoftwareRegisterAccessDaemon_CP_2867_elements(130);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_122 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(122), clk => clk, reset => reset); --
    end block;
    -- CP-element group 123:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	121 
    -- CP-element group 123: successors 
    -- CP-element group 123: marked-successors 
    -- CP-element group 123: 	18 
    -- CP-element group 123: 	121 
    -- CP-element group 123: 	54 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_1950_sample_completed_
      -- CP-element group 123: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_1950_Sample/$exit
      -- CP-element group 123: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_1950_Sample/ack
      -- 
    ack_3317_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 123_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_update_free_q_pipe_1900_delayed_5_0_1948_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(123)); -- 
    -- CP-element group 124:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: 	122 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	129 
    -- CP-element group 124: 	125 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_1950_update_completed_
      -- CP-element group 124: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_1950_Update/$exit
      -- CP-element group 124: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_1950_Update/ack
      -- 
    ack_3322_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 124_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_update_free_q_pipe_1900_delayed_5_0_1948_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(124)); -- 
    -- CP-element group 125:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	120 
    -- CP-element group 125: 	124 
    -- CP-element group 125: marked-predecessors 
    -- CP-element group 125: 	127 
    -- CP-element group 125: successors 
    -- CP-element group 125: 	127 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1954_sample_start_
      -- CP-element group 125: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1954_Sample/$entry
      -- CP-element group 125: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1954_Sample/rr
      -- 
    rr_3330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(125), ack => type_cast_1954_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_125: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_125"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(120) & SoftwareRegisterAccessDaemon_CP_2867_elements(124) & SoftwareRegisterAccessDaemon_CP_2867_elements(127);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_125 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(125), clk => clk, reset => reset); --
    end block;
    -- CP-element group 126:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: marked-predecessors 
    -- CP-element group 126: 	130 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	128 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1954_update_start_
      -- CP-element group 126: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1954_Update/$entry
      -- CP-element group 126: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1954_Update/cr
      -- 
    cr_3335_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3335_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(126), ack => type_cast_1954_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_126: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_126"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2867_elements(130);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_126 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(126), clk => clk, reset => reset); --
    end block;
    -- CP-element group 127:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	125 
    -- CP-element group 127: successors 
    -- CP-element group 127: marked-successors 
    -- CP-element group 127: 	118 
    -- CP-element group 127: 	122 
    -- CP-element group 127: 	125 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1954_sample_completed_
      -- CP-element group 127: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1954_Sample/$exit
      -- CP-element group 127: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1954_Sample/ra
      -- 
    ra_3331_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 127_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1954_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(127)); -- 
    -- CP-element group 128:  transition  input  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: 	126 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	129 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1954_update_completed_
      -- CP-element group 128: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1954_Update/$exit
      -- CP-element group 128: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/type_cast_1954_Update/ca
      -- 
    ca_3336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 128_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => type_cast_1954_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(128)); -- 
    -- CP-element group 129:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	128 
    -- CP-element group 129: 	124 
    -- CP-element group 129: marked-predecessors 
    -- CP-element group 129: 	131 
    -- CP-element group 129: successors 
    -- CP-element group 129: 	130 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_FREE_Q_1952_sample_start_
      -- CP-element group 129: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_FREE_Q_1952_Sample/$entry
      -- CP-element group 129: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_FREE_Q_1952_Sample/req
      -- 
    req_3344_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3344_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(129), ack => WPIPE_FREE_Q_1952_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_129: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_129"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(128) & SoftwareRegisterAccessDaemon_CP_2867_elements(124) & SoftwareRegisterAccessDaemon_CP_2867_elements(131);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_129 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(129), clk => clk, reset => reset); --
    end block;
    -- CP-element group 130:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	129 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130: marked-successors 
    -- CP-element group 130: 	122 
    -- CP-element group 130: 	126 
    -- CP-element group 130:  members (6) 
      -- CP-element group 130: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_FREE_Q_1952_sample_completed_
      -- CP-element group 130: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_FREE_Q_1952_update_start_
      -- CP-element group 130: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_FREE_Q_1952_Sample/$exit
      -- CP-element group 130: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_FREE_Q_1952_Sample/ack
      -- CP-element group 130: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_FREE_Q_1952_Update/$entry
      -- CP-element group 130: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_FREE_Q_1952_Update/req
      -- 
    ack_3345_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_FREE_Q_1952_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(130)); -- 
    req_3349_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3349_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(130), ack => WPIPE_FREE_Q_1952_inst_req_1); -- 
    -- CP-element group 131:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	130 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	181 
    -- CP-element group 131: marked-successors 
    -- CP-element group 131: 	129 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_FREE_Q_1952_update_completed_
      -- CP-element group 131: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_FREE_Q_1952_Update/$exit
      -- CP-element group 131: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_FREE_Q_1952_Update/ack
      -- 
    ack_3350_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 131_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_FREE_Q_1952_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(131)); -- 
    -- CP-element group 132:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: 	11 
    -- CP-element group 132: 	20 
    -- CP-element group 132: 	77 
    -- CP-element group 132: marked-predecessors 
    -- CP-element group 132: 	166 
    -- CP-element group 132: 	134 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (5) 
      -- CP-element group 132: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1959_sample_start_
      -- CP-element group 132: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1959_Sample/$entry
      -- CP-element group 132: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1959_Sample/word_access_start/$entry
      -- CP-element group 132: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1959_Sample/word_access_start/word_0/$entry
      -- CP-element group 132: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1959_Sample/word_access_start/word_0/rr
      -- 
    rr_3367_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3367_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(132), ack => array_obj_ref_1959_load_0_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 31,1 => 31,2 => 31,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 1,4 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(11) & SoftwareRegisterAccessDaemon_CP_2867_elements(20) & SoftwareRegisterAccessDaemon_CP_2867_elements(77) & SoftwareRegisterAccessDaemon_CP_2867_elements(166) & SoftwareRegisterAccessDaemon_CP_2867_elements(134);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: marked-predecessors 
    -- CP-element group 133: 	137 
    -- CP-element group 133: successors 
    -- CP-element group 133: 	135 
    -- CP-element group 133:  members (5) 
      -- CP-element group 133: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1959_update_start_
      -- CP-element group 133: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1959_Update/$entry
      -- CP-element group 133: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1959_Update/word_access_complete/$entry
      -- CP-element group 133: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1959_Update/word_access_complete/word_0/$entry
      -- CP-element group 133: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1959_Update/word_access_complete/word_0/cr
      -- 
    cr_3378_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3378_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(133), ack => array_obj_ref_1959_load_0_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_133: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_133"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2867_elements(137);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_133 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(133), clk => clk, reset => reset); --
    end block;
    -- CP-element group 134:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	179 
    -- CP-element group 134: marked-successors 
    -- CP-element group 134: 	18 
    -- CP-element group 134: 	132 
    -- CP-element group 134: 	73 
    -- CP-element group 134:  members (5) 
      -- CP-element group 134: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1959_sample_completed_
      -- CP-element group 134: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1959_Sample/$exit
      -- CP-element group 134: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1959_Sample/word_access_start/$exit
      -- CP-element group 134: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1959_Sample/word_access_start/word_0/$exit
      -- CP-element group 134: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1959_Sample/word_access_start/word_0/ra
      -- 
    ra_3368_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1959_load_0_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(134)); -- 
    -- CP-element group 135:  transition  input  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	133 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	136 
    -- CP-element group 135:  members (9) 
      -- CP-element group 135: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1959_update_completed_
      -- CP-element group 135: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1959_Update/$exit
      -- CP-element group 135: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1959_Update/word_access_complete/$exit
      -- CP-element group 135: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1959_Update/word_access_complete/word_0/$exit
      -- CP-element group 135: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1959_Update/word_access_complete/word_0/ca
      -- CP-element group 135: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1959_Update/array_obj_ref_1959_Merge/$entry
      -- CP-element group 135: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1959_Update/array_obj_ref_1959_Merge/$exit
      -- CP-element group 135: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1959_Update/array_obj_ref_1959_Merge/merge_req
      -- CP-element group 135: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1959_Update/array_obj_ref_1959_Merge/merge_ack
      -- 
    ca_3379_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 135_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_1959_load_0_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(135)); -- 
    -- CP-element group 136:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: 	20 
    -- CP-element group 136: 	135 
    -- CP-element group 136: 	77 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	138 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	137 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_NUMBER_OF_SERVERS_1957_sample_start_
      -- CP-element group 136: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_NUMBER_OF_SERVERS_1957_Sample/$entry
      -- CP-element group 136: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_NUMBER_OF_SERVERS_1957_Sample/req
      -- 
    req_3392_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3392_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(136), ack => WPIPE_NUMBER_OF_SERVERS_1957_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 1,2 => 31,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(20) & SoftwareRegisterAccessDaemon_CP_2867_elements(135) & SoftwareRegisterAccessDaemon_CP_2867_elements(77) & SoftwareRegisterAccessDaemon_CP_2867_elements(138);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	136 
    -- CP-element group 137: successors 
    -- CP-element group 137: 	138 
    -- CP-element group 137: marked-successors 
    -- CP-element group 137: 	18 
    -- CP-element group 137: 	133 
    -- CP-element group 137: 	73 
    -- CP-element group 137:  members (6) 
      -- CP-element group 137: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_NUMBER_OF_SERVERS_1957_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_NUMBER_OF_SERVERS_1957_update_start_
      -- CP-element group 137: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_NUMBER_OF_SERVERS_1957_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_NUMBER_OF_SERVERS_1957_Sample/ack
      -- CP-element group 137: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_NUMBER_OF_SERVERS_1957_Update/$entry
      -- CP-element group 137: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_NUMBER_OF_SERVERS_1957_Update/req
      -- 
    ack_3393_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NUMBER_OF_SERVERS_1957_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(137)); -- 
    req_3397_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3397_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(137), ack => WPIPE_NUMBER_OF_SERVERS_1957_inst_req_1); -- 
    -- CP-element group 138:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	137 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	181 
    -- CP-element group 138: marked-successors 
    -- CP-element group 138: 	136 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_NUMBER_OF_SERVERS_1957_update_completed_
      -- CP-element group 138: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_NUMBER_OF_SERVERS_1957_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_NUMBER_OF_SERVERS_1957_Update/ack
      -- 
    ack_3398_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NUMBER_OF_SERVERS_1957_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(138)); -- 
    -- CP-element group 139:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	11 
    -- CP-element group 139: marked-predecessors 
    -- CP-element group 139: 	142 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	141 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/RPIPE_AFB_NIC_REQUEST_1962_sample_start_
      -- CP-element group 139: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/RPIPE_AFB_NIC_REQUEST_1962_Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/RPIPE_AFB_NIC_REQUEST_1962_Sample/rr
      -- 
    rr_3406_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3406_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(139), ack => RPIPE_AFB_NIC_REQUEST_1962_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_139: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_139"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(11) & SoftwareRegisterAccessDaemon_CP_2867_elements(142);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_139 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(139), clk => clk, reset => reset); --
    end block;
    -- CP-element group 140:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: 	14 
    -- CP-element group 140: 	141 
    -- CP-element group 140: marked-predecessors 
    -- CP-element group 140: 	145 
    -- CP-element group 140: 	149 
    -- CP-element group 140: 	153 
    -- CP-element group 140: 	157 
    -- CP-element group 140: 	161 
    -- CP-element group 140: 	169 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	142 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/RPIPE_AFB_NIC_REQUEST_1962_update_start_
      -- CP-element group 140: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/RPIPE_AFB_NIC_REQUEST_1962_Update/$entry
      -- CP-element group 140: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/RPIPE_AFB_NIC_REQUEST_1962_Update/cr
      -- 
    cr_3411_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3411_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(140), ack => RPIPE_AFB_NIC_REQUEST_1962_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_140: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 31,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_140"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(14) & SoftwareRegisterAccessDaemon_CP_2867_elements(141) & SoftwareRegisterAccessDaemon_CP_2867_elements(145) & SoftwareRegisterAccessDaemon_CP_2867_elements(149) & SoftwareRegisterAccessDaemon_CP_2867_elements(153) & SoftwareRegisterAccessDaemon_CP_2867_elements(157) & SoftwareRegisterAccessDaemon_CP_2867_elements(161) & SoftwareRegisterAccessDaemon_CP_2867_elements(169);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_140 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(140), clk => clk, reset => reset); --
    end block;
    -- CP-element group 141:  transition  input  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	139 
    -- CP-element group 141: successors 
    -- CP-element group 141: 	140 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/RPIPE_AFB_NIC_REQUEST_1962_sample_completed_
      -- CP-element group 141: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/RPIPE_AFB_NIC_REQUEST_1962_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/RPIPE_AFB_NIC_REQUEST_1962_Sample/ra
      -- 
    ra_3407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_AFB_NIC_REQUEST_1962_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(141)); -- 
    -- CP-element group 142:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	140 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	147 
    -- CP-element group 142: 	151 
    -- CP-element group 142: 	155 
    -- CP-element group 142: 	159 
    -- CP-element group 142: 	167 
    -- CP-element group 142: 	143 
    -- CP-element group 142: marked-successors 
    -- CP-element group 142: 	139 
    -- CP-element group 142: 	34 
    -- CP-element group 142: 	53 
    -- CP-element group 142: 	72 
    -- CP-element group 142:  members (29) 
      -- CP-element group 142: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/RPIPE_AFB_NIC_REQUEST_1962_update_completed_
      -- CP-element group 142: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/RPIPE_AFB_NIC_REQUEST_1962_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/RPIPE_AFB_NIC_REQUEST_1962_Update/ca
      -- CP-element group 142: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_word_address_calculated
      -- CP-element group 142: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_root_address_calculated
      -- CP-element group 142: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_offset_calculated
      -- CP-element group 142: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_index_resized_0
      -- CP-element group 142: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_index_scaled_0
      -- CP-element group 142: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_index_computed_0
      -- CP-element group 142: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_index_resize_0/$entry
      -- CP-element group 142: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_index_resize_0/$exit
      -- CP-element group 142: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_index_resize_0/index_resize_req
      -- CP-element group 142: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_index_resize_0/index_resize_ack
      -- CP-element group 142: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_index_scale_0/$entry
      -- CP-element group 142: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_index_scale_0/$exit
      -- CP-element group 142: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_index_scale_0/scale_rename_req
      -- CP-element group 142: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_index_scale_0/scale_rename_ack
      -- CP-element group 142: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_final_index_sum_regn/$entry
      -- CP-element group 142: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_final_index_sum_regn/$exit
      -- CP-element group 142: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_final_index_sum_regn/req
      -- CP-element group 142: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_final_index_sum_regn/ack
      -- CP-element group 142: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_base_plus_offset/$entry
      -- CP-element group 142: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_base_plus_offset/$exit
      -- CP-element group 142: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_base_plus_offset/sum_rename_req
      -- CP-element group 142: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_base_plus_offset/sum_rename_ack
      -- CP-element group 142: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_word_addrgen/$entry
      -- CP-element group 142: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_word_addrgen/$exit
      -- CP-element group 142: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_word_addrgen/root_register_req
      -- CP-element group 142: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_word_addrgen/root_register_ack
      -- 
    ca_3412_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_AFB_NIC_REQUEST_1962_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(142)); -- 
    -- CP-element group 143:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	142 
    -- CP-element group 143: marked-predecessors 
    -- CP-element group 143: 	145 
    -- CP-element group 143: 	166 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	145 
    -- CP-element group 143:  members (5) 
      -- CP-element group 143: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_Sample/word_access_start/$entry
      -- CP-element group 143: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_Sample/word_access_start/word_0/$entry
      -- CP-element group 143: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_Sample/word_access_start/word_0/rr
      -- 
    rr_3458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(143), ack => array_obj_ref_2015_load_0_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_143: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_143"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(142) & SoftwareRegisterAccessDaemon_CP_2867_elements(145) & SoftwareRegisterAccessDaemon_CP_2867_elements(166);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_143 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(143), clk => clk, reset => reset); --
    end block;
    -- CP-element group 144:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: marked-predecessors 
    -- CP-element group 144: 	165 
    -- CP-element group 144: 	172 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	146 
    -- CP-element group 144:  members (5) 
      -- CP-element group 144: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_update_start_
      -- CP-element group 144: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_Update/$entry
      -- CP-element group 144: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_Update/word_access_complete/$entry
      -- CP-element group 144: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_Update/word_access_complete/word_0/$entry
      -- CP-element group 144: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_Update/word_access_complete/word_0/cr
      -- 
    cr_3469_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3469_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(144), ack => array_obj_ref_2015_load_0_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_144: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_144"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(165) & SoftwareRegisterAccessDaemon_CP_2867_elements(172);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_144 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(144), clk => clk, reset => reset); --
    end block;
    -- CP-element group 145:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	143 
    -- CP-element group 145: successors 
    -- CP-element group 145: 	180 
    -- CP-element group 145: marked-successors 
    -- CP-element group 145: 	140 
    -- CP-element group 145: 	143 
    -- CP-element group 145:  members (5) 
      -- CP-element group 145: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_sample_completed_
      -- CP-element group 145: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_Sample/word_access_start/$exit
      -- CP-element group 145: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_Sample/word_access_start/word_0/$exit
      -- CP-element group 145: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_Sample/word_access_start/word_0/ra
      -- 
    ra_3459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2015_load_0_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(145)); -- 
    -- CP-element group 146:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	144 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	163 
    -- CP-element group 146: 	171 
    -- CP-element group 146:  members (9) 
      -- CP-element group 146: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_update_completed_
      -- CP-element group 146: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_Update/word_access_complete/$exit
      -- CP-element group 146: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_Update/word_access_complete/word_0/$exit
      -- CP-element group 146: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_Update/word_access_complete/word_0/ca
      -- CP-element group 146: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_Update/array_obj_ref_2015_Merge/$entry
      -- CP-element group 146: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_Update/array_obj_ref_2015_Merge/$exit
      -- CP-element group 146: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_Update/array_obj_ref_2015_Merge/merge_req
      -- CP-element group 146: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_Update/array_obj_ref_2015_Merge/merge_ack
      -- 
    ca_3470_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_2015_load_0_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(146)); -- 
    -- CP-element group 147:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	142 
    -- CP-element group 147: marked-predecessors 
    -- CP-element group 147: 	149 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2019_sample_start_
      -- CP-element group 147: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2019_Sample/$entry
      -- CP-element group 147: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2019_Sample/req
      -- 
    req_3483_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3483_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(147), ack => W_rwbar_1966_delayed_5_0_2017_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_147: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_147"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(142) & SoftwareRegisterAccessDaemon_CP_2867_elements(149);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_147 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(147), clk => clk, reset => reset); --
    end block;
    -- CP-element group 148:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: marked-predecessors 
    -- CP-element group 148: 	165 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	150 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2019_update_start_
      -- CP-element group 148: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2019_Update/$entry
      -- CP-element group 148: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2019_Update/req
      -- 
    req_3488_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3488_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(148), ack => W_rwbar_1966_delayed_5_0_2017_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_148: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_148"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2867_elements(165);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_148 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(148), clk => clk, reset => reset); --
    end block;
    -- CP-element group 149:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: marked-successors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: 	140 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2019_sample_completed_
      -- CP-element group 149: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2019_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2019_Sample/ack
      -- 
    ack_3484_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_1966_delayed_5_0_2017_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(149)); -- 
    -- CP-element group 150:  transition  input  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	148 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	163 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2019_update_completed_
      -- CP-element group 150: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2019_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2019_Update/ack
      -- 
    ack_3489_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_1966_delayed_5_0_2017_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(150)); -- 
    -- CP-element group 151:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	142 
    -- CP-element group 151: marked-predecessors 
    -- CP-element group 151: 	153 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2022_sample_start_
      -- CP-element group 151: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2022_Sample/$entry
      -- CP-element group 151: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2022_Sample/req
      -- 
    req_3497_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3497_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(151), ack => W_bmask_1967_delayed_5_0_2020_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(142) & SoftwareRegisterAccessDaemon_CP_2867_elements(153);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_151 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: marked-predecessors 
    -- CP-element group 152: 	165 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	154 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2022_update_start_
      -- CP-element group 152: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2022_Update/$entry
      -- CP-element group 152: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2022_Update/req
      -- 
    req_3502_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3502_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(152), ack => W_bmask_1967_delayed_5_0_2020_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_152: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_152"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2867_elements(165);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_152 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(152), clk => clk, reset => reset); --
    end block;
    -- CP-element group 153:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153: marked-successors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: 	140 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2022_sample_completed_
      -- CP-element group 153: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2022_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2022_Sample/ack
      -- 
    ack_3498_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bmask_1967_delayed_5_0_2020_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(153)); -- 
    -- CP-element group 154:  transition  input  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	152 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	163 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2022_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2022_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2022_Update/ack
      -- 
    ack_3503_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bmask_1967_delayed_5_0_2020_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(154)); -- 
    -- CP-element group 155:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	142 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	157 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2025_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2025_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2025_Sample/req
      -- 
    req_3511_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3511_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(155), ack => W_wdata_1969_delayed_5_0_2023_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(142) & SoftwareRegisterAccessDaemon_CP_2867_elements(157);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: marked-predecessors 
    -- CP-element group 156: 	165 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2025_update_start_
      -- CP-element group 156: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2025_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2025_Update/req
      -- 
    req_3516_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3516_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(156), ack => W_wdata_1969_delayed_5_0_2023_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2867_elements(165);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157: marked-successors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: 	140 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2025_sample_completed_
      -- CP-element group 157: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2025_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2025_Sample/ack
      -- 
    ack_3512_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_wdata_1969_delayed_5_0_2023_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(157)); -- 
    -- CP-element group 158:  transition  input  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	163 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2025_update_completed_
      -- CP-element group 158: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2025_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2025_Update/ack
      -- 
    ack_3517_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_wdata_1969_delayed_5_0_2023_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(158)); -- 
    -- CP-element group 159:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	142 
    -- CP-element group 159: marked-predecessors 
    -- CP-element group 159: 	161 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	161 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2028_sample_start_
      -- CP-element group 159: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2028_Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2028_Sample/req
      -- 
    req_3525_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3525_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(159), ack => W_index_1970_delayed_5_0_2026_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_159: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_159"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(142) & SoftwareRegisterAccessDaemon_CP_2867_elements(161);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_159 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(159), clk => clk, reset => reset); --
    end block;
    -- CP-element group 160:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: marked-predecessors 
    -- CP-element group 160: 	165 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	162 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2028_update_start_
      -- CP-element group 160: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2028_Update/$entry
      -- CP-element group 160: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2028_Update/req
      -- 
    req_3530_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3530_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(160), ack => W_index_1970_delayed_5_0_2026_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2867_elements(165);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: successors 
    -- CP-element group 161: marked-successors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: 	140 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2028_sample_completed_
      -- CP-element group 161: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2028_Sample/$exit
      -- CP-element group 161: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2028_Sample/ack
      -- 
    ack_3526_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_index_1970_delayed_5_0_2026_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(161)); -- 
    -- CP-element group 162:  transition  input  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	160 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	163 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2028_update_completed_
      -- CP-element group 162: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2028_Update/$exit
      -- CP-element group 162: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2028_Update/ack
      -- 
    ack_3531_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_index_1970_delayed_5_0_2026_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(162)); -- 
    -- CP-element group 163:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	146 
    -- CP-element group 163: 	150 
    -- CP-element group 163: 	154 
    -- CP-element group 163: 	158 
    -- CP-element group 163: 	162 
    -- CP-element group 163: 	175 
    -- CP-element group 163: 	176 
    -- CP-element group 163: 	177 
    -- CP-element group 163: 	178 
    -- CP-element group 163: 	179 
    -- CP-element group 163: 	180 
    -- CP-element group 163: marked-predecessors 
    -- CP-element group 163: 	165 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	165 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/call_stmt_2035_sample_start_
      -- CP-element group 163: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/call_stmt_2035_Sample/$entry
      -- CP-element group 163: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/call_stmt_2035_Sample/crr
      -- 
    crr_3539_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3539_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(163), ack => call_stmt_2035_call_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 31,6 => 31,7 => 31,8 => 31,9 => 31,10 => 31,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 1);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(146) & SoftwareRegisterAccessDaemon_CP_2867_elements(150) & SoftwareRegisterAccessDaemon_CP_2867_elements(154) & SoftwareRegisterAccessDaemon_CP_2867_elements(158) & SoftwareRegisterAccessDaemon_CP_2867_elements(162) & SoftwareRegisterAccessDaemon_CP_2867_elements(175) & SoftwareRegisterAccessDaemon_CP_2867_elements(176) & SoftwareRegisterAccessDaemon_CP_2867_elements(177) & SoftwareRegisterAccessDaemon_CP_2867_elements(178) & SoftwareRegisterAccessDaemon_CP_2867_elements(179) & SoftwareRegisterAccessDaemon_CP_2867_elements(180) & SoftwareRegisterAccessDaemon_CP_2867_elements(165);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: marked-predecessors 
    -- CP-element group 164: 	166 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/call_stmt_2035_update_start_
      -- CP-element group 164: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/call_stmt_2035_Update/$entry
      -- CP-element group 164: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/call_stmt_2035_Update/ccr
      -- 
    ccr_3544_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3544_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(164), ack => call_stmt_2035_call_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2867_elements(166);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: successors 
    -- CP-element group 165: marked-successors 
    -- CP-element group 165: 	148 
    -- CP-element group 165: 	152 
    -- CP-element group 165: 	156 
    -- CP-element group 165: 	160 
    -- CP-element group 165: 	163 
    -- CP-element group 165: 	144 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/call_stmt_2035_sample_completed_
      -- CP-element group 165: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/call_stmt_2035_Sample/$exit
      -- CP-element group 165: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/call_stmt_2035_Sample/cra
      -- 
    cra_3540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2035_call_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(165)); -- 
    -- CP-element group 166:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	181 
    -- CP-element group 166: marked-successors 
    -- CP-element group 166: 	95 
    -- CP-element group 166: 	117 
    -- CP-element group 166: 	164 
    -- CP-element group 166: 	132 
    -- CP-element group 166: 	143 
    -- CP-element group 166: 	91 
    -- CP-element group 166: 	108 
    -- CP-element group 166:  members (4) 
      -- CP-element group 166: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/call_stmt_2035_update_completed_
      -- CP-element group 166: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/call_stmt_2035_Update/$exit
      -- CP-element group 166: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/call_stmt_2035_Update/cca
      -- CP-element group 166: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/ring_reenable_memory_space_2
      -- 
    cca_3545_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_2035_call_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(166)); -- 
    -- CP-element group 167:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	142 
    -- CP-element group 167: marked-predecessors 
    -- CP-element group 167: 	169 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	169 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2038_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2038_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2038_Sample/req
      -- 
    req_3553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(167), ack => W_rwbar_1974_delayed_5_0_2036_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_167: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_167"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(142) & SoftwareRegisterAccessDaemon_CP_2867_elements(169);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_167 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(167), clk => clk, reset => reset); --
    end block;
    -- CP-element group 168:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: marked-predecessors 
    -- CP-element group 168: 	172 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	170 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2038_update_start_
      -- CP-element group 168: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2038_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2038_Update/req
      -- 
    req_3558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(168), ack => W_rwbar_1974_delayed_5_0_2036_inst_req_1); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_168: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_168"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= SoftwareRegisterAccessDaemon_CP_2867_elements(172);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_168 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(168), clk => clk, reset => reset); --
    end block;
    -- CP-element group 169:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: successors 
    -- CP-element group 169: marked-successors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: 	140 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2038_sample_completed_
      -- CP-element group 169: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2038_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2038_Sample/ack
      -- 
    ack_3554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_1974_delayed_5_0_2036_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(169)); -- 
    -- CP-element group 170:  transition  input  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	168 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	171 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2038_update_completed_
      -- CP-element group 170: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2038_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/assign_stmt_2038_Update/ack
      -- 
    ack_3559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_1974_delayed_5_0_2036_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(170)); -- 
    -- CP-element group 171:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	146 
    -- CP-element group 171: 	170 
    -- CP-element group 171: marked-predecessors 
    -- CP-element group 171: 	173 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	172 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_AFB_NIC_RESPONSE_2052_sample_start_
      -- CP-element group 171: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_AFB_NIC_RESPONSE_2052_Sample/$entry
      -- CP-element group 171: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_AFB_NIC_RESPONSE_2052_Sample/req
      -- 
    req_3567_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3567_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(171), ack => WPIPE_AFB_NIC_RESPONSE_2052_inst_req_0); -- 
    SoftwareRegisterAccessDaemon_cp_element_group_171: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_171"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(146) & SoftwareRegisterAccessDaemon_CP_2867_elements(170) & SoftwareRegisterAccessDaemon_CP_2867_elements(173);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_171 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(171), clk => clk, reset => reset); --
    end block;
    -- CP-element group 172:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: 	171 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	173 
    -- CP-element group 172: marked-successors 
    -- CP-element group 172: 	168 
    -- CP-element group 172: 	144 
    -- CP-element group 172:  members (6) 
      -- CP-element group 172: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_AFB_NIC_RESPONSE_2052_sample_completed_
      -- CP-element group 172: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_AFB_NIC_RESPONSE_2052_update_start_
      -- CP-element group 172: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_AFB_NIC_RESPONSE_2052_Sample/$exit
      -- CP-element group 172: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_AFB_NIC_RESPONSE_2052_Sample/ack
      -- CP-element group 172: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_AFB_NIC_RESPONSE_2052_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_AFB_NIC_RESPONSE_2052_Update/req
      -- 
    ack_3568_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 172_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_AFB_NIC_RESPONSE_2052_inst_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(172)); -- 
    req_3572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(172), ack => WPIPE_AFB_NIC_RESPONSE_2052_inst_req_1); -- 
    -- CP-element group 173:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	172 
    -- CP-element group 173: successors 
    -- CP-element group 173: 	181 
    -- CP-element group 173: marked-successors 
    -- CP-element group 173: 	171 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_AFB_NIC_RESPONSE_2052_update_completed_
      -- CP-element group 173: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_AFB_NIC_RESPONSE_2052_Update/$exit
      -- CP-element group 173: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/WPIPE_AFB_NIC_RESPONSE_2052_Update/ack
      -- 
    ack_3573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_AFB_NIC_RESPONSE_2052_inst_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(173)); -- 
    -- CP-element group 174:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	11 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	12 
    -- CP-element group 174:  members (1) 
      -- CP-element group 174: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(174) is a control-delay.
    cp_element_174_delay: control_delay_element  generic map(name => " 174_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2867_elements(11), ack => SoftwareRegisterAccessDaemon_CP_2867_elements(174), clk => clk, reset =>reset);
    -- CP-element group 175:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	93 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	163 
    -- CP-element group 175:  members (1) 
      -- CP-element group 175: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1899_call_stmt_2035_delay
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(175) is a control-delay.
    cp_element_175_delay: control_delay_element  generic map(name => " 175_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2867_elements(93), ack => SoftwareRegisterAccessDaemon_CP_2867_elements(175), clk => clk, reset =>reset);
    -- CP-element group 176:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: 	97 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	163 
    -- CP-element group 176:  members (1) 
      -- CP-element group 176: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1930_call_stmt_2035_delay
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(176) is a control-delay.
    cp_element_176_delay: control_delay_element  generic map(name => " 176_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2867_elements(97), ack => SoftwareRegisterAccessDaemon_CP_2867_elements(176), clk => clk, reset =>reset);
    -- CP-element group 177:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	110 
    -- CP-element group 177: successors 
    -- CP-element group 177: 	163 
    -- CP-element group 177:  members (1) 
      -- CP-element group 177: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1938_call_stmt_2035_delay
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(177) is a control-delay.
    cp_element_177_delay: control_delay_element  generic map(name => " 177_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2867_elements(110), ack => SoftwareRegisterAccessDaemon_CP_2867_elements(177), clk => clk, reset =>reset);
    -- CP-element group 178:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	119 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	163 
    -- CP-element group 178:  members (1) 
      -- CP-element group 178: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1946_call_stmt_2035_delay
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(178) is a control-delay.
    cp_element_178_delay: control_delay_element  generic map(name => " 178_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2867_elements(119), ack => SoftwareRegisterAccessDaemon_CP_2867_elements(178), clk => clk, reset =>reset);
    -- CP-element group 179:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	134 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	163 
    -- CP-element group 179:  members (1) 
      -- CP-element group 179: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_1959_call_stmt_2035_delay
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(179) is a control-delay.
    cp_element_179_delay: control_delay_element  generic map(name => " 179_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2867_elements(134), ack => SoftwareRegisterAccessDaemon_CP_2867_elements(179), clk => clk, reset =>reset);
    -- CP-element group 180:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: 	145 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	163 
    -- CP-element group 180:  members (1) 
      -- CP-element group 180: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/array_obj_ref_2015_call_stmt_2035_delay
      -- 
    -- Element group SoftwareRegisterAccessDaemon_CP_2867_elements(180) is a control-delay.
    cp_element_180_delay: control_delay_element  generic map(name => " 180_delay", delay_value => 1)  port map(req => SoftwareRegisterAccessDaemon_CP_2867_elements(145), ack => SoftwareRegisterAccessDaemon_CP_2867_elements(180), clk => clk, reset =>reset);
    -- CP-element group 181:  join  transition  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	14 
    -- CP-element group 181: 	94 
    -- CP-element group 181: 	116 
    -- CP-element group 181: 	166 
    -- CP-element group 181: 	131 
    -- CP-element group 181: 	173 
    -- CP-element group 181: 	138 
    -- CP-element group 181: 	101 
    -- CP-element group 181: successors 
    -- CP-element group 181: 	8 
    -- CP-element group 181:  members (1) 
      -- CP-element group 181: 	 branch_block_stmt_1862/do_while_stmt_1872/do_while_stmt_1872_loop_body/$exit
      -- 
    SoftwareRegisterAccessDaemon_cp_element_group_181: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 31,1 => 31,2 => 31,3 => 31,4 => 31,5 => 31,6 => 31,7 => 31);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 49) := "SoftwareRegisterAccessDaemon_cp_element_group_181"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= SoftwareRegisterAccessDaemon_CP_2867_elements(14) & SoftwareRegisterAccessDaemon_CP_2867_elements(94) & SoftwareRegisterAccessDaemon_CP_2867_elements(116) & SoftwareRegisterAccessDaemon_CP_2867_elements(166) & SoftwareRegisterAccessDaemon_CP_2867_elements(131) & SoftwareRegisterAccessDaemon_CP_2867_elements(173) & SoftwareRegisterAccessDaemon_CP_2867_elements(138) & SoftwareRegisterAccessDaemon_CP_2867_elements(101);
      gj_SoftwareRegisterAccessDaemon_cp_element_group_181 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(181), clk => clk, reset => reset); --
    end block;
    -- CP-element group 182:  transition  input  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	7 
    -- CP-element group 182: successors 
    -- CP-element group 182:  members (2) 
      -- CP-element group 182: 	 branch_block_stmt_1862/do_while_stmt_1872/loop_exit/$exit
      -- CP-element group 182: 	 branch_block_stmt_1862/do_while_stmt_1872/loop_exit/ack
      -- 
    ack_3585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1872_branch_ack_0, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(182)); -- 
    -- CP-element group 183:  transition  input  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	7 
    -- CP-element group 183: successors 
    -- CP-element group 183:  members (2) 
      -- CP-element group 183: 	 branch_block_stmt_1862/do_while_stmt_1872/loop_taken/$exit
      -- CP-element group 183: 	 branch_block_stmt_1862/do_while_stmt_1872/loop_taken/ack
      -- 
    ack_3589_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 183_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1872_branch_ack_1, ack => SoftwareRegisterAccessDaemon_CP_2867_elements(183)); -- 
    -- CP-element group 184:  transition  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: 	5 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	1 
    -- CP-element group 184:  members (1) 
      -- CP-element group 184: 	 branch_block_stmt_1862/do_while_stmt_1872/$exit
      -- 
    SoftwareRegisterAccessDaemon_CP_2867_elements(184) <= SoftwareRegisterAccessDaemon_CP_2867_elements(5);
    -- CP-element group 185:  merge  branch  transition  place  output  bypass 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	2 
    -- CP-element group 185: 	0 
    -- CP-element group 185: successors 
    -- CP-element group 185: 	2 
    -- CP-element group 185: 	3 
    -- CP-element group 185:  members (37) 
      -- CP-element group 185: 	 branch_block_stmt_1862/merge_stmt_1863__exit__
      -- CP-element group 185: 	 branch_block_stmt_1862/if_stmt_1866__entry__
      -- CP-element group 185: 	 branch_block_stmt_1862/if_stmt_1866_dead_link/$entry
      -- CP-element group 185: 	 branch_block_stmt_1862/if_stmt_1866_eval_test/$entry
      -- CP-element group 185: 	 branch_block_stmt_1862/if_stmt_1866_eval_test/$exit
      -- CP-element group 185: 	 branch_block_stmt_1862/if_stmt_1866_eval_test/EQ_u1_u1_1869/$entry
      -- CP-element group 185: 	 branch_block_stmt_1862/if_stmt_1866_eval_test/EQ_u1_u1_1869/$exit
      -- CP-element group 185: 	 branch_block_stmt_1862/if_stmt_1866_eval_test/EQ_u1_u1_1869/EQ_u1_u1_1869_inputs/$entry
      -- CP-element group 185: 	 branch_block_stmt_1862/if_stmt_1866_eval_test/EQ_u1_u1_1869/EQ_u1_u1_1869_inputs/$exit
      -- CP-element group 185: 	 branch_block_stmt_1862/if_stmt_1866_eval_test/EQ_u1_u1_1869/EQ_u1_u1_1869_inputs/RPIPE_MAC_ENABLE_1867/$entry
      -- CP-element group 185: 	 branch_block_stmt_1862/if_stmt_1866_eval_test/EQ_u1_u1_1869/EQ_u1_u1_1869_inputs/RPIPE_MAC_ENABLE_1867/$exit
      -- CP-element group 185: 	 branch_block_stmt_1862/if_stmt_1866_eval_test/EQ_u1_u1_1869/EQ_u1_u1_1869_inputs/RPIPE_MAC_ENABLE_1867/Sample/$entry
      -- CP-element group 185: 	 branch_block_stmt_1862/if_stmt_1866_eval_test/EQ_u1_u1_1869/EQ_u1_u1_1869_inputs/RPIPE_MAC_ENABLE_1867/Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_1862/if_stmt_1866_eval_test/EQ_u1_u1_1869/EQ_u1_u1_1869_inputs/RPIPE_MAC_ENABLE_1867/Sample/req
      -- CP-element group 185: 	 branch_block_stmt_1862/if_stmt_1866_eval_test/EQ_u1_u1_1869/EQ_u1_u1_1869_inputs/RPIPE_MAC_ENABLE_1867/Sample/ack
      -- CP-element group 185: 	 branch_block_stmt_1862/if_stmt_1866_eval_test/EQ_u1_u1_1869/EQ_u1_u1_1869_inputs/RPIPE_MAC_ENABLE_1867/Update/$entry
      -- CP-element group 185: 	 branch_block_stmt_1862/if_stmt_1866_eval_test/EQ_u1_u1_1869/EQ_u1_u1_1869_inputs/RPIPE_MAC_ENABLE_1867/Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_1862/if_stmt_1866_eval_test/EQ_u1_u1_1869/EQ_u1_u1_1869_inputs/RPIPE_MAC_ENABLE_1867/Update/req
      -- CP-element group 185: 	 branch_block_stmt_1862/if_stmt_1866_eval_test/EQ_u1_u1_1869/EQ_u1_u1_1869_inputs/RPIPE_MAC_ENABLE_1867/Update/ack
      -- CP-element group 185: 	 branch_block_stmt_1862/if_stmt_1866_eval_test/EQ_u1_u1_1869/SplitProtocol/$entry
      -- CP-element group 185: 	 branch_block_stmt_1862/if_stmt_1866_eval_test/EQ_u1_u1_1869/SplitProtocol/$exit
      -- CP-element group 185: 	 branch_block_stmt_1862/if_stmt_1866_eval_test/EQ_u1_u1_1869/SplitProtocol/Sample/$entry
      -- CP-element group 185: 	 branch_block_stmt_1862/if_stmt_1866_eval_test/EQ_u1_u1_1869/SplitProtocol/Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_1862/if_stmt_1866_eval_test/EQ_u1_u1_1869/SplitProtocol/Sample/rr
      -- CP-element group 185: 	 branch_block_stmt_1862/if_stmt_1866_eval_test/EQ_u1_u1_1869/SplitProtocol/Sample/ra
      -- CP-element group 185: 	 branch_block_stmt_1862/if_stmt_1866_eval_test/EQ_u1_u1_1869/SplitProtocol/Update/$entry
      -- CP-element group 185: 	 branch_block_stmt_1862/if_stmt_1866_eval_test/EQ_u1_u1_1869/SplitProtocol/Update/$exit
      -- CP-element group 185: 	 branch_block_stmt_1862/if_stmt_1866_eval_test/EQ_u1_u1_1869/SplitProtocol/Update/cr
      -- CP-element group 185: 	 branch_block_stmt_1862/if_stmt_1866_eval_test/EQ_u1_u1_1869/SplitProtocol/Update/ca
      -- CP-element group 185: 	 branch_block_stmt_1862/if_stmt_1866_eval_test/branch_req
      -- CP-element group 185: 	 branch_block_stmt_1862/EQ_u1_u1_1869_place
      -- CP-element group 185: 	 branch_block_stmt_1862/if_stmt_1866_if_link/$entry
      -- CP-element group 185: 	 branch_block_stmt_1862/if_stmt_1866_else_link/$entry
      -- CP-element group 185: 	 branch_block_stmt_1862/merge_stmt_1863_PhiReqMerge
      -- CP-element group 185: 	 branch_block_stmt_1862/merge_stmt_1863_PhiAck/$entry
      -- CP-element group 185: 	 branch_block_stmt_1862/merge_stmt_1863_PhiAck/$exit
      -- CP-element group 185: 	 branch_block_stmt_1862/merge_stmt_1863_PhiAck/dummy
      -- 
    branch_req_2920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SoftwareRegisterAccessDaemon_CP_2867_elements(185), ack => if_stmt_1866_branch_req_0); -- 
    SoftwareRegisterAccessDaemon_CP_2867_elements(185) <= OrReduce(SoftwareRegisterAccessDaemon_CP_2867_elements(2) & SoftwareRegisterAccessDaemon_CP_2867_elements(0));
    SoftwareRegisterAccessDaemon_do_while_stmt_1872_terminator_3590: loop_terminator -- 
      generic map (name => " SoftwareRegisterAccessDaemon_do_while_stmt_1872_terminator_3590", max_iterations_in_flight =>31) 
      port map(loop_body_exit => SoftwareRegisterAccessDaemon_CP_2867_elements(8),loop_continue => SoftwareRegisterAccessDaemon_CP_2867_elements(183),loop_terminate => SoftwareRegisterAccessDaemon_CP_2867_elements(182),loop_back => SoftwareRegisterAccessDaemon_CP_2867_elements(6),loop_exit => SoftwareRegisterAccessDaemon_CP_2867_elements(5),clk => clk, reset => reset); -- 
    phi_stmt_1874_phi_seq_2984_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= SoftwareRegisterAccessDaemon_CP_2867_elements(23);
      SoftwareRegisterAccessDaemon_CP_2867_elements(26)<= src_sample_reqs(0);
      src_sample_acks(0)  <= SoftwareRegisterAccessDaemon_CP_2867_elements(26);
      SoftwareRegisterAccessDaemon_CP_2867_elements(27)<= src_update_reqs(0);
      src_update_acks(0)  <= SoftwareRegisterAccessDaemon_CP_2867_elements(28);
      SoftwareRegisterAccessDaemon_CP_2867_elements(24) <= phi_mux_reqs(0);
      triggers(1)  <= SoftwareRegisterAccessDaemon_CP_2867_elements(21);
      SoftwareRegisterAccessDaemon_CP_2867_elements(30)<= src_sample_reqs(1);
      src_sample_acks(1)  <= SoftwareRegisterAccessDaemon_CP_2867_elements(30);
      SoftwareRegisterAccessDaemon_CP_2867_elements(31)<= src_update_reqs(1);
      src_update_acks(1)  <= SoftwareRegisterAccessDaemon_CP_2867_elements(32);
      SoftwareRegisterAccessDaemon_CP_2867_elements(22) <= phi_mux_reqs(1);
      phi_stmt_1874_phi_seq_2984 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_1874_phi_seq_2984") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => SoftwareRegisterAccessDaemon_CP_2867_elements(13), 
          phi_sample_ack => SoftwareRegisterAccessDaemon_CP_2867_elements(19), 
          phi_update_req => SoftwareRegisterAccessDaemon_CP_2867_elements(15), 
          phi_update_ack => SoftwareRegisterAccessDaemon_CP_2867_elements(20), 
          phi_mux_ack => SoftwareRegisterAccessDaemon_CP_2867_elements(25), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1880_phi_seq_3028_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= SoftwareRegisterAccessDaemon_CP_2867_elements(40);
      SoftwareRegisterAccessDaemon_CP_2867_elements(45)<= src_sample_reqs(0);
      src_sample_acks(0)  <= SoftwareRegisterAccessDaemon_CP_2867_elements(47);
      SoftwareRegisterAccessDaemon_CP_2867_elements(46)<= src_update_reqs(0);
      src_update_acks(0)  <= SoftwareRegisterAccessDaemon_CP_2867_elements(48);
      SoftwareRegisterAccessDaemon_CP_2867_elements(41) <= phi_mux_reqs(0);
      triggers(1)  <= SoftwareRegisterAccessDaemon_CP_2867_elements(42);
      SoftwareRegisterAccessDaemon_CP_2867_elements(49)<= src_sample_reqs(1);
      src_sample_acks(1)  <= SoftwareRegisterAccessDaemon_CP_2867_elements(49);
      SoftwareRegisterAccessDaemon_CP_2867_elements(50)<= src_update_reqs(1);
      src_update_acks(1)  <= SoftwareRegisterAccessDaemon_CP_2867_elements(51);
      SoftwareRegisterAccessDaemon_CP_2867_elements(43) <= phi_mux_reqs(1);
      phi_stmt_1880_phi_seq_3028 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_1880_phi_seq_3028") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => SoftwareRegisterAccessDaemon_CP_2867_elements(36), 
          phi_sample_ack => SoftwareRegisterAccessDaemon_CP_2867_elements(37), 
          phi_update_req => SoftwareRegisterAccessDaemon_CP_2867_elements(38), 
          phi_update_ack => SoftwareRegisterAccessDaemon_CP_2867_elements(39), 
          phi_mux_ack => SoftwareRegisterAccessDaemon_CP_2867_elements(44), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1885_phi_seq_3072_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= SoftwareRegisterAccessDaemon_CP_2867_elements(61);
      SoftwareRegisterAccessDaemon_CP_2867_elements(64)<= src_sample_reqs(0);
      src_sample_acks(0)  <= SoftwareRegisterAccessDaemon_CP_2867_elements(64);
      SoftwareRegisterAccessDaemon_CP_2867_elements(65)<= src_update_reqs(0);
      src_update_acks(0)  <= SoftwareRegisterAccessDaemon_CP_2867_elements(66);
      SoftwareRegisterAccessDaemon_CP_2867_elements(62) <= phi_mux_reqs(0);
      triggers(1)  <= SoftwareRegisterAccessDaemon_CP_2867_elements(59);
      SoftwareRegisterAccessDaemon_CP_2867_elements(68)<= src_sample_reqs(1);
      src_sample_acks(1)  <= SoftwareRegisterAccessDaemon_CP_2867_elements(70);
      SoftwareRegisterAccessDaemon_CP_2867_elements(69)<= src_update_reqs(1);
      src_update_acks(1)  <= SoftwareRegisterAccessDaemon_CP_2867_elements(71);
      SoftwareRegisterAccessDaemon_CP_2867_elements(60) <= phi_mux_reqs(1);
      phi_stmt_1885_phi_seq_3072 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_1885_phi_seq_3072") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => SoftwareRegisterAccessDaemon_CP_2867_elements(55), 
          phi_sample_ack => SoftwareRegisterAccessDaemon_CP_2867_elements(56), 
          phi_update_req => SoftwareRegisterAccessDaemon_CP_2867_elements(57), 
          phi_update_ack => SoftwareRegisterAccessDaemon_CP_2867_elements(58), 
          phi_mux_ack => SoftwareRegisterAccessDaemon_CP_2867_elements(63), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1890_phi_seq_3116_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= SoftwareRegisterAccessDaemon_CP_2867_elements(80);
      SoftwareRegisterAccessDaemon_CP_2867_elements(83)<= src_sample_reqs(0);
      src_sample_acks(0)  <= SoftwareRegisterAccessDaemon_CP_2867_elements(83);
      SoftwareRegisterAccessDaemon_CP_2867_elements(84)<= src_update_reqs(0);
      src_update_acks(0)  <= SoftwareRegisterAccessDaemon_CP_2867_elements(85);
      SoftwareRegisterAccessDaemon_CP_2867_elements(81) <= phi_mux_reqs(0);
      triggers(1)  <= SoftwareRegisterAccessDaemon_CP_2867_elements(78);
      SoftwareRegisterAccessDaemon_CP_2867_elements(87)<= src_sample_reqs(1);
      src_sample_acks(1)  <= SoftwareRegisterAccessDaemon_CP_2867_elements(89);
      SoftwareRegisterAccessDaemon_CP_2867_elements(88)<= src_update_reqs(1);
      src_update_acks(1)  <= SoftwareRegisterAccessDaemon_CP_2867_elements(90);
      SoftwareRegisterAccessDaemon_CP_2867_elements(79) <= phi_mux_reqs(1);
      phi_stmt_1890_phi_seq_3116 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_1890_phi_seq_3116") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => SoftwareRegisterAccessDaemon_CP_2867_elements(74), 
          phi_sample_ack => SoftwareRegisterAccessDaemon_CP_2867_elements(75), 
          phi_update_req => SoftwareRegisterAccessDaemon_CP_2867_elements(76), 
          phi_update_ack => SoftwareRegisterAccessDaemon_CP_2867_elements(77), 
          phi_mux_ack => SoftwareRegisterAccessDaemon_CP_2867_elements(82), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_2946_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= SoftwareRegisterAccessDaemon_CP_2867_elements(9);
        preds(1)  <= SoftwareRegisterAccessDaemon_CP_2867_elements(10);
        entry_tmerge_2946 : transition_merge -- 
          generic map(name => " entry_tmerge_2946")
          port map (preds => preds, symbol_out => SoftwareRegisterAccessDaemon_CP_2867_elements(11));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_1908_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_1916_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_1924_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_1869_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_1992_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_2001_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_2010_wire : std_logic_vector(0 downto 0);
    signal EQ_u32_u1_1941_wire : std_logic_vector(0 downto 0);
    signal EQ_u6_u1_1989_wire : std_logic_vector(0 downto 0);
    signal EQ_u6_u1_1998_wire : std_logic_vector(0 downto 0);
    signal EQ_u6_u1_2007_wire : std_logic_vector(0 downto 0);
    signal FREE_Q_32_1947 : std_logic_vector(31 downto 0);
    signal INIT_1874 : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1905_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1913_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1921_wire : std_logic_vector(0 downto 0);
    signal RPIPE_MAC_ENABLE_1867_wire : std_logic_vector(0 downto 0);
    signal R_index_2014_resized : std_logic_vector(5 downto 0);
    signal R_index_2014_scaled : std_logic_vector(5 downto 0);
    signal addr_1977 : std_logic_vector(35 downto 0);
    signal array_obj_ref_1899_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1899_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_1930_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1930_wire : std_logic_vector(31 downto 0);
    signal array_obj_ref_1930_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_1938_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1938_wire : std_logic_vector(31 downto 0);
    signal array_obj_ref_1938_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_1946_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1946_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_1959_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_1959_wire : std_logic_vector(31 downto 0);
    signal array_obj_ref_1959_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_2015_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_2015_final_offset : std_logic_vector(5 downto 0);
    signal array_obj_ref_2015_offset_scale_factor_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_2015_resized_base_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_2015_root_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_2015_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_2015_word_offset_0 : std_logic_vector(5 downto 0);
    signal bmask_1967_delayed_5_0_2022 : std_logic_vector(3 downto 0);
    signal bmask_1973 : std_logic_vector(3 downto 0);
    signal check_control_regsiter_1994 : std_logic_vector(0 downto 0);
    signal check_control_regsiter_1994_1882_buffered : std_logic_vector(0 downto 0);
    signal check_free_q_2003 : std_logic_vector(0 downto 0);
    signal check_free_q_2003_1889_buffered : std_logic_vector(0 downto 0);
    signal check_num_server_2012 : std_logic_vector(0 downto 0);
    signal check_num_server_2012_1894_buffered : std_logic_vector(0 downto 0);
    signal control_data_1900 : std_logic_vector(31 downto 0);
    signal control_register_1880 : std_logic_vector(0 downto 0);
    signal free_q_1885 : std_logic_vector(0 downto 0);
    signal index_1970_delayed_5_0_2028 : std_logic_vector(5 downto 0);
    signal index_1985 : std_logic_vector(5 downto 0);
    signal konst_1868_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1988_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1991_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1997_wire_constant : std_logic_vector(5 downto 0);
    signal konst_2000_wire_constant : std_logic_vector(0 downto 0);
    signal konst_2006_wire_constant : std_logic_vector(5 downto 0);
    signal konst_2009_wire_constant : std_logic_vector(0 downto 0);
    signal konst_2056_wire_constant : std_logic_vector(0 downto 0);
    signal num_server_1890 : std_logic_vector(0 downto 0);
    signal rdata_2045 : std_logic_vector(31 downto 0);
    signal req_1963 : std_logic_vector(73 downto 0);
    signal resp_2051 : std_logic_vector(32 downto 0);
    signal rval_2016 : std_logic_vector(31 downto 0);
    signal rwbar_1966_delayed_5_0_2019 : std_logic_vector(0 downto 0);
    signal rwbar_1969 : std_logic_vector(0 downto 0);
    signal rwbar_1974_delayed_5_0_2038 : std_logic_vector(0 downto 0);
    signal type_cast_1877_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1879_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1884_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1888_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1893_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1940_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1954_wire : std_logic_vector(35 downto 0);
    signal type_cast_2043_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_2048_wire_constant : std_logic_vector(0 downto 0);
    signal update_control_register_pipe_1887_delayed_5_0_1934 : std_logic_vector(0 downto 0);
    signal update_control_register_pipe_1910 : std_logic_vector(0 downto 0);
    signal update_free_q_pipe_1900_delayed_5_0_1950 : std_logic_vector(0 downto 0);
    signal update_free_q_pipe_1918 : std_logic_vector(0 downto 0);
    signal update_server_num_1926 : std_logic_vector(0 downto 0);
    signal wdata_1969_delayed_5_0_2025 : std_logic_vector(31 downto 0);
    signal wdata_1981 : std_logic_vector(31 downto 0);
    signal wval_2035 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    array_obj_ref_1899_word_address_0 <= "000000";
    array_obj_ref_1930_word_address_0 <= "000000";
    array_obj_ref_1938_word_address_0 <= "000000";
    array_obj_ref_1946_word_address_0 <= "010010";
    array_obj_ref_1959_word_address_0 <= "000001";
    array_obj_ref_2015_offset_scale_factor_0 <= "000001";
    array_obj_ref_2015_resized_base_address <= "000000";
    array_obj_ref_2015_word_offset_0 <= "000000";
    konst_1868_wire_constant <= "0";
    konst_1988_wire_constant <= "000000";
    konst_1991_wire_constant <= "0";
    konst_1997_wire_constant <= "010010";
    konst_2000_wire_constant <= "0";
    konst_2006_wire_constant <= "000001";
    konst_2009_wire_constant <= "0";
    konst_2056_wire_constant <= "1";
    type_cast_1877_wire_constant <= "0";
    type_cast_1879_wire_constant <= "1";
    type_cast_1884_wire_constant <= "0";
    type_cast_1888_wire_constant <= "0";
    type_cast_1893_wire_constant <= "0";
    type_cast_1940_wire_constant <= "00000000000000000000000000000001";
    type_cast_2043_wire_constant <= "00000000000000000000000000000000";
    type_cast_2048_wire_constant <= "0";
    phi_stmt_1874: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1877_wire_constant & type_cast_1879_wire_constant;
      req <= phi_stmt_1874_req_0 & phi_stmt_1874_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1874",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1874_ack_0,
          idata => idata,
          odata => INIT_1874,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1874
    phi_stmt_1880: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= check_control_regsiter_1994_1882_buffered & type_cast_1884_wire_constant;
      req <= phi_stmt_1880_req_0 & phi_stmt_1880_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1880",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1880_ack_0,
          idata => idata,
          odata => control_register_1880,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1880
    phi_stmt_1885: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1888_wire_constant & check_free_q_2003_1889_buffered;
      req <= phi_stmt_1885_req_0 & phi_stmt_1885_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1885",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1885_ack_0,
          idata => idata,
          odata => free_q_1885,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1885
    phi_stmt_1890: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1893_wire_constant & check_num_server_2012_1894_buffered;
      req <= phi_stmt_1890_req_0 & phi_stmt_1890_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1890",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1890_ack_0,
          idata => idata,
          odata => num_server_1890,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1890
    -- flow-through select operator MUX_2044_inst
    rdata_2045 <= rval_2016 when (rwbar_1974_delayed_5_0_2038(0) /=  '0') else type_cast_2043_wire_constant;
    -- flow-through slice operator slice_1968_inst
    rwbar_1969 <= req_1963(72 downto 72);
    -- flow-through slice operator slice_1972_inst
    bmask_1973 <= req_1963(71 downto 68);
    -- flow-through slice operator slice_1976_inst
    addr_1977 <= req_1963(67 downto 32);
    -- flow-through slice operator slice_1980_inst
    wdata_1981 <= req_1963(31 downto 0);
    -- flow-through slice operator slice_1984_inst
    index_1985 <= addr_1977(7 downto 2);
    W_bmask_1967_delayed_5_0_2020_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_bmask_1967_delayed_5_0_2020_inst_req_0;
      W_bmask_1967_delayed_5_0_2020_inst_ack_0<= wack(0);
      rreq(0) <= W_bmask_1967_delayed_5_0_2020_inst_req_1;
      W_bmask_1967_delayed_5_0_2020_inst_ack_1<= rack(0);
      W_bmask_1967_delayed_5_0_2020_inst : InterlockBuffer generic map ( -- 
        name => "W_bmask_1967_delayed_5_0_2020_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 4,
        out_data_width => 4,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => bmask_1973,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => bmask_1967_delayed_5_0_2022,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_index_1970_delayed_5_0_2026_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_index_1970_delayed_5_0_2026_inst_req_0;
      W_index_1970_delayed_5_0_2026_inst_ack_0<= wack(0);
      rreq(0) <= W_index_1970_delayed_5_0_2026_inst_req_1;
      W_index_1970_delayed_5_0_2026_inst_ack_1<= rack(0);
      W_index_1970_delayed_5_0_2026_inst : InterlockBuffer generic map ( -- 
        name => "W_index_1970_delayed_5_0_2026_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 6,
        out_data_width => 6,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => index_1985,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => index_1970_delayed_5_0_2028,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rwbar_1966_delayed_5_0_2017_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rwbar_1966_delayed_5_0_2017_inst_req_0;
      W_rwbar_1966_delayed_5_0_2017_inst_ack_0<= wack(0);
      rreq(0) <= W_rwbar_1966_delayed_5_0_2017_inst_req_1;
      W_rwbar_1966_delayed_5_0_2017_inst_ack_1<= rack(0);
      W_rwbar_1966_delayed_5_0_2017_inst : InterlockBuffer generic map ( -- 
        name => "W_rwbar_1966_delayed_5_0_2017_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rwbar_1969,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rwbar_1966_delayed_5_0_2019,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rwbar_1974_delayed_5_0_2036_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rwbar_1974_delayed_5_0_2036_inst_req_0;
      W_rwbar_1974_delayed_5_0_2036_inst_ack_0<= wack(0);
      rreq(0) <= W_rwbar_1974_delayed_5_0_2036_inst_req_1;
      W_rwbar_1974_delayed_5_0_2036_inst_ack_1<= rack(0);
      W_rwbar_1974_delayed_5_0_2036_inst : InterlockBuffer generic map ( -- 
        name => "W_rwbar_1974_delayed_5_0_2036_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rwbar_1969,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rwbar_1974_delayed_5_0_2038,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_update_control_register_pipe_1887_delayed_5_0_1932_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_update_control_register_pipe_1887_delayed_5_0_1932_inst_req_0;
      W_update_control_register_pipe_1887_delayed_5_0_1932_inst_ack_0<= wack(0);
      rreq(0) <= W_update_control_register_pipe_1887_delayed_5_0_1932_inst_req_1;
      W_update_control_register_pipe_1887_delayed_5_0_1932_inst_ack_1<= rack(0);
      W_update_control_register_pipe_1887_delayed_5_0_1932_inst : InterlockBuffer generic map ( -- 
        name => "W_update_control_register_pipe_1887_delayed_5_0_1932_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => update_control_register_pipe_1910,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => update_control_register_pipe_1887_delayed_5_0_1934,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_update_free_q_pipe_1900_delayed_5_0_1948_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_update_free_q_pipe_1900_delayed_5_0_1948_inst_req_0;
      W_update_free_q_pipe_1900_delayed_5_0_1948_inst_ack_0<= wack(0);
      rreq(0) <= W_update_free_q_pipe_1900_delayed_5_0_1948_inst_req_1;
      W_update_free_q_pipe_1900_delayed_5_0_1948_inst_ack_1<= rack(0);
      W_update_free_q_pipe_1900_delayed_5_0_1948_inst : InterlockBuffer generic map ( -- 
        name => "W_update_free_q_pipe_1900_delayed_5_0_1948_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => update_free_q_pipe_1918,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => update_free_q_pipe_1900_delayed_5_0_1950,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_wdata_1969_delayed_5_0_2023_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_wdata_1969_delayed_5_0_2023_inst_req_0;
      W_wdata_1969_delayed_5_0_2023_inst_ack_0<= wack(0);
      rreq(0) <= W_wdata_1969_delayed_5_0_2023_inst_req_1;
      W_wdata_1969_delayed_5_0_2023_inst_ack_1<= rack(0);
      W_wdata_1969_delayed_5_0_2023_inst : InterlockBuffer generic map ( -- 
        name => "W_wdata_1969_delayed_5_0_2023_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => wdata_1981,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => wdata_1969_delayed_5_0_2025,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    check_control_regsiter_1994_1882_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= check_control_regsiter_1994_1882_buf_req_0;
      check_control_regsiter_1994_1882_buf_ack_0<= wack(0);
      rreq(0) <= check_control_regsiter_1994_1882_buf_req_1;
      check_control_regsiter_1994_1882_buf_ack_1<= rack(0);
      check_control_regsiter_1994_1882_buf : InterlockBuffer generic map ( -- 
        name => "check_control_regsiter_1994_1882_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => check_control_regsiter_1994,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => check_control_regsiter_1994_1882_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    check_free_q_2003_1889_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= check_free_q_2003_1889_buf_req_0;
      check_free_q_2003_1889_buf_ack_0<= wack(0);
      rreq(0) <= check_free_q_2003_1889_buf_req_1;
      check_free_q_2003_1889_buf_ack_1<= rack(0);
      check_free_q_2003_1889_buf : InterlockBuffer generic map ( -- 
        name => "check_free_q_2003_1889_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => check_free_q_2003,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => check_free_q_2003_1889_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    check_num_server_2012_1894_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= check_num_server_2012_1894_buf_req_0;
      check_num_server_2012_1894_buf_ack_0<= wack(0);
      rreq(0) <= check_num_server_2012_1894_buf_req_1;
      check_num_server_2012_1894_buf_ack_1<= rack(0);
      check_num_server_2012_1894_buf : InterlockBuffer generic map ( -- 
        name => "check_num_server_2012_1894_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => check_num_server_2012,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => check_num_server_2012_1894_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    type_cast_1954_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= type_cast_1954_inst_req_0;
      type_cast_1954_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= type_cast_1954_inst_req_1;
      type_cast_1954_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  update_free_q_pipe_1900_delayed_5_0_1950(0);
      type_cast_1954_inst_gI: SplitGuardInterface generic map(name => "type_cast_1954_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      type_cast_1954_inst : InterlockBuffer generic map ( -- 
        name => "type_cast_1954_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 36,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => FREE_Q_32_1947,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => type_cast_1954_wire,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- equivalence array_obj_ref_1899_gather_scatter
    process(array_obj_ref_1899_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1899_data_0;
      ov(31 downto 0) := iv;
      control_data_1900 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1930_gather_scatter
    process(array_obj_ref_1930_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1930_data_0;
      ov(31 downto 0) := iv;
      array_obj_ref_1930_wire <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1938_gather_scatter
    process(array_obj_ref_1938_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1938_data_0;
      ov(31 downto 0) := iv;
      array_obj_ref_1938_wire <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1946_gather_scatter
    process(array_obj_ref_1946_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1946_data_0;
      ov(31 downto 0) := iv;
      FREE_Q_32_1947 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_1959_gather_scatter
    process(array_obj_ref_1959_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_1959_data_0;
      ov(31 downto 0) := iv;
      array_obj_ref_1959_wire <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2015_addr_0
    process(array_obj_ref_2015_root_address) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2015_root_address;
      ov(5 downto 0) := iv;
      array_obj_ref_2015_word_address_0 <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2015_gather_scatter
    process(array_obj_ref_2015_data_0) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2015_data_0;
      ov(31 downto 0) := iv;
      rval_2016 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2015_index_0_rename
    process(R_index_2014_resized) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_2014_resized;
      ov(5 downto 0) := iv;
      R_index_2014_scaled <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2015_index_0_resize
    process(index_1985) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := index_1985;
      ov(5 downto 0) := iv;
      R_index_2014_resized <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2015_index_offset
    process(R_index_2014_scaled) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_2014_scaled;
      ov(5 downto 0) := iv;
      array_obj_ref_2015_final_offset <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_2015_root_address_inst
    process(array_obj_ref_2015_final_offset) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_2015_final_offset;
      ov(5 downto 0) := iv;
      array_obj_ref_2015_root_address <= ov(5 downto 0);
      --
    end process;
    do_while_stmt_1872_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_2056_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1872_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1872_branch_req_0,
          ack0 => do_while_stmt_1872_branch_ack_0,
          ack1 => do_while_stmt_1872_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1866_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= EQ_u1_u1_1869_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1866_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1866_branch_req_0,
          ack0 => if_stmt_1866_branch_ack_0,
          ack1 => if_stmt_1866_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator AND_u1_u1_1908_inst
    process(INIT_1874, control_register_1880) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(INIT_1874, control_register_1880, tmp_var);
      AND_u1_u1_1908_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1916_inst
    process(INIT_1874, free_q_1885) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(INIT_1874, free_q_1885, tmp_var);
      AND_u1_u1_1916_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1924_inst
    process(INIT_1874, num_server_1890) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(INIT_1874, num_server_1890, tmp_var);
      AND_u1_u1_1924_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1993_inst
    process(EQ_u6_u1_1989_wire, EQ_u1_u1_1992_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u6_u1_1989_wire, EQ_u1_u1_1992_wire, tmp_var);
      check_control_regsiter_1994 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2002_inst
    process(EQ_u6_u1_1998_wire, EQ_u1_u1_2001_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u6_u1_1998_wire, EQ_u1_u1_2001_wire, tmp_var);
      check_free_q_2003 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2011_inst
    process(EQ_u6_u1_2007_wire, EQ_u1_u1_2010_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u6_u1_2007_wire, EQ_u1_u1_2010_wire, tmp_var);
      check_num_server_2012 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u33_2050_inst
    process(type_cast_2048_wire_constant, rdata_2045) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_2048_wire_constant, rdata_2045, tmp_var);
      resp_2051 <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_1869_inst
    process(RPIPE_MAC_ENABLE_1867_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(RPIPE_MAC_ENABLE_1867_wire, konst_1868_wire_constant, tmp_var);
      EQ_u1_u1_1869_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_1992_inst
    process(rwbar_1969) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(rwbar_1969, konst_1991_wire_constant, tmp_var);
      EQ_u1_u1_1992_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_2001_inst
    process(rwbar_1969) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(rwbar_1969, konst_2000_wire_constant, tmp_var);
      EQ_u1_u1_2001_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_2010_inst
    process(rwbar_1969) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(rwbar_1969, konst_2009_wire_constant, tmp_var);
      EQ_u1_u1_2010_wire <= tmp_var; --
    end process;
    -- shared split operator group (11) : EQ_u32_u1_1941_inst 
    ApIntEq_group_11: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= array_obj_ref_1938_wire;
      EQ_u32_u1_1941_wire <= data_out(0 downto 0);
      guard_vector(0)  <= update_control_register_pipe_1887_delayed_5_0_1934(0);
      reqL_unguarded(0) <= EQ_u32_u1_1941_inst_req_0;
      EQ_u32_u1_1941_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u32_u1_1941_inst_req_1;
      EQ_u32_u1_1941_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_11_gI: SplitGuardInterface generic map(name => "ApIntEq_group_11_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_11",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 11
    -- binary operator EQ_u6_u1_1989_inst
    process(index_1985) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(index_1985, konst_1988_wire_constant, tmp_var);
      EQ_u6_u1_1989_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u6_u1_1998_inst
    process(index_1985) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(index_1985, konst_1997_wire_constant, tmp_var);
      EQ_u6_u1_1998_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u6_u1_2007_inst
    process(index_1985) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(index_1985, konst_2006_wire_constant, tmp_var);
      EQ_u6_u1_2007_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1905_inst
    process(INIT_1874) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", INIT_1874, tmp_var);
      NOT_u1_u1_1905_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1913_inst
    process(INIT_1874) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", INIT_1874, tmp_var);
      NOT_u1_u1_1913_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1921_inst
    process(INIT_1874) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", INIT_1874, tmp_var);
      NOT_u1_u1_1921_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_1909_inst
    process(NOT_u1_u1_1905_wire, AND_u1_u1_1908_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1905_wire, AND_u1_u1_1908_wire, tmp_var);
      update_control_register_pipe_1910 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1917_inst
    process(NOT_u1_u1_1913_wire, AND_u1_u1_1916_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1913_wire, AND_u1_u1_1916_wire, tmp_var);
      update_free_q_pipe_1918 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1925_inst
    process(NOT_u1_u1_1921_wire, AND_u1_u1_1924_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_1921_wire, AND_u1_u1_1924_wire, tmp_var);
      update_server_num_1926 <= tmp_var; --
    end process;
    -- shared load operator group (0) : array_obj_ref_1946_load_0 array_obj_ref_1959_load_0 array_obj_ref_2015_load_0 array_obj_ref_1938_load_0 array_obj_ref_1930_load_0 array_obj_ref_1899_load_0 
    LoadGroup0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(191 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 5 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 5 downto 0);
      signal reqL_unregulated, ackL_unregulated: BooleanArray( 5 downto 0);
      signal guard_vector : std_logic_vector( 5 downto 0);
      constant inBUFs : IntegerArray(5 downto 0) := (5 => 2, 4 => 2, 3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant outBUFs : IntegerArray(5 downto 0) := (5 => 2, 4 => 2, 3 => 2, 2 => 2, 1 => 2, 0 => 2);
      constant guardFlags : BooleanArray(5 downto 0) := (0 => false, 1 => true, 2 => true, 3 => false, 4 => true, 5 => true);
      constant guardBuffering: IntegerArray(5 downto 0)  := (0 => 5, 1 => 5, 2 => 5, 3 => 5, 4 => 5, 5 => 5);
      -- 
    begin -- 
      reqL_unguarded(5) <= array_obj_ref_1946_load_0_req_0;
      reqL_unguarded(4) <= array_obj_ref_1959_load_0_req_0;
      reqL_unguarded(3) <= array_obj_ref_2015_load_0_req_0;
      reqL_unguarded(2) <= array_obj_ref_1938_load_0_req_0;
      reqL_unguarded(1) <= array_obj_ref_1930_load_0_req_0;
      reqL_unguarded(0) <= array_obj_ref_1899_load_0_req_0;
      array_obj_ref_1946_load_0_ack_0 <= ackL_unguarded(5);
      array_obj_ref_1959_load_0_ack_0 <= ackL_unguarded(4);
      array_obj_ref_2015_load_0_ack_0 <= ackL_unguarded(3);
      array_obj_ref_1938_load_0_ack_0 <= ackL_unguarded(2);
      array_obj_ref_1930_load_0_ack_0 <= ackL_unguarded(1);
      array_obj_ref_1899_load_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(5) <= array_obj_ref_1946_load_0_req_1;
      reqR_unguarded(4) <= array_obj_ref_1959_load_0_req_1;
      reqR_unguarded(3) <= array_obj_ref_2015_load_0_req_1;
      reqR_unguarded(2) <= array_obj_ref_1938_load_0_req_1;
      reqR_unguarded(1) <= array_obj_ref_1930_load_0_req_1;
      reqR_unguarded(0) <= array_obj_ref_1899_load_0_req_1;
      array_obj_ref_1946_load_0_ack_1 <= ackR_unguarded(5);
      array_obj_ref_1959_load_0_ack_1 <= ackR_unguarded(4);
      array_obj_ref_2015_load_0_ack_1 <= ackR_unguarded(3);
      array_obj_ref_1938_load_0_ack_1 <= ackR_unguarded(2);
      array_obj_ref_1930_load_0_ack_1 <= ackR_unguarded(1);
      array_obj_ref_1899_load_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <= update_control_register_pipe_1910(0);
      guard_vector(2)  <= update_control_register_pipe_1887_delayed_5_0_1934(0);
      guard_vector(3)  <=  '1';
      guard_vector(4)  <= update_server_num_1926(0);
      guard_vector(5)  <= update_free_q_pipe_1918(0);
      LoadGroup0_accessRegulator_0: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_1: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_2: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_3: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_4: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_4", num_slots => 1) -- 
        port map (req => reqL_unregulated(4), -- 
          ack => ackL_unregulated(4),
          regulated_req => reqL(4),
          regulated_ack => ackL(4),
          release_req => reqR(4),
          release_ack => ackR(4),
          clk => clk, reset => reset); -- 
      LoadGroup0_accessRegulator_5: access_regulator_base generic map (name => "LoadGroup0_accessRegulator_5", num_slots => 1) -- 
        port map (req => reqL_unregulated(5), -- 
          ack => ackL_unregulated(5),
          regulated_req => reqL(5),
          regulated_ack => ackL(5),
          release_req => reqR(5),
          release_ack => ackR(5),
          clk => clk, reset => reset); -- 
      LoadGroup0_gI: SplitGuardInterface generic map(name => "LoadGroup0_gI", nreqs => 6, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= array_obj_ref_1946_word_address_0 & array_obj_ref_1959_word_address_0 & array_obj_ref_2015_word_address_0 & array_obj_ref_1938_word_address_0 & array_obj_ref_1930_word_address_0 & array_obj_ref_1899_word_address_0;
      array_obj_ref_1946_data_0 <= data_out(191 downto 160);
      array_obj_ref_1959_data_0 <= data_out(159 downto 128);
      array_obj_ref_2015_data_0 <= data_out(127 downto 96);
      array_obj_ref_1938_data_0 <= data_out(95 downto 64);
      array_obj_ref_1930_data_0 <= data_out(63 downto 32);
      array_obj_ref_1899_data_0 <= data_out(31 downto 0);
      LoadReq: LoadReqSharedWithInputBuffers -- 
        generic map ( name => "LoadGroup0", addr_width => 6,
        num_reqs => 6,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          mreq => memory_space_2_lr_req(0),
          mack => memory_space_2_lr_ack(0),
          maddr => memory_space_2_lr_addr(5 downto 0),
          mtag => memory_space_2_lr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      LoadComplete: LoadCompleteShared -- 
        generic map ( name => "LoadGroup0 load-complete ",
        data_width => 32,
        num_reqs => 6,
        tag_length => 3,
        detailed_buffering_per_output => outBUFs, 
        no_arbitration => false)
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          mreq => memory_space_2_lc_req(0),
          mack => memory_space_2_lc_ack(0),
          mdata => memory_space_2_lc_data(31 downto 0),
          mtag => memory_space_2_lc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- load group 0
    -- shared inport operator group (0) : RPIPE_AFB_NIC_REQUEST_1962_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(73 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_AFB_NIC_REQUEST_1962_inst_req_0;
      RPIPE_AFB_NIC_REQUEST_1962_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_AFB_NIC_REQUEST_1962_inst_req_1;
      RPIPE_AFB_NIC_REQUEST_1962_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      req_1963 <= data_out(73 downto 0);
      AFB_NIC_REQUEST_read_0_gI: SplitGuardInterface generic map(name => "AFB_NIC_REQUEST_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      AFB_NIC_REQUEST_read_0: InputPortRevised -- 
        generic map ( name => "AFB_NIC_REQUEST_read_0", data_width => 74,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => AFB_NIC_REQUEST_pipe_read_req(0),
          oack => AFB_NIC_REQUEST_pipe_read_ack(0),
          odata => AFB_NIC_REQUEST_pipe_read_data(73 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- read from input-signal MAC_ENABLE
    RPIPE_MAC_ENABLE_1867_wire <= MAC_ENABLE;
    -- shared outport operator group (0) : WPIPE_AFB_NIC_RESPONSE_2052_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(32 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_AFB_NIC_RESPONSE_2052_inst_req_0;
      WPIPE_AFB_NIC_RESPONSE_2052_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_AFB_NIC_RESPONSE_2052_inst_req_1;
      WPIPE_AFB_NIC_RESPONSE_2052_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= resp_2051;
      AFB_NIC_RESPONSE_write_0_gI: SplitGuardInterface generic map(name => "AFB_NIC_RESPONSE_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      AFB_NIC_RESPONSE_write_0: OutputPortRevised -- 
        generic map ( name => "AFB_NIC_RESPONSE", data_width => 33, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => AFB_NIC_RESPONSE_pipe_write_req(0),
          oack => AFB_NIC_RESPONSE_pipe_write_ack(0),
          odata => AFB_NIC_RESPONSE_pipe_write_data(32 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_CONTROL_REGISTER_1928_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_CONTROL_REGISTER_1928_inst_req_0;
      WPIPE_CONTROL_REGISTER_1928_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_CONTROL_REGISTER_1928_inst_req_1;
      WPIPE_CONTROL_REGISTER_1928_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= update_control_register_pipe_1910(0);
      data_in <= array_obj_ref_1930_wire;
      CONTROL_REGISTER_write_1_gI: SplitGuardInterface generic map(name => "CONTROL_REGISTER_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      CONTROL_REGISTER_write_1: OutputPortRevised -- 
        generic map ( name => "CONTROL_REGISTER", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => CONTROL_REGISTER_pipe_write_req(0),
          oack => CONTROL_REGISTER_pipe_write_ack(0),
          odata => CONTROL_REGISTER_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_FREE_Q_1952_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_FREE_Q_1952_inst_req_0;
      WPIPE_FREE_Q_1952_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_FREE_Q_1952_inst_req_1;
      WPIPE_FREE_Q_1952_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= update_free_q_pipe_1900_delayed_5_0_1950(0);
      data_in <= type_cast_1954_wire;
      FREE_Q_write_2_gI: SplitGuardInterface generic map(name => "FREE_Q_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      FREE_Q_write_2: OutputPortRevised -- 
        generic map ( name => "FREE_Q", data_width => 36, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => FREE_Q_pipe_write_req(0),
          oack => FREE_Q_pipe_write_ack(0),
          odata => FREE_Q_pipe_write_data(35 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_NUMBER_OF_SERVERS_1957_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_NUMBER_OF_SERVERS_1957_inst_req_0;
      WPIPE_NUMBER_OF_SERVERS_1957_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_NUMBER_OF_SERVERS_1957_inst_req_1;
      WPIPE_NUMBER_OF_SERVERS_1957_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= update_server_num_1926(0);
      data_in <= array_obj_ref_1959_wire;
      NUMBER_OF_SERVERS_write_3_gI: SplitGuardInterface generic map(name => "NUMBER_OF_SERVERS_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      NUMBER_OF_SERVERS_write_3: OutputPortRevised -- 
        generic map ( name => "NUMBER_OF_SERVERS", data_width => 32, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => NUMBER_OF_SERVERS_pipe_write_req(0),
          oack => NUMBER_OF_SERVERS_pipe_write_ack(0),
          odata => NUMBER_OF_SERVERS_pipe_write_data(31 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    -- shared outport operator group (4) : WPIPE_enable_mac_1936_inst 
    OutportGroup_4: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_enable_mac_1936_inst_req_0;
      WPIPE_enable_mac_1936_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_enable_mac_1936_inst_req_1;
      WPIPE_enable_mac_1936_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= update_control_register_pipe_1887_delayed_5_0_1934(0);
      data_in <= EQ_u32_u1_1941_wire;
      enable_mac_write_4_gI: SplitGuardInterface generic map(name => "enable_mac_write_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      enable_mac_write_4: OutputPortRevised -- 
        generic map ( name => "enable_mac", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => enable_mac_pipe_write_req(0),
          oack => enable_mac_pipe_write_ack(0),
          odata => enable_mac_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 4
    -- shared call operator group (0) : call_stmt_2035_call 
    UpdateRegister_call_group_0: Block -- 
      signal data_in: std_logic_vector(73 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_2035_call_req_0;
      call_stmt_2035_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_2035_call_req_1;
      call_stmt_2035_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not rwbar_1966_delayed_5_0_2019(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      UpdateRegister_call_group_0_gI: SplitGuardInterface generic map(name => "UpdateRegister_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= bmask_1967_delayed_5_0_2022 & rval_2016 & wdata_1969_delayed_5_0_2025 & index_1970_delayed_5_0_2028;
      wval_2035 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 74,
        owidth => 74,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => UpdateRegister_call_reqs(0),
          ackR => UpdateRegister_call_acks(0),
          dataR => UpdateRegister_call_data(73 downto 0),
          tagR => UpdateRegister_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => UpdateRegister_return_acks(0), -- cross-over
          ackL => UpdateRegister_return_reqs(0), -- cross-over
          dataL => UpdateRegister_return_data(31 downto 0),
          tagL => UpdateRegister_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end SoftwareRegisterAccessDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.nic_system_global_package.all;
entity UpdateRegister is -- 
  generic (tag_length : integer); 
  port ( -- 
    bmask : in  std_logic_vector(3 downto 0);
    rval : in  std_logic_vector(31 downto 0);
    wdata : in  std_logic_vector(31 downto 0);
    index : in  std_logic_vector(5 downto 0);
    wval : out  std_logic_vector(31 downto 0);
    memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sr_addr : out  std_logic_vector(5 downto 0);
    memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
    memory_space_2_sr_tag :  out  std_logic_vector(20 downto 0);
    memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
    memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
    memory_space_2_sc_tag :  in  std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity UpdateRegister;
architecture UpdateRegister_arch of UpdateRegister is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 74)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal bmask_buffer :  std_logic_vector(3 downto 0);
  signal bmask_update_enable: Boolean;
  signal rval_buffer :  std_logic_vector(31 downto 0);
  signal rval_update_enable: Boolean;
  signal wdata_buffer :  std_logic_vector(31 downto 0);
  signal wdata_update_enable: Boolean;
  signal index_buffer :  std_logic_vector(5 downto 0);
  signal index_update_enable: Boolean;
  -- output port buffer signals
  signal wval_buffer :  std_logic_vector(31 downto 0);
  signal wval_update_enable: Boolean;
  signal UpdateRegister_CP_434_start: Boolean;
  signal UpdateRegister_CP_434_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal CONCAT_u16_u32_395_inst_req_0 : boolean;
  signal CONCAT_u16_u32_395_inst_ack_0 : boolean;
  signal CONCAT_u16_u32_395_inst_req_1 : boolean;
  signal CONCAT_u16_u32_395_inst_ack_1 : boolean;
  signal array_obj_ref_398_store_0_req_0 : boolean;
  signal array_obj_ref_398_store_0_ack_0 : boolean;
  signal array_obj_ref_398_store_0_req_1 : boolean;
  signal array_obj_ref_398_store_0_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "UpdateRegister_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 74) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(3 downto 0) <= bmask;
  bmask_buffer <= in_buffer_data_out(3 downto 0);
  in_buffer_data_in(35 downto 4) <= rval;
  rval_buffer <= in_buffer_data_out(35 downto 4);
  in_buffer_data_in(67 downto 36) <= wdata;
  wdata_buffer <= in_buffer_data_out(67 downto 36);
  in_buffer_data_in(73 downto 68) <= index;
  index_buffer <= in_buffer_data_out(73 downto 68);
  in_buffer_data_in(tag_length + 73 downto 74) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 73 downto 74);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  UpdateRegister_CP_434_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "UpdateRegister_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= wval_buffer;
  wval <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= UpdateRegister_CP_434_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= UpdateRegister_CP_434_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= UpdateRegister_CP_434_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  UpdateRegister_CP_434: Block -- control-path 
    signal UpdateRegister_CP_434_elements: BooleanArray(5 downto 0);
    -- 
  begin -- 
    UpdateRegister_CP_434_elements(0) <= UpdateRegister_CP_434_start;
    UpdateRegister_CP_434_symbol <= UpdateRegister_CP_434_elements(5);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	3 
    -- CP-element group 0: 	5 
    -- CP-element group 0:  members (39) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/$entry
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/CONCAT_u16_u32_395_sample_start_
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/CONCAT_u16_u32_395_update_start_
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/CONCAT_u16_u32_395_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/CONCAT_u16_u32_395_Sample/rr
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/CONCAT_u16_u32_395_Update/$entry
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/CONCAT_u16_u32_395_Update/cr
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_update_start_
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_word_address_calculated
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_root_address_calculated
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_offset_calculated
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_index_resized_0
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_index_scaled_0
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_index_computed_0
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_index_resize_0/$entry
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_index_resize_0/$exit
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_index_resize_0/index_resize_req
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_index_resize_0/index_resize_ack
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_index_scale_0/$entry
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_index_scale_0/$exit
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_index_scale_0/scale_rename_req
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_index_scale_0/scale_rename_ack
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_final_index_sum_regn/$entry
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_final_index_sum_regn/$exit
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_final_index_sum_regn/req
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_final_index_sum_regn/ack
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_base_plus_offset/$entry
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_base_plus_offset/$exit
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_base_plus_offset/sum_rename_req
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_base_plus_offset/sum_rename_ack
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_word_addrgen/$entry
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_word_addrgen/$exit
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_word_addrgen/root_register_req
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_word_addrgen/root_register_ack
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_Update/$entry
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_Update/word_access_complete/$entry
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_Update/word_access_complete/word_0/$entry
      -- CP-element group 0: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_Update/word_access_complete/word_0/cr
      -- 
    rr_447_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_447_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UpdateRegister_CP_434_elements(0), ack => CONCAT_u16_u32_395_inst_req_0); -- 
    cr_452_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_452_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UpdateRegister_CP_434_elements(0), ack => CONCAT_u16_u32_395_inst_req_1); -- 
    cr_514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UpdateRegister_CP_434_elements(0), ack => array_obj_ref_398_store_0_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_331_to_assign_stmt_400/CONCAT_u16_u32_395_sample_completed_
      -- CP-element group 1: 	 assign_stmt_331_to_assign_stmt_400/CONCAT_u16_u32_395_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_331_to_assign_stmt_400/CONCAT_u16_u32_395_Sample/ra
      -- 
    ra_448_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u16_u32_395_inst_ack_0, ack => UpdateRegister_CP_434_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 assign_stmt_331_to_assign_stmt_400/CONCAT_u16_u32_395_update_completed_
      -- CP-element group 2: 	 assign_stmt_331_to_assign_stmt_400/CONCAT_u16_u32_395_Update/$exit
      -- CP-element group 2: 	 assign_stmt_331_to_assign_stmt_400/CONCAT_u16_u32_395_Update/ca
      -- 
    ca_453_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u16_u32_395_inst_ack_1, ack => UpdateRegister_CP_434_elements(2)); -- 
    -- CP-element group 3:  join  transition  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (9) 
      -- CP-element group 3: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_sample_start_
      -- CP-element group 3: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_Sample/$entry
      -- CP-element group 3: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_Sample/array_obj_ref_398_Split/$entry
      -- CP-element group 3: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_Sample/array_obj_ref_398_Split/$exit
      -- CP-element group 3: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_Sample/array_obj_ref_398_Split/split_req
      -- CP-element group 3: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_Sample/array_obj_ref_398_Split/split_ack
      -- CP-element group 3: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_Sample/word_access_start/$entry
      -- CP-element group 3: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_Sample/word_access_start/word_0/$entry
      -- CP-element group 3: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_Sample/word_access_start/word_0/rr
      -- 
    rr_503_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_503_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => UpdateRegister_CP_434_elements(3), ack => array_obj_ref_398_store_0_req_0); -- 
    UpdateRegister_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "UpdateRegister_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= UpdateRegister_CP_434_elements(0) & UpdateRegister_CP_434_elements(2);
      gj_UpdateRegister_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => UpdateRegister_CP_434_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_sample_completed_
      -- CP-element group 4: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_Sample/$exit
      -- CP-element group 4: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_Sample/word_access_start/$exit
      -- CP-element group 4: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_Sample/word_access_start/word_0/$exit
      -- CP-element group 4: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_Sample/word_access_start/word_0/ra
      -- 
    ra_504_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_398_store_0_ack_0, ack => UpdateRegister_CP_434_elements(4)); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	0 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (7) 
      -- CP-element group 5: 	 $exit
      -- CP-element group 5: 	 assign_stmt_331_to_assign_stmt_400/$exit
      -- CP-element group 5: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_update_completed_
      -- CP-element group 5: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_Update/$exit
      -- CP-element group 5: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_Update/word_access_complete/$exit
      -- CP-element group 5: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_Update/word_access_complete/word_0/$exit
      -- CP-element group 5: 	 assign_stmt_331_to_assign_stmt_400/array_obj_ref_398_Update/word_access_complete/word_0/ca
      -- 
    ca_515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => array_obj_ref_398_store_0_ack_1, ack => UpdateRegister_CP_434_elements(5)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u8_u16_385_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_394_wire : std_logic_vector(15 downto 0);
    signal MUX_380_wire : std_logic_vector(7 downto 0);
    signal MUX_384_wire : std_logic_vector(7 downto 0);
    signal MUX_389_wire : std_logic_vector(7 downto 0);
    signal MUX_393_wire : std_logic_vector(7 downto 0);
    signal R_index_397_resized : std_logic_vector(5 downto 0);
    signal R_index_397_scaled : std_logic_vector(5 downto 0);
    signal array_obj_ref_398_data_0 : std_logic_vector(31 downto 0);
    signal array_obj_ref_398_final_offset : std_logic_vector(5 downto 0);
    signal array_obj_ref_398_offset_scale_factor_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_398_resized_base_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_398_root_address : std_logic_vector(5 downto 0);
    signal array_obj_ref_398_word_address_0 : std_logic_vector(5 downto 0);
    signal array_obj_ref_398_word_offset_0 : std_logic_vector(5 downto 0);
    signal b0_331 : std_logic_vector(0 downto 0);
    signal b1_335 : std_logic_vector(0 downto 0);
    signal b2_339 : std_logic_vector(0 downto 0);
    signal b3_343 : std_logic_vector(0 downto 0);
    signal r0_347 : std_logic_vector(7 downto 0);
    signal r1_351 : std_logic_vector(7 downto 0);
    signal r2_355 : std_logic_vector(7 downto 0);
    signal r3_359 : std_logic_vector(7 downto 0);
    signal w0_363 : std_logic_vector(7 downto 0);
    signal w1_367 : std_logic_vector(7 downto 0);
    signal w2_371 : std_logic_vector(7 downto 0);
    signal w3_375 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    array_obj_ref_398_offset_scale_factor_0 <= "000001";
    array_obj_ref_398_resized_base_address <= "000000";
    array_obj_ref_398_word_offset_0 <= "000000";
    -- flow-through select operator MUX_380_inst
    MUX_380_wire <= w0_363 when (b0_331(0) /=  '0') else r0_347;
    -- flow-through select operator MUX_384_inst
    MUX_384_wire <= w1_367 when (b1_335(0) /=  '0') else r1_351;
    -- flow-through select operator MUX_389_inst
    MUX_389_wire <= w2_371 when (b2_339(0) /=  '0') else r2_355;
    -- flow-through select operator MUX_393_inst
    MUX_393_wire <= w3_375 when (b3_343(0) /=  '0') else r3_359;
    -- flow-through slice operator slice_330_inst
    b0_331 <= bmask_buffer(3 downto 3);
    -- flow-through slice operator slice_334_inst
    b1_335 <= bmask_buffer(2 downto 2);
    -- flow-through slice operator slice_338_inst
    b2_339 <= bmask_buffer(1 downto 1);
    -- flow-through slice operator slice_342_inst
    b3_343 <= bmask_buffer(0 downto 0);
    -- flow-through slice operator slice_346_inst
    r0_347 <= rval_buffer(31 downto 24);
    -- flow-through slice operator slice_350_inst
    r1_351 <= rval_buffer(23 downto 16);
    -- flow-through slice operator slice_354_inst
    r2_355 <= rval_buffer(15 downto 8);
    -- flow-through slice operator slice_358_inst
    r3_359 <= rval_buffer(7 downto 0);
    -- flow-through slice operator slice_362_inst
    w0_363 <= wdata_buffer(31 downto 24);
    -- flow-through slice operator slice_366_inst
    w1_367 <= wdata_buffer(23 downto 16);
    -- flow-through slice operator slice_370_inst
    w2_371 <= wdata_buffer(15 downto 8);
    -- flow-through slice operator slice_374_inst
    w3_375 <= wdata_buffer(7 downto 0);
    -- equivalence array_obj_ref_398_addr_0
    process(array_obj_ref_398_root_address) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_398_root_address;
      ov(5 downto 0) := iv;
      array_obj_ref_398_word_address_0 <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_398_gather_scatter
    process(wval_buffer) --
      variable iv : std_logic_vector(31 downto 0);
      variable ov : std_logic_vector(31 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := wval_buffer;
      ov(31 downto 0) := iv;
      array_obj_ref_398_data_0 <= ov(31 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_398_index_0_rename
    process(R_index_397_resized) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_397_resized;
      ov(5 downto 0) := iv;
      R_index_397_scaled <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_398_index_0_resize
    process(index_buffer) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := index_buffer;
      ov(5 downto 0) := iv;
      R_index_397_resized <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_398_index_offset
    process(R_index_397_scaled) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := R_index_397_scaled;
      ov(5 downto 0) := iv;
      array_obj_ref_398_final_offset <= ov(5 downto 0);
      --
    end process;
    -- equivalence array_obj_ref_398_root_address_inst
    process(array_obj_ref_398_final_offset) --
      variable iv : std_logic_vector(5 downto 0);
      variable ov : std_logic_vector(5 downto 0);
      -- 
    begin -- 
      ov := (others => '0');
      iv := array_obj_ref_398_final_offset;
      ov(5 downto 0) := iv;
      array_obj_ref_398_root_address <= ov(5 downto 0);
      --
    end process;
    -- shared split operator group (0) : CONCAT_u16_u32_395_inst 
    ApConcat_group_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u8_u16_385_wire & CONCAT_u8_u16_394_wire;
      wval_buffer <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u16_u32_395_inst_req_0;
      CONCAT_u16_u32_395_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u16_u32_395_inst_req_1;
      CONCAT_u16_u32_395_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_0_gI: SplitGuardInterface generic map(name => "ApConcat_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 16,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 16, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- binary operator CONCAT_u8_u16_385_inst
    process(MUX_380_wire, MUX_384_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_380_wire, MUX_384_wire, tmp_var);
      CONCAT_u8_u16_385_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u16_394_inst
    process(MUX_389_wire, MUX_393_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_389_wire, MUX_393_wire, tmp_var);
      CONCAT_u8_u16_394_wire <= tmp_var; --
    end process;
    -- shared store operator group (0) : array_obj_ref_398_store_0 
    StoreGroup0: Block -- 
      signal addr_in: std_logic_vector(5 downto 0);
      signal data_in: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= array_obj_ref_398_store_0_req_0;
      array_obj_ref_398_store_0_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= array_obj_ref_398_store_0_req_1;
      array_obj_ref_398_store_0_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      StoreGroup0_gI: SplitGuardInterface generic map(name => "StoreGroup0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      addr_in <= array_obj_ref_398_word_address_0;
      data_in <= array_obj_ref_398_data_0;
      StoreReq: StoreReqSharedWithInputBuffers -- 
        generic map ( name => "StoreGroup0 Req ", addr_width => 6,
        data_width => 32,
        num_reqs => 1,
        tag_length => 3,
        time_stamp_width => 18,
        min_clock_period => false,
        input_buffering => inBUFs, 
        no_arbitration => false)
        port map (--
          reqL => reqL , 
          ackL => ackL , 
          addr => addr_in, 
          data => data_in, 
          mreq => memory_space_2_sr_req(0),
          mack => memory_space_2_sr_ack(0),
          maddr => memory_space_2_sr_addr(5 downto 0),
          mdata => memory_space_2_sr_data(31 downto 0),
          mtag => memory_space_2_sr_tag(20 downto 0),
          clk => clk, reset => reset -- 
        );--
      StoreComplete: StoreCompleteShared -- 
        generic map ( -- 
          name => "StoreGroup0 Complete ",
          num_reqs => 1,
          detailed_buffering_per_output => outBUFs,
          tag_length => 3 -- 
        )
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          mreq => memory_space_2_sc_req(0),
          mack => memory_space_2_sc_ack(0),
          mtag => memory_space_2_sc_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- store group 0
    -- 
  end Block; -- data_path
  -- 
end UpdateRegister_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.nic_system_global_package.all;
entity accessMemory is -- 
  generic (tag_length : integer); 
  port ( -- 
    lock : in  std_logic_vector(0 downto 0);
    rwbar : in  std_logic_vector(0 downto 0);
    bmask : in  std_logic_vector(7 downto 0);
    addr : in  std_logic_vector(35 downto 0);
    wdata : in  std_logic_vector(63 downto 0);
    rdata : out  std_logic_vector(63 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity accessMemory;
architecture accessMemory_arch of accessMemory is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 110)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal lock_buffer :  std_logic_vector(0 downto 0);
  signal lock_update_enable: Boolean;
  signal rwbar_buffer :  std_logic_vector(0 downto 0);
  signal rwbar_update_enable: Boolean;
  signal bmask_buffer :  std_logic_vector(7 downto 0);
  signal bmask_update_enable: Boolean;
  signal addr_buffer :  std_logic_vector(35 downto 0);
  signal addr_update_enable: Boolean;
  signal wdata_buffer :  std_logic_vector(63 downto 0);
  signal wdata_update_enable: Boolean;
  -- output port buffer signals
  signal rdata_buffer :  std_logic_vector(63 downto 0);
  signal rdata_update_enable: Boolean;
  signal accessMemory_CP_913_start: Boolean;
  signal accessMemory_CP_913_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_518_branch_ack_1 : boolean;
  signal WPIPE_NIC_TO_MEMORY_REQUEST_531_inst_ack_0 : boolean;
  signal do_while_stmt_518_branch_req_0 : boolean;
  signal WPIPE_NIC_TO_MEMORY_REQUEST_531_inst_req_0 : boolean;
  signal WPIPE_NIC_TO_MEMORY_REQUEST_531_inst_req_1 : boolean;
  signal WPIPE_NIC_TO_MEMORY_REQUEST_531_inst_ack_1 : boolean;
  signal RPIPE_MEMORY_TO_NIC_RESPONSE_535_inst_req_0 : boolean;
  signal RPIPE_MEMORY_TO_NIC_RESPONSE_535_inst_ack_0 : boolean;
  signal RPIPE_MEMORY_TO_NIC_RESPONSE_535_inst_req_1 : boolean;
  signal RPIPE_MEMORY_TO_NIC_RESPONSE_535_inst_ack_1 : boolean;
  signal do_while_stmt_518_branch_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "accessMemory_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 110) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= lock;
  lock_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(1 downto 1) <= rwbar;
  rwbar_buffer <= in_buffer_data_out(1 downto 1);
  in_buffer_data_in(9 downto 2) <= bmask;
  bmask_buffer <= in_buffer_data_out(9 downto 2);
  in_buffer_data_in(45 downto 10) <= addr;
  addr_buffer <= in_buffer_data_out(45 downto 10);
  in_buffer_data_in(109 downto 46) <= wdata;
  wdata_buffer <= in_buffer_data_out(109 downto 46);
  in_buffer_data_in(tag_length + 109 downto 110) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 109 downto 110);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  accessMemory_CP_913_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "accessMemory_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= rdata_buffer;
  rdata <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMemory_CP_913_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= accessMemory_CP_913_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessMemory_CP_913_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  accessMemory_CP_913: Block -- control-path 
    signal accessMemory_CP_913_elements: BooleanArray(20 downto 0);
    -- 
  begin -- 
    accessMemory_CP_913_elements(0) <= accessMemory_CP_913_start;
    accessMemory_CP_913_symbol <= accessMemory_CP_913_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_517/do_while_stmt_518__entry__
      -- CP-element group 0: 	 branch_block_stmt_517/branch_block_stmt_517__entry__
      -- CP-element group 0: 	 branch_block_stmt_517/$entry
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	20 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_517/do_while_stmt_518__exit__
      -- CP-element group 1: 	 branch_block_stmt_517/branch_block_stmt_517__exit__
      -- CP-element group 1: 	 branch_block_stmt_517/$exit
      -- CP-element group 1: 	 $exit
      -- 
    accessMemory_CP_913_elements(1) <= accessMemory_CP_913_elements(20);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_517/do_while_stmt_518/do_while_stmt_518__entry__
      -- CP-element group 2: 	 branch_block_stmt_517/do_while_stmt_518/$entry
      -- 
    accessMemory_CP_913_elements(2) <= accessMemory_CP_913_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	20 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_517/do_while_stmt_518/do_while_stmt_518__exit__
      -- 
    -- Element group accessMemory_CP_913_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_517/do_while_stmt_518/loop_back
      -- 
    -- Element group accessMemory_CP_913_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	18 
    -- CP-element group 5: 	19 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_517/do_while_stmt_518/condition_done
      -- CP-element group 5: 	 branch_block_stmt_517/do_while_stmt_518/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_517/do_while_stmt_518/loop_taken/$entry
      -- 
    accessMemory_CP_913_elements(5) <= accessMemory_CP_913_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	13 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_517/do_while_stmt_518/loop_body_done
      -- 
    accessMemory_CP_913_elements(6) <= accessMemory_CP_913_elements(13);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_517/do_while_stmt_518/do_while_stmt_518_loop_body/back_edge_to_loop_body
      -- 
    accessMemory_CP_913_elements(7) <= accessMemory_CP_913_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_517/do_while_stmt_518/do_while_stmt_518_loop_body/first_time_through_loop_body
      -- 
    accessMemory_CP_913_elements(8) <= accessMemory_CP_913_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	17 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	14 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_517/do_while_stmt_518/do_while_stmt_518_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_517/do_while_stmt_518/do_while_stmt_518_loop_body/loop_body_start
      -- 
    -- Element group accessMemory_CP_913_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	16 
    -- CP-element group 10: 	17 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_517/do_while_stmt_518/do_while_stmt_518_loop_body/condition_evaluated
      -- 
    condition_evaluated_937_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_937_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemory_CP_913_elements(10), ack => do_while_stmt_518_branch_req_0); -- 
    accessMemory_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "accessMemory_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemory_CP_913_elements(16) & accessMemory_CP_913_elements(17);
      gj_accessMemory_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_913_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	13 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_517/do_while_stmt_518/do_while_stmt_518_loop_body/WPIPE_NIC_TO_MEMORY_REQUEST_531_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_517/do_while_stmt_518/do_while_stmt_518_loop_body/WPIPE_NIC_TO_MEMORY_REQUEST_531_Sample/$entry
      -- CP-element group 11: 	 branch_block_stmt_517/do_while_stmt_518/do_while_stmt_518_loop_body/WPIPE_NIC_TO_MEMORY_REQUEST_531_Sample/req
      -- 
    req_946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemory_CP_913_elements(11), ack => WPIPE_NIC_TO_MEMORY_REQUEST_531_inst_req_0); -- 
    accessMemory_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "accessMemory_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemory_CP_913_elements(9) & accessMemory_CP_913_elements(13);
      gj_accessMemory_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_913_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_517/do_while_stmt_518/do_while_stmt_518_loop_body/WPIPE_NIC_TO_MEMORY_REQUEST_531_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_517/do_while_stmt_518/do_while_stmt_518_loop_body/WPIPE_NIC_TO_MEMORY_REQUEST_531_update_start_
      -- CP-element group 12: 	 branch_block_stmt_517/do_while_stmt_518/do_while_stmt_518_loop_body/WPIPE_NIC_TO_MEMORY_REQUEST_531_Sample/ack
      -- CP-element group 12: 	 branch_block_stmt_517/do_while_stmt_518/do_while_stmt_518_loop_body/WPIPE_NIC_TO_MEMORY_REQUEST_531_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_517/do_while_stmt_518/do_while_stmt_518_loop_body/WPIPE_NIC_TO_MEMORY_REQUEST_531_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_517/do_while_stmt_518/do_while_stmt_518_loop_body/WPIPE_NIC_TO_MEMORY_REQUEST_531_Update/req
      -- 
    ack_947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_TO_MEMORY_REQUEST_531_inst_ack_0, ack => accessMemory_CP_913_elements(12)); -- 
    req_951_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_951_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemory_CP_913_elements(12), ack => WPIPE_NIC_TO_MEMORY_REQUEST_531_inst_req_1); -- 
    -- CP-element group 13:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	6 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	11 
    -- CP-element group 13:  members (4) 
      -- CP-element group 13: 	 branch_block_stmt_517/do_while_stmt_518/do_while_stmt_518_loop_body/$exit
      -- CP-element group 13: 	 branch_block_stmt_517/do_while_stmt_518/do_while_stmt_518_loop_body/WPIPE_NIC_TO_MEMORY_REQUEST_531_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_517/do_while_stmt_518/do_while_stmt_518_loop_body/WPIPE_NIC_TO_MEMORY_REQUEST_531_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_517/do_while_stmt_518/do_while_stmt_518_loop_body/WPIPE_NIC_TO_MEMORY_REQUEST_531_Update/ack
      -- 
    ack_952_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NIC_TO_MEMORY_REQUEST_531_inst_ack_1, ack => accessMemory_CP_913_elements(13)); -- 
    -- CP-element group 14:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	9 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	16 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_517/do_while_stmt_518/do_while_stmt_518_loop_body/RPIPE_MEMORY_TO_NIC_RESPONSE_535_sample_start_
      -- CP-element group 14: 	 branch_block_stmt_517/do_while_stmt_518/do_while_stmt_518_loop_body/RPIPE_MEMORY_TO_NIC_RESPONSE_535_Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_517/do_while_stmt_518/do_while_stmt_518_loop_body/RPIPE_MEMORY_TO_NIC_RESPONSE_535_Sample/rr
      -- 
    rr_960_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_960_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemory_CP_913_elements(14), ack => RPIPE_MEMORY_TO_NIC_RESPONSE_535_inst_req_0); -- 
    accessMemory_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "accessMemory_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessMemory_CP_913_elements(9) & accessMemory_CP_913_elements(16);
      gj_accessMemory_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessMemory_CP_913_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	16 
    -- CP-element group 15:  members (6) 
      -- CP-element group 15: 	 branch_block_stmt_517/do_while_stmt_518/do_while_stmt_518_loop_body/RPIPE_MEMORY_TO_NIC_RESPONSE_535_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_517/do_while_stmt_518/do_while_stmt_518_loop_body/RPIPE_MEMORY_TO_NIC_RESPONSE_535_update_start_
      -- CP-element group 15: 	 branch_block_stmt_517/do_while_stmt_518/do_while_stmt_518_loop_body/RPIPE_MEMORY_TO_NIC_RESPONSE_535_Update/$entry
      -- CP-element group 15: 	 branch_block_stmt_517/do_while_stmt_518/do_while_stmt_518_loop_body/RPIPE_MEMORY_TO_NIC_RESPONSE_535_Sample/$exit
      -- CP-element group 15: 	 branch_block_stmt_517/do_while_stmt_518/do_while_stmt_518_loop_body/RPIPE_MEMORY_TO_NIC_RESPONSE_535_Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_517/do_while_stmt_518/do_while_stmt_518_loop_body/RPIPE_MEMORY_TO_NIC_RESPONSE_535_Update/cr
      -- 
    ra_961_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_MEMORY_TO_NIC_RESPONSE_535_inst_ack_0, ack => accessMemory_CP_913_elements(15)); -- 
    cr_965_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_965_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessMemory_CP_913_elements(15), ack => RPIPE_MEMORY_TO_NIC_RESPONSE_535_inst_req_1); -- 
    -- CP-element group 16:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	10 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	14 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_517/do_while_stmt_518/do_while_stmt_518_loop_body/RPIPE_MEMORY_TO_NIC_RESPONSE_535_update_completed_
      -- CP-element group 16: 	 branch_block_stmt_517/do_while_stmt_518/do_while_stmt_518_loop_body/RPIPE_MEMORY_TO_NIC_RESPONSE_535_Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_517/do_while_stmt_518/do_while_stmt_518_loop_body/RPIPE_MEMORY_TO_NIC_RESPONSE_535_Update/ca
      -- 
    ca_966_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_MEMORY_TO_NIC_RESPONSE_535_inst_ack_1, ack => accessMemory_CP_913_elements(16)); -- 
    -- CP-element group 17:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	9 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	10 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_517/do_while_stmt_518/do_while_stmt_518_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group accessMemory_CP_913_elements(17) is a control-delay.
    cp_element_17_delay: control_delay_element  generic map(name => " 17_delay", delay_value => 1)  port map(req => accessMemory_CP_913_elements(9), ack => accessMemory_CP_913_elements(17), clk => clk, reset =>reset);
    -- CP-element group 18:  transition  input  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	5 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_517/do_while_stmt_518/loop_exit/$exit
      -- CP-element group 18: 	 branch_block_stmt_517/do_while_stmt_518/loop_exit/ack
      -- 
    ack_971_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_518_branch_ack_0, ack => accessMemory_CP_913_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	5 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_517/do_while_stmt_518/loop_taken/ack
      -- CP-element group 19: 	 branch_block_stmt_517/do_while_stmt_518/loop_taken/$exit
      -- 
    ack_975_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_518_branch_ack_1, ack => accessMemory_CP_913_elements(19)); -- 
    -- CP-element group 20:  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	3 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	1 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_517/do_while_stmt_518/$exit
      -- 
    accessMemory_CP_913_elements(20) <= accessMemory_CP_913_elements(3);
    accessMemory_do_while_stmt_518_terminator_976: loop_terminator -- 
      generic map (name => " accessMemory_do_while_stmt_518_terminator_976", max_iterations_in_flight =>15) 
      port map(loop_body_exit => accessMemory_CP_913_elements(6),loop_continue => accessMemory_CP_913_elements(19),loop_terminate => accessMemory_CP_913_elements(18),loop_back => accessMemory_CP_913_elements(4),loop_exit => accessMemory_CP_913_elements(3),clk => clk, reset => reset); -- 
    entry_tmerge_938_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= accessMemory_CP_913_elements(7);
        preds(1)  <= accessMemory_CP_913_elements(8);
        entry_tmerge_938 : transition_merge -- 
          generic map(name => " entry_tmerge_938")
          port map (preds => preds, symbol_out => accessMemory_CP_913_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u1_u2_523_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u2_u10_525_wire : std_logic_vector(9 downto 0);
    signal CONCAT_u36_u100_528_wire : std_logic_vector(99 downto 0);
    signal EQ_u1_u1_554_wire : std_logic_vector(0 downto 0);
    signal err_540 : std_logic_vector(0 downto 0);
    signal konst_553_wire_constant : std_logic_vector(0 downto 0);
    signal request_530 : std_logic_vector(109 downto 0);
    signal response_536 : std_logic_vector(64 downto 0);
    -- 
  begin -- 
    konst_553_wire_constant <= "1";
    -- flow-through slice operator slice_539_inst
    err_540 <= response_536(64 downto 64);
    -- flow-through slice operator slice_543_inst
    rdata_buffer <= response_536(63 downto 0);
    do_while_stmt_518_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= EQ_u1_u1_554_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_518_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_518_branch_req_0,
          ack0 => do_while_stmt_518_branch_ack_0,
          ack1 => do_while_stmt_518_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator CONCAT_u10_u110_529_inst
    process(CONCAT_u2_u10_525_wire, CONCAT_u36_u100_528_wire) -- 
      variable tmp_var : std_logic_vector(109 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u2_u10_525_wire, CONCAT_u36_u100_528_wire, tmp_var);
      request_530 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_523_inst
    process(lock_buffer, rwbar_buffer) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(lock_buffer, rwbar_buffer, tmp_var);
      CONCAT_u1_u2_523_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u2_u10_525_inst
    process(CONCAT_u1_u2_523_wire, bmask_buffer) -- 
      variable tmp_var : std_logic_vector(9 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_523_wire, bmask_buffer, tmp_var);
      CONCAT_u2_u10_525_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u36_u100_528_inst
    process(addr_buffer, wdata_buffer) -- 
      variable tmp_var : std_logic_vector(99 downto 0); -- 
    begin -- 
      ApConcat_proc(addr_buffer, wdata_buffer, tmp_var);
      CONCAT_u36_u100_528_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_554_inst
    process(err_540) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(err_540, konst_553_wire_constant, tmp_var);
      EQ_u1_u1_554_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_MEMORY_TO_NIC_RESPONSE_535_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(64 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_MEMORY_TO_NIC_RESPONSE_535_inst_req_0;
      RPIPE_MEMORY_TO_NIC_RESPONSE_535_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_MEMORY_TO_NIC_RESPONSE_535_inst_req_1;
      RPIPE_MEMORY_TO_NIC_RESPONSE_535_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      response_536 <= data_out(64 downto 0);
      MEMORY_TO_NIC_RESPONSE_read_0_gI: SplitGuardInterface generic map(name => "MEMORY_TO_NIC_RESPONSE_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      MEMORY_TO_NIC_RESPONSE_read_0: InputPortRevised -- 
        generic map ( name => "MEMORY_TO_NIC_RESPONSE_read_0", data_width => 65,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => MEMORY_TO_NIC_RESPONSE_pipe_read_req(0),
          oack => MEMORY_TO_NIC_RESPONSE_pipe_read_ack(0),
          odata => MEMORY_TO_NIC_RESPONSE_pipe_read_data(64 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_NIC_TO_MEMORY_REQUEST_531_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_NIC_TO_MEMORY_REQUEST_531_inst_req_0;
      WPIPE_NIC_TO_MEMORY_REQUEST_531_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_NIC_TO_MEMORY_REQUEST_531_inst_req_1;
      WPIPE_NIC_TO_MEMORY_REQUEST_531_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= request_530;
      NIC_TO_MEMORY_REQUEST_write_0_gI: SplitGuardInterface generic map(name => "NIC_TO_MEMORY_REQUEST_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      NIC_TO_MEMORY_REQUEST_write_0: OutputPortRevised -- 
        generic map ( name => "NIC_TO_MEMORY_REQUEST", data_width => 110, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => NIC_TO_MEMORY_REQUEST_pipe_write_req(0),
          oack => NIC_TO_MEMORY_REQUEST_pipe_write_ack(0),
          odata => NIC_TO_MEMORY_REQUEST_pipe_write_data(109 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end accessMemory_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.nic_system_global_package.all;
entity acquireLock is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    m_ok : out  std_logic_vector(0 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity acquireLock;
architecture acquireLock_arch of acquireLock is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 1)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  -- output port buffer signals
  signal m_ok_buffer :  std_logic_vector(0 downto 0);
  signal acquireLock_CP_977_start: Boolean;
  signal acquireLock_CP_977_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_734_call_ack_0 : boolean;
  signal call_stmt_603_call_ack_0 : boolean;
  signal call_stmt_807_call_req_0 : boolean;
  signal call_stmt_734_call_req_1 : boolean;
  signal call_stmt_734_call_ack_1 : boolean;
  signal if_stmt_717_branch_req_0 : boolean;
  signal call_stmt_603_call_req_0 : boolean;
  signal call_stmt_734_call_req_0 : boolean;
  signal if_stmt_717_branch_ack_0 : boolean;
  signal call_stmt_579_call_ack_1 : boolean;
  signal call_stmt_579_call_req_1 : boolean;
  signal call_stmt_807_call_ack_1 : boolean;
  signal call_stmt_603_call_ack_1 : boolean;
  signal if_stmt_717_branch_ack_1 : boolean;
  signal call_stmt_603_call_req_1 : boolean;
  signal call_stmt_807_call_req_1 : boolean;
  signal call_stmt_579_call_ack_0 : boolean;
  signal call_stmt_579_call_req_0 : boolean;
  signal call_stmt_807_call_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "acquireLock_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  acquireLock_CP_977_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "acquireLock_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 1) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  m_ok_buffer <= "1";
  out_buffer_data_in(0 downto 0) <= m_ok_buffer;
  m_ok <= out_buffer_data_out(0 downto 0);
  out_buffer_data_in(tag_length + 0 downto 1) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 0 downto 1);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= acquireLock_CP_977_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= acquireLock_CP_977_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= acquireLock_CP_977_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  acquireLock_CP_977: Block -- control-path 
    signal acquireLock_CP_977_elements: BooleanArray(11 downto 0);
    -- 
  begin -- 
    acquireLock_CP_977_elements(0) <= acquireLock_CP_977_start;
    acquireLock_CP_977_symbol <= acquireLock_CP_977_elements(10);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	11 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 branch_block_stmt_560/assign_stmt_566/$entry
      -- CP-element group 0: 	 branch_block_stmt_560/assign_stmt_566/$exit
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_560/$entry
      -- CP-element group 0: 	 branch_block_stmt_560/branch_block_stmt_560__entry__
      -- CP-element group 0: 	 branch_block_stmt_560/assign_stmt_566__entry__
      -- CP-element group 0: 	 branch_block_stmt_560/merge_stmt_567_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_560/assign_stmt_566__exit__
      -- CP-element group 0: 	 branch_block_stmt_560/merge_stmt_567__entry__
      -- CP-element group 0: 	 branch_block_stmt_560/merge_stmt_567__entry___PhiReq/$entry
      -- CP-element group 0: 	 branch_block_stmt_560/merge_stmt_567__entry___PhiReq/$exit
      -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	11 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 branch_block_stmt_560/call_stmt_579_to_assign_stmt_716/call_stmt_579_sample_completed_
      -- CP-element group 1: 	 branch_block_stmt_560/call_stmt_579_to_assign_stmt_716/call_stmt_579_Sample/cra
      -- CP-element group 1: 	 branch_block_stmt_560/call_stmt_579_to_assign_stmt_716/call_stmt_579_Sample/$exit
      -- 
    cra_1009_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_579_call_ack_0, ack => acquireLock_CP_977_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	11 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 branch_block_stmt_560/call_stmt_579_to_assign_stmt_716/call_stmt_603_sample_start_
      -- CP-element group 2: 	 branch_block_stmt_560/call_stmt_579_to_assign_stmt_716/call_stmt_603_Sample/$entry
      -- CP-element group 2: 	 branch_block_stmt_560/call_stmt_579_to_assign_stmt_716/call_stmt_603_Sample/crr
      -- CP-element group 2: 	 branch_block_stmt_560/call_stmt_579_to_assign_stmt_716/call_stmt_579_update_completed_
      -- CP-element group 2: 	 branch_block_stmt_560/call_stmt_579_to_assign_stmt_716/call_stmt_579_Update/cca
      -- CP-element group 2: 	 branch_block_stmt_560/call_stmt_579_to_assign_stmt_716/call_stmt_579_Update/$exit
      -- 
    cca_1014_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_579_call_ack_1, ack => acquireLock_CP_977_elements(2)); -- 
    crr_1022_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1022_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireLock_CP_977_elements(2), ack => call_stmt_603_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_560/call_stmt_579_to_assign_stmt_716/call_stmt_603_Sample/cra
      -- CP-element group 3: 	 branch_block_stmt_560/call_stmt_579_to_assign_stmt_716/call_stmt_603_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_560/call_stmt_579_to_assign_stmt_716/call_stmt_603_Sample/$exit
      -- 
    cra_1023_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_603_call_ack_0, ack => acquireLock_CP_977_elements(3)); -- 
    -- CP-element group 4:  branch  transition  place  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	11 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4: 	6 
    -- CP-element group 4:  members (27) 
      -- CP-element group 4: 	 branch_block_stmt_560/if_stmt_717_dead_link/$entry
      -- CP-element group 4: 	 branch_block_stmt_560/call_stmt_579_to_assign_stmt_716__exit__
      -- CP-element group 4: 	 branch_block_stmt_560/if_stmt_717_eval_test/EQ_u8_u1_722/$entry
      -- CP-element group 4: 	 branch_block_stmt_560/if_stmt_717_eval_test/$entry
      -- CP-element group 4: 	 branch_block_stmt_560/if_stmt_717_eval_test/$exit
      -- CP-element group 4: 	 branch_block_stmt_560/call_stmt_579_to_assign_stmt_716/$exit
      -- CP-element group 4: 	 branch_block_stmt_560/if_stmt_717_eval_test/EQ_u8_u1_722/$exit
      -- CP-element group 4: 	 branch_block_stmt_560/if_stmt_717_eval_test/EQ_u8_u1_722/EQ_u8_u1_722_inputs/$entry
      -- CP-element group 4: 	 branch_block_stmt_560/if_stmt_717_eval_test/EQ_u8_u1_722/SplitProtocol/Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_560/if_stmt_717_eval_test/EQ_u8_u1_722/EQ_u8_u1_722_inputs/$exit
      -- CP-element group 4: 	 branch_block_stmt_560/if_stmt_717_eval_test/EQ_u8_u1_722/SplitProtocol/Update/cr
      -- CP-element group 4: 	 branch_block_stmt_560/if_stmt_717_eval_test/EQ_u8_u1_722/SplitProtocol/$entry
      -- CP-element group 4: 	 branch_block_stmt_560/if_stmt_717_eval_test/EQ_u8_u1_722/SplitProtocol/$exit
      -- CP-element group 4: 	 branch_block_stmt_560/if_stmt_717_eval_test/EQ_u8_u1_722/SplitProtocol/Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_560/if_stmt_717_eval_test/branch_req
      -- CP-element group 4: 	 branch_block_stmt_560/if_stmt_717_eval_test/EQ_u8_u1_722/SplitProtocol/Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_560/if_stmt_717_eval_test/EQ_u8_u1_722/SplitProtocol/Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_560/call_stmt_579_to_assign_stmt_716/call_stmt_603_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_560/if_stmt_717_eval_test/EQ_u8_u1_722/SplitProtocol/Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_560/EQ_u8_u1_722_place
      -- CP-element group 4: 	 branch_block_stmt_560/if_stmt_717__entry__
      -- CP-element group 4: 	 branch_block_stmt_560/if_stmt_717_eval_test/EQ_u8_u1_722/SplitProtocol/Update/ca
      -- CP-element group 4: 	 branch_block_stmt_560/if_stmt_717_else_link/$entry
      -- CP-element group 4: 	 branch_block_stmt_560/call_stmt_579_to_assign_stmt_716/call_stmt_603_Update/cca
      -- CP-element group 4: 	 branch_block_stmt_560/if_stmt_717_eval_test/EQ_u8_u1_722/SplitProtocol/Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_560/call_stmt_579_to_assign_stmt_716/call_stmt_603_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_560/if_stmt_717_if_link/$entry
      -- 
    cca_1028_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_603_call_ack_1, ack => acquireLock_CP_977_elements(4)); -- 
    branch_req_1055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_1055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireLock_CP_977_elements(4), ack => if_stmt_717_branch_req_0); -- 
    -- CP-element group 5:  fork  transition  place  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	7 
    -- CP-element group 5: 	8 
    -- CP-element group 5:  members (10) 
      -- CP-element group 5: 	 branch_block_stmt_560/call_stmt_734__entry__
      -- CP-element group 5: 	 branch_block_stmt_560/call_stmt_734/call_stmt_734_Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_560/call_stmt_734/call_stmt_734_Update/ccr
      -- CP-element group 5: 	 branch_block_stmt_560/call_stmt_734/call_stmt_734_Sample/crr
      -- CP-element group 5: 	 branch_block_stmt_560/call_stmt_734/call_stmt_734_Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_560/call_stmt_734/call_stmt_734_update_start_
      -- CP-element group 5: 	 branch_block_stmt_560/call_stmt_734/call_stmt_734_sample_start_
      -- CP-element group 5: 	 branch_block_stmt_560/if_stmt_717_if_link/if_choice_transition
      -- CP-element group 5: 	 branch_block_stmt_560/call_stmt_734/$entry
      -- CP-element group 5: 	 branch_block_stmt_560/if_stmt_717_if_link/$exit
      -- 
    if_choice_transition_1060_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_717_branch_ack_1, ack => acquireLock_CP_977_elements(5)); -- 
    ccr_1083_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1083_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireLock_CP_977_elements(5), ack => call_stmt_734_call_req_1); -- 
    crr_1078_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1078_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireLock_CP_977_elements(5), ack => call_stmt_734_call_req_0); -- 
    -- CP-element group 6:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	4 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6: 	10 
    -- CP-element group 6:  members (11) 
      -- CP-element group 6: 	 branch_block_stmt_560/if_stmt_717__exit__
      -- CP-element group 6: 	 branch_block_stmt_560/assign_stmt_793_to_call_stmt_807/call_stmt_807_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_560/assign_stmt_793_to_call_stmt_807__entry__
      -- CP-element group 6: 	 branch_block_stmt_560/assign_stmt_793_to_call_stmt_807/call_stmt_807_Sample/crr
      -- CP-element group 6: 	 branch_block_stmt_560/assign_stmt_793_to_call_stmt_807/call_stmt_807_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_560/assign_stmt_793_to_call_stmt_807/call_stmt_807_update_start_
      -- CP-element group 6: 	 branch_block_stmt_560/assign_stmt_793_to_call_stmt_807/$entry
      -- CP-element group 6: 	 branch_block_stmt_560/if_stmt_717_else_link/else_choice_transition
      -- CP-element group 6: 	 branch_block_stmt_560/if_stmt_717_else_link/$exit
      -- CP-element group 6: 	 branch_block_stmt_560/assign_stmt_793_to_call_stmt_807/call_stmt_807_Update/ccr
      -- CP-element group 6: 	 branch_block_stmt_560/assign_stmt_793_to_call_stmt_807/call_stmt_807_Update/$entry
      -- 
    else_choice_transition_1064_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_717_branch_ack_0, ack => acquireLock_CP_977_elements(6)); -- 
    crr_1095_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1095_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireLock_CP_977_elements(6), ack => call_stmt_807_call_req_0); -- 
    ccr_1100_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1100_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireLock_CP_977_elements(6), ack => call_stmt_807_call_req_1); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	5 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_560/call_stmt_734/call_stmt_734_Sample/cra
      -- CP-element group 7: 	 branch_block_stmt_560/call_stmt_734/call_stmt_734_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_560/call_stmt_734/call_stmt_734_sample_completed_
      -- 
    cra_1079_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_734_call_ack_0, ack => acquireLock_CP_977_elements(7)); -- 
    -- CP-element group 8:  transition  place  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	5 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	11 
    -- CP-element group 8:  members (8) 
      -- CP-element group 8: 	 branch_block_stmt_560/loopback_PhiReq/$exit
      -- CP-element group 8: 	 branch_block_stmt_560/call_stmt_734__exit__
      -- CP-element group 8: 	 branch_block_stmt_560/call_stmt_734/call_stmt_734_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_560/call_stmt_734/call_stmt_734_Update/cca
      -- CP-element group 8: 	 branch_block_stmt_560/call_stmt_734/call_stmt_734_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_560/call_stmt_734/$exit
      -- CP-element group 8: 	 branch_block_stmt_560/loopback
      -- CP-element group 8: 	 branch_block_stmt_560/loopback_PhiReq/$entry
      -- 
    cca_1084_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_734_call_ack_1, ack => acquireLock_CP_977_elements(8)); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_560/assign_stmt_793_to_call_stmt_807/call_stmt_807_Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_560/assign_stmt_793_to_call_stmt_807/call_stmt_807_sample_completed_
      -- CP-element group 9: 	 branch_block_stmt_560/assign_stmt_793_to_call_stmt_807/call_stmt_807_Sample/cra
      -- 
    cra_1096_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_807_call_ack_0, ack => acquireLock_CP_977_elements(9)); -- 
    -- CP-element group 10:  transition  place  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	6 
    -- CP-element group 10: successors 
    -- CP-element group 10:  members (10) 
      -- CP-element group 10: 	 assign_stmt_812/$entry
      -- CP-element group 10: 	 branch_block_stmt_560/assign_stmt_793_to_call_stmt_807/call_stmt_807_update_completed_
      -- CP-element group 10: 	 branch_block_stmt_560/assign_stmt_793_to_call_stmt_807/$exit
      -- CP-element group 10: 	 assign_stmt_812/$exit
      -- CP-element group 10: 	 $exit
      -- CP-element group 10: 	 branch_block_stmt_560/$exit
      -- CP-element group 10: 	 branch_block_stmt_560/branch_block_stmt_560__exit__
      -- CP-element group 10: 	 branch_block_stmt_560/assign_stmt_793_to_call_stmt_807__exit__
      -- CP-element group 10: 	 branch_block_stmt_560/assign_stmt_793_to_call_stmt_807/call_stmt_807_Update/cca
      -- CP-element group 10: 	 branch_block_stmt_560/assign_stmt_793_to_call_stmt_807/call_stmt_807_Update/$exit
      -- 
    cca_1101_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_807_call_ack_1, ack => acquireLock_CP_977_elements(10)); -- 
    -- CP-element group 11:  merge  fork  transition  place  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	8 
    -- CP-element group 11: 	0 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	4 
    -- CP-element group 11: 	1 
    -- CP-element group 11: 	2 
    -- CP-element group 11:  members (16) 
      -- CP-element group 11: 	 branch_block_stmt_560/merge_stmt_567_PhiReqMerge
      -- CP-element group 11: 	 branch_block_stmt_560/call_stmt_579_to_assign_stmt_716__entry__
      -- CP-element group 11: 	 branch_block_stmt_560/call_stmt_579_to_assign_stmt_716/$entry
      -- CP-element group 11: 	 branch_block_stmt_560/merge_stmt_567_PhiAck/$exit
      -- CP-element group 11: 	 branch_block_stmt_560/merge_stmt_567_PhiAck/dummy
      -- CP-element group 11: 	 branch_block_stmt_560/call_stmt_579_to_assign_stmt_716/call_stmt_579_sample_start_
      -- CP-element group 11: 	 branch_block_stmt_560/merge_stmt_567__exit__
      -- CP-element group 11: 	 branch_block_stmt_560/call_stmt_579_to_assign_stmt_716/call_stmt_603_update_start_
      -- CP-element group 11: 	 branch_block_stmt_560/call_stmt_579_to_assign_stmt_716/call_stmt_579_update_start_
      -- CP-element group 11: 	 branch_block_stmt_560/merge_stmt_567_PhiAck/$entry
      -- CP-element group 11: 	 branch_block_stmt_560/call_stmt_579_to_assign_stmt_716/call_stmt_579_Update/ccr
      -- CP-element group 11: 	 branch_block_stmt_560/call_stmt_579_to_assign_stmt_716/call_stmt_579_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_560/call_stmt_579_to_assign_stmt_716/call_stmt_603_Update/ccr
      -- CP-element group 11: 	 branch_block_stmt_560/call_stmt_579_to_assign_stmt_716/call_stmt_603_Update/$entry
      -- CP-element group 11: 	 branch_block_stmt_560/call_stmt_579_to_assign_stmt_716/call_stmt_579_Sample/crr
      -- CP-element group 11: 	 branch_block_stmt_560/call_stmt_579_to_assign_stmt_716/call_stmt_579_Sample/$entry
      -- 
    ccr_1013_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1013_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireLock_CP_977_elements(11), ack => call_stmt_579_call_req_1); -- 
    ccr_1027_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1027_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireLock_CP_977_elements(11), ack => call_stmt_603_call_req_1); -- 
    crr_1008_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1008_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => acquireLock_CP_977_elements(11), ack => call_stmt_579_call_req_0); -- 
    acquireLock_CP_977_elements(11) <= OrReduce(acquireLock_CP_977_elements(8) & acquireLock_CP_977_elements(0));
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u1_u2_750_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_763_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_777_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_790_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u2_u4_764_wire : std_logic_vector(3 downto 0);
    signal CONCAT_u2_u4_791_wire : std_logic_vector(3 downto 0);
    signal CONCAT_u4_u36_599_wire : std_logic_vector(35 downto 0);
    signal CONCAT_u4_u36_802_wire : std_logic_vector(35 downto 0);
    signal EQ_u8_u1_722_wire : std_logic_vector(0 downto 0);
    signal MUX_680_wire : std_logic_vector(7 downto 0);
    signal MUX_684_wire : std_logic_vector(7 downto 0);
    signal MUX_689_wire : std_logic_vector(7 downto 0);
    signal MUX_693_wire : std_logic_vector(7 downto 0);
    signal MUX_699_wire : std_logic_vector(7 downto 0);
    signal MUX_703_wire : std_logic_vector(7 downto 0);
    signal MUX_708_wire : std_logic_vector(7 downto 0);
    signal MUX_712_wire : std_logic_vector(7 downto 0);
    signal MUX_743_wire : std_logic_vector(0 downto 0);
    signal MUX_749_wire : std_logic_vector(0 downto 0);
    signal MUX_756_wire : std_logic_vector(0 downto 0);
    signal MUX_762_wire : std_logic_vector(0 downto 0);
    signal MUX_770_wire : std_logic_vector(0 downto 0);
    signal MUX_776_wire : std_logic_vector(0 downto 0);
    signal MUX_783_wire : std_logic_vector(0 downto 0);
    signal MUX_789_wire : std_logic_vector(0 downto 0);
    signal NOT_u64_u64_805_wire_constant : std_logic_vector(63 downto 0);
    signal NOT_u8_u8_574_wire_constant : std_logic_vector(7 downto 0);
    signal NOT_u8_u8_595_wire_constant : std_logic_vector(7 downto 0);
    signal NOT_u8_u8_721_wire_constant : std_logic_vector(7 downto 0);
    signal NOT_u8_u8_729_wire_constant : std_logic_vector(7 downto 0);
    signal OR_u8_u8_685_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_694_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_695_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_704_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_713_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_714_wire : std_logic_vector(7 downto 0);
    signal err_734 : std_logic_vector(63 downto 0);
    signal ignore_807 : std_logic_vector(63 downto 0);
    signal konst_638_wire_constant : std_logic_vector(2 downto 0);
    signal konst_643_wire_constant : std_logic_vector(2 downto 0);
    signal konst_648_wire_constant : std_logic_vector(2 downto 0);
    signal konst_653_wire_constant : std_logic_vector(2 downto 0);
    signal konst_658_wire_constant : std_logic_vector(2 downto 0);
    signal konst_663_wire_constant : std_logic_vector(2 downto 0);
    signal konst_668_wire_constant : std_logic_vector(2 downto 0);
    signal konst_673_wire_constant : std_logic_vector(2 downto 0);
    signal konst_679_wire_constant : std_logic_vector(7 downto 0);
    signal konst_683_wire_constant : std_logic_vector(7 downto 0);
    signal konst_688_wire_constant : std_logic_vector(7 downto 0);
    signal konst_692_wire_constant : std_logic_vector(7 downto 0);
    signal konst_698_wire_constant : std_logic_vector(7 downto 0);
    signal konst_702_wire_constant : std_logic_vector(7 downto 0);
    signal konst_707_wire_constant : std_logic_vector(7 downto 0);
    signal konst_711_wire_constant : std_logic_vector(7 downto 0);
    signal l0_607 : std_logic_vector(7 downto 0);
    signal l1_611 : std_logic_vector(7 downto 0);
    signal l2_615 : std_logic_vector(7 downto 0);
    signal l3_619 : std_logic_vector(7 downto 0);
    signal l4_623 : std_logic_vector(7 downto 0);
    signal l5_627 : std_logic_vector(7 downto 0);
    signal l6_631 : std_logic_vector(7 downto 0);
    signal l7_635 : std_logic_vector(7 downto 0);
    signal lock_addr_32_583 : std_logic_vector(31 downto 0);
    signal lock_address_pointer_566 : std_logic_vector(35 downto 0);
    signal lock_val_716 : std_logic_vector(7 downto 0);
    signal lock_values_603 : std_logic_vector(63 downto 0);
    signal msg_size_plus_lock_579 : std_logic_vector(63 downto 0);
    signal new_bmask_793 : std_logic_vector(7 downto 0);
    signal s0_640 : std_logic_vector(0 downto 0);
    signal s1_645 : std_logic_vector(0 downto 0);
    signal s2_650 : std_logic_vector(0 downto 0);
    signal s3_655 : std_logic_vector(0 downto 0);
    signal s4_660 : std_logic_vector(0 downto 0);
    signal s5_665 : std_logic_vector(0 downto 0);
    signal s6_670 : std_logic_vector(0 downto 0);
    signal s7_675 : std_logic_vector(0 downto 0);
    signal sel_588 : std_logic_vector(2 downto 0);
    signal type_cast_564_wire_constant : std_logic_vector(35 downto 0);
    signal type_cast_569_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_571_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_577_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_590_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_592_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_597_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_601_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_724_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_726_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_732_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_740_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_742_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_746_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_748_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_753_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_755_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_759_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_761_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_767_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_769_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_773_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_775_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_780_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_782_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_786_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_788_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_795_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_797_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_800_wire_constant : std_logic_vector(3 downto 0);
    -- 
  begin -- 
    NOT_u64_u64_805_wire_constant <= "1111111111111111111111111111111111111111111111111111111111111111";
    NOT_u8_u8_574_wire_constant <= "11111111";
    NOT_u8_u8_595_wire_constant <= "11111111";
    NOT_u8_u8_721_wire_constant <= "11111111";
    NOT_u8_u8_729_wire_constant <= "11111111";
    konst_638_wire_constant <= "000";
    konst_643_wire_constant <= "001";
    konst_648_wire_constant <= "010";
    konst_653_wire_constant <= "011";
    konst_658_wire_constant <= "100";
    konst_663_wire_constant <= "101";
    konst_668_wire_constant <= "110";
    konst_673_wire_constant <= "111";
    konst_679_wire_constant <= "00000000";
    konst_683_wire_constant <= "00000000";
    konst_688_wire_constant <= "00000000";
    konst_692_wire_constant <= "00000000";
    konst_698_wire_constant <= "00000000";
    konst_702_wire_constant <= "00000000";
    konst_707_wire_constant <= "00000000";
    konst_711_wire_constant <= "00000000";
    type_cast_564_wire_constant <= "000000000000000000000000000000010000";
    type_cast_569_wire_constant <= "1";
    type_cast_571_wire_constant <= "1";
    type_cast_577_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_590_wire_constant <= "1";
    type_cast_592_wire_constant <= "1";
    type_cast_597_wire_constant <= "0000";
    type_cast_601_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_724_wire_constant <= "0";
    type_cast_726_wire_constant <= "1";
    type_cast_732_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_740_wire_constant <= "1";
    type_cast_742_wire_constant <= "0";
    type_cast_746_wire_constant <= "1";
    type_cast_748_wire_constant <= "0";
    type_cast_753_wire_constant <= "1";
    type_cast_755_wire_constant <= "0";
    type_cast_759_wire_constant <= "1";
    type_cast_761_wire_constant <= "0";
    type_cast_767_wire_constant <= "1";
    type_cast_769_wire_constant <= "0";
    type_cast_773_wire_constant <= "1";
    type_cast_775_wire_constant <= "0";
    type_cast_780_wire_constant <= "1";
    type_cast_782_wire_constant <= "0";
    type_cast_786_wire_constant <= "1";
    type_cast_788_wire_constant <= "0";
    type_cast_795_wire_constant <= "0";
    type_cast_797_wire_constant <= "0";
    type_cast_800_wire_constant <= "0000";
    -- flow-through select operator MUX_680_inst
    MUX_680_wire <= l0_607 when (s0_640(0) /=  '0') else konst_679_wire_constant;
    -- flow-through select operator MUX_684_inst
    MUX_684_wire <= l1_611 when (s1_645(0) /=  '0') else konst_683_wire_constant;
    -- flow-through select operator MUX_689_inst
    MUX_689_wire <= l2_615 when (s2_650(0) /=  '0') else konst_688_wire_constant;
    -- flow-through select operator MUX_693_inst
    MUX_693_wire <= l3_619 when (s3_655(0) /=  '0') else konst_692_wire_constant;
    -- flow-through select operator MUX_699_inst
    MUX_699_wire <= l4_623 when (s4_660(0) /=  '0') else konst_698_wire_constant;
    -- flow-through select operator MUX_703_inst
    MUX_703_wire <= l5_627 when (s5_665(0) /=  '0') else konst_702_wire_constant;
    -- flow-through select operator MUX_708_inst
    MUX_708_wire <= l6_631 when (s6_670(0) /=  '0') else konst_707_wire_constant;
    -- flow-through select operator MUX_712_inst
    MUX_712_wire <= l7_635 when (s7_675(0) /=  '0') else konst_711_wire_constant;
    -- flow-through select operator MUX_743_inst
    MUX_743_wire <= type_cast_740_wire_constant when (s0_640(0) /=  '0') else type_cast_742_wire_constant;
    -- flow-through select operator MUX_749_inst
    MUX_749_wire <= type_cast_746_wire_constant when (s1_645(0) /=  '0') else type_cast_748_wire_constant;
    -- flow-through select operator MUX_756_inst
    MUX_756_wire <= type_cast_753_wire_constant when (s2_650(0) /=  '0') else type_cast_755_wire_constant;
    -- flow-through select operator MUX_762_inst
    MUX_762_wire <= type_cast_759_wire_constant when (s3_655(0) /=  '0') else type_cast_761_wire_constant;
    -- flow-through select operator MUX_770_inst
    MUX_770_wire <= type_cast_767_wire_constant when (s4_660(0) /=  '0') else type_cast_769_wire_constant;
    -- flow-through select operator MUX_776_inst
    MUX_776_wire <= type_cast_773_wire_constant when (s5_665(0) /=  '0') else type_cast_775_wire_constant;
    -- flow-through select operator MUX_783_inst
    MUX_783_wire <= type_cast_780_wire_constant when (s6_670(0) /=  '0') else type_cast_782_wire_constant;
    -- flow-through select operator MUX_789_inst
    MUX_789_wire <= type_cast_786_wire_constant when (s7_675(0) /=  '0') else type_cast_788_wire_constant;
    -- flow-through slice operator slice_582_inst
    lock_addr_32_583 <= msg_size_plus_lock_579(31 downto 0);
    -- flow-through slice operator slice_587_inst
    sel_588 <= lock_addr_32_583(2 downto 0);
    -- flow-through slice operator slice_606_inst
    l0_607 <= lock_values_603(63 downto 56);
    -- flow-through slice operator slice_610_inst
    l1_611 <= lock_values_603(55 downto 48);
    -- flow-through slice operator slice_614_inst
    l2_615 <= lock_values_603(47 downto 40);
    -- flow-through slice operator slice_618_inst
    l3_619 <= lock_values_603(39 downto 32);
    -- flow-through slice operator slice_622_inst
    l4_623 <= lock_values_603(31 downto 24);
    -- flow-through slice operator slice_626_inst
    l5_627 <= lock_values_603(23 downto 16);
    -- flow-through slice operator slice_630_inst
    l6_631 <= lock_values_603(15 downto 8);
    -- flow-through slice operator slice_634_inst
    l7_635 <= lock_values_603(7 downto 0);
    if_stmt_717_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= EQ_u8_u1_722_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_717_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_717_branch_req_0,
          ack0 => if_stmt_717_branch_ack_0,
          ack1 => if_stmt_717_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u36_u36_565_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, type_cast_564_wire_constant, tmp_var);
      lock_address_pointer_566 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_750_inst
    process(MUX_743_wire, MUX_749_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_743_wire, MUX_749_wire, tmp_var);
      CONCAT_u1_u2_750_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_763_inst
    process(MUX_756_wire, MUX_762_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_756_wire, MUX_762_wire, tmp_var);
      CONCAT_u1_u2_763_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_777_inst
    process(MUX_770_wire, MUX_776_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_770_wire, MUX_776_wire, tmp_var);
      CONCAT_u1_u2_777_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_790_inst
    process(MUX_783_wire, MUX_789_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_783_wire, MUX_789_wire, tmp_var);
      CONCAT_u1_u2_790_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u2_u4_764_inst
    process(CONCAT_u1_u2_750_wire, CONCAT_u1_u2_763_wire) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_750_wire, CONCAT_u1_u2_763_wire, tmp_var);
      CONCAT_u2_u4_764_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u2_u4_791_inst
    process(CONCAT_u1_u2_777_wire, CONCAT_u1_u2_790_wire) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_777_wire, CONCAT_u1_u2_790_wire, tmp_var);
      CONCAT_u2_u4_791_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u4_u36_599_inst
    process(type_cast_597_wire_constant, lock_addr_32_583) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_597_wire_constant, lock_addr_32_583, tmp_var);
      CONCAT_u4_u36_599_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u4_u36_802_inst
    process(type_cast_800_wire_constant, lock_addr_32_583) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_800_wire_constant, lock_addr_32_583, tmp_var);
      CONCAT_u4_u36_802_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u4_u8_792_inst
    process(CONCAT_u2_u4_764_wire, CONCAT_u2_u4_791_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u2_u4_764_wire, CONCAT_u2_u4_791_wire, tmp_var);
      new_bmask_793 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_639_inst
    process(sel_588) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_588, konst_638_wire_constant, tmp_var);
      s0_640 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_644_inst
    process(sel_588) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_588, konst_643_wire_constant, tmp_var);
      s1_645 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_649_inst
    process(sel_588) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_588, konst_648_wire_constant, tmp_var);
      s2_650 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_654_inst
    process(sel_588) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_588, konst_653_wire_constant, tmp_var);
      s3_655 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_659_inst
    process(sel_588) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_588, konst_658_wire_constant, tmp_var);
      s4_660 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_664_inst
    process(sel_588) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_588, konst_663_wire_constant, tmp_var);
      s5_665 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_669_inst
    process(sel_588) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_588, konst_668_wire_constant, tmp_var);
      s6_670 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_674_inst
    process(sel_588) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_588, konst_673_wire_constant, tmp_var);
      s7_675 <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_722_inst
    process(lock_val_716) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(lock_val_716, NOT_u8_u8_721_wire_constant, tmp_var);
      EQ_u8_u1_722_wire <= tmp_var; --
    end process;
    -- binary operator OR_u8_u8_685_inst
    process(MUX_680_wire, MUX_684_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_680_wire, MUX_684_wire, tmp_var);
      OR_u8_u8_685_wire <= tmp_var; --
    end process;
    -- binary operator OR_u8_u8_694_inst
    process(MUX_689_wire, MUX_693_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_689_wire, MUX_693_wire, tmp_var);
      OR_u8_u8_694_wire <= tmp_var; --
    end process;
    -- binary operator OR_u8_u8_695_inst
    process(OR_u8_u8_685_wire, OR_u8_u8_694_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u8_u8_685_wire, OR_u8_u8_694_wire, tmp_var);
      OR_u8_u8_695_wire <= tmp_var; --
    end process;
    -- binary operator OR_u8_u8_704_inst
    process(MUX_699_wire, MUX_703_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_699_wire, MUX_703_wire, tmp_var);
      OR_u8_u8_704_wire <= tmp_var; --
    end process;
    -- binary operator OR_u8_u8_713_inst
    process(MUX_708_wire, MUX_712_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_708_wire, MUX_712_wire, tmp_var);
      OR_u8_u8_713_wire <= tmp_var; --
    end process;
    -- binary operator OR_u8_u8_714_inst
    process(OR_u8_u8_704_wire, OR_u8_u8_713_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u8_u8_704_wire, OR_u8_u8_713_wire, tmp_var);
      OR_u8_u8_714_wire <= tmp_var; --
    end process;
    -- binary operator OR_u8_u8_715_inst
    process(OR_u8_u8_695_wire, OR_u8_u8_714_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u8_u8_695_wire, OR_u8_u8_714_wire, tmp_var);
      lock_val_716 <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_579_call call_stmt_603_call call_stmt_734_call call_stmt_807_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(439 downto 0);
      signal data_out: std_logic_vector(255 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 3 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 3 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 3 downto 0);
      signal guard_vector : std_logic_vector( 3 downto 0);
      constant inBUFs : IntegerArray(3 downto 0) := (3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(3 downto 0) := (3 => 1, 2 => 1, 1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(3 downto 0) := (0 => false, 1 => false, 2 => false, 3 => false);
      constant guardBuffering: IntegerArray(3 downto 0)  := (0 => 2, 1 => 2, 2 => 2, 3 => 2);
      -- 
    begin -- 
      reqL_unguarded(3) <= call_stmt_579_call_req_0;
      reqL_unguarded(2) <= call_stmt_603_call_req_0;
      reqL_unguarded(1) <= call_stmt_734_call_req_0;
      reqL_unguarded(0) <= call_stmt_807_call_req_0;
      call_stmt_579_call_ack_0 <= ackL_unguarded(3);
      call_stmt_603_call_ack_0 <= ackL_unguarded(2);
      call_stmt_734_call_ack_0 <= ackL_unguarded(1);
      call_stmt_807_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(3) <= call_stmt_579_call_req_1;
      reqR_unguarded(2) <= call_stmt_603_call_req_1;
      reqR_unguarded(1) <= call_stmt_734_call_req_1;
      reqR_unguarded(0) <= call_stmt_807_call_req_1;
      call_stmt_579_call_ack_1 <= ackR_unguarded(3);
      call_stmt_603_call_ack_1 <= ackR_unguarded(2);
      call_stmt_734_call_ack_1 <= ackR_unguarded(1);
      call_stmt_807_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      guard_vector(2)  <=  '1';
      guard_vector(3)  <=  '1';
      accessMemory_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_accessRegulator_2: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_2", num_slots => 1) -- 
        port map (req => reqL_unregulated(2), -- 
          ack => ackL_unregulated(2),
          regulated_req => reqL(2),
          regulated_ack => ackL(2),
          release_req => reqR(2),
          release_ack => ackR(2),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_accessRegulator_3: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_3", num_slots => 1) -- 
        port map (req => reqL_unregulated(3), -- 
          ack => ackL_unregulated(3),
          regulated_req => reqL(3),
          regulated_ack => ackL(3),
          release_req => reqR(3),
          release_ack => ackR(3),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 4, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_569_wire_constant & type_cast_571_wire_constant & NOT_u8_u8_574_wire_constant & lock_address_pointer_566 & type_cast_577_wire_constant & type_cast_590_wire_constant & type_cast_592_wire_constant & NOT_u8_u8_595_wire_constant & CONCAT_u4_u36_599_wire & type_cast_601_wire_constant & type_cast_724_wire_constant & type_cast_726_wire_constant & NOT_u8_u8_729_wire_constant & lock_address_pointer_566 & type_cast_732_wire_constant & type_cast_795_wire_constant & type_cast_797_wire_constant & new_bmask_793 & CONCAT_u4_u36_802_wire & NOT_u64_u64_805_wire_constant;
      msg_size_plus_lock_579 <= data_out(255 downto 192);
      lock_values_603 <= data_out(191 downto 128);
      err_734 <= data_out(127 downto 64);
      ignore_807 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 440,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 4,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 256,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 4) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end acquireLock_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.nic_system_global_package.all;
entity delay_time_Operator is -- 
  port ( -- 
    sample_req: in boolean;
    sample_ack: out boolean;
    update_req: in boolean;
    update_ack: out boolean;
    T : in  std_logic_vector(31 downto 0);
    delay_done : out  std_logic_vector(0 downto 0);
    clk, reset: in std_logic
    -- 
  );
  -- 
end entity delay_time_Operator;
architecture delay_time_Operator_arch of delay_time_Operator is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal update_ack_symbol: Boolean;
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal T_buffer :  std_logic_vector(31 downto 0);
  signal T_update_enable: Boolean;
  signal T_update_enable_unmarked: Boolean;
  -- output port buffer signals
  signal delay_done_buffer :  std_logic_vector(0 downto 0);
  signal delay_time_CP_2100_start: Boolean;
  signal delay_time_CP_2100_symbol: Boolean;
  signal cp_all_inputs_sampled: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal do_while_stmt_1610_branch_req_0 : boolean;
  signal phi_stmt_1612_req_0 : boolean;
  signal phi_stmt_1612_req_1 : boolean;
  signal phi_stmt_1612_ack_0 : boolean;
  signal nR_1621_1614_buf_req_0 : boolean;
  signal nR_1621_1614_buf_ack_0 : boolean;
  signal nR_1621_1614_buf_req_1 : boolean;
  signal nR_1621_1614_buf_ack_1 : boolean;
  signal T_1615_buf_req_0 : boolean;
  signal T_1615_buf_ack_0 : boolean;
  signal T_1615_buf_req_1 : boolean;
  signal T_1615_buf_ack_1 : boolean;
  signal do_while_stmt_1610_branch_ack_0 : boolean;
  signal do_while_stmt_1610_branch_ack_1 : boolean;
  -- 
begin --  
  sample_ack <= delay_time_CP_2100_symbol;
  -- input handling ------------------------------------------------
  T_buffer <= T;
  -- join of sample-req and update-req.. used to trigger CP.
  delay_time_CP_2100_start_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
    constant joinName: string(1 to 29) := "delay_time_CP_2100_start_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= sample_req & update_req;
    gj_delay_time_CP_2100_start_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => delay_time_CP_2100_start, clk => clk, reset => reset); --
  end block;
  -- output handling  -------------------------------------------------------
  delay_done_buffer <= "1";
  delay_done <= delay_done_buffer;
  update_ack_symbol <= delay_time_CP_2100_symbol;
  update_ack <= update_ack_symbol;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  delay_time_CP_2100: Block -- control-path 
    signal delay_time_CP_2100_elements: BooleanArray(32 downto 0);
    -- 
  begin -- 
    delay_time_CP_2100_elements(0) <= delay_time_CP_2100_start;
    delay_time_CP_2100_symbol <= delay_time_CP_2100_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1609/$entry
      -- CP-element group 0: 	 branch_block_stmt_1609/branch_block_stmt_1609__entry__
      -- CP-element group 0: 	 branch_block_stmt_1609/do_while_stmt_1610__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	32 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (8) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1609/$exit
      -- CP-element group 1: 	 branch_block_stmt_1609/branch_block_stmt_1609__exit__
      -- CP-element group 1: 	 branch_block_stmt_1609/do_while_stmt_1610__exit__
      -- CP-element group 1: 	 branch_block_stmt_1609/assign_stmt_1628__entry__
      -- CP-element group 1: 	 branch_block_stmt_1609/assign_stmt_1628__exit__
      -- CP-element group 1: 	 branch_block_stmt_1609/assign_stmt_1628/$entry
      -- CP-element group 1: 	 branch_block_stmt_1609/assign_stmt_1628/$exit
      -- 
    delay_time_CP_2100_elements(1) <= delay_time_CP_2100_elements(32);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1609/do_while_stmt_1610/$entry
      -- CP-element group 2: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610__entry__
      -- 
    delay_time_CP_2100_elements(2) <= delay_time_CP_2100_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	32 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610__exit__
      -- 
    -- Element group delay_time_CP_2100_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1609/do_while_stmt_1610/loop_back
      -- 
    -- Element group delay_time_CP_2100_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	30 
    -- CP-element group 5: 	31 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1609/do_while_stmt_1610/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1609/do_while_stmt_1610/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1609/do_while_stmt_1610/loop_taken/$entry
      -- 
    delay_time_CP_2100_elements(5) <= delay_time_CP_2100_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	14 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1609/do_while_stmt_1610/loop_body_done
      -- 
    delay_time_CP_2100_elements(6) <= delay_time_CP_2100_elements(14);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	16 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/back_edge_to_loop_body
      -- 
    delay_time_CP_2100_elements(7) <= delay_time_CP_2100_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	18 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/first_time_through_loop_body
      -- 
    delay_time_CP_2100_elements(8) <= delay_time_CP_2100_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9: 	13 
    -- CP-element group 9: 	29 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/loop_body_start
      -- 
    -- Element group delay_time_CP_2100_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	29 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/condition_evaluated
      -- 
    condition_evaluated_2126_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2126_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_2100_elements(10), ack => do_while_stmt_1610_branch_req_0); -- 
    delay_time_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "delay_time_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= delay_time_CP_2100_elements(15) & delay_time_CP_2100_elements(29);
      gj_delay_time_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => delay_time_CP_2100_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/phi_stmt_1612_sample_start__ps
      -- 
    delay_time_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "delay_time_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= delay_time_CP_2100_elements(12) & delay_time_CP_2100_elements(15);
      gj_delay_time_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => delay_time_CP_2100_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	11 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/phi_stmt_1612_sample_start_
      -- 
    delay_time_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "delay_time_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= delay_time_CP_2100_elements(9) & delay_time_CP_2100_elements(14);
      gj_delay_time_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => delay_time_CP_2100_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	9 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	15 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/phi_stmt_1612_update_start_
      -- CP-element group 13: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/phi_stmt_1612_update_start__ps
      -- 
    delay_time_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "delay_time_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= delay_time_CP_2100_elements(9) & delay_time_CP_2100_elements(15);
      gj_delay_time_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => delay_time_CP_2100_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	6 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (4) 
      -- CP-element group 14: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/$exit
      -- CP-element group 14: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/aggregated_phi_sample_ack
      -- CP-element group 14: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/phi_stmt_1612_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/phi_stmt_1612_sample_completed__ps
      -- 
    -- Element group delay_time_CP_2100_elements(14) is bound as output of CP function.
    -- CP-element group 15:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15: 	13 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/aggregated_phi_update_ack
      -- CP-element group 15: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/phi_stmt_1612_update_completed_
      -- CP-element group 15: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/phi_stmt_1612_update_completed__ps
      -- 
    -- Element group delay_time_CP_2100_elements(15) is bound as output of CP function.
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	7 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/phi_stmt_1612_loopback_trigger
      -- 
    delay_time_CP_2100_elements(16) <= delay_time_CP_2100_elements(7);
    -- CP-element group 17:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/phi_stmt_1612_loopback_sample_req
      -- CP-element group 17: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/phi_stmt_1612_loopback_sample_req_ps
      -- 
    phi_stmt_1612_loopback_sample_req_2141_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1612_loopback_sample_req_2141_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_2100_elements(17), ack => phi_stmt_1612_req_0); -- 
    -- Element group delay_time_CP_2100_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	8 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/phi_stmt_1612_entry_trigger
      -- 
    delay_time_CP_2100_elements(18) <= delay_time_CP_2100_elements(8);
    -- CP-element group 19:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/phi_stmt_1612_entry_sample_req
      -- CP-element group 19: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/phi_stmt_1612_entry_sample_req_ps
      -- 
    phi_stmt_1612_entry_sample_req_2144_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1612_entry_sample_req_2144_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_2100_elements(19), ack => phi_stmt_1612_req_1); -- 
    -- Element group delay_time_CP_2100_elements(19) is bound as output of CP function.
    -- CP-element group 20:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/phi_stmt_1612_phi_mux_ack
      -- CP-element group 20: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/phi_stmt_1612_phi_mux_ack_ps
      -- 
    phi_stmt_1612_phi_mux_ack_2147_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1612_ack_0, ack => delay_time_CP_2100_elements(20)); -- 
    -- CP-element group 21:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (4) 
      -- CP-element group 21: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/R_nR_1614_sample_start__ps
      -- CP-element group 21: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/R_nR_1614_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/R_nR_1614_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/R_nR_1614_Sample/req
      -- 
    req_2160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_2100_elements(21), ack => nR_1621_1614_buf_req_0); -- 
    -- Element group delay_time_CP_2100_elements(21) is bound as output of CP function.
    -- CP-element group 22:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (4) 
      -- CP-element group 22: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/R_nR_1614_update_start__ps
      -- CP-element group 22: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/R_nR_1614_update_start_
      -- CP-element group 22: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/R_nR_1614_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/R_nR_1614_Update/req
      -- 
    req_2165_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2165_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_2100_elements(22), ack => nR_1621_1614_buf_req_1); -- 
    -- Element group delay_time_CP_2100_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (4) 
      -- CP-element group 23: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/R_nR_1614_sample_completed__ps
      -- CP-element group 23: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/R_nR_1614_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/R_nR_1614_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/R_nR_1614_Sample/ack
      -- 
    ack_2161_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nR_1621_1614_buf_ack_0, ack => delay_time_CP_2100_elements(23)); -- 
    -- CP-element group 24:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/R_nR_1614_update_completed__ps
      -- CP-element group 24: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/R_nR_1614_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/R_nR_1614_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/R_nR_1614_Update/ack
      -- 
    ack_2166_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nR_1621_1614_buf_ack_1, ack => delay_time_CP_2100_elements(24)); -- 
    -- CP-element group 25:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/R_T_1615_sample_start__ps
      -- CP-element group 25: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/R_T_1615_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/R_T_1615_Sample/$entry
      -- CP-element group 25: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/R_T_1615_Sample/req
      -- 
    req_2178_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2178_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_2100_elements(25), ack => T_1615_buf_req_0); -- 
    -- Element group delay_time_CP_2100_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/R_T_1615_update_start__ps
      -- CP-element group 26: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/R_T_1615_update_start_
      -- CP-element group 26: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/R_T_1615_Update/$entry
      -- CP-element group 26: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/R_T_1615_Update/req
      -- 
    req_2183_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2183_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => delay_time_CP_2100_elements(26), ack => T_1615_buf_req_1); -- 
    -- Element group delay_time_CP_2100_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/R_T_1615_sample_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/R_T_1615_sample_completed_
      -- CP-element group 27: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/R_T_1615_Sample/$exit
      -- CP-element group 27: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/R_T_1615_Sample/ack
      -- 
    ack_2179_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => T_1615_buf_ack_0, ack => delay_time_CP_2100_elements(27)); -- 
    -- CP-element group 28:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/R_T_1615_update_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/R_T_1615_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/R_T_1615_Update/$exit
      -- CP-element group 28: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/R_T_1615_Update/ack
      -- 
    ack_2184_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 28_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => T_1615_buf_ack_1, ack => delay_time_CP_2100_elements(28)); -- 
    -- CP-element group 29:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	9 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	10 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_1609/do_while_stmt_1610/do_while_stmt_1610_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group delay_time_CP_2100_elements(29) is a control-delay.
    cp_element_29_delay: control_delay_element  generic map(name => " 29_delay", delay_value => 1)  port map(req => delay_time_CP_2100_elements(9), ack => delay_time_CP_2100_elements(29), clk => clk, reset =>reset);
    -- CP-element group 30:  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	5 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_1609/do_while_stmt_1610/loop_exit/$exit
      -- CP-element group 30: 	 branch_block_stmt_1609/do_while_stmt_1610/loop_exit/ack
      -- 
    ack_2190_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1610_branch_ack_0, ack => delay_time_CP_2100_elements(30)); -- 
    -- CP-element group 31:  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	5 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (2) 
      -- CP-element group 31: 	 branch_block_stmt_1609/do_while_stmt_1610/loop_taken/$exit
      -- CP-element group 31: 	 branch_block_stmt_1609/do_while_stmt_1610/loop_taken/ack
      -- 
    ack_2194_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1610_branch_ack_1, ack => delay_time_CP_2100_elements(31)); -- 
    -- CP-element group 32:  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	3 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	1 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_1609/do_while_stmt_1610/$exit
      -- 
    delay_time_CP_2100_elements(32) <= delay_time_CP_2100_elements(3);
    delay_time_do_while_stmt_1610_terminator_2195: loop_terminator -- 
      generic map (name => " delay_time_do_while_stmt_1610_terminator_2195", max_iterations_in_flight =>7) 
      port map(loop_body_exit => delay_time_CP_2100_elements(6),loop_continue => delay_time_CP_2100_elements(31),loop_terminate => delay_time_CP_2100_elements(30),loop_back => delay_time_CP_2100_elements(4),loop_exit => delay_time_CP_2100_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1612_phi_seq_2185_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= delay_time_CP_2100_elements(16);
      delay_time_CP_2100_elements(21)<= src_sample_reqs(0);
      src_sample_acks(0)  <= delay_time_CP_2100_elements(23);
      delay_time_CP_2100_elements(22)<= src_update_reqs(0);
      src_update_acks(0)  <= delay_time_CP_2100_elements(24);
      delay_time_CP_2100_elements(17) <= phi_mux_reqs(0);
      triggers(1)  <= delay_time_CP_2100_elements(18);
      delay_time_CP_2100_elements(25)<= src_sample_reqs(1);
      src_sample_acks(1)  <= delay_time_CP_2100_elements(27);
      delay_time_CP_2100_elements(26)<= src_update_reqs(1);
      src_update_acks(1)  <= delay_time_CP_2100_elements(28);
      delay_time_CP_2100_elements(19) <= phi_mux_reqs(1);
      phi_stmt_1612_phi_seq_2185 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_1612_phi_seq_2185") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => delay_time_CP_2100_elements(11), 
          phi_sample_ack => delay_time_CP_2100_elements(14), 
          phi_update_req => delay_time_CP_2100_elements(13), 
          phi_update_ack => delay_time_CP_2100_elements(15), 
          phi_mux_ack => delay_time_CP_2100_elements(20), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_2127_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= delay_time_CP_2100_elements(7);
        preds(1)  <= delay_time_CP_2100_elements(8);
        entry_tmerge_2127 : transition_merge -- 
          generic map(name => " entry_tmerge_2127")
          port map (preds => preds, symbol_out => delay_time_CP_2100_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal R_1612 : std_logic_vector(31 downto 0);
    signal T_1615_buffered : std_logic_vector(31 downto 0);
    signal UGT_u32_u1_1625_wire : std_logic_vector(0 downto 0);
    signal konst_1619_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1624_wire_constant : std_logic_vector(31 downto 0);
    signal nR_1621 : std_logic_vector(31 downto 0);
    signal nR_1621_1614_buffered : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    konst_1619_wire_constant <= "00000000000000000000000000000001";
    konst_1624_wire_constant <= "00000000000000000000000000000000";
    phi_stmt_1612: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nR_1621_1614_buffered & T_1615_buffered;
      req <= phi_stmt_1612_req_0 & phi_stmt_1612_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1612",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1612_ack_0,
          idata => idata,
          odata => R_1612,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1612
    T_1615_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= T_1615_buf_req_0;
      T_1615_buf_ack_0<= wack(0);
      rreq(0) <= T_1615_buf_req_1;
      T_1615_buf_ack_1<= rack(0);
      T_1615_buf : InterlockBuffer generic map ( -- 
        name => "T_1615_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => T_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => T_1615_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nR_1621_1614_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nR_1621_1614_buf_req_0;
      nR_1621_1614_buf_ack_0<= wack(0);
      rreq(0) <= nR_1621_1614_buf_req_1;
      nR_1621_1614_buf_ack_1<= rack(0);
      nR_1621_1614_buf : InterlockBuffer generic map ( -- 
        name => "nR_1621_1614_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nR_1621,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nR_1621_1614_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_1610_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= UGT_u32_u1_1625_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1610_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1610_branch_req_0,
          ack0 => do_while_stmt_1610_branch_ack_0,
          ack1 => do_while_stmt_1610_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator SUB_u32_u32_1620_inst
    process(R_1612) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(R_1612, konst_1619_wire_constant, tmp_var);
      nR_1621 <= tmp_var; --
    end process;
    -- binary operator UGT_u32_u1_1625_inst
    process(R_1612) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(R_1612, konst_1624_wire_constant, tmp_var);
      UGT_u32_u1_1625_wire <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end delay_time_Operator_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.nic_system_global_package.all;
entity getQueueElement is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    read_index : in  std_logic_vector(31 downto 0);
    q_r_data : out  std_logic_vector(31 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity getQueueElement;
architecture getQueueElement_arch of getQueueElement is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 68)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  signal read_index_buffer :  std_logic_vector(31 downto 0);
  signal read_index_update_enable: Boolean;
  -- output port buffer signals
  signal q_r_data_buffer :  std_logic_vector(31 downto 0);
  signal q_r_data_update_enable: Boolean;
  signal getQueueElement_CP_1222_start: Boolean;
  signal getQueueElement_CP_1222_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_932_call_ack_0 : boolean;
  signal MUX_947_inst_req_1 : boolean;
  signal call_stmt_932_call_req_0 : boolean;
  signal MUX_947_inst_ack_0 : boolean;
  signal MUX_947_inst_req_0 : boolean;
  signal MUX_947_inst_ack_1 : boolean;
  signal call_stmt_932_call_req_1 : boolean;
  signal call_stmt_932_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "getQueueElement_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 68) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(67 downto 36) <= read_index;
  read_index_buffer <= in_buffer_data_out(67 downto 36);
  in_buffer_data_in(tag_length + 67 downto 68) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 67 downto 68);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  getQueueElement_CP_1222_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "getQueueElement_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= q_r_data_buffer;
  q_r_data <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueueElement_CP_1222_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= getQueueElement_CP_1222_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueueElement_CP_1222_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  getQueueElement_CP_1222: Block -- control-path 
    signal getQueueElement_CP_1222_elements: BooleanArray(4 downto 0);
    -- 
  begin -- 
    getQueueElement_CP_1222_elements(0) <= getQueueElement_CP_1222_start;
    getQueueElement_CP_1222_symbol <= getQueueElement_CP_1222_elements(4);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 assign_stmt_908_to_assign_stmt_948/call_stmt_932_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_908_to_assign_stmt_948/call_stmt_932_update_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_908_to_assign_stmt_948/MUX_947_complete/req
      -- CP-element group 0: 	 assign_stmt_908_to_assign_stmt_948/call_stmt_932_Update/$entry
      -- CP-element group 0: 	 assign_stmt_908_to_assign_stmt_948/call_stmt_932_sample_start_
      -- CP-element group 0: 	 assign_stmt_908_to_assign_stmt_948/call_stmt_932_Sample/crr
      -- CP-element group 0: 	 assign_stmt_908_to_assign_stmt_948/$entry
      -- CP-element group 0: 	 assign_stmt_908_to_assign_stmt_948/MUX_947_update_start_
      -- CP-element group 0: 	 assign_stmt_908_to_assign_stmt_948/MUX_947_complete/$entry
      -- CP-element group 0: 	 assign_stmt_908_to_assign_stmt_948/call_stmt_932_Update/ccr
      -- 
    crr_1235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueElement_CP_1222_elements(0), ack => call_stmt_932_call_req_0); -- 
    ccr_1240_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1240_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueElement_CP_1222_elements(0), ack => call_stmt_932_call_req_1); -- 
    req_1254_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1254_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueElement_CP_1222_elements(0), ack => MUX_947_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_908_to_assign_stmt_948/call_stmt_932_sample_completed_
      -- CP-element group 1: 	 assign_stmt_908_to_assign_stmt_948/call_stmt_932_Sample/cra
      -- CP-element group 1: 	 assign_stmt_908_to_assign_stmt_948/call_stmt_932_Sample/$exit
      -- 
    cra_1236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_932_call_ack_0, ack => getQueueElement_CP_1222_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 assign_stmt_908_to_assign_stmt_948/call_stmt_932_update_completed_
      -- CP-element group 2: 	 assign_stmt_908_to_assign_stmt_948/call_stmt_932_Update/$exit
      -- CP-element group 2: 	 assign_stmt_908_to_assign_stmt_948/MUX_947_start/req
      -- CP-element group 2: 	 assign_stmt_908_to_assign_stmt_948/MUX_947_start/$entry
      -- CP-element group 2: 	 assign_stmt_908_to_assign_stmt_948/call_stmt_932_Update/cca
      -- CP-element group 2: 	 assign_stmt_908_to_assign_stmt_948/MUX_947_sample_start_
      -- 
    cca_1241_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_932_call_ack_1, ack => getQueueElement_CP_1222_elements(2)); -- 
    req_1249_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1249_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueElement_CP_1222_elements(2), ack => MUX_947_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_908_to_assign_stmt_948/MUX_947_sample_completed_
      -- CP-element group 3: 	 assign_stmt_908_to_assign_stmt_948/MUX_947_start/ack
      -- CP-element group 3: 	 assign_stmt_908_to_assign_stmt_948/MUX_947_start/$exit
      -- 
    ack_1250_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_947_inst_ack_0, ack => getQueueElement_CP_1222_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 assign_stmt_908_to_assign_stmt_948/MUX_947_update_completed_
      -- CP-element group 4: 	 assign_stmt_908_to_assign_stmt_948/$exit
      -- CP-element group 4: 	 $exit
      -- CP-element group 4: 	 assign_stmt_908_to_assign_stmt_948/MUX_947_complete/$exit
      -- CP-element group 4: 	 assign_stmt_908_to_assign_stmt_948/MUX_947_complete/ack
      -- 
    ack_1255_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_947_inst_ack_1, ack => getQueueElement_CP_1222_elements(4)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u32_u1_944_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u31_u34_916_wire : std_logic_vector(33 downto 0);
    signal NOT_u8_u8_927_wire_constant : std_logic_vector(7 downto 0);
    signal buffer_address_908 : std_logic_vector(35 downto 0);
    signal e0_936 : std_logic_vector(31 downto 0);
    signal e1_940 : std_logic_vector(31 downto 0);
    signal element_pair_932 : std_logic_vector(63 downto 0);
    signal element_pair_address_920 : std_logic_vector(35 downto 0);
    signal konst_943_wire_constant : std_logic_vector(31 downto 0);
    signal slice_913_wire : std_logic_vector(30 downto 0);
    signal type_cast_906_wire_constant : std_logic_vector(35 downto 0);
    signal type_cast_915_wire_constant : std_logic_vector(2 downto 0);
    signal type_cast_918_wire : std_logic_vector(35 downto 0);
    signal type_cast_922_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_924_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_930_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    NOT_u8_u8_927_wire_constant <= "11111111";
    konst_943_wire_constant <= "00000000000000000000000000000000";
    type_cast_906_wire_constant <= "000000000000000000000000000000100000";
    type_cast_915_wire_constant <= "000";
    type_cast_922_wire_constant <= "0";
    type_cast_924_wire_constant <= "1";
    type_cast_930_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    MUX_947_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= MUX_947_inst_req_0;
      MUX_947_inst_ack_0<= sample_ack(0);
      update_req(0) <= MUX_947_inst_req_1;
      MUX_947_inst_ack_1<= update_ack(0);
      MUX_947_inst: SelectSplitProtocol generic map(name => "MUX_947_inst", data_width => 32, buffering => 1, flow_through => false, full_rate => false) -- 
        port map( x => e1_940, y => e0_936, sel => BITSEL_u32_u1_944_wire, z => q_r_data_buffer, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through slice operator slice_913_inst
    slice_913_wire <= read_index_buffer(31 downto 1);
    -- flow-through slice operator slice_935_inst
    e0_936 <= element_pair_932(63 downto 32);
    -- flow-through slice operator slice_939_inst
    e1_940 <= element_pair_932(31 downto 0);
    -- interlock type_cast_918_inst
    process(CONCAT_u31_u34_916_wire) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 33 downto 0) := CONCAT_u31_u34_916_wire(33 downto 0);
      type_cast_918_wire <= tmp_var; -- 
    end process;
    -- binary operator ADD_u36_u36_907_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, type_cast_906_wire_constant, tmp_var);
      buffer_address_908 <= tmp_var; --
    end process;
    -- binary operator ADD_u36_u36_919_inst
    process(buffer_address_908, type_cast_918_wire) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(buffer_address_908, type_cast_918_wire, tmp_var);
      element_pair_address_920 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_944_inst
    process(read_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(read_index_buffer, konst_943_wire_constant, tmp_var);
      BITSEL_u32_u1_944_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u31_u34_916_inst
    process(slice_913_wire) -- 
      variable tmp_var : std_logic_vector(33 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_913_wire, type_cast_915_wire_constant, tmp_var);
      CONCAT_u31_u34_916_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_932_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_932_call_req_0;
      call_stmt_932_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_932_call_req_1;
      call_stmt_932_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_922_wire_constant & type_cast_924_wire_constant & NOT_u8_u8_927_wire_constant & element_pair_address_920 & type_cast_930_wire_constant;
      element_pair_932 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end getQueueElement_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.nic_system_global_package.all;
entity getQueueLength is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    Queue_Length : out  std_logic_vector(31 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity getQueueLength;
architecture getQueueLength_arch of getQueueLength is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  -- output port buffer signals
  signal Queue_Length_buffer :  std_logic_vector(31 downto 0);
  signal Queue_Length_update_enable: Boolean;
  signal getQueueLength_CP_1154_start: Boolean;
  signal getQueueLength_CP_1154_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_873_call_ack_1 : boolean;
  signal call_stmt_873_call_req_1 : boolean;
  signal slice_876_inst_req_1 : boolean;
  signal slice_876_inst_ack_1 : boolean;
  signal call_stmt_873_call_req_0 : boolean;
  signal call_stmt_873_call_ack_0 : boolean;
  signal slice_876_inst_req_0 : boolean;
  signal slice_876_inst_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "getQueueLength_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  getQueueLength_CP_1154_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "getQueueLength_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= Queue_Length_buffer;
  Queue_Length <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueueLength_CP_1154_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= getQueueLength_CP_1154_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueueLength_CP_1154_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  getQueueLength_CP_1154: Block -- control-path 
    signal getQueueLength_CP_1154_elements: BooleanArray(4 downto 0);
    -- 
  begin -- 
    getQueueLength_CP_1154_elements(0) <= getQueueLength_CP_1154_start;
    getQueueLength_CP_1154_symbol <= getQueueLength_CP_1154_elements(4);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 call_stmt_873_to_assign_stmt_877/call_stmt_873_Sample/$entry
      -- CP-element group 0: 	 call_stmt_873_to_assign_stmt_877/call_stmt_873_Update/ccr
      -- CP-element group 0: 	 call_stmt_873_to_assign_stmt_877/slice_876_update_start_
      -- CP-element group 0: 	 call_stmt_873_to_assign_stmt_877/call_stmt_873_Update/$entry
      -- CP-element group 0: 	 call_stmt_873_to_assign_stmt_877/slice_876_Update/cr
      -- CP-element group 0: 	 call_stmt_873_to_assign_stmt_877/call_stmt_873_Sample/crr
      -- CP-element group 0: 	 call_stmt_873_to_assign_stmt_877/slice_876_Update/$entry
      -- CP-element group 0: 	 call_stmt_873_to_assign_stmt_877/call_stmt_873_update_start_
      -- CP-element group 0: 	 call_stmt_873_to_assign_stmt_877/call_stmt_873_sample_start_
      -- CP-element group 0: 	 call_stmt_873_to_assign_stmt_877/$entry
      -- CP-element group 0: 	 $entry
      -- 
    cr_1186_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1186_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueLength_CP_1154_elements(0), ack => slice_876_inst_req_1); -- 
    crr_1167_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1167_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueLength_CP_1154_elements(0), ack => call_stmt_873_call_req_0); -- 
    ccr_1172_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1172_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueLength_CP_1154_elements(0), ack => call_stmt_873_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_873_to_assign_stmt_877/call_stmt_873_Sample/$exit
      -- CP-element group 1: 	 call_stmt_873_to_assign_stmt_877/call_stmt_873_Sample/cra
      -- CP-element group 1: 	 call_stmt_873_to_assign_stmt_877/call_stmt_873_sample_completed_
      -- 
    cra_1168_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_873_call_ack_0, ack => getQueueLength_CP_1154_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 call_stmt_873_to_assign_stmt_877/call_stmt_873_Update/$exit
      -- CP-element group 2: 	 call_stmt_873_to_assign_stmt_877/call_stmt_873_Update/cca
      -- CP-element group 2: 	 call_stmt_873_to_assign_stmt_877/slice_876_sample_start_
      -- CP-element group 2: 	 call_stmt_873_to_assign_stmt_877/slice_876_Sample/$entry
      -- CP-element group 2: 	 call_stmt_873_to_assign_stmt_877/slice_876_Sample/rr
      -- CP-element group 2: 	 call_stmt_873_to_assign_stmt_877/call_stmt_873_update_completed_
      -- 
    cca_1173_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_873_call_ack_1, ack => getQueueLength_CP_1154_elements(2)); -- 
    rr_1181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueueLength_CP_1154_elements(2), ack => slice_876_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 call_stmt_873_to_assign_stmt_877/slice_876_sample_completed_
      -- CP-element group 3: 	 call_stmt_873_to_assign_stmt_877/slice_876_Sample/$exit
      -- CP-element group 3: 	 call_stmt_873_to_assign_stmt_877/slice_876_Sample/ra
      -- 
    ra_1182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_876_inst_ack_0, ack => getQueueLength_CP_1154_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 call_stmt_873_to_assign_stmt_877/slice_876_Update/$exit
      -- CP-element group 4: 	 call_stmt_873_to_assign_stmt_877/slice_876_Update/ca
      -- CP-element group 4: 	 call_stmt_873_to_assign_stmt_877/slice_876_update_completed_
      -- CP-element group 4: 	 call_stmt_873_to_assign_stmt_877/$exit
      -- CP-element group 4: 	 $exit
      -- 
    ca_1187_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_876_inst_ack_1, ack => getQueueLength_CP_1154_elements(4)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u36_u36_869_wire : std_logic_vector(35 downto 0);
    signal NOT_u8_u8_866_wire_constant : std_logic_vector(7 downto 0);
    signal konst_868_wire_constant : std_logic_vector(35 downto 0);
    signal type_cast_861_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_863_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_871_wire_constant : std_logic_vector(63 downto 0);
    signal wi_and_len_873 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    NOT_u8_u8_866_wire_constant <= "11111111";
    konst_868_wire_constant <= "000000000000000000000000000000001000";
    type_cast_861_wire_constant <= "0";
    type_cast_863_wire_constant <= "1";
    type_cast_871_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    slice_876_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_876_inst_req_0;
      slice_876_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_876_inst_req_1;
      slice_876_inst_ack_1<= update_ack(0);
      slice_876_inst: SliceSplitProtocol generic map(name => "slice_876_inst", in_data_width => 64, high_index => 31, low_index => 0, buffering => 1, flow_through => false,  full_rate => false) -- 
        port map( din => wi_and_len_873, dout => Queue_Length_buffer, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- binary operator ADD_u36_u36_869_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, konst_868_wire_constant, tmp_var);
      ADD_u36_u36_869_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_873_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_873_call_req_0;
      call_stmt_873_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_873_call_req_1;
      call_stmt_873_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_861_wire_constant & type_cast_863_wire_constant & NOT_u8_u8_866_wire_constant & ADD_u36_u36_869_wire & type_cast_871_wire_constant;
      wi_and_len_873 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end getQueueLength_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.nic_system_global_package.all;
entity getQueuePointers is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    wp : out  std_logic_vector(31 downto 0);
    rp : out  std_logic_vector(31 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity getQueuePointers;
architecture getQueuePointers_arch of getQueuePointers is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  -- output port buffer signals
  signal wp_buffer :  std_logic_vector(31 downto 0);
  signal wp_update_enable: Boolean;
  signal rp_buffer :  std_logic_vector(31 downto 0);
  signal rp_update_enable: Boolean;
  signal getQueuePointers_CP_1120_start: Boolean;
  signal getQueuePointers_CP_1120_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_829_call_req_0 : boolean;
  signal call_stmt_829_call_ack_0 : boolean;
  signal call_stmt_829_call_req_1 : boolean;
  signal call_stmt_829_call_ack_1 : boolean;
  signal call_stmt_843_call_req_0 : boolean;
  signal call_stmt_843_call_ack_0 : boolean;
  signal call_stmt_843_call_req_1 : boolean;
  signal call_stmt_843_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "getQueuePointers_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  getQueuePointers_CP_1120_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "getQueuePointers_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= wp_buffer;
  wp <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(63 downto 32) <= rp_buffer;
  rp <= out_buffer_data_out(63 downto 32);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueuePointers_CP_1120_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= getQueuePointers_CP_1120_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getQueuePointers_CP_1120_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  getQueuePointers_CP_1120: Block -- control-path 
    signal getQueuePointers_CP_1120_elements: BooleanArray(4 downto 0);
    -- 
  begin -- 
    getQueuePointers_CP_1120_elements(0) <= getQueuePointers_CP_1120_start;
    getQueuePointers_CP_1120_symbol <= getQueuePointers_CP_1120_elements(4);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_829_to_assign_stmt_851/$entry
      -- CP-element group 0: 	 call_stmt_829_to_assign_stmt_851/call_stmt_829_sample_start_
      -- CP-element group 0: 	 call_stmt_829_to_assign_stmt_851/call_stmt_829_update_start_
      -- CP-element group 0: 	 call_stmt_829_to_assign_stmt_851/call_stmt_829_Sample/$entry
      -- CP-element group 0: 	 call_stmt_829_to_assign_stmt_851/call_stmt_829_Sample/crr
      -- CP-element group 0: 	 call_stmt_829_to_assign_stmt_851/call_stmt_829_Update/$entry
      -- CP-element group 0: 	 call_stmt_829_to_assign_stmt_851/call_stmt_829_Update/ccr
      -- CP-element group 0: 	 call_stmt_829_to_assign_stmt_851/call_stmt_843_update_start_
      -- CP-element group 0: 	 call_stmt_829_to_assign_stmt_851/call_stmt_843_Update/$entry
      -- CP-element group 0: 	 call_stmt_829_to_assign_stmt_851/call_stmt_843_Update/ccr
      -- 
    crr_1133_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1133_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueuePointers_CP_1120_elements(0), ack => call_stmt_829_call_req_0); -- 
    ccr_1138_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1138_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueuePointers_CP_1120_elements(0), ack => call_stmt_829_call_req_1); -- 
    ccr_1152_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1152_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueuePointers_CP_1120_elements(0), ack => call_stmt_843_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_829_to_assign_stmt_851/call_stmt_829_sample_completed_
      -- CP-element group 1: 	 call_stmt_829_to_assign_stmt_851/call_stmt_829_Sample/$exit
      -- CP-element group 1: 	 call_stmt_829_to_assign_stmt_851/call_stmt_829_Sample/cra
      -- 
    cra_1134_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_829_call_ack_0, ack => getQueuePointers_CP_1120_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 call_stmt_829_to_assign_stmt_851/call_stmt_829_update_completed_
      -- CP-element group 2: 	 call_stmt_829_to_assign_stmt_851/call_stmt_829_Update/$exit
      -- CP-element group 2: 	 call_stmt_829_to_assign_stmt_851/call_stmt_829_Update/cca
      -- CP-element group 2: 	 call_stmt_829_to_assign_stmt_851/call_stmt_843_sample_start_
      -- CP-element group 2: 	 call_stmt_829_to_assign_stmt_851/call_stmt_843_Sample/$entry
      -- CP-element group 2: 	 call_stmt_829_to_assign_stmt_851/call_stmt_843_Sample/crr
      -- 
    cca_1139_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_829_call_ack_1, ack => getQueuePointers_CP_1120_elements(2)); -- 
    crr_1147_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1147_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getQueuePointers_CP_1120_elements(2), ack => call_stmt_843_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 call_stmt_829_to_assign_stmt_851/call_stmt_843_sample_completed_
      -- CP-element group 3: 	 call_stmt_829_to_assign_stmt_851/call_stmt_843_Sample/$exit
      -- CP-element group 3: 	 call_stmt_829_to_assign_stmt_851/call_stmt_843_Sample/cra
      -- 
    cra_1148_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_843_call_ack_0, ack => getQueuePointers_CP_1120_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 $exit
      -- CP-element group 4: 	 call_stmt_829_to_assign_stmt_851/$exit
      -- CP-element group 4: 	 call_stmt_829_to_assign_stmt_851/call_stmt_843_update_completed_
      -- CP-element group 4: 	 call_stmt_829_to_assign_stmt_851/call_stmt_843_Update/$exit
      -- CP-element group 4: 	 call_stmt_829_to_assign_stmt_851/call_stmt_843_Update/cca
      -- 
    cca_1153_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_843_call_ack_1, ack => getQueuePointers_CP_1120_elements(4)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u36_u36_839_wire : std_logic_vector(35 downto 0);
    signal NOT_u8_u8_824_wire_constant : std_logic_vector(7 downto 0);
    signal NOT_u8_u8_836_wire_constant : std_logic_vector(7 downto 0);
    signal konst_838_wire_constant : std_logic_vector(35 downto 0);
    signal msgs_rp_829 : std_logic_vector(63 downto 0);
    signal type_cast_819_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_821_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_827_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_831_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_833_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_841_wire_constant : std_logic_vector(63 downto 0);
    signal wp_len_843 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    NOT_u8_u8_824_wire_constant <= "11111111";
    NOT_u8_u8_836_wire_constant <= "11111111";
    konst_838_wire_constant <= "000000000000000000000000000000001000";
    type_cast_819_wire_constant <= "0";
    type_cast_821_wire_constant <= "1";
    type_cast_827_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_831_wire_constant <= "0";
    type_cast_833_wire_constant <= "1";
    type_cast_841_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    -- flow-through slice operator slice_846_inst
    rp_buffer <= msgs_rp_829(31 downto 0);
    -- flow-through slice operator slice_850_inst
    wp_buffer <= wp_len_843(63 downto 32);
    -- binary operator ADD_u36_u36_839_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, konst_838_wire_constant, tmp_var);
      ADD_u36_u36_839_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_843_call call_stmt_829_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(219 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_843_call_req_0;
      reqL_unguarded(0) <= call_stmt_829_call_req_0;
      call_stmt_843_call_ack_0 <= ackL_unguarded(1);
      call_stmt_829_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_843_call_req_1;
      reqR_unguarded(0) <= call_stmt_829_call_req_1;
      call_stmt_843_call_ack_1 <= ackR_unguarded(1);
      call_stmt_829_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      accessMemory_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_831_wire_constant & type_cast_833_wire_constant & NOT_u8_u8_836_wire_constant & ADD_u36_u36_839_wire & type_cast_841_wire_constant & type_cast_819_wire_constant & type_cast_821_wire_constant & NOT_u8_u8_824_wire_constant & q_base_address_buffer & type_cast_827_wire_constant;
      wp_len_843 <= data_out(127 downto 64);
      msgs_rp_829 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 220,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end getQueuePointers_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.nic_system_global_package.all;
entity getTotalMessages is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    total_msgs : out  std_logic_vector(31 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity getTotalMessages;
architecture getTotalMessages_arch of getTotalMessages is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  -- output port buffer signals
  signal total_msgs_buffer :  std_logic_vector(31 downto 0);
  signal total_msgs_update_enable: Boolean;
  signal getTotalMessages_CP_1188_start: Boolean;
  signal getTotalMessages_CP_1188_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal slice_896_inst_req_1 : boolean;
  signal slice_896_inst_ack_0 : boolean;
  signal slice_896_inst_ack_1 : boolean;
  signal slice_896_inst_req_0 : boolean;
  signal call_stmt_893_call_ack_1 : boolean;
  signal call_stmt_893_call_req_1 : boolean;
  signal call_stmt_893_call_ack_0 : boolean;
  signal call_stmt_893_call_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "getTotalMessages_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  getTotalMessages_CP_1188_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "getTotalMessages_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 32) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= total_msgs_buffer;
  total_msgs <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(tag_length + 31 downto 32) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 31 downto 32);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getTotalMessages_CP_1188_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= getTotalMessages_CP_1188_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getTotalMessages_CP_1188_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  getTotalMessages_CP_1188: Block -- control-path 
    signal getTotalMessages_CP_1188_elements: BooleanArray(4 downto 0);
    -- 
  begin -- 
    getTotalMessages_CP_1188_elements(0) <= getTotalMessages_CP_1188_start;
    getTotalMessages_CP_1188_symbol <= getTotalMessages_CP_1188_elements(4);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 call_stmt_893_to_assign_stmt_897/call_stmt_893_sample_start_
      -- CP-element group 0: 	 call_stmt_893_to_assign_stmt_897/$entry
      -- CP-element group 0: 	 call_stmt_893_to_assign_stmt_897/slice_896_Update/cr
      -- CP-element group 0: 	 call_stmt_893_to_assign_stmt_897/call_stmt_893_update_start_
      -- CP-element group 0: 	 call_stmt_893_to_assign_stmt_897/call_stmt_893_Sample/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_893_to_assign_stmt_897/slice_896_Update/$entry
      -- CP-element group 0: 	 call_stmt_893_to_assign_stmt_897/slice_896_update_start_
      -- CP-element group 0: 	 call_stmt_893_to_assign_stmt_897/call_stmt_893_Update/ccr
      -- CP-element group 0: 	 call_stmt_893_to_assign_stmt_897/call_stmt_893_Update/$entry
      -- CP-element group 0: 	 call_stmt_893_to_assign_stmt_897/call_stmt_893_Sample/crr
      -- 
    crr_1201_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1201_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTotalMessages_CP_1188_elements(0), ack => call_stmt_893_call_req_0); -- 
    ccr_1206_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1206_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTotalMessages_CP_1188_elements(0), ack => call_stmt_893_call_req_1); -- 
    cr_1220_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1220_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTotalMessages_CP_1188_elements(0), ack => slice_896_inst_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_893_to_assign_stmt_897/call_stmt_893_sample_completed_
      -- CP-element group 1: 	 call_stmt_893_to_assign_stmt_897/call_stmt_893_Sample/cra
      -- CP-element group 1: 	 call_stmt_893_to_assign_stmt_897/call_stmt_893_Sample/$exit
      -- 
    cra_1202_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_893_call_ack_0, ack => getTotalMessages_CP_1188_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 call_stmt_893_to_assign_stmt_897/slice_896_Sample/$entry
      -- CP-element group 2: 	 call_stmt_893_to_assign_stmt_897/call_stmt_893_update_completed_
      -- CP-element group 2: 	 call_stmt_893_to_assign_stmt_897/slice_896_Sample/rr
      -- CP-element group 2: 	 call_stmt_893_to_assign_stmt_897/slice_896_sample_start_
      -- CP-element group 2: 	 call_stmt_893_to_assign_stmt_897/call_stmt_893_Update/cca
      -- CP-element group 2: 	 call_stmt_893_to_assign_stmt_897/call_stmt_893_Update/$exit
      -- 
    cca_1207_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_893_call_ack_1, ack => getTotalMessages_CP_1188_elements(2)); -- 
    rr_1215_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1215_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTotalMessages_CP_1188_elements(2), ack => slice_896_inst_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 call_stmt_893_to_assign_stmt_897/slice_896_Sample/ra
      -- CP-element group 3: 	 call_stmt_893_to_assign_stmt_897/slice_896_Sample/$exit
      -- CP-element group 3: 	 call_stmt_893_to_assign_stmt_897/slice_896_sample_completed_
      -- 
    ra_1216_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_896_inst_ack_0, ack => getTotalMessages_CP_1188_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 call_stmt_893_to_assign_stmt_897/slice_896_Update/$exit
      -- CP-element group 4: 	 call_stmt_893_to_assign_stmt_897/$exit
      -- CP-element group 4: 	 $exit
      -- CP-element group 4: 	 call_stmt_893_to_assign_stmt_897/slice_896_Update/ca
      -- CP-element group 4: 	 call_stmt_893_to_assign_stmt_897/slice_896_update_completed_
      -- 
    ca_1221_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => slice_896_inst_ack_1, ack => getTotalMessages_CP_1188_elements(4)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal NOT_u8_u8_888_wire_constant : std_logic_vector(7 downto 0);
    signal rdata_893 : std_logic_vector(63 downto 0);
    signal type_cast_883_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_885_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_891_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    NOT_u8_u8_888_wire_constant <= "11111111";
    type_cast_883_wire_constant <= "0";
    type_cast_885_wire_constant <= "1";
    type_cast_891_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    slice_896_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= slice_896_inst_req_0;
      slice_896_inst_ack_0<= sample_ack(0);
      update_req(0) <= slice_896_inst_req_1;
      slice_896_inst_ack_1<= update_ack(0);
      slice_896_inst: SliceSplitProtocol generic map(name => "slice_896_inst", in_data_width => 64, high_index => 63, low_index => 32, buffering => 1, flow_through => false,  full_rate => false) -- 
        port map( din => rdata_893, dout => total_msgs_buffer, sample_req => sample_req(0) , sample_ack => sample_ack(0) , update_req => update_req(0) , update_ack => update_ack(0) , clk => clk, reset => reset); -- 
      -- 
    end block;
    -- shared call operator group (0) : call_stmt_893_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_893_call_req_0;
      call_stmt_893_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_893_call_req_1;
      call_stmt_893_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_883_wire_constant & type_cast_885_wire_constant & NOT_u8_u8_888_wire_constant & q_base_address_buffer & type_cast_891_wire_constant;
      rdata_893 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end getTotalMessages_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.nic_system_global_package.all;
entity getTxPacketPointerFromServer is -- 
  generic (tag_length : integer); 
  port ( -- 
    queue_index : in  std_logic_vector(5 downto 0);
    pkt_pointer : out  std_logic_vector(31 downto 0);
    status : out  std_logic_vector(0 downto 0);
    AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_call_data : out  std_logic_vector(42 downto 0);
    AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
    AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_return_data : in   std_logic_vector(31 downto 0);
    AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
    popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
    popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
    popFromQueue_call_data : out  std_logic_vector(36 downto 0);
    popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
    popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
    popFromQueue_return_data : in   std_logic_vector(32 downto 0);
    popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity getTxPacketPointerFromServer;
architecture getTxPacketPointerFromServer_arch of getTxPacketPointerFromServer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 6)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 33)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal queue_index_buffer :  std_logic_vector(5 downto 0);
  signal queue_index_update_enable: Boolean;
  -- output port buffer signals
  signal pkt_pointer_buffer :  std_logic_vector(31 downto 0);
  signal pkt_pointer_update_enable: Boolean;
  signal status_buffer :  std_logic_vector(0 downto 0);
  signal status_update_enable: Boolean;
  signal getTxPacketPointerFromServer_CP_30524_start: Boolean;
  signal getTxPacketPointerFromServer_CP_30524_symbol: Boolean;
  -- volatile/operator module components. 
  component AccessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      register_index : in  std_logic_vector(5 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component popFromQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_r_data : out  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_call_acks : in   std_logic_vector(0 downto 0);
      releaseLock_call_data : out  std_logic_vector(35 downto 0);
      releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_return_acks : in   std_logic_vector(0 downto 0);
      releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_call_acks : in   std_logic_vector(0 downto 0);
      acquireLock_call_data : out  std_logic_vector(35 downto 0);
      acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_return_acks : in   std_logic_vector(0 downto 0);
      acquireLock_return_data : in   std_logic_vector(0 downto 0);
      acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      updateTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_data : out  std_logic_vector(67 downto 0);
      updateTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_call_data : out  std_logic_vector(67 downto 0);
      getQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_return_data : in   std_logic_vector(31 downto 0);
      getQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_call_data : out  std_logic_vector(35 downto 0);
      getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
      getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_call_data : out  std_logic_vector(35 downto 0);
      getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_return_data : in   std_logic_vector(31 downto 0);
      getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_15844_call_req_0 : boolean;
  signal call_stmt_15844_call_ack_0 : boolean;
  signal call_stmt_15832_call_ack_1 : boolean;
  signal call_stmt_15832_call_req_1 : boolean;
  signal call_stmt_15832_call_ack_0 : boolean;
  signal call_stmt_15832_call_req_0 : boolean;
  signal call_stmt_15844_call_ack_1 : boolean;
  signal call_stmt_15844_call_req_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "getTxPacketPointerFromServer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 6) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(5 downto 0) <= queue_index;
  queue_index_buffer <= in_buffer_data_out(5 downto 0);
  in_buffer_data_in(tag_length + 5 downto 6) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 5 downto 6);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 7);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= queue_index_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  getTxPacketPointerFromServer_CP_30524_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "getTxPacketPointerFromServer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 33) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= pkt_pointer_buffer;
  pkt_pointer <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(32 downto 32) <= status_buffer;
  status <= out_buffer_data_out(32 downto 32);
  out_buffer_data_in(tag_length + 32 downto 33) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 32 downto 33);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getTxPacketPointerFromServer_CP_30524_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  pkt_pointer_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 30) := "pkt_pointer_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_pkt_pointer_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => pkt_pointer_update_enable, clk => clk, reset => reset); --
  end block;
  status_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 25) := "status_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_status_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => status_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 7,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= getTxPacketPointerFromServer_CP_30524_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= getTxPacketPointerFromServer_CP_30524_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  getTxPacketPointerFromServer_CP_30524: Block -- control-path 
    signal getTxPacketPointerFromServer_CP_30524_elements: BooleanArray(16 downto 0);
    -- 
  begin -- 
    getTxPacketPointerFromServer_CP_30524_elements(0) <= getTxPacketPointerFromServer_CP_30524_start;
    getTxPacketPointerFromServer_CP_30524_symbol <= getTxPacketPointerFromServer_CP_30524_elements(16);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	5 
    -- CP-element group 1:  members (1) 
      -- CP-element group 1: 	 assign_stmt_15822_to_stmt_15849/$entry
      -- 
    getTxPacketPointerFromServer_CP_30524_elements(1) <= getTxPacketPointerFromServer_CP_30524_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	7 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	13 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_15822_to_stmt_15849/queue_index_update_enable
      -- CP-element group 2: 	 assign_stmt_15822_to_stmt_15849/queue_index_update_enable_out
      -- 
    getTxPacketPointerFromServer_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 47) := "getTxPacketPointerFromServer_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= getTxPacketPointerFromServer_CP_30524_elements(7);
      gj_getTxPacketPointerFromServer_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getTxPacketPointerFromServer_CP_30524_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	14 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	10 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_15822_to_stmt_15849/pkt_pointer_update_enable_in
      -- CP-element group 3: 	 assign_stmt_15822_to_stmt_15849/pkt_pointer_update_enable
      -- 
    getTxPacketPointerFromServer_CP_30524_elements(3) <= getTxPacketPointerFromServer_CP_30524_elements(14);
    -- CP-element group 4:  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	15 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	10 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_15822_to_stmt_15849/status_update_enable_in
      -- CP-element group 4: 	 assign_stmt_15822_to_stmt_15849/status_update_enable
      -- 
    getTxPacketPointerFromServer_CP_30524_elements(4) <= getTxPacketPointerFromServer_CP_30524_elements(15);
    -- CP-element group 5:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	1 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	7 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	7 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 assign_stmt_15822_to_stmt_15849/call_stmt_15832_Sample/crr
      -- CP-element group 5: 	 assign_stmt_15822_to_stmt_15849/call_stmt_15832_Sample/$entry
      -- CP-element group 5: 	 assign_stmt_15822_to_stmt_15849/call_stmt_15832_sample_start_
      -- 
    crr_30543_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_30543_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTxPacketPointerFromServer_CP_30524_elements(5), ack => call_stmt_15832_call_req_0); -- 
    getTxPacketPointerFromServer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 47) := "getTxPacketPointerFromServer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= getTxPacketPointerFromServer_CP_30524_elements(1) & getTxPacketPointerFromServer_CP_30524_elements(7);
      gj_getTxPacketPointerFromServer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getTxPacketPointerFromServer_CP_30524_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: marked-predecessors 
    -- CP-element group 6: 	8 
    -- CP-element group 6: 	11 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	8 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 assign_stmt_15822_to_stmt_15849/call_stmt_15832_Update/ccr
      -- CP-element group 6: 	 assign_stmt_15822_to_stmt_15849/call_stmt_15832_Update/$entry
      -- CP-element group 6: 	 assign_stmt_15822_to_stmt_15849/call_stmt_15832_update_start_
      -- 
    ccr_30548_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_30548_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTxPacketPointerFromServer_CP_30524_elements(6), ack => call_stmt_15832_call_req_1); -- 
    getTxPacketPointerFromServer_cp_element_group_6: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 47) := "getTxPacketPointerFromServer_cp_element_group_6"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= getTxPacketPointerFromServer_CP_30524_elements(8) & getTxPacketPointerFromServer_CP_30524_elements(11);
      gj_getTxPacketPointerFromServer_cp_element_group_6 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getTxPacketPointerFromServer_CP_30524_elements(6), clk => clk, reset => reset); --
    end block;
    -- CP-element group 7:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	5 
    -- CP-element group 7: successors 
    -- CP-element group 7: marked-successors 
    -- CP-element group 7: 	2 
    -- CP-element group 7: 	5 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 assign_stmt_15822_to_stmt_15849/call_stmt_15832_Sample/cra
      -- CP-element group 7: 	 assign_stmt_15822_to_stmt_15849/call_stmt_15832_Sample/$exit
      -- CP-element group 7: 	 assign_stmt_15822_to_stmt_15849/call_stmt_15832_sample_completed_
      -- 
    cra_30544_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_15832_call_ack_0, ack => getTxPacketPointerFromServer_CP_30524_elements(7)); -- 
    -- CP-element group 8:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	6 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8: marked-successors 
    -- CP-element group 8: 	6 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 assign_stmt_15822_to_stmt_15849/call_stmt_15832_Update/cca
      -- CP-element group 8: 	 assign_stmt_15822_to_stmt_15849/call_stmt_15832_Update/$exit
      -- CP-element group 8: 	 assign_stmt_15822_to_stmt_15849/call_stmt_15832_update_completed_
      -- 
    cca_30549_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_15832_call_ack_1, ack => getTxPacketPointerFromServer_CP_30524_elements(8)); -- 
    -- CP-element group 9:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: marked-predecessors 
    -- CP-element group 9: 	11 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 assign_stmt_15822_to_stmt_15849/call_stmt_15844_Sample/crr
      -- CP-element group 9: 	 assign_stmt_15822_to_stmt_15849/call_stmt_15844_Sample/$entry
      -- CP-element group 9: 	 assign_stmt_15822_to_stmt_15849/call_stmt_15844_sample_start_
      -- 
    crr_30557_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_30557_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTxPacketPointerFromServer_CP_30524_elements(9), ack => call_stmt_15844_call_req_0); -- 
    getTxPacketPointerFromServer_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 47) := "getTxPacketPointerFromServer_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= getTxPacketPointerFromServer_CP_30524_elements(8) & getTxPacketPointerFromServer_CP_30524_elements(11);
      gj_getTxPacketPointerFromServer_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getTxPacketPointerFromServer_CP_30524_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	3 
    -- CP-element group 10: 	4 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	12 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_15822_to_stmt_15849/call_stmt_15844_update_start_
      -- CP-element group 10: 	 assign_stmt_15822_to_stmt_15849/call_stmt_15844_Update/ccr
      -- CP-element group 10: 	 assign_stmt_15822_to_stmt_15849/call_stmt_15844_Update/$entry
      -- 
    ccr_30562_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_30562_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => getTxPacketPointerFromServer_CP_30524_elements(10), ack => call_stmt_15844_call_req_1); -- 
    getTxPacketPointerFromServer_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 7,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 48) := "getTxPacketPointerFromServer_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= getTxPacketPointerFromServer_CP_30524_elements(3) & getTxPacketPointerFromServer_CP_30524_elements(4) & getTxPacketPointerFromServer_CP_30524_elements(12);
      gj_getTxPacketPointerFromServer_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => getTxPacketPointerFromServer_CP_30524_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: marked-successors 
    -- CP-element group 11: 	6 
    -- CP-element group 11: 	9 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 assign_stmt_15822_to_stmt_15849/call_stmt_15844_Sample/$exit
      -- CP-element group 11: 	 assign_stmt_15822_to_stmt_15849/call_stmt_15844_sample_completed_
      -- CP-element group 11: 	 assign_stmt_15822_to_stmt_15849/call_stmt_15844_Sample/cra
      -- 
    cra_30558_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_15844_call_ack_0, ack => getTxPacketPointerFromServer_CP_30524_elements(11)); -- 
    -- CP-element group 12:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	16 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	10 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 assign_stmt_15822_to_stmt_15849/$exit
      -- CP-element group 12: 	 assign_stmt_15822_to_stmt_15849/call_stmt_15844_update_completed_
      -- CP-element group 12: 	 assign_stmt_15822_to_stmt_15849/call_stmt_15844_Update/cca
      -- CP-element group 12: 	 assign_stmt_15822_to_stmt_15849/call_stmt_15844_Update/$exit
      -- 
    cca_30563_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_15844_call_ack_1, ack => getTxPacketPointerFromServer_CP_30524_elements(12)); -- 
    -- CP-element group 13:  place  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	2 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 queue_index_update_enable
      -- 
    getTxPacketPointerFromServer_CP_30524_elements(13) <= getTxPacketPointerFromServer_CP_30524_elements(2);
    -- CP-element group 14:  place  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	3 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 pkt_pointer_update_enable
      -- 
    -- CP-element group 15:  place  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	4 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 status_update_enable
      -- 
    -- CP-element group 16:  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	12 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 $exit
      -- 
    getTxPacketPointerFromServer_CP_30524_elements(16) <= getTxPacketPointerFromServer_CP_30524_elements(12);
    --  hookup: inputs to control-path 
    getTxPacketPointerFromServer_CP_30524_elements(15) <= status_update_enable;
    getTxPacketPointerFromServer_CP_30524_elements(14) <= pkt_pointer_update_enable;
    -- hookup: output from control-path 
    queue_index_update_enable <= getTxPacketPointerFromServer_CP_30524_elements(13);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u6_u6_15820_wire : std_logic_vector(5 downto 0);
    signal NOT_u4_u4_15827_wire_constant : std_logic_vector(3 downto 0);
    signal R_TX_QUEUES_REG_START_OFFSET_15819_wire_constant : std_logic_vector(5 downto 0);
    signal register_index_15822 : std_logic_vector(5 downto 0);
    signal tx_queue_pointer_32_15832 : std_logic_vector(31 downto 0);
    signal tx_queue_pointer_36_15838 : std_logic_vector(35 downto 0);
    signal type_cast_15824_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_15830_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_15835_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_15840_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    NOT_u4_u4_15827_wire_constant <= "1111";
    R_TX_QUEUES_REG_START_OFFSET_15819_wire_constant <= "001010";
    type_cast_15824_wire_constant <= "1";
    type_cast_15830_wire_constant <= "00000000000000000000000000000000";
    type_cast_15835_wire_constant <= "0000";
    type_cast_15840_wire_constant <= "1";
    -- interlock type_cast_15821_inst
    process(ADD_u6_u6_15820_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := ADD_u6_u6_15820_wire(5 downto 0);
      register_index_15822 <= tmp_var; -- 
    end process;
    -- binary operator ADD_u6_u6_15820_inst
    process(queue_index_buffer) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(queue_index_buffer, R_TX_QUEUES_REG_START_OFFSET_15819_wire_constant, tmp_var);
      ADD_u6_u6_15820_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u4_u36_15837_inst
    process(type_cast_15835_wire_constant, tx_queue_pointer_32_15832) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_15835_wire_constant, tx_queue_pointer_32_15832, tmp_var);
      tx_queue_pointer_36_15838 <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_15832_call 
    AccessRegister_call_group_0: Block -- 
      signal data_in: std_logic_vector(42 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_15832_call_req_0;
      call_stmt_15832_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_15832_call_req_1;
      call_stmt_15832_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      AccessRegister_call_group_0_gI: SplitGuardInterface generic map(name => "AccessRegister_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_15824_wire_constant & NOT_u4_u4_15827_wire_constant & register_index_15822 & type_cast_15830_wire_constant;
      tx_queue_pointer_32_15832 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 43,
        owidth => 43,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => AccessRegister_call_reqs(0),
          ackR => AccessRegister_call_acks(0),
          dataR => AccessRegister_call_data(42 downto 0),
          tagR => AccessRegister_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => AccessRegister_return_acks(0), -- cross-over
          ackL => AccessRegister_return_reqs(0), -- cross-over
          dataL => AccessRegister_return_data(31 downto 0),
          tagL => AccessRegister_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_15844_call 
    popFromQueue_call_group_1: Block -- 
      signal data_in: std_logic_vector(36 downto 0);
      signal data_out: std_logic_vector(32 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_15844_call_req_0;
      call_stmt_15844_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_15844_call_req_1;
      call_stmt_15844_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      popFromQueue_call_group_1_gI: SplitGuardInterface generic map(name => "popFromQueue_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_15840_wire_constant & tx_queue_pointer_36_15838;
      pkt_pointer_buffer <= data_out(32 downto 1);
      status_buffer <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 37,
        owidth => 37,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => popFromQueue_call_reqs(0),
          ackR => popFromQueue_call_acks(0),
          dataR => popFromQueue_call_data(36 downto 0),
          tagR => popFromQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 33,
          owidth => 33,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => popFromQueue_return_acks(0), -- cross-over
          ackL => popFromQueue_return_reqs(0), -- cross-over
          dataL => popFromQueue_return_data(32 downto 0),
          tagL => popFromQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- 
  end Block; -- data_path
  -- 
end getTxPacketPointerFromServer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.nic_system_global_package.all;
entity loadBuffer is -- 
  generic (tag_length : integer); 
  port ( -- 
    rx_buffer_pointer : in  std_logic_vector(35 downto 0);
    bad_packet_identifier : out  std_logic_vector(0 downto 0);
    writePayloadToMem_call_reqs : out  std_logic_vector(0 downto 0);
    writePayloadToMem_call_acks : in   std_logic_vector(0 downto 0);
    writePayloadToMem_call_data : out  std_logic_vector(71 downto 0);
    writePayloadToMem_call_tag  :  out  std_logic_vector(0 downto 0);
    writePayloadToMem_return_reqs : out  std_logic_vector(0 downto 0);
    writePayloadToMem_return_acks : in   std_logic_vector(0 downto 0);
    writePayloadToMem_return_data : in   std_logic_vector(19 downto 0);
    writePayloadToMem_return_tag :  in   std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_call_reqs : out  std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_call_acks : in   std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_call_data : out  std_logic_vector(35 downto 0);
    writeEthernetHeaderToMem_call_tag  :  out  std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_return_reqs : out  std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_return_acks : in   std_logic_vector(0 downto 0);
    writeEthernetHeaderToMem_return_data : in   std_logic_vector(35 downto 0);
    writeEthernetHeaderToMem_return_tag :  in   std_logic_vector(0 downto 0);
    writeControlInformationToMem_call_reqs : out  std_logic_vector(0 downto 0);
    writeControlInformationToMem_call_acks : in   std_logic_vector(0 downto 0);
    writeControlInformationToMem_call_data : out  std_logic_vector(54 downto 0);
    writeControlInformationToMem_call_tag  :  out  std_logic_vector(0 downto 0);
    writeControlInformationToMem_return_reqs : out  std_logic_vector(0 downto 0);
    writeControlInformationToMem_return_acks : in   std_logic_vector(0 downto 0);
    writeControlInformationToMem_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity loadBuffer;
architecture loadBuffer_arch of loadBuffer is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 1)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rx_buffer_pointer_buffer :  std_logic_vector(35 downto 0);
  signal rx_buffer_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal bad_packet_identifier_buffer :  std_logic_vector(0 downto 0);
  signal bad_packet_identifier_update_enable: Boolean;
  signal loadBuffer_CP_1832_start: Boolean;
  signal loadBuffer_CP_1832_symbol: Boolean;
  -- volatile/operator module components. 
  component writePayloadToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      base_buf_pointer : in  std_logic_vector(35 downto 0);
      buf_pointer : in  std_logic_vector(35 downto 0);
      packet_size_32 : out  std_logic_vector(10 downto 0);
      bad_packet_identifier : out  std_logic_vector(0 downto 0);
      last_keep : out  std_logic_vector(7 downto 0);
      nic_rx_to_packet_pipe_read_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_read_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_read_data : in   std_logic_vector(72 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component writeEthernetHeaderToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      buf_pointer : in  std_logic_vector(35 downto 0);
      buf_position_out : out  std_logic_vector(35 downto 0);
      nic_rx_to_header_pipe_read_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_read_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_read_data : in   std_logic_vector(72 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component writeControlInformationToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      base_buffer_pointer : in  std_logic_vector(35 downto 0);
      packet_size : in  std_logic_vector(10 downto 0);
      last_keep : in  std_logic_vector(7 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1438_call_req_0 : boolean;
  signal call_stmt_1438_call_ack_1 : boolean;
  signal call_stmt_1438_call_req_1 : boolean;
  signal W_bad_packet_identifier_1410_delayed_8_0_1431_inst_ack_1 : boolean;
  signal call_stmt_1438_call_ack_0 : boolean;
  signal W_bad_packet_identifier_1410_delayed_8_0_1431_inst_req_1 : boolean;
  signal call_stmt_1418_call_req_0 : boolean;
  signal call_stmt_1418_call_ack_0 : boolean;
  signal call_stmt_1418_call_req_1 : boolean;
  signal call_stmt_1418_call_ack_1 : boolean;
  signal W_rx_buffer_pointer_1404_delayed_4_0_1419_inst_req_0 : boolean;
  signal W_rx_buffer_pointer_1404_delayed_4_0_1419_inst_ack_0 : boolean;
  signal W_rx_buffer_pointer_1404_delayed_4_0_1419_inst_req_1 : boolean;
  signal W_rx_buffer_pointer_1404_delayed_4_0_1419_inst_ack_1 : boolean;
  signal call_stmt_1427_call_req_0 : boolean;
  signal call_stmt_1427_call_ack_0 : boolean;
  signal call_stmt_1427_call_req_1 : boolean;
  signal call_stmt_1427_call_ack_1 : boolean;
  signal W_rx_buffer_pointer_1411_delayed_8_0_1428_inst_req_0 : boolean;
  signal W_rx_buffer_pointer_1411_delayed_8_0_1428_inst_ack_0 : boolean;
  signal W_rx_buffer_pointer_1411_delayed_8_0_1428_inst_req_1 : boolean;
  signal W_rx_buffer_pointer_1411_delayed_8_0_1428_inst_ack_1 : boolean;
  signal W_bad_packet_identifier_1410_delayed_8_0_1431_inst_req_0 : boolean;
  signal W_bad_packet_identifier_1410_delayed_8_0_1431_inst_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "loadBuffer_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= rx_buffer_pointer;
  rx_buffer_pointer_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 31);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 31);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= rx_buffer_pointer_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  loadBuffer_CP_1832_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "loadBuffer_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 1) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(0 downto 0) <= bad_packet_identifier_buffer;
  bad_packet_identifier <= out_buffer_data_out(0 downto 0);
  out_buffer_data_in(tag_length + 0 downto 1) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 0 downto 1);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 31);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadBuffer_CP_1832_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  bad_packet_identifier_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 40) := "bad_packet_identifier_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_bad_packet_identifier_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => bad_packet_identifier_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 31,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= loadBuffer_CP_1832_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= loadBuffer_CP_1832_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  loadBuffer_CP_1832: Block -- control-path 
    signal loadBuffer_CP_1832_elements: BooleanArray(30 downto 0);
    -- 
  begin -- 
    loadBuffer_CP_1832_elements(0) <= loadBuffer_CP_1832_start;
    loadBuffer_CP_1832_symbol <= loadBuffer_CP_1832_elements(30);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	16 
    -- CP-element group 1: 	4 
    -- CP-element group 1: 	8 
    -- CP-element group 1:  members (1) 
      -- CP-element group 1: 	 call_stmt_1418_to_call_stmt_1438/$entry
      -- 
    loadBuffer_CP_1832_elements(1) <= loadBuffer_CP_1832_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	18 
    -- CP-element group 2: 	6 
    -- CP-element group 2: 	10 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	28 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 call_stmt_1418_to_call_stmt_1438/rx_buffer_pointer_update_enable
      -- CP-element group 2: 	 call_stmt_1418_to_call_stmt_1438/rx_buffer_pointer_update_enable_out
      -- 
    loadBuffer_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_1832_elements(18) & loadBuffer_CP_1832_elements(6) & loadBuffer_CP_1832_elements(10);
      gj_loadBuffer_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1832_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	29 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	13 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 call_stmt_1418_to_call_stmt_1438/bad_packet_identifier_update_enable
      -- CP-element group 3: 	 call_stmt_1418_to_call_stmt_1438/bad_packet_identifier_update_enable_in
      -- 
    loadBuffer_CP_1832_elements(3) <= loadBuffer_CP_1832_elements(29);
    -- CP-element group 4:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	1 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	27 
    -- CP-element group 4: 	6 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	6 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1418_sample_start_
      -- CP-element group 4: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1418_Sample/$entry
      -- CP-element group 4: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1418_Sample/crr
      -- 
    crr_1849_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1849_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1832_elements(4), ack => call_stmt_1418_call_req_0); -- 
    loadBuffer_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_1832_elements(1) & loadBuffer_CP_1832_elements(27) & loadBuffer_CP_1832_elements(6);
      gj_loadBuffer_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1832_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	27 
    -- CP-element group 5: 	14 
    -- CP-element group 5: 	7 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	7 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1418_update_start_
      -- CP-element group 5: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1418_Update/$entry
      -- CP-element group 5: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1418_Update/ccr
      -- 
    ccr_1854_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1854_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1832_elements(5), ack => call_stmt_1418_call_req_1); -- 
    loadBuffer_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_1832_elements(27) & loadBuffer_CP_1832_elements(14) & loadBuffer_CP_1832_elements(7);
      gj_loadBuffer_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1832_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	4 
    -- CP-element group 6: successors 
    -- CP-element group 6: marked-successors 
    -- CP-element group 6: 	4 
    -- CP-element group 6: 	2 
    -- CP-element group 6:  members (3) 
      -- CP-element group 6: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1418_sample_completed_
      -- CP-element group 6: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1418_Sample/$exit
      -- CP-element group 6: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1418_Sample/cra
      -- 
    cra_1850_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1418_call_ack_0, ack => loadBuffer_CP_1832_elements(6)); -- 
    -- CP-element group 7:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	5 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	12 
    -- CP-element group 7: marked-successors 
    -- CP-element group 7: 	5 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1418_update_completed_
      -- CP-element group 7: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1418_Update/$exit
      -- CP-element group 7: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1418_Update/cca
      -- 
    cca_1855_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1418_call_ack_1, ack => loadBuffer_CP_1832_elements(7)); -- 
    -- CP-element group 8:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	1 
    -- CP-element group 8: marked-predecessors 
    -- CP-element group 8: 	10 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	10 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1421_sample_start_
      -- CP-element group 8: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1421_Sample/$entry
      -- CP-element group 8: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1421_Sample/req
      -- 
    req_1863_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1863_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1832_elements(8), ack => W_rx_buffer_pointer_1404_delayed_4_0_1419_inst_req_0); -- 
    loadBuffer_cp_element_group_8: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_8"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_1832_elements(1) & loadBuffer_CP_1832_elements(10);
      gj_loadBuffer_cp_element_group_8 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1832_elements(8), clk => clk, reset => reset); --
    end block;
    -- CP-element group 9:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: marked-predecessors 
    -- CP-element group 9: 	14 
    -- CP-element group 9: 	11 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1421_update_start_
      -- CP-element group 9: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1421_Update/$entry
      -- CP-element group 9: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1421_Update/req
      -- 
    req_1868_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1868_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1832_elements(9), ack => W_rx_buffer_pointer_1404_delayed_4_0_1419_inst_req_1); -- 
    loadBuffer_cp_element_group_9: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 29) := "loadBuffer_cp_element_group_9"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_1832_elements(14) & loadBuffer_CP_1832_elements(11);
      gj_loadBuffer_cp_element_group_9 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1832_elements(9), clk => clk, reset => reset); --
    end block;
    -- CP-element group 10:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	8 
    -- CP-element group 10: successors 
    -- CP-element group 10: marked-successors 
    -- CP-element group 10: 	8 
    -- CP-element group 10: 	2 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1421_sample_completed_
      -- CP-element group 10: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1421_Sample/$exit
      -- CP-element group 10: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1421_Sample/ack
      -- 
    ack_1864_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_1404_delayed_4_0_1419_inst_ack_0, ack => loadBuffer_CP_1832_elements(10)); -- 
    -- CP-element group 11:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11: marked-successors 
    -- CP-element group 11: 	9 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1421_update_completed_
      -- CP-element group 11: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1421_Update/$exit
      -- CP-element group 11: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1421_Update/ack
      -- 
    ack_1869_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_1404_delayed_4_0_1419_inst_ack_1, ack => loadBuffer_CP_1832_elements(11)); -- 
    -- CP-element group 12:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	7 
    -- CP-element group 12: 	11 
    -- CP-element group 12: marked-predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	14 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1427_sample_start_
      -- CP-element group 12: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1427_Sample/$entry
      -- CP-element group 12: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1427_Sample/crr
      -- 
    crr_1877_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1877_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1832_elements(12), ack => call_stmt_1427_call_req_0); -- 
    loadBuffer_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= loadBuffer_CP_1832_elements(7) & loadBuffer_CP_1832_elements(11) & loadBuffer_CP_1832_elements(14);
      gj_loadBuffer_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1832_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	3 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	22 
    -- CP-element group 13: 	26 
    -- CP-element group 13: 	15 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	15 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1427_update_start_
      -- CP-element group 13: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1427_Update/$entry
      -- CP-element group 13: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1427_Update/ccr
      -- 
    ccr_1882_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1882_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1832_elements(13), ack => call_stmt_1427_call_req_1); -- 
    loadBuffer_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= loadBuffer_CP_1832_elements(3) & loadBuffer_CP_1832_elements(22) & loadBuffer_CP_1832_elements(26) & loadBuffer_CP_1832_elements(15);
      gj_loadBuffer_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1832_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	12 
    -- CP-element group 14: successors 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	5 
    -- CP-element group 14: 	9 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1427_sample_completed_
      -- CP-element group 14: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1427_Sample/$exit
      -- CP-element group 14: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1427_Sample/cra
      -- 
    cra_1878_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 14_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1427_call_ack_0, ack => loadBuffer_CP_1832_elements(14)); -- 
    -- CP-element group 15:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	13 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	24 
    -- CP-element group 15: 	20 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	13 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1427_update_completed_
      -- CP-element group 15: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1427_Update/$exit
      -- CP-element group 15: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1427_Update/cca
      -- 
    cca_1883_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1427_call_ack_1, ack => loadBuffer_CP_1832_elements(15)); -- 
    -- CP-element group 16:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	1 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	18 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	18 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1430_sample_start_
      -- CP-element group 16: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1430_Sample/$entry
      -- CP-element group 16: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1430_Sample/req
      -- 
    req_1891_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1891_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1832_elements(16), ack => W_rx_buffer_pointer_1411_delayed_8_0_1428_inst_req_0); -- 
    loadBuffer_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_1832_elements(1) & loadBuffer_CP_1832_elements(18);
      gj_loadBuffer_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1832_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	26 
    -- CP-element group 17: 	19 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	19 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1430_update_start_
      -- CP-element group 17: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1430_Update/$entry
      -- CP-element group 17: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1430_Update/req
      -- 
    req_1896_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1896_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1832_elements(17), ack => W_rx_buffer_pointer_1411_delayed_8_0_1428_inst_req_1); -- 
    loadBuffer_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_1832_elements(26) & loadBuffer_CP_1832_elements(19);
      gj_loadBuffer_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1832_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	16 
    -- CP-element group 18: successors 
    -- CP-element group 18: marked-successors 
    -- CP-element group 18: 	16 
    -- CP-element group 18: 	2 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1430_sample_completed_
      -- CP-element group 18: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1430_Sample/$exit
      -- CP-element group 18: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1430_Sample/ack
      -- 
    ack_1892_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_1411_delayed_8_0_1428_inst_ack_0, ack => loadBuffer_CP_1832_elements(18)); -- 
    -- CP-element group 19:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	17 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	24 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	17 
    -- CP-element group 19:  members (3) 
      -- CP-element group 19: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1430_update_completed_
      -- CP-element group 19: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1430_Update/$exit
      -- CP-element group 19: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1430_Update/ack
      -- 
    ack_1897_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rx_buffer_pointer_1411_delayed_8_0_1428_inst_ack_1, ack => loadBuffer_CP_1832_elements(19)); -- 
    -- CP-element group 20:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	15 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	22 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	22 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1433_sample_start_
      -- CP-element group 20: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1433_Sample/$entry
      -- CP-element group 20: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1433_Sample/req
      -- 
    req_1905_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1905_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1832_elements(20), ack => W_bad_packet_identifier_1410_delayed_8_0_1431_inst_req_0); -- 
    loadBuffer_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_1832_elements(15) & loadBuffer_CP_1832_elements(22);
      gj_loadBuffer_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1832_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	23 
    -- CP-element group 21: 	26 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1433_Update/req
      -- CP-element group 21: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1433_update_start_
      -- CP-element group 21: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1433_Update/$entry
      -- 
    req_1910_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1910_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1832_elements(21), ack => W_bad_packet_identifier_1410_delayed_8_0_1431_inst_req_1); -- 
    loadBuffer_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= loadBuffer_CP_1832_elements(23) & loadBuffer_CP_1832_elements(26);
      gj_loadBuffer_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1832_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	20 
    -- CP-element group 22: successors 
    -- CP-element group 22: marked-successors 
    -- CP-element group 22: 	13 
    -- CP-element group 22: 	20 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1433_sample_completed_
      -- CP-element group 22: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1433_Sample/$exit
      -- CP-element group 22: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1433_Sample/ack
      -- 
    ack_1906_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bad_packet_identifier_1410_delayed_8_0_1431_inst_ack_0, ack => loadBuffer_CP_1832_elements(22)); -- 
    -- CP-element group 23:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	21 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1433_Update/ack
      -- CP-element group 23: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1433_update_completed_
      -- CP-element group 23: 	 call_stmt_1418_to_call_stmt_1438/assign_stmt_1433_Update/$exit
      -- 
    ack_1911_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_bad_packet_identifier_1410_delayed_8_0_1431_inst_ack_1, ack => loadBuffer_CP_1832_elements(23)); -- 
    -- CP-element group 24:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	23 
    -- CP-element group 24: 	15 
    -- CP-element group 24: 	19 
    -- CP-element group 24: marked-predecessors 
    -- CP-element group 24: 	26 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (3) 
      -- CP-element group 24: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1438_Sample/crr
      -- CP-element group 24: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1438_sample_start_
      -- CP-element group 24: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1438_Sample/$entry
      -- 
    crr_1919_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1919_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1832_elements(24), ack => call_stmt_1438_call_req_0); -- 
    loadBuffer_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= loadBuffer_CP_1832_elements(23) & loadBuffer_CP_1832_elements(15) & loadBuffer_CP_1832_elements(19) & loadBuffer_CP_1832_elements(26);
      gj_loadBuffer_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1832_elements(24), clk => clk, reset => reset); --
    end block;
    -- CP-element group 25:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	27 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (3) 
      -- CP-element group 25: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1438_update_start_
      -- CP-element group 25: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1438_Update/ccr
      -- CP-element group 25: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1438_Update/$entry
      -- 
    ccr_1924_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1924_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => loadBuffer_CP_1832_elements(25), ack => call_stmt_1438_call_req_1); -- 
    loadBuffer_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 30) := "loadBuffer_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= loadBuffer_CP_1832_elements(27);
      gj_loadBuffer_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => loadBuffer_CP_1832_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26: marked-successors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: 	13 
    -- CP-element group 26: 	17 
    -- CP-element group 26: 	21 
    -- CP-element group 26:  members (3) 
      -- CP-element group 26: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1438_sample_completed_
      -- CP-element group 26: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1438_Sample/$exit
      -- CP-element group 26: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1438_Sample/cra
      -- 
    cra_1920_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1438_call_ack_0, ack => loadBuffer_CP_1832_elements(26)); -- 
    -- CP-element group 27:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	30 
    -- CP-element group 27: marked-successors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: 	4 
    -- CP-element group 27: 	5 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1438_Update/cca
      -- CP-element group 27: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1438_update_completed_
      -- CP-element group 27: 	 call_stmt_1418_to_call_stmt_1438/call_stmt_1438_Update/$exit
      -- CP-element group 27: 	 call_stmt_1418_to_call_stmt_1438/$exit
      -- 
    cca_1925_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1438_call_ack_1, ack => loadBuffer_CP_1832_elements(27)); -- 
    -- CP-element group 28:  place  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	2 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 rx_buffer_pointer_update_enable
      -- 
    loadBuffer_CP_1832_elements(28) <= loadBuffer_CP_1832_elements(2);
    -- CP-element group 29:  place  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	3 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 bad_packet_identifier_update_enable
      -- 
    -- CP-element group 30:  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	27 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 $exit
      -- 
    loadBuffer_CP_1832_elements(30) <= loadBuffer_CP_1832_elements(27);
    --  hookup: inputs to control-path 
    loadBuffer_CP_1832_elements(29) <= bad_packet_identifier_update_enable;
    -- hookup: output from control-path 
    rx_buffer_pointer_update_enable <= loadBuffer_CP_1832_elements(28);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal bad_packet_identifier_1410_delayed_8_0_1433 : std_logic_vector(0 downto 0);
    signal last_keep_1427 : std_logic_vector(7 downto 0);
    signal new_buf_pointer_1418 : std_logic_vector(35 downto 0);
    signal packet_size_1427 : std_logic_vector(10 downto 0);
    signal rx_buffer_pointer_1404_delayed_4_0_1421 : std_logic_vector(35 downto 0);
    signal rx_buffer_pointer_1411_delayed_8_0_1430 : std_logic_vector(35 downto 0);
    -- 
  begin -- 
    W_bad_packet_identifier_1410_delayed_8_0_1431_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_bad_packet_identifier_1410_delayed_8_0_1431_inst_req_0;
      W_bad_packet_identifier_1410_delayed_8_0_1431_inst_ack_0<= wack(0);
      rreq(0) <= W_bad_packet_identifier_1410_delayed_8_0_1431_inst_req_1;
      W_bad_packet_identifier_1410_delayed_8_0_1431_inst_ack_1<= rack(0);
      W_bad_packet_identifier_1410_delayed_8_0_1431_inst : InterlockBuffer generic map ( -- 
        name => "W_bad_packet_identifier_1410_delayed_8_0_1431_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => bad_packet_identifier_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => bad_packet_identifier_1410_delayed_8_0_1433,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rx_buffer_pointer_1404_delayed_4_0_1419_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rx_buffer_pointer_1404_delayed_4_0_1419_inst_req_0;
      W_rx_buffer_pointer_1404_delayed_4_0_1419_inst_ack_0<= wack(0);
      rreq(0) <= W_rx_buffer_pointer_1404_delayed_4_0_1419_inst_req_1;
      W_rx_buffer_pointer_1404_delayed_4_0_1419_inst_ack_1<= rack(0);
      W_rx_buffer_pointer_1404_delayed_4_0_1419_inst : InterlockBuffer generic map ( -- 
        name => "W_rx_buffer_pointer_1404_delayed_4_0_1419_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rx_buffer_pointer_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rx_buffer_pointer_1404_delayed_4_0_1421,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rx_buffer_pointer_1411_delayed_8_0_1428_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rx_buffer_pointer_1411_delayed_8_0_1428_inst_req_0;
      W_rx_buffer_pointer_1411_delayed_8_0_1428_inst_ack_0<= wack(0);
      rreq(0) <= W_rx_buffer_pointer_1411_delayed_8_0_1428_inst_req_1;
      W_rx_buffer_pointer_1411_delayed_8_0_1428_inst_ack_1<= rack(0);
      W_rx_buffer_pointer_1411_delayed_8_0_1428_inst : InterlockBuffer generic map ( -- 
        name => "W_rx_buffer_pointer_1411_delayed_8_0_1428_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rx_buffer_pointer_buffer,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rx_buffer_pointer_1411_delayed_8_0_1430,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- shared call operator group (0) : call_stmt_1418_call 
    writeEthernetHeaderToMem_call_group_0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1418_call_req_0;
      call_stmt_1418_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1418_call_req_1;
      call_stmt_1418_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      writeEthernetHeaderToMem_call_group_0_gI: SplitGuardInterface generic map(name => "writeEthernetHeaderToMem_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_buffer_pointer_buffer;
      new_buf_pointer_1418 <= data_out(35 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => writeEthernetHeaderToMem_call_reqs(0),
          ackR => writeEthernetHeaderToMem_call_acks(0),
          dataR => writeEthernetHeaderToMem_call_data(35 downto 0),
          tagR => writeEthernetHeaderToMem_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 36,
          owidth => 36,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => writeEthernetHeaderToMem_return_acks(0), -- cross-over
          ackL => writeEthernetHeaderToMem_return_reqs(0), -- cross-over
          dataL => writeEthernetHeaderToMem_return_data(35 downto 0),
          tagL => writeEthernetHeaderToMem_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1427_call 
    writePayloadToMem_call_group_1: Block -- 
      signal data_in: std_logic_vector(71 downto 0);
      signal data_out: std_logic_vector(19 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1427_call_req_0;
      call_stmt_1427_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1427_call_req_1;
      call_stmt_1427_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      writePayloadToMem_call_group_1_gI: SplitGuardInterface generic map(name => "writePayloadToMem_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_buffer_pointer_1404_delayed_4_0_1421 & new_buf_pointer_1418;
      packet_size_1427 <= data_out(19 downto 9);
      bad_packet_identifier_buffer <= data_out(8 downto 8);
      last_keep_1427 <= data_out(7 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 72,
        owidth => 72,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => writePayloadToMem_call_reqs(0),
          ackR => writePayloadToMem_call_acks(0),
          dataR => writePayloadToMem_call_data(71 downto 0),
          tagR => writePayloadToMem_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 20,
          owidth => 20,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => writePayloadToMem_return_acks(0), -- cross-over
          ackL => writePayloadToMem_return_reqs(0), -- cross-over
          dataL => writePayloadToMem_return_data(19 downto 0),
          tagL => writePayloadToMem_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1438_call 
    writeControlInformationToMem_call_group_2: Block -- 
      signal data_in: std_logic_vector(54 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1438_call_req_0;
      call_stmt_1438_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1438_call_req_1;
      call_stmt_1438_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not bad_packet_identifier_1410_delayed_8_0_1433(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      writeControlInformationToMem_call_group_2_gI: SplitGuardInterface generic map(name => "writeControlInformationToMem_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= rx_buffer_pointer_1411_delayed_8_0_1430 & packet_size_1427 & last_keep_1427;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 55,
        owidth => 55,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => writeControlInformationToMem_call_reqs(0),
          ackR => writeControlInformationToMem_call_acks(0),
          dataR => writeControlInformationToMem_call_data(54 downto 0),
          tagR => writeControlInformationToMem_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => writeControlInformationToMem_return_acks(0), -- cross-over
          ackL => writeControlInformationToMem_return_reqs(0), -- cross-over
          tagL => writeControlInformationToMem_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end loadBuffer_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.nic_system_global_package.all;
entity nextLSTATE_Volatile is -- 
  port ( -- 
    RX : in  std_logic_vector(72 downto 0);
    LSTATE : in  std_logic_vector(1 downto 0);
    nLSTATE : out  std_logic_vector(1 downto 0)-- 
  );
  -- 
end entity nextLSTATE_Volatile;
architecture nextLSTATE_Volatile_arch of nextLSTATE_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(75-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal RX_buffer :  std_logic_vector(72 downto 0);
  signal LSTATE_buffer :  std_logic_vector(1 downto 0);
  -- output port buffer signals
  signal nLSTATE_buffer :  std_logic_vector(1 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  RX_buffer <= RX;
  LSTATE_buffer <= LSTATE;
  -- output handling  -------------------------------------------------------
  nLSTATE <= nLSTATE_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_15911_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_15919_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_15875_wire : std_logic_vector(0 downto 0);
    signal EQ_u1_u1_15893_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_15884_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_15890_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_15901_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_15908_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_15917_wire : std_logic_vector(0 downto 0);
    signal MUX_15887_wire : std_logic_vector(1 downto 0);
    signal MUX_15897_wire : std_logic_vector(1 downto 0);
    signal MUX_15904_wire : std_logic_vector(1 downto 0);
    signal MUX_15914_wire : std_logic_vector(1 downto 0);
    signal MUX_15922_wire : std_logic_vector(1 downto 0);
    signal NEQ_u2_u1_15878_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_15910_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_15894_wire : std_logic_vector(0 downto 0);
    signal OR_u2_u2_15898_wire : std_logic_vector(1 downto 0);
    signal OR_u2_u2_15905_wire : std_logic_vector(1 downto 0);
    signal OR_u2_u2_15923_wire : std_logic_vector(1 downto 0);
    signal R_S0_15883_wire_constant : std_logic_vector(1 downto 0);
    signal R_S0_15895_wire_constant : std_logic_vector(1 downto 0);
    signal R_S0_15920_wire_constant : std_logic_vector(1 downto 0);
    signal R_S1_15885_wire_constant : std_logic_vector(1 downto 0);
    signal R_S1_15900_wire_constant : std_logic_vector(1 downto 0);
    signal R_S2_15877_wire_constant : std_logic_vector(1 downto 0);
    signal R_S2_15902_wire_constant : std_logic_vector(1 downto 0);
    signal R_S2_15907_wire_constant : std_logic_vector(1 downto 0);
    signal R_S2_15912_wire_constant : std_logic_vector(1 downto 0);
    signal R_S2_15916_wire_constant : std_logic_vector(1 downto 0);
    signal R_S3_15889_wire_constant : std_logic_vector(1 downto 0);
    signal go_to_s0_15880 : std_logic_vector(0 downto 0);
    signal konst_15869_wire_constant : std_logic_vector(0 downto 0);
    signal konst_15874_wire_constant : std_logic_vector(0 downto 0);
    signal konst_15886_wire_constant : std_logic_vector(1 downto 0);
    signal konst_15892_wire_constant : std_logic_vector(0 downto 0);
    signal konst_15896_wire_constant : std_logic_vector(1 downto 0);
    signal konst_15903_wire_constant : std_logic_vector(1 downto 0);
    signal konst_15913_wire_constant : std_logic_vector(1 downto 0);
    signal konst_15921_wire_constant : std_logic_vector(1 downto 0);
    signal last_word_15871 : std_logic_vector(0 downto 0);
    signal tlast_15866 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_S0_15883_wire_constant <= "00";
    R_S0_15895_wire_constant <= "00";
    R_S0_15920_wire_constant <= "00";
    R_S1_15885_wire_constant <= "01";
    R_S1_15900_wire_constant <= "01";
    R_S2_15877_wire_constant <= "10";
    R_S2_15902_wire_constant <= "10";
    R_S2_15907_wire_constant <= "10";
    R_S2_15912_wire_constant <= "10";
    R_S2_15916_wire_constant <= "10";
    R_S3_15889_wire_constant <= "11";
    konst_15869_wire_constant <= "1";
    konst_15874_wire_constant <= "1";
    konst_15886_wire_constant <= "00";
    konst_15892_wire_constant <= "1";
    konst_15896_wire_constant <= "00";
    konst_15903_wire_constant <= "00";
    konst_15913_wire_constant <= "00";
    konst_15921_wire_constant <= "00";
    -- flow-through select operator MUX_15887_inst
    MUX_15887_wire <= R_S1_15885_wire_constant when (EQ_u2_u1_15884_wire(0) /=  '0') else konst_15886_wire_constant;
    -- flow-through select operator MUX_15897_inst
    MUX_15897_wire <= R_S0_15895_wire_constant when (OR_u1_u1_15894_wire(0) /=  '0') else konst_15896_wire_constant;
    -- flow-through select operator MUX_15904_inst
    MUX_15904_wire <= R_S2_15902_wire_constant when (EQ_u2_u1_15901_wire(0) /=  '0') else konst_15903_wire_constant;
    -- flow-through select operator MUX_15914_inst
    MUX_15914_wire <= R_S2_15912_wire_constant when (AND_u1_u1_15911_wire(0) /=  '0') else konst_15913_wire_constant;
    -- flow-through select operator MUX_15922_inst
    MUX_15922_wire <= R_S0_15920_wire_constant when (AND_u1_u1_15919_wire(0) /=  '0') else konst_15921_wire_constant;
    -- flow-through slice operator slice_15865_inst
    tlast_15866 <= RX_buffer(72 downto 72);
    -- binary operator AND_u1_u1_15879_inst
    process(EQ_u1_u1_15875_wire, NEQ_u2_u1_15878_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u1_u1_15875_wire, NEQ_u2_u1_15878_wire, tmp_var);
      go_to_s0_15880 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_15911_inst
    process(EQ_u2_u1_15908_wire, NOT_u1_u1_15910_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_15908_wire, NOT_u1_u1_15910_wire, tmp_var);
      AND_u1_u1_15911_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_15919_inst
    process(EQ_u2_u1_15917_wire, last_word_15871) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u2_u1_15917_wire, last_word_15871, tmp_var);
      AND_u1_u1_15919_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_15870_inst
    process(tlast_15866) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(tlast_15866, konst_15869_wire_constant, tmp_var);
      last_word_15871 <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_15875_inst
    process(last_word_15871) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(last_word_15871, konst_15874_wire_constant, tmp_var);
      EQ_u1_u1_15875_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_15893_inst
    process(go_to_s0_15880) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(go_to_s0_15880, konst_15892_wire_constant, tmp_var);
      EQ_u1_u1_15893_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_15884_inst
    process(LSTATE_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_buffer, R_S0_15883_wire_constant, tmp_var);
      EQ_u2_u1_15884_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_15890_inst
    process(LSTATE_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_buffer, R_S3_15889_wire_constant, tmp_var);
      EQ_u2_u1_15890_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_15901_inst
    process(LSTATE_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_buffer, R_S1_15900_wire_constant, tmp_var);
      EQ_u2_u1_15901_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_15908_inst
    process(LSTATE_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_buffer, R_S2_15907_wire_constant, tmp_var);
      EQ_u2_u1_15908_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_15917_inst
    process(LSTATE_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_buffer, R_S2_15916_wire_constant, tmp_var);
      EQ_u2_u1_15917_wire <= tmp_var; --
    end process;
    -- binary operator NEQ_u2_u1_15878_inst
    process(LSTATE_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(LSTATE_buffer, R_S2_15877_wire_constant, tmp_var);
      NEQ_u2_u1_15878_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_15910_inst
    process(last_word_15871) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", last_word_15871, tmp_var);
      NOT_u1_u1_15910_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_15894_inst
    process(EQ_u2_u1_15890_wire, EQ_u1_u1_15893_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u2_u1_15890_wire, EQ_u1_u1_15893_wire, tmp_var);
      OR_u1_u1_15894_wire <= tmp_var; --
    end process;
    -- binary operator OR_u2_u2_15898_inst
    process(MUX_15887_wire, MUX_15897_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_15887_wire, MUX_15897_wire, tmp_var);
      OR_u2_u2_15898_wire <= tmp_var; --
    end process;
    -- binary operator OR_u2_u2_15905_inst
    process(OR_u2_u2_15898_wire, MUX_15904_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u2_u2_15898_wire, MUX_15904_wire, tmp_var);
      OR_u2_u2_15905_wire <= tmp_var; --
    end process;
    -- binary operator OR_u2_u2_15923_inst
    process(MUX_15914_wire, MUX_15922_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_15914_wire, MUX_15922_wire, tmp_var);
      OR_u2_u2_15923_wire <= tmp_var; --
    end process;
    -- binary operator OR_u2_u2_15924_inst
    process(OR_u2_u2_15905_wire, OR_u2_u2_15923_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u2_u2_15905_wire, OR_u2_u2_15923_wire, tmp_var);
      nLSTATE_buffer <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end nextLSTATE_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.nic_system_global_package.all;
entity nicRxFromMacDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    mac_to_nic_data_pipe_read_req : out  std_logic_vector(0 downto 0);
    mac_to_nic_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
    mac_to_nic_data_pipe_read_data : in   std_logic_vector(72 downto 0);
    CONTROL_REGISTER : in std_logic_vector(31 downto 0);
    nic_rx_to_header_pipe_write_req : out  std_logic_vector(0 downto 0);
    nic_rx_to_header_pipe_write_ack : in   std_logic_vector(0 downto 0);
    nic_rx_to_header_pipe_write_data : out  std_logic_vector(72 downto 0);
    nic_rx_to_packet_pipe_write_req : out  std_logic_vector(0 downto 0);
    nic_rx_to_packet_pipe_write_ack : in   std_logic_vector(0 downto 0);
    nic_rx_to_packet_pipe_write_data : out  std_logic_vector(72 downto 0);
    AccessRegister_call_reqs : out  std_logic_vector(1 downto 0);
    AccessRegister_call_acks : in   std_logic_vector(1 downto 0);
    AccessRegister_call_data : out  std_logic_vector(85 downto 0);
    AccessRegister_call_tag  :  out  std_logic_vector(3 downto 0);
    AccessRegister_return_reqs : out  std_logic_vector(1 downto 0);
    AccessRegister_return_acks : in   std_logic_vector(1 downto 0);
    AccessRegister_return_data : in   std_logic_vector(63 downto 0);
    AccessRegister_return_tag :  in   std_logic_vector(3 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity nicRxFromMacDaemon;
architecture nicRxFromMacDaemon_arch of nicRxFromMacDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal nicRxFromMacDaemon_CP_30596_start: Boolean;
  signal nicRxFromMacDaemon_CP_30596_symbol: Boolean;
  -- volatile/operator module components. 
  component AccessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      register_index : in  std_logic_vector(5 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component nextLSTATE_Volatile is -- 
    port ( -- 
      RX : in  std_logic_vector(72 downto 0);
      LSTATE : in  std_logic_vector(1 downto 0);
      nLSTATE : out  std_logic_vector(1 downto 0)-- 
    );
    -- 
  end component; 
  -- links between control-path and data-path
  signal call_stmt_15940_call_req_0 : boolean;
  signal call_stmt_15940_call_ack_0 : boolean;
  signal call_stmt_15940_call_req_1 : boolean;
  signal call_stmt_15940_call_ack_1 : boolean;
  signal if_stmt_15941_branch_req_0 : boolean;
  signal if_stmt_15941_branch_ack_1 : boolean;
  signal if_stmt_15941_branch_ack_0 : boolean;
  signal call_stmt_15958_call_req_0 : boolean;
  signal call_stmt_15958_call_ack_0 : boolean;
  signal call_stmt_15958_call_req_1 : boolean;
  signal call_stmt_15958_call_ack_1 : boolean;
  signal do_while_stmt_15959_branch_req_0 : boolean;
  signal phi_stmt_15961_req_1 : boolean;
  signal phi_stmt_15961_req_0 : boolean;
  signal phi_stmt_15961_ack_0 : boolean;
  signal nLSTATE_15980_15964_buf_req_0 : boolean;
  signal nLSTATE_15980_15964_buf_ack_0 : boolean;
  signal nLSTATE_15980_15964_buf_req_1 : boolean;
  signal nLSTATE_15980_15964_buf_ack_1 : boolean;
  signal RPIPE_mac_to_nic_data_15967_inst_req_0 : boolean;
  signal RPIPE_mac_to_nic_data_15967_inst_ack_0 : boolean;
  signal RPIPE_mac_to_nic_data_15967_inst_req_1 : boolean;
  signal RPIPE_mac_to_nic_data_15967_inst_ack_1 : boolean;
  signal phi_stmt_15968_req_1 : boolean;
  signal phi_stmt_15968_req_0 : boolean;
  signal phi_stmt_15968_ack_0 : boolean;
  signal npkt_cnt_16018_15972_buf_req_0 : boolean;
  signal npkt_cnt_16018_15972_buf_ack_0 : boolean;
  signal npkt_cnt_16018_15972_buf_req_1 : boolean;
  signal npkt_cnt_16018_15972_buf_ack_1 : boolean;
  signal MUX_16000_inst_req_0 : boolean;
  signal MUX_16000_inst_ack_0 : boolean;
  signal MUX_16000_inst_req_1 : boolean;
  signal MUX_16000_inst_ack_1 : boolean;
  signal WPIPE_nic_rx_to_header_15991_inst_req_0 : boolean;
  signal WPIPE_nic_rx_to_header_15991_inst_ack_0 : boolean;
  signal WPIPE_nic_rx_to_header_15991_inst_req_1 : boolean;
  signal WPIPE_nic_rx_to_header_15991_inst_ack_1 : boolean;
  signal WPIPE_nic_rx_to_packet_16002_inst_req_0 : boolean;
  signal WPIPE_nic_rx_to_packet_16002_inst_ack_0 : boolean;
  signal WPIPE_nic_rx_to_packet_16002_inst_req_1 : boolean;
  signal WPIPE_nic_rx_to_packet_16002_inst_ack_1 : boolean;
  signal call_stmt_16028_call_req_0 : boolean;
  signal call_stmt_16028_call_ack_0 : boolean;
  signal call_stmt_16028_call_req_1 : boolean;
  signal call_stmt_16028_call_ack_1 : boolean;
  signal do_while_stmt_15959_branch_ack_0 : boolean;
  signal do_while_stmt_15959_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "nicRxFromMacDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  nicRxFromMacDaemon_CP_30596_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "nicRxFromMacDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= nicRxFromMacDaemon_CP_30596_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= nicRxFromMacDaemon_CP_30596_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= nicRxFromMacDaemon_CP_30596_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  nicRxFromMacDaemon_CP_30596: Block -- control-path 
    signal nicRxFromMacDaemon_CP_30596_elements: BooleanArray(82 downto 0);
    -- 
  begin -- 
    nicRxFromMacDaemon_CP_30596_elements(0) <= nicRxFromMacDaemon_CP_30596_start;
    nicRxFromMacDaemon_CP_30596_symbol <= nicRxFromMacDaemon_CP_30596_elements(1);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	82 
    -- CP-element group 0:  members (7) 
      -- CP-element group 0: 	 branch_block_stmt_15928/merge_stmt_15930__entry___PhiReq/$entry
      -- CP-element group 0: 	 branch_block_stmt_15928/merge_stmt_15930__entry___PhiReq/$exit
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_15928/$entry
      -- CP-element group 0: 	 branch_block_stmt_15928/branch_block_stmt_15928__entry__
      -- CP-element group 0: 	 branch_block_stmt_15928/merge_stmt_15930__entry__
      -- CP-element group 0: 	 branch_block_stmt_15928/merge_stmt_15930_dead_link/$entry
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_15928/$exit
      -- CP-element group 1: 	 branch_block_stmt_15928/branch_block_stmt_15928__exit__
      -- 
    nicRxFromMacDaemon_CP_30596_elements(1) <= false; 
    -- CP-element group 2:  transition  place  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	81 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	82 
    -- CP-element group 2:  members (4) 
      -- CP-element group 2: 	 branch_block_stmt_15928/disable_loopback_PhiReq/$entry
      -- CP-element group 2: 	 branch_block_stmt_15928/disable_loopback_PhiReq/$exit
      -- CP-element group 2: 	 branch_block_stmt_15928/do_while_stmt_15959__exit__
      -- CP-element group 2: 	 branch_block_stmt_15928/disable_loopback
      -- 
    nicRxFromMacDaemon_CP_30596_elements(2) <= nicRxFromMacDaemon_CP_30596_elements(81);
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	82 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 branch_block_stmt_15928/call_stmt_15940/call_stmt_15940_sample_completed_
      -- CP-element group 3: 	 branch_block_stmt_15928/call_stmt_15940/call_stmt_15940_Sample/$exit
      -- CP-element group 3: 	 branch_block_stmt_15928/call_stmt_15940/call_stmt_15940_Sample/cra
      -- 
    cra_30626_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_15940_call_ack_0, ack => nicRxFromMacDaemon_CP_30596_elements(3)); -- 
    -- CP-element group 4:  branch  transition  place  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	82 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4: 	6 
    -- CP-element group 4:  members (49) 
      -- CP-element group 4: 	 branch_block_stmt_15928/call_stmt_15940__exit__
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941__entry__
      -- CP-element group 4: 	 branch_block_stmt_15928/call_stmt_15940/$exit
      -- CP-element group 4: 	 branch_block_stmt_15928/call_stmt_15940/call_stmt_15940_update_completed_
      -- CP-element group 4: 	 branch_block_stmt_15928/call_stmt_15940/call_stmt_15940_Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_15928/call_stmt_15940/call_stmt_15940_Update/cca
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_dead_link/$entry
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/$entry
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/$exit
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/$entry
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/$exit
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/BITSEL_u32_u1_15944/$entry
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/BITSEL_u32_u1_15944/$exit
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/BITSEL_u32_u1_15944/BITSEL_u32_u1_15944_inputs/$entry
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/BITSEL_u32_u1_15944/BITSEL_u32_u1_15944_inputs/$exit
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/BITSEL_u32_u1_15944/BITSEL_u32_u1_15944_inputs/RPIPE_CONTROL_REGISTER_15942/$entry
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/BITSEL_u32_u1_15944/BITSEL_u32_u1_15944_inputs/RPIPE_CONTROL_REGISTER_15942/$exit
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/BITSEL_u32_u1_15944/BITSEL_u32_u1_15944_inputs/RPIPE_CONTROL_REGISTER_15942/Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/BITSEL_u32_u1_15944/BITSEL_u32_u1_15944_inputs/RPIPE_CONTROL_REGISTER_15942/Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/BITSEL_u32_u1_15944/BITSEL_u32_u1_15944_inputs/RPIPE_CONTROL_REGISTER_15942/Sample/req
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/BITSEL_u32_u1_15944/BITSEL_u32_u1_15944_inputs/RPIPE_CONTROL_REGISTER_15942/Sample/ack
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/BITSEL_u32_u1_15944/BITSEL_u32_u1_15944_inputs/RPIPE_CONTROL_REGISTER_15942/Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/BITSEL_u32_u1_15944/BITSEL_u32_u1_15944_inputs/RPIPE_CONTROL_REGISTER_15942/Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/BITSEL_u32_u1_15944/BITSEL_u32_u1_15944_inputs/RPIPE_CONTROL_REGISTER_15942/Update/req
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/BITSEL_u32_u1_15944/BITSEL_u32_u1_15944_inputs/RPIPE_CONTROL_REGISTER_15942/Update/ack
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/BITSEL_u32_u1_15944/SplitProtocol/$entry
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/BITSEL_u32_u1_15944/SplitProtocol/$exit
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/BITSEL_u32_u1_15944/SplitProtocol/Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/BITSEL_u32_u1_15944/SplitProtocol/Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/BITSEL_u32_u1_15944/SplitProtocol/Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/BITSEL_u32_u1_15944/SplitProtocol/Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/BITSEL_u32_u1_15944/SplitProtocol/Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/BITSEL_u32_u1_15944/SplitProtocol/Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/BITSEL_u32_u1_15944/SplitProtocol/Update/cr
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/BITSEL_u32_u1_15944/SplitProtocol/Update/ca
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/SplitProtocol/$entry
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/SplitProtocol/$exit
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/SplitProtocol/Sample/$entry
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/SplitProtocol/Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/SplitProtocol/Sample/rr
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/SplitProtocol/Sample/ra
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/SplitProtocol/Update/$entry
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/SplitProtocol/Update/$exit
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/SplitProtocol/Update/cr
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/NOT_u1_u1_15945/SplitProtocol/Update/ca
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_eval_test/branch_req
      -- CP-element group 4: 	 branch_block_stmt_15928/NOT_u1_u1_15945_place
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_if_link/$entry
      -- CP-element group 4: 	 branch_block_stmt_15928/if_stmt_15941_else_link/$entry
      -- 
    cca_30631_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_15940_call_ack_1, ack => nicRxFromMacDaemon_CP_30596_elements(4)); -- 
    branch_req_30687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_30687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_30596_elements(4), ack => if_stmt_15941_branch_req_0); -- 
    -- CP-element group 5:  transition  place  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	82 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_15928/not_enabled_yet_loopback_PhiReq/$entry
      -- CP-element group 5: 	 branch_block_stmt_15928/not_enabled_yet_loopback_PhiReq/$exit
      -- CP-element group 5: 	 branch_block_stmt_15928/if_stmt_15941_if_link/$exit
      -- CP-element group 5: 	 branch_block_stmt_15928/if_stmt_15941_if_link/if_choice_transition
      -- CP-element group 5: 	 branch_block_stmt_15928/not_enabled_yet_loopback
      -- 
    if_choice_transition_30692_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_15941_branch_ack_1, ack => nicRxFromMacDaemon_CP_30596_elements(5)); -- 
    -- CP-element group 6:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	4 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	8 
    -- CP-element group 6:  members (11) 
      -- CP-element group 6: 	 branch_block_stmt_15928/if_stmt_15941__exit__
      -- CP-element group 6: 	 branch_block_stmt_15928/call_stmt_15958__entry__
      -- CP-element group 6: 	 branch_block_stmt_15928/if_stmt_15941_else_link/$exit
      -- CP-element group 6: 	 branch_block_stmt_15928/if_stmt_15941_else_link/else_choice_transition
      -- CP-element group 6: 	 branch_block_stmt_15928/call_stmt_15958/$entry
      -- CP-element group 6: 	 branch_block_stmt_15928/call_stmt_15958/call_stmt_15958_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_15928/call_stmt_15958/call_stmt_15958_update_start_
      -- CP-element group 6: 	 branch_block_stmt_15928/call_stmt_15958/call_stmt_15958_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_15928/call_stmt_15958/call_stmt_15958_Sample/crr
      -- CP-element group 6: 	 branch_block_stmt_15928/call_stmt_15958/call_stmt_15958_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_15928/call_stmt_15958/call_stmt_15958_Update/ccr
      -- 
    else_choice_transition_30696_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_15941_branch_ack_0, ack => nicRxFromMacDaemon_CP_30596_elements(6)); -- 
    crr_30708_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_30708_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_30596_elements(6), ack => call_stmt_15958_call_req_0); -- 
    ccr_30713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_30713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_30596_elements(6), ack => call_stmt_15958_call_req_1); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_15928/call_stmt_15958/call_stmt_15958_sample_completed_
      -- CP-element group 7: 	 branch_block_stmt_15928/call_stmt_15958/call_stmt_15958_Sample/$exit
      -- CP-element group 7: 	 branch_block_stmt_15928/call_stmt_15958/call_stmt_15958_Sample/cra
      -- 
    cra_30709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_15958_call_ack_0, ack => nicRxFromMacDaemon_CP_30596_elements(7)); -- 
    -- CP-element group 8:  transition  place  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	6 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 branch_block_stmt_15928/call_stmt_15958__exit__
      -- CP-element group 8: 	 branch_block_stmt_15928/do_while_stmt_15959__entry__
      -- CP-element group 8: 	 branch_block_stmt_15928/call_stmt_15958/$exit
      -- CP-element group 8: 	 branch_block_stmt_15928/call_stmt_15958/call_stmt_15958_update_completed_
      -- CP-element group 8: 	 branch_block_stmt_15928/call_stmt_15958/call_stmt_15958_Update/$exit
      -- CP-element group 8: 	 branch_block_stmt_15928/call_stmt_15958/call_stmt_15958_Update/cca
      -- 
    cca_30714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_15958_call_ack_1, ack => nicRxFromMacDaemon_CP_30596_elements(8)); -- 
    -- CP-element group 9:  transition  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	15 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_15928/do_while_stmt_15959/$entry
      -- CP-element group 9: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959__entry__
      -- 
    nicRxFromMacDaemon_CP_30596_elements(9) <= nicRxFromMacDaemon_CP_30596_elements(8);
    -- CP-element group 10:  merge  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	81 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959__exit__
      -- 
    -- Element group nicRxFromMacDaemon_CP_30596_elements(10) is bound as output of CP function.
    -- CP-element group 11:  merge  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	14 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_15928/do_while_stmt_15959/loop_back
      -- 
    -- Element group nicRxFromMacDaemon_CP_30596_elements(11) is bound as output of CP function.
    -- CP-element group 12:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	17 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	79 
    -- CP-element group 12: 	80 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_15928/do_while_stmt_15959/condition_done
      -- CP-element group 12: 	 branch_block_stmt_15928/do_while_stmt_15959/loop_exit/$entry
      -- CP-element group 12: 	 branch_block_stmt_15928/do_while_stmt_15959/loop_taken/$entry
      -- 
    nicRxFromMacDaemon_CP_30596_elements(12) <= nicRxFromMacDaemon_CP_30596_elements(17);
    -- CP-element group 13:  branch  place  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	78 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_15928/do_while_stmt_15959/loop_body_done
      -- 
    nicRxFromMacDaemon_CP_30596_elements(13) <= nicRxFromMacDaemon_CP_30596_elements(78);
    -- CP-element group 14:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	11 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	26 
    -- CP-element group 14: 	50 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/back_edge_to_loop_body
      -- 
    nicRxFromMacDaemon_CP_30596_elements(14) <= nicRxFromMacDaemon_CP_30596_elements(11);
    -- CP-element group 15:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	28 
    -- CP-element group 15: 	52 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/first_time_through_loop_body
      -- 
    nicRxFromMacDaemon_CP_30596_elements(15) <= nicRxFromMacDaemon_CP_30596_elements(9);
    -- CP-element group 16:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	39 
    -- CP-element group 16: 	23 
    -- CP-element group 16: 	44 
    -- CP-element group 16: 	45 
    -- CP-element group 16: 	18 
    -- CP-element group 16: 	22 
    -- CP-element group 16: 	77 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/$entry
      -- CP-element group 16: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/loop_body_start
      -- CP-element group 16: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15965_sample_start_
      -- 
    -- Element group nicRxFromMacDaemon_CP_30596_elements(16) is bound as output of CP function.
    -- CP-element group 17:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	21 
    -- CP-element group 17: 	77 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/condition_evaluated
      -- 
    condition_evaluated_30729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_30729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_30596_elements(17), ack => do_while_stmt_15959_branch_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 7);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_30596_elements(21) & nicRxFromMacDaemon_CP_30596_elements(77);
      gj_nicRxFromMacDaemon_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_30596_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	44 
    -- CP-element group 18: 	16 
    -- CP-element group 18: 	22 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	21 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	40 
    -- CP-element group 18: 	46 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/aggregated_phi_sample_req
      -- CP-element group 18: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15961_sample_start__ps
      -- 
    nicRxFromMacDaemon_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 7,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_30596_elements(44) & nicRxFromMacDaemon_CP_30596_elements(16) & nicRxFromMacDaemon_CP_30596_elements(22) & nicRxFromMacDaemon_CP_30596_elements(21);
      gj_nicRxFromMacDaemon_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_30596_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	42 
    -- CP-element group 19: 	24 
    -- CP-element group 19: 	47 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	78 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	44 
    -- CP-element group 19: 	22 
    -- CP-element group 19:  members (4) 
      -- CP-element group 19: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/aggregated_phi_sample_ack
      -- CP-element group 19: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15961_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15965_sample_completed_
      -- CP-element group 19: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15968_sample_completed_
      -- 
    nicRxFromMacDaemon_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 7,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_30596_elements(42) & nicRxFromMacDaemon_CP_30596_elements(24) & nicRxFromMacDaemon_CP_30596_elements(47);
      gj_nicRxFromMacDaemon_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_30596_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	39 
    -- CP-element group 20: 	23 
    -- CP-element group 20: 	45 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	41 
    -- CP-element group 20: 	48 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/aggregated_phi_update_req
      -- CP-element group 20: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15961_update_start__ps
      -- 
    nicRxFromMacDaemon_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_30596_elements(39) & nicRxFromMacDaemon_CP_30596_elements(23) & nicRxFromMacDaemon_CP_30596_elements(45);
      gj_nicRxFromMacDaemon_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_30596_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	25 
    -- CP-element group 21: 	43 
    -- CP-element group 21: 	49 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	17 
    -- CP-element group 21: marked-successors 
    -- CP-element group 21: 	18 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/aggregated_phi_update_ack
      -- 
    nicRxFromMacDaemon_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 7);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_30596_elements(25) & nicRxFromMacDaemon_CP_30596_elements(43) & nicRxFromMacDaemon_CP_30596_elements(49);
      gj_nicRxFromMacDaemon_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_30596_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	16 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	18 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15961_sample_start_
      -- 
    nicRxFromMacDaemon_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_30596_elements(16) & nicRxFromMacDaemon_CP_30596_elements(19);
      gj_nicRxFromMacDaemon_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_30596_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  join  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	16 
    -- CP-element group 23: marked-predecessors 
    -- CP-element group 23: 	65 
    -- CP-element group 23: 	25 
    -- CP-element group 23: 	68 
    -- CP-element group 23: 	75 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	20 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15961_update_start_
      -- 
    nicRxFromMacDaemon_cp_element_group_23: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 7,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_23"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_30596_elements(16) & nicRxFromMacDaemon_CP_30596_elements(65) & nicRxFromMacDaemon_CP_30596_elements(25) & nicRxFromMacDaemon_CP_30596_elements(68) & nicRxFromMacDaemon_CP_30596_elements(75);
      gj_nicRxFromMacDaemon_cp_element_group_23 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_30596_elements(23), clk => clk, reset => reset); --
    end block;
    -- CP-element group 24:  join  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	19 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15961_sample_completed__ps
      -- 
    -- Element group nicRxFromMacDaemon_CP_30596_elements(24) is bound as output of CP function.
    -- CP-element group 25:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	63 
    -- CP-element group 25: 	21 
    -- CP-element group 25: 	67 
    -- CP-element group 25: 	73 
    -- CP-element group 25: marked-successors 
    -- CP-element group 25: 	23 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15961_update_completed_
      -- CP-element group 25: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15961_update_completed__ps
      -- 
    -- Element group nicRxFromMacDaemon_CP_30596_elements(25) is bound as output of CP function.
    -- CP-element group 26:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	14 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15961_loopback_trigger
      -- 
    nicRxFromMacDaemon_CP_30596_elements(26) <= nicRxFromMacDaemon_CP_30596_elements(14);
    -- CP-element group 27:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15961_loopback_sample_req
      -- CP-element group 27: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15961_loopback_sample_req_ps
      -- 
    phi_stmt_15961_loopback_sample_req_30744_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_15961_loopback_sample_req_30744_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_30596_elements(27), ack => phi_stmt_15961_req_1); -- 
    -- Element group nicRxFromMacDaemon_CP_30596_elements(27) is bound as output of CP function.
    -- CP-element group 28:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	15 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15961_entry_trigger
      -- 
    nicRxFromMacDaemon_CP_30596_elements(28) <= nicRxFromMacDaemon_CP_30596_elements(15);
    -- CP-element group 29:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15961_entry_sample_req
      -- CP-element group 29: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15961_entry_sample_req_ps
      -- 
    phi_stmt_15961_entry_sample_req_30747_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_15961_entry_sample_req_30747_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_30596_elements(29), ack => phi_stmt_15961_req_0); -- 
    -- Element group nicRxFromMacDaemon_CP_30596_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15961_phi_mux_ack
      -- CP-element group 30: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15961_phi_mux_ack_ps
      -- 
    phi_stmt_15961_phi_mux_ack_30750_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_15961_ack_0, ack => nicRxFromMacDaemon_CP_30596_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_S0_15963_sample_start__ps
      -- CP-element group 31: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_S0_15963_sample_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_S0_15963_sample_start_
      -- CP-element group 31: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_S0_15963_sample_completed_
      -- 
    -- Element group nicRxFromMacDaemon_CP_30596_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_S0_15963_update_start__ps
      -- CP-element group 32: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_S0_15963_update_start_
      -- 
    -- Element group nicRxFromMacDaemon_CP_30596_elements(32) is bound as output of CP function.
    -- CP-element group 33:  join  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	34 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (1) 
      -- CP-element group 33: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_S0_15963_update_completed__ps
      -- 
    nicRxFromMacDaemon_CP_30596_elements(33) <= nicRxFromMacDaemon_CP_30596_elements(34);
    -- CP-element group 34:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	33 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_S0_15963_update_completed_
      -- 
    -- Element group nicRxFromMacDaemon_CP_30596_elements(34) is a control-delay.
    cp_element_34_delay: control_delay_element  generic map(name => " 34_delay", delay_value => 1)  port map(req => nicRxFromMacDaemon_CP_30596_elements(32), ack => nicRxFromMacDaemon_CP_30596_elements(34), clk => clk, reset =>reset);
    -- CP-element group 35:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_nLSTATE_15964_sample_start__ps
      -- CP-element group 35: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_nLSTATE_15964_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_nLSTATE_15964_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_nLSTATE_15964_Sample/req
      -- 
    req_30771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_30771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_30596_elements(35), ack => nLSTATE_15980_15964_buf_req_0); -- 
    -- Element group nicRxFromMacDaemon_CP_30596_elements(35) is bound as output of CP function.
    -- CP-element group 36:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_nLSTATE_15964_update_start__ps
      -- CP-element group 36: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_nLSTATE_15964_update_start_
      -- CP-element group 36: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_nLSTATE_15964_Update/$entry
      -- CP-element group 36: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_nLSTATE_15964_Update/req
      -- 
    req_30776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_30776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_30596_elements(36), ack => nLSTATE_15980_15964_buf_req_1); -- 
    -- Element group nicRxFromMacDaemon_CP_30596_elements(36) is bound as output of CP function.
    -- CP-element group 37:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (4) 
      -- CP-element group 37: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_nLSTATE_15964_sample_completed__ps
      -- CP-element group 37: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_nLSTATE_15964_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_nLSTATE_15964_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_nLSTATE_15964_Sample/ack
      -- 
    ack_30772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nLSTATE_15980_15964_buf_ack_0, ack => nicRxFromMacDaemon_CP_30596_elements(37)); -- 
    -- CP-element group 38:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_nLSTATE_15964_update_completed__ps
      -- CP-element group 38: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_nLSTATE_15964_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_nLSTATE_15964_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_nLSTATE_15964_Update/ack
      -- 
    ack_30777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nLSTATE_15980_15964_buf_ack_1, ack => nicRxFromMacDaemon_CP_30596_elements(38)); -- 
    -- CP-element group 39:  join  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	16 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	65 
    -- CP-element group 39: 	71 
    -- CP-element group 39: 	75 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	20 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15965_update_start_
      -- 
    nicRxFromMacDaemon_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_30596_elements(16) & nicRxFromMacDaemon_CP_30596_elements(65) & nicRxFromMacDaemon_CP_30596_elements(71) & nicRxFromMacDaemon_CP_30596_elements(75);
      gj_nicRxFromMacDaemon_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_30596_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	18 
    -- CP-element group 40: marked-predecessors 
    -- CP-element group 40: 	43 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	42 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/RPIPE_mac_to_nic_data_15967_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/RPIPE_mac_to_nic_data_15967_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/RPIPE_mac_to_nic_data_15967_Sample/rr
      -- 
    rr_30790_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_30790_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_30596_elements(40), ack => RPIPE_mac_to_nic_data_15967_inst_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_40: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_40"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_30596_elements(18) & nicRxFromMacDaemon_CP_30596_elements(43);
      gj_nicRxFromMacDaemon_cp_element_group_40 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_30596_elements(40), clk => clk, reset => reset); --
    end block;
    -- CP-element group 41:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	42 
    -- CP-element group 41: 	20 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	43 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/RPIPE_mac_to_nic_data_15967_update_start_
      -- CP-element group 41: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/RPIPE_mac_to_nic_data_15967_Update/$entry
      -- CP-element group 41: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/RPIPE_mac_to_nic_data_15967_Update/cr
      -- 
    cr_30795_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_30795_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_30596_elements(41), ack => RPIPE_mac_to_nic_data_15967_inst_req_1); -- 
    nicRxFromMacDaemon_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_30596_elements(42) & nicRxFromMacDaemon_CP_30596_elements(20);
      gj_nicRxFromMacDaemon_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_30596_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	40 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	41 
    -- CP-element group 42: 	19 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/RPIPE_mac_to_nic_data_15967_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/RPIPE_mac_to_nic_data_15967_Sample/$exit
      -- CP-element group 42: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/RPIPE_mac_to_nic_data_15967_Sample/ra
      -- 
    ra_30791_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_mac_to_nic_data_15967_inst_ack_0, ack => nicRxFromMacDaemon_CP_30596_elements(42)); -- 
    -- CP-element group 43:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	63 
    -- CP-element group 43: 	21 
    -- CP-element group 43: 	70 
    -- CP-element group 43: 	73 
    -- CP-element group 43: marked-successors 
    -- CP-element group 43: 	40 
    -- CP-element group 43:  members (4) 
      -- CP-element group 43: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15965_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/RPIPE_mac_to_nic_data_15967_update_completed_
      -- CP-element group 43: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/RPIPE_mac_to_nic_data_15967_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/RPIPE_mac_to_nic_data_15967_Update/ca
      -- 
    ca_30796_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_mac_to_nic_data_15967_inst_ack_1, ack => nicRxFromMacDaemon_CP_30596_elements(43)); -- 
    -- CP-element group 44:  join  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	16 
    -- CP-element group 44: marked-predecessors 
    -- CP-element group 44: 	19 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	18 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15968_sample_start_
      -- 
    nicRxFromMacDaemon_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 7,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_30596_elements(16) & nicRxFromMacDaemon_CP_30596_elements(19);
      gj_nicRxFromMacDaemon_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_30596_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  join  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	16 
    -- CP-element group 45: marked-predecessors 
    -- CP-element group 45: 	49 
    -- CP-element group 45: 	75 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	20 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15968_update_start_
      -- 
    nicRxFromMacDaemon_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_30596_elements(16) & nicRxFromMacDaemon_CP_30596_elements(49) & nicRxFromMacDaemon_CP_30596_elements(75);
      gj_nicRxFromMacDaemon_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_30596_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	18 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (1) 
      -- CP-element group 46: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15968_sample_start__ps
      -- 
    nicRxFromMacDaemon_CP_30596_elements(46) <= nicRxFromMacDaemon_CP_30596_elements(18);
    -- CP-element group 47:  join  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	19 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15968_sample_completed__ps
      -- 
    -- Element group nicRxFromMacDaemon_CP_30596_elements(47) is bound as output of CP function.
    -- CP-element group 48:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	20 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15968_update_start__ps
      -- 
    nicRxFromMacDaemon_CP_30596_elements(48) <= nicRxFromMacDaemon_CP_30596_elements(20);
    -- CP-element group 49:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	21 
    -- CP-element group 49: 	73 
    -- CP-element group 49: marked-successors 
    -- CP-element group 49: 	45 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15968_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15968_update_completed__ps
      -- 
    -- Element group nicRxFromMacDaemon_CP_30596_elements(49) is bound as output of CP function.
    -- CP-element group 50:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	14 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15968_loopback_trigger
      -- 
    nicRxFromMacDaemon_CP_30596_elements(50) <= nicRxFromMacDaemon_CP_30596_elements(14);
    -- CP-element group 51:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (2) 
      -- CP-element group 51: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15968_loopback_sample_req
      -- CP-element group 51: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15968_loopback_sample_req_ps
      -- 
    phi_stmt_15968_loopback_sample_req_30806_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_15968_loopback_sample_req_30806_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_30596_elements(51), ack => phi_stmt_15968_req_1); -- 
    -- Element group nicRxFromMacDaemon_CP_30596_elements(51) is bound as output of CP function.
    -- CP-element group 52:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	15 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15968_entry_trigger
      -- 
    nicRxFromMacDaemon_CP_30596_elements(52) <= nicRxFromMacDaemon_CP_30596_elements(15);
    -- CP-element group 53:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (2) 
      -- CP-element group 53: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15968_entry_sample_req
      -- CP-element group 53: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15968_entry_sample_req_ps
      -- 
    phi_stmt_15968_entry_sample_req_30809_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_15968_entry_sample_req_30809_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_30596_elements(53), ack => phi_stmt_15968_req_0); -- 
    -- Element group nicRxFromMacDaemon_CP_30596_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (2) 
      -- CP-element group 54: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15968_phi_mux_ack
      -- CP-element group 54: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/phi_stmt_15968_phi_mux_ack_ps
      -- 
    phi_stmt_15968_phi_mux_ack_30812_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_15968_ack_0, ack => nicRxFromMacDaemon_CP_30596_elements(54)); -- 
    -- CP-element group 55:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/type_cast_15971_sample_start__ps
      -- CP-element group 55: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/type_cast_15971_sample_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/type_cast_15971_sample_start_
      -- CP-element group 55: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/type_cast_15971_sample_completed_
      -- 
    -- Element group nicRxFromMacDaemon_CP_30596_elements(55) is bound as output of CP function.
    -- CP-element group 56:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (2) 
      -- CP-element group 56: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/type_cast_15971_update_start__ps
      -- CP-element group 56: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/type_cast_15971_update_start_
      -- 
    -- Element group nicRxFromMacDaemon_CP_30596_elements(56) is bound as output of CP function.
    -- CP-element group 57:  join  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: successors 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/type_cast_15971_update_completed__ps
      -- 
    nicRxFromMacDaemon_CP_30596_elements(57) <= nicRxFromMacDaemon_CP_30596_elements(58);
    -- CP-element group 58:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	57 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/type_cast_15971_update_completed_
      -- 
    -- Element group nicRxFromMacDaemon_CP_30596_elements(58) is a control-delay.
    cp_element_58_delay: control_delay_element  generic map(name => " 58_delay", delay_value => 1)  port map(req => nicRxFromMacDaemon_CP_30596_elements(56), ack => nicRxFromMacDaemon_CP_30596_elements(58), clk => clk, reset =>reset);
    -- CP-element group 59:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (4) 
      -- CP-element group 59: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_npkt_cnt_15972_sample_start__ps
      -- CP-element group 59: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_npkt_cnt_15972_sample_start_
      -- CP-element group 59: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_npkt_cnt_15972_Sample/$entry
      -- CP-element group 59: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_npkt_cnt_15972_Sample/req
      -- 
    req_30833_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_30833_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_30596_elements(59), ack => npkt_cnt_16018_15972_buf_req_0); -- 
    -- Element group nicRxFromMacDaemon_CP_30596_elements(59) is bound as output of CP function.
    -- CP-element group 60:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (4) 
      -- CP-element group 60: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_npkt_cnt_15972_update_start__ps
      -- CP-element group 60: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_npkt_cnt_15972_update_start_
      -- CP-element group 60: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_npkt_cnt_15972_Update/$entry
      -- CP-element group 60: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_npkt_cnt_15972_Update/req
      -- 
    req_30838_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_30838_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_30596_elements(60), ack => npkt_cnt_16018_15972_buf_req_1); -- 
    -- Element group nicRxFromMacDaemon_CP_30596_elements(60) is bound as output of CP function.
    -- CP-element group 61:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (4) 
      -- CP-element group 61: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_npkt_cnt_15972_sample_completed__ps
      -- CP-element group 61: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_npkt_cnt_15972_sample_completed_
      -- CP-element group 61: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_npkt_cnt_15972_Sample/$exit
      -- CP-element group 61: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_npkt_cnt_15972_Sample/ack
      -- 
    ack_30834_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => npkt_cnt_16018_15972_buf_ack_0, ack => nicRxFromMacDaemon_CP_30596_elements(61)); -- 
    -- CP-element group 62:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (4) 
      -- CP-element group 62: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_npkt_cnt_15972_update_completed__ps
      -- CP-element group 62: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_npkt_cnt_15972_update_completed_
      -- CP-element group 62: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_npkt_cnt_15972_Update/$exit
      -- CP-element group 62: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/R_npkt_cnt_15972_Update/ack
      -- 
    ack_30839_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => npkt_cnt_16018_15972_buf_ack_1, ack => nicRxFromMacDaemon_CP_30596_elements(62)); -- 
    -- CP-element group 63:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	25 
    -- CP-element group 63: 	43 
    -- CP-element group 63: marked-predecessors 
    -- CP-element group 63: 	65 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/MUX_16000_sample_start_
      -- CP-element group 63: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/MUX_16000_start/$entry
      -- CP-element group 63: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/MUX_16000_start/req
      -- 
    req_30848_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_30848_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_30596_elements(63), ack => MUX_16000_inst_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_30596_elements(25) & nicRxFromMacDaemon_CP_30596_elements(43) & nicRxFromMacDaemon_CP_30596_elements(65);
      gj_nicRxFromMacDaemon_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_30596_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: marked-predecessors 
    -- CP-element group 64: 	66 
    -- CP-element group 64: 	68 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/MUX_16000_update_start_
      -- CP-element group 64: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/MUX_16000_complete/$entry
      -- CP-element group 64: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/MUX_16000_complete/req
      -- 
    req_30853_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_30853_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_30596_elements(64), ack => MUX_16000_inst_req_1); -- 
    nicRxFromMacDaemon_cp_element_group_64: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_64"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_30596_elements(66) & nicRxFromMacDaemon_CP_30596_elements(68);
      gj_nicRxFromMacDaemon_cp_element_group_64 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_30596_elements(64), clk => clk, reset => reset); --
    end block;
    -- CP-element group 65:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: marked-successors 
    -- CP-element group 65: 	39 
    -- CP-element group 65: 	63 
    -- CP-element group 65: 	23 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/MUX_16000_sample_completed_
      -- CP-element group 65: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/MUX_16000_start/$exit
      -- CP-element group 65: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/MUX_16000_start/ack
      -- 
    ack_30849_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_16000_inst_ack_0, ack => nicRxFromMacDaemon_CP_30596_elements(65)); -- 
    -- CP-element group 66:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	64 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/MUX_16000_update_completed_
      -- CP-element group 66: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/MUX_16000_complete/$exit
      -- CP-element group 66: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/MUX_16000_complete/ack
      -- 
    ack_30854_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => MUX_16000_inst_ack_1, ack => nicRxFromMacDaemon_CP_30596_elements(66)); -- 
    -- CP-element group 67:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	25 
    -- CP-element group 67: 	66 
    -- CP-element group 67: marked-predecessors 
    -- CP-element group 67: 	69 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	68 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/WPIPE_nic_rx_to_header_15991_sample_start_
      -- CP-element group 67: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/WPIPE_nic_rx_to_header_15991_Sample/$entry
      -- CP-element group 67: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/WPIPE_nic_rx_to_header_15991_Sample/req
      -- 
    req_30862_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_30862_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_30596_elements(67), ack => WPIPE_nic_rx_to_header_15991_inst_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 7,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_30596_elements(25) & nicRxFromMacDaemon_CP_30596_elements(66) & nicRxFromMacDaemon_CP_30596_elements(69);
      gj_nicRxFromMacDaemon_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_30596_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	67 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	69 
    -- CP-element group 68: marked-successors 
    -- CP-element group 68: 	64 
    -- CP-element group 68: 	23 
    -- CP-element group 68:  members (6) 
      -- CP-element group 68: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/WPIPE_nic_rx_to_header_15991_sample_completed_
      -- CP-element group 68: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/WPIPE_nic_rx_to_header_15991_update_start_
      -- CP-element group 68: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/WPIPE_nic_rx_to_header_15991_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/WPIPE_nic_rx_to_header_15991_Sample/ack
      -- CP-element group 68: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/WPIPE_nic_rx_to_header_15991_Update/$entry
      -- CP-element group 68: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/WPIPE_nic_rx_to_header_15991_Update/req
      -- 
    ack_30863_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_rx_to_header_15991_inst_ack_0, ack => nicRxFromMacDaemon_CP_30596_elements(68)); -- 
    req_30867_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_30867_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_30596_elements(68), ack => WPIPE_nic_rx_to_header_15991_inst_req_1); -- 
    -- CP-element group 69:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	68 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	78 
    -- CP-element group 69: marked-successors 
    -- CP-element group 69: 	67 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/WPIPE_nic_rx_to_header_15991_update_completed_
      -- CP-element group 69: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/WPIPE_nic_rx_to_header_15991_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/WPIPE_nic_rx_to_header_15991_Update/ack
      -- 
    ack_30868_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_rx_to_header_15991_inst_ack_1, ack => nicRxFromMacDaemon_CP_30596_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	43 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	72 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	71 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/WPIPE_nic_rx_to_packet_16002_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/WPIPE_nic_rx_to_packet_16002_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/WPIPE_nic_rx_to_packet_16002_Sample/req
      -- 
    req_30876_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_30876_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_30596_elements(70), ack => WPIPE_nic_rx_to_packet_16002_inst_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_30596_elements(43) & nicRxFromMacDaemon_CP_30596_elements(72);
      gj_nicRxFromMacDaemon_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_30596_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	70 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71: marked-successors 
    -- CP-element group 71: 	39 
    -- CP-element group 71:  members (6) 
      -- CP-element group 71: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/WPIPE_nic_rx_to_packet_16002_sample_completed_
      -- CP-element group 71: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/WPIPE_nic_rx_to_packet_16002_update_start_
      -- CP-element group 71: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/WPIPE_nic_rx_to_packet_16002_Sample/$exit
      -- CP-element group 71: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/WPIPE_nic_rx_to_packet_16002_Sample/ack
      -- CP-element group 71: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/WPIPE_nic_rx_to_packet_16002_Update/$entry
      -- CP-element group 71: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/WPIPE_nic_rx_to_packet_16002_Update/req
      -- 
    ack_30877_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_rx_to_packet_16002_inst_ack_0, ack => nicRxFromMacDaemon_CP_30596_elements(71)); -- 
    req_30881_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_30881_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_30596_elements(71), ack => WPIPE_nic_rx_to_packet_16002_inst_req_1); -- 
    -- CP-element group 72:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	71 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	78 
    -- CP-element group 72: marked-successors 
    -- CP-element group 72: 	70 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/WPIPE_nic_rx_to_packet_16002_update_completed_
      -- CP-element group 72: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/WPIPE_nic_rx_to_packet_16002_Update/$exit
      -- CP-element group 72: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/WPIPE_nic_rx_to_packet_16002_Update/ack
      -- 
    ack_30882_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_rx_to_packet_16002_inst_ack_1, ack => nicRxFromMacDaemon_CP_30596_elements(72)); -- 
    -- CP-element group 73:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	25 
    -- CP-element group 73: 	43 
    -- CP-element group 73: 	49 
    -- CP-element group 73: marked-predecessors 
    -- CP-element group 73: 	75 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/call_stmt_16028_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/call_stmt_16028_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/call_stmt_16028_Sample/crr
      -- 
    crr_30890_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_30890_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_30596_elements(73), ack => call_stmt_16028_call_req_0); -- 
    nicRxFromMacDaemon_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 1,2 => 7,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_30596_elements(25) & nicRxFromMacDaemon_CP_30596_elements(43) & nicRxFromMacDaemon_CP_30596_elements(49) & nicRxFromMacDaemon_CP_30596_elements(75);
      gj_nicRxFromMacDaemon_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_30596_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	76 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/call_stmt_16028_update_start_
      -- CP-element group 74: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/call_stmt_16028_Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/call_stmt_16028_Update/ccr
      -- 
    ccr_30895_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_30895_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_30596_elements(74), ack => call_stmt_16028_call_req_1); -- 
    nicRxFromMacDaemon_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= nicRxFromMacDaemon_CP_30596_elements(76);
      gj_nicRxFromMacDaemon_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_30596_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	39 
    -- CP-element group 75: 	23 
    -- CP-element group 75: 	45 
    -- CP-element group 75: 	73 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/call_stmt_16028_sample_completed_
      -- CP-element group 75: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/call_stmt_16028_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/call_stmt_16028_Sample/cra
      -- 
    cra_30891_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_16028_call_ack_0, ack => nicRxFromMacDaemon_CP_30596_elements(75)); -- 
    -- CP-element group 76:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76: marked-successors 
    -- CP-element group 76: 	74 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/call_stmt_16028_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/call_stmt_16028_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/call_stmt_16028_Update/cca
      -- 
    cca_30896_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_16028_call_ack_1, ack => nicRxFromMacDaemon_CP_30596_elements(76)); -- 
    -- CP-element group 77:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	16 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	17 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group nicRxFromMacDaemon_CP_30596_elements(77) is a control-delay.
    cp_element_77_delay: control_delay_element  generic map(name => " 77_delay", delay_value => 1)  port map(req => nicRxFromMacDaemon_CP_30596_elements(16), ack => nicRxFromMacDaemon_CP_30596_elements(77), clk => clk, reset =>reset);
    -- CP-element group 78:  join  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	19 
    -- CP-element group 78: 	69 
    -- CP-element group 78: 	72 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	13 
    -- CP-element group 78:  members (1) 
      -- CP-element group 78: 	 branch_block_stmt_15928/do_while_stmt_15959/do_while_stmt_15959_loop_body/$exit
      -- 
    nicRxFromMacDaemon_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 7,1 => 7,2 => 7,3 => 7);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 38) := "nicRxFromMacDaemon_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= nicRxFromMacDaemon_CP_30596_elements(19) & nicRxFromMacDaemon_CP_30596_elements(69) & nicRxFromMacDaemon_CP_30596_elements(72) & nicRxFromMacDaemon_CP_30596_elements(76);
      gj_nicRxFromMacDaemon_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => nicRxFromMacDaemon_CP_30596_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  transition  input  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	12 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (2) 
      -- CP-element group 79: 	 branch_block_stmt_15928/do_while_stmt_15959/loop_exit/$exit
      -- CP-element group 79: 	 branch_block_stmt_15928/do_while_stmt_15959/loop_exit/ack
      -- 
    ack_30901_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_15959_branch_ack_0, ack => nicRxFromMacDaemon_CP_30596_elements(79)); -- 
    -- CP-element group 80:  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	12 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_15928/do_while_stmt_15959/loop_taken/$exit
      -- CP-element group 80: 	 branch_block_stmt_15928/do_while_stmt_15959/loop_taken/ack
      -- 
    ack_30905_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_15959_branch_ack_1, ack => nicRxFromMacDaemon_CP_30596_elements(80)); -- 
    -- CP-element group 81:  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	10 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	2 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_15928/do_while_stmt_15959/$exit
      -- 
    nicRxFromMacDaemon_CP_30596_elements(81) <= nicRxFromMacDaemon_CP_30596_elements(10);
    -- CP-element group 82:  merge  fork  transition  place  output  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	5 
    -- CP-element group 82: 	0 
    -- CP-element group 82: 	2 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	3 
    -- CP-element group 82: 	4 
    -- CP-element group 82:  members (13) 
      -- CP-element group 82: 	 branch_block_stmt_15928/merge_stmt_15930_PhiAck/$entry
      -- CP-element group 82: 	 branch_block_stmt_15928/merge_stmt_15930_PhiAck/$exit
      -- CP-element group 82: 	 branch_block_stmt_15928/merge_stmt_15930__exit__
      -- CP-element group 82: 	 branch_block_stmt_15928/call_stmt_15940__entry__
      -- CP-element group 82: 	 branch_block_stmt_15928/call_stmt_15940/$entry
      -- CP-element group 82: 	 branch_block_stmt_15928/call_stmt_15940/call_stmt_15940_sample_start_
      -- CP-element group 82: 	 branch_block_stmt_15928/call_stmt_15940/call_stmt_15940_update_start_
      -- CP-element group 82: 	 branch_block_stmt_15928/call_stmt_15940/call_stmt_15940_Sample/$entry
      -- CP-element group 82: 	 branch_block_stmt_15928/call_stmt_15940/call_stmt_15940_Sample/crr
      -- CP-element group 82: 	 branch_block_stmt_15928/call_stmt_15940/call_stmt_15940_Update/$entry
      -- CP-element group 82: 	 branch_block_stmt_15928/call_stmt_15940/call_stmt_15940_Update/ccr
      -- CP-element group 82: 	 branch_block_stmt_15928/merge_stmt_15930_PhiAck/dummy
      -- CP-element group 82: 	 branch_block_stmt_15928/merge_stmt_15930_PhiReqMerge
      -- 
    crr_30625_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_30625_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_30596_elements(82), ack => call_stmt_15940_call_req_0); -- 
    ccr_30630_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_30630_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nicRxFromMacDaemon_CP_30596_elements(82), ack => call_stmt_15940_call_req_1); -- 
    nicRxFromMacDaemon_CP_30596_elements(82) <= OrReduce(nicRxFromMacDaemon_CP_30596_elements(5) & nicRxFromMacDaemon_CP_30596_elements(0) & nicRxFromMacDaemon_CP_30596_elements(2));
    nicRxFromMacDaemon_do_while_stmt_15959_terminator_30906: loop_terminator -- 
      generic map (name => " nicRxFromMacDaemon_do_while_stmt_15959_terminator_30906", max_iterations_in_flight =>7) 
      port map(loop_body_exit => nicRxFromMacDaemon_CP_30596_elements(13),loop_continue => nicRxFromMacDaemon_CP_30596_elements(80),loop_terminate => nicRxFromMacDaemon_CP_30596_elements(79),loop_back => nicRxFromMacDaemon_CP_30596_elements(11),loop_exit => nicRxFromMacDaemon_CP_30596_elements(10),clk => clk, reset => reset); -- 
    phi_stmt_15961_phi_seq_30778_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= nicRxFromMacDaemon_CP_30596_elements(28);
      nicRxFromMacDaemon_CP_30596_elements(31)<= src_sample_reqs(0);
      src_sample_acks(0)  <= nicRxFromMacDaemon_CP_30596_elements(31);
      nicRxFromMacDaemon_CP_30596_elements(32)<= src_update_reqs(0);
      src_update_acks(0)  <= nicRxFromMacDaemon_CP_30596_elements(33);
      nicRxFromMacDaemon_CP_30596_elements(29) <= phi_mux_reqs(0);
      triggers(1)  <= nicRxFromMacDaemon_CP_30596_elements(26);
      nicRxFromMacDaemon_CP_30596_elements(35)<= src_sample_reqs(1);
      src_sample_acks(1)  <= nicRxFromMacDaemon_CP_30596_elements(37);
      nicRxFromMacDaemon_CP_30596_elements(36)<= src_update_reqs(1);
      src_update_acks(1)  <= nicRxFromMacDaemon_CP_30596_elements(38);
      nicRxFromMacDaemon_CP_30596_elements(27) <= phi_mux_reqs(1);
      phi_stmt_15961_phi_seq_30778 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_15961_phi_seq_30778") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => nicRxFromMacDaemon_CP_30596_elements(18), 
          phi_sample_ack => nicRxFromMacDaemon_CP_30596_elements(24), 
          phi_update_req => nicRxFromMacDaemon_CP_30596_elements(20), 
          phi_update_ack => nicRxFromMacDaemon_CP_30596_elements(25), 
          phi_mux_ack => nicRxFromMacDaemon_CP_30596_elements(30), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_15968_phi_seq_30840_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= nicRxFromMacDaemon_CP_30596_elements(52);
      nicRxFromMacDaemon_CP_30596_elements(55)<= src_sample_reqs(0);
      src_sample_acks(0)  <= nicRxFromMacDaemon_CP_30596_elements(55);
      nicRxFromMacDaemon_CP_30596_elements(56)<= src_update_reqs(0);
      src_update_acks(0)  <= nicRxFromMacDaemon_CP_30596_elements(57);
      nicRxFromMacDaemon_CP_30596_elements(53) <= phi_mux_reqs(0);
      triggers(1)  <= nicRxFromMacDaemon_CP_30596_elements(50);
      nicRxFromMacDaemon_CP_30596_elements(59)<= src_sample_reqs(1);
      src_sample_acks(1)  <= nicRxFromMacDaemon_CP_30596_elements(61);
      nicRxFromMacDaemon_CP_30596_elements(60)<= src_update_reqs(1);
      src_update_acks(1)  <= nicRxFromMacDaemon_CP_30596_elements(62);
      nicRxFromMacDaemon_CP_30596_elements(51) <= phi_mux_reqs(1);
      phi_stmt_15968_phi_seq_30840 : phi_sequencer_v2-- 
        generic map (place_capacity => 7, ntriggers => 2, name => "phi_stmt_15968_phi_seq_30840") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => nicRxFromMacDaemon_CP_30596_elements(46), 
          phi_sample_ack => nicRxFromMacDaemon_CP_30596_elements(47), 
          phi_update_req => nicRxFromMacDaemon_CP_30596_elements(48), 
          phi_update_ack => nicRxFromMacDaemon_CP_30596_elements(49), 
          phi_mux_ack => nicRxFromMacDaemon_CP_30596_elements(54), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_30730_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= nicRxFromMacDaemon_CP_30596_elements(14);
        preds(1)  <= nicRxFromMacDaemon_CP_30596_elements(15);
        entry_tmerge_30730 : transition_merge -- 
          generic map(name => " entry_tmerge_30730")
          port map (preds => preds, symbol_out => nicRxFromMacDaemon_CP_30596_elements(16));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_16015_wire : std_logic_vector(31 downto 0);
    signal BITSEL_u32_u1_15944_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_16035_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u65_u73_15998_wire : std_logic_vector(72 downto 0);
    signal EQ_u2_u1_15984_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_15987_wire : std_logic_vector(0 downto 0);
    signal EQ_u2_u1_15994_wire : std_logic_vector(0 downto 0);
    signal LSTATE_15961 : std_logic_vector(1 downto 0);
    signal MUX_16000_wire : std_logic_vector(72 downto 0);
    signal NOT_u1_u1_15945_wire : std_logic_vector(0 downto 0);
    signal NOT_u4_u4_15935_wire_constant : std_logic_vector(3 downto 0);
    signal NOT_u4_u4_15953_wire_constant : std_logic_vector(3 downto 0);
    signal NOT_u4_u4_16024_wire_constant : std_logic_vector(3 downto 0);
    signal RPIPE_CONTROL_REGISTER_15942_wire : std_logic_vector(31 downto 0);
    signal RPIPE_CONTROL_REGISTER_16033_wire : std_logic_vector(31 downto 0);
    signal RPIPE_mac_to_nic_data_15967_wire : std_logic_vector(72 downto 0);
    signal RX_15965 : std_logic_vector(72 downto 0);
    signal R_HEADER_TKEEP_15997_wire_constant : std_logic_vector(7 downto 0);
    signal R_S0_15963_wire_constant : std_logic_vector(1 downto 0);
    signal R_S0_15983_wire_constant : std_logic_vector(1 downto 0);
    signal R_S0_16007_wire_constant : std_logic_vector(1 downto 0);
    signal R_S1_15986_wire_constant : std_logic_vector(1 downto 0);
    signal R_S1_15993_wire_constant : std_logic_vector(1 downto 0);
    signal ignore_resp0_15940 : std_logic_vector(31 downto 0);
    signal ignore_resp1_15958 : std_logic_vector(31 downto 0);
    signal ignore_resp2_16028 : std_logic_vector(31 downto 0);
    signal konst_15936_wire_constant : std_logic_vector(5 downto 0);
    signal konst_15943_wire_constant : std_logic_vector(31 downto 0);
    signal konst_15954_wire_constant : std_logic_vector(5 downto 0);
    signal konst_16025_wire_constant : std_logic_vector(5 downto 0);
    signal konst_16034_wire_constant : std_logic_vector(31 downto 0);
    signal nLSTATE_15980 : std_logic_vector(1 downto 0);
    signal nLSTATE_15980_15964_buffered : std_logic_vector(1 downto 0);
    signal npkt_cnt_16018 : std_logic_vector(31 downto 0);
    signal npkt_cnt_16018_15972_buffered : std_logic_vector(31 downto 0);
    signal pkt_cnt_15968 : std_logic_vector(31 downto 0);
    signal pkt_complete_16009 : std_logic_vector(0 downto 0);
    signal slice_15996_wire : std_logic_vector(64 downto 0);
    signal type_cast_15932_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_15938_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_15950_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_15956_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_15971_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_16014_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_16021_wire_constant : std_logic_vector(0 downto 0);
    signal write_to_header_15989 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    NOT_u4_u4_15935_wire_constant <= "1111";
    NOT_u4_u4_15953_wire_constant <= "1111";
    NOT_u4_u4_16024_wire_constant <= "1111";
    R_HEADER_TKEEP_15997_wire_constant <= "00111111";
    R_S0_15963_wire_constant <= "00";
    R_S0_15983_wire_constant <= "00";
    R_S0_16007_wire_constant <= "00";
    R_S1_15986_wire_constant <= "01";
    R_S1_15993_wire_constant <= "01";
    konst_15936_wire_constant <= "010110";
    konst_15943_wire_constant <= "00000000000000000000000000000000";
    konst_15954_wire_constant <= "010110";
    konst_16025_wire_constant <= "010111";
    konst_16034_wire_constant <= "00000000000000000000000000000000";
    type_cast_15932_wire_constant <= "0";
    type_cast_15938_wire_constant <= "00000000000000000000000000000000";
    type_cast_15950_wire_constant <= "0";
    type_cast_15956_wire_constant <= "00000000000000000000000000000001";
    type_cast_15971_wire_constant <= "00000000000000000000000000000000";
    type_cast_16014_wire_constant <= "00000000000000000000000000000001";
    type_cast_16021_wire_constant <= "0";
    phi_stmt_15961: Block -- phi operator 
      signal idata: std_logic_vector(3 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= R_S0_15963_wire_constant & nLSTATE_15980_15964_buffered;
      req <= phi_stmt_15961_req_0 & phi_stmt_15961_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_15961",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 2) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_15961_ack_0,
          idata => idata,
          odata => LSTATE_15961,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_15961
    phi_stmt_15968: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_15971_wire_constant & npkt_cnt_16018_15972_buffered;
      req <= phi_stmt_15968_req_0 & phi_stmt_15968_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_15968",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_15968_ack_0,
          idata => idata,
          odata => pkt_cnt_15968,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_15968
    MUX_16000_inst_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      signal sample_req_ug, sample_ack_ug, update_req_ug, update_ack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      sample_req_ug(0) <= MUX_16000_inst_req_0;
      MUX_16000_inst_ack_0<= sample_ack_ug(0);
      update_req_ug(0) <= MUX_16000_inst_req_1;
      MUX_16000_inst_ack_1<= update_ack_ug(0);
      guard_vector(0) <=  write_to_header_15989(0);
      MUX_16000_inst_gI: SplitGuardInterface generic map(name => "MUX_16000_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_ug,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_ug,
        cr_in => update_req_ug,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_ug,
        guards => guard_vector); -- 
      MUX_16000_inst: SelectSplitProtocol generic map(name => "MUX_16000_inst", data_width => 73, buffering => 1, flow_through => false, full_rate => true) -- 
        port map( x => CONCAT_u65_u73_15998_wire, y => RX_15965, sel => EQ_u2_u1_15994_wire, z => MUX_16000_wire, sample_req => sample_req(0), sample_ack => sample_ack(0), update_req => update_req(0), update_ack => update_ack(0), clk => clk, reset => reset); -- 
      -- 
    end block;
    -- flow-through select operator MUX_16017_inst
    npkt_cnt_16018 <= ADD_u32_u32_16015_wire when (pkt_complete_16009(0) /=  '0') else pkt_cnt_15968;
    -- flow-through slice operator slice_15996_inst
    slice_15996_wire <= RX_15965(72 downto 8);
    nLSTATE_15980_15964_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nLSTATE_15980_15964_buf_req_0;
      nLSTATE_15980_15964_buf_ack_0<= wack(0);
      rreq(0) <= nLSTATE_15980_15964_buf_req_1;
      nLSTATE_15980_15964_buf_ack_1<= rack(0);
      nLSTATE_15980_15964_buf : InterlockBuffer generic map ( -- 
        name => "nLSTATE_15980_15964_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 2,
        out_data_width => 2,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nLSTATE_15980,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nLSTATE_15980_15964_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    npkt_cnt_16018_15972_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= npkt_cnt_16018_15972_buf_req_0;
      npkt_cnt_16018_15972_buf_ack_0<= wack(0);
      rreq(0) <= npkt_cnt_16018_15972_buf_req_1;
      npkt_cnt_16018_15972_buf_ack_1<= rack(0);
      npkt_cnt_16018_15972_buf : InterlockBuffer generic map ( -- 
        name => "npkt_cnt_16018_15972_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => npkt_cnt_16018,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => npkt_cnt_16018_15972_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_15965
    process(RPIPE_mac_to_nic_data_15967_wire) -- 
      variable tmp_var : std_logic_vector(72 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 72 downto 0) := RPIPE_mac_to_nic_data_15967_wire(72 downto 0);
      RX_15965 <= tmp_var; -- 
    end process;
    do_while_stmt_15959_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= BITSEL_u32_u1_16035_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_15959_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_15959_branch_req_0,
          ack0 => do_while_stmt_15959_branch_ack_0,
          ack1 => do_while_stmt_15959_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_15941_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_15945_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_15941_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_15941_branch_req_0,
          ack0 => if_stmt_15941_branch_ack_0,
          ack1 => if_stmt_15941_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u32_u32_16015_inst
    process(pkt_cnt_15968) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(pkt_cnt_15968, type_cast_16014_wire_constant, tmp_var);
      ADD_u32_u32_16015_wire <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_15944_inst
    process(RPIPE_CONTROL_REGISTER_15942_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_CONTROL_REGISTER_15942_wire, konst_15943_wire_constant, tmp_var);
      BITSEL_u32_u1_15944_wire <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_16035_inst
    process(RPIPE_CONTROL_REGISTER_16033_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_CONTROL_REGISTER_16033_wire, konst_16034_wire_constant, tmp_var);
      BITSEL_u32_u1_16035_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u65_u73_15998_inst
    process(slice_15996_wire) -- 
      variable tmp_var : std_logic_vector(72 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_15996_wire, R_HEADER_TKEEP_15997_wire_constant, tmp_var);
      CONCAT_u65_u73_15998_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_15984_inst
    process(LSTATE_15961) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_15961, R_S0_15983_wire_constant, tmp_var);
      EQ_u2_u1_15984_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_15987_inst
    process(LSTATE_15961) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_15961, R_S1_15986_wire_constant, tmp_var);
      EQ_u2_u1_15987_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_15994_inst
    process(LSTATE_15961) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(LSTATE_15961, R_S1_15993_wire_constant, tmp_var);
      EQ_u2_u1_15994_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u2_u1_16008_inst
    process(nLSTATE_15980) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(nLSTATE_15980, R_S0_16007_wire_constant, tmp_var);
      pkt_complete_16009 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_15945_inst
    process(BITSEL_u32_u1_15944_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", BITSEL_u32_u1_15944_wire, tmp_var);
      NOT_u1_u1_15945_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_15988_inst
    process(EQ_u2_u1_15984_wire, EQ_u2_u1_15987_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u2_u1_15984_wire, EQ_u2_u1_15987_wire, tmp_var);
      write_to_header_15989 <= tmp_var; --
    end process;
    -- read from input-signal CONTROL_REGISTER
    RPIPE_CONTROL_REGISTER_15942_wire <= CONTROL_REGISTER;
    -- read from input-signal CONTROL_REGISTER
    RPIPE_CONTROL_REGISTER_16033_wire <= CONTROL_REGISTER;
    -- shared inport operator group (2) : RPIPE_mac_to_nic_data_15967_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(72 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_mac_to_nic_data_15967_inst_req_0;
      RPIPE_mac_to_nic_data_15967_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_mac_to_nic_data_15967_inst_req_1;
      RPIPE_mac_to_nic_data_15967_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_mac_to_nic_data_15967_wire <= data_out(72 downto 0);
      mac_to_nic_data_read_2_gI: SplitGuardInterface generic map(name => "mac_to_nic_data_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      mac_to_nic_data_read_2: InputPortRevised -- 
        generic map ( name => "mac_to_nic_data_read_2", data_width => 73,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => mac_to_nic_data_pipe_read_req(0),
          oack => mac_to_nic_data_pipe_read_ack(0),
          odata => mac_to_nic_data_pipe_read_data(72 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared outport operator group (0) : WPIPE_nic_rx_to_header_15991_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_nic_rx_to_header_15991_inst_req_0;
      WPIPE_nic_rx_to_header_15991_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_nic_rx_to_header_15991_inst_req_1;
      WPIPE_nic_rx_to_header_15991_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= write_to_header_15989(0);
      data_in <= MUX_16000_wire;
      nic_rx_to_header_write_0_gI: SplitGuardInterface generic map(name => "nic_rx_to_header_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      nic_rx_to_header_write_0: OutputPortRevised -- 
        generic map ( name => "nic_rx_to_header", data_width => 73, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => nic_rx_to_header_pipe_write_req(0),
          oack => nic_rx_to_header_pipe_write_ack(0),
          odata => nic_rx_to_header_pipe_write_data(72 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_nic_rx_to_packet_16002_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_nic_rx_to_packet_16002_inst_req_0;
      WPIPE_nic_rx_to_packet_16002_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_nic_rx_to_packet_16002_inst_req_1;
      WPIPE_nic_rx_to_packet_16002_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= RX_15965;
      nic_rx_to_packet_write_1_gI: SplitGuardInterface generic map(name => "nic_rx_to_packet_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      nic_rx_to_packet_write_1: OutputPortRevised -- 
        generic map ( name => "nic_rx_to_packet", data_width => 73, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => nic_rx_to_packet_pipe_write_req(0),
          oack => nic_rx_to_packet_pipe_write_ack(0),
          odata => nic_rx_to_packet_pipe_write_data(72 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_15958_call call_stmt_15940_call 
    AccessRegister_call_group_0: Block -- 
      signal data_in: std_logic_vector(85 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_15958_call_req_0;
      reqL_unguarded(0) <= call_stmt_15940_call_req_0;
      call_stmt_15958_call_ack_0 <= ackL_unguarded(1);
      call_stmt_15940_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_15958_call_req_1;
      reqR_unguarded(0) <= call_stmt_15940_call_req_1;
      call_stmt_15958_call_ack_1 <= ackR_unguarded(1);
      call_stmt_15940_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      AccessRegister_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "AccessRegister_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      AccessRegister_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "AccessRegister_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      AccessRegister_call_group_0_gI: SplitGuardInterface generic map(name => "AccessRegister_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_15950_wire_constant & NOT_u4_u4_15953_wire_constant & konst_15954_wire_constant & type_cast_15956_wire_constant & type_cast_15932_wire_constant & NOT_u4_u4_15935_wire_constant & konst_15936_wire_constant & type_cast_15938_wire_constant;
      ignore_resp1_15958 <= data_out(63 downto 32);
      ignore_resp0_15940 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 86,
        owidth => 43,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => AccessRegister_call_reqs(1),
          ackR => AccessRegister_call_acks(1),
          dataR => AccessRegister_call_data(85 downto 43),
          tagR => AccessRegister_call_tag(3 downto 2),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => AccessRegister_return_acks(1), -- cross-over
          ackL => AccessRegister_return_reqs(1), -- cross-over
          dataL => AccessRegister_return_data(63 downto 32),
          tagL => AccessRegister_return_tag(3 downto 2),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    volatile_operator_nextLSTATE_43052: nextLSTATE_Volatile port map(RX => RX_15965, LSTATE => LSTATE_15961, nLSTATE => nLSTATE_15980); 
    -- shared call operator group (2) : call_stmt_16028_call 
    AccessRegister_call_group_2: Block -- 
      signal data_in: std_logic_vector(42 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_16028_call_req_0;
      call_stmt_16028_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_16028_call_req_1;
      call_stmt_16028_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= pkt_complete_16009(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      AccessRegister_call_group_2_gI: SplitGuardInterface generic map(name => "AccessRegister_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_16021_wire_constant & NOT_u4_u4_16024_wire_constant & konst_16025_wire_constant & pkt_cnt_15968;
      ignore_resp2_16028 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 43,
        owidth => 43,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => AccessRegister_call_reqs(0),
          ackR => AccessRegister_call_acks(0),
          dataR => AccessRegister_call_data(42 downto 0),
          tagR => AccessRegister_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => AccessRegister_return_acks(0), -- cross-over
          ackL => AccessRegister_return_reqs(0), -- cross-over
          dataL => AccessRegister_return_data(31 downto 0),
          tagL => AccessRegister_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end nicRxFromMacDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.nic_system_global_package.all;
entity popFromQueue is -- 
  generic (tag_length : integer); 
  port ( -- 
    lock : in  std_logic_vector(0 downto 0);
    q_base_address : in  std_logic_vector(35 downto 0);
    q_r_data : out  std_logic_vector(31 downto 0);
    status : out  std_logic_vector(0 downto 0);
    releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
    releaseLock_call_acks : in   std_logic_vector(0 downto 0);
    releaseLock_call_data : out  std_logic_vector(35 downto 0);
    releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
    releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
    releaseLock_return_acks : in   std_logic_vector(0 downto 0);
    releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
    setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
    setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
    setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
    setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
    setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
    setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
    setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
    acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
    acquireLock_call_acks : in   std_logic_vector(0 downto 0);
    acquireLock_call_data : out  std_logic_vector(35 downto 0);
    acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
    acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
    acquireLock_return_acks : in   std_logic_vector(0 downto 0);
    acquireLock_return_data : in   std_logic_vector(0 downto 0);
    acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    updateTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
    updateTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
    updateTotalMessages_call_data : out  std_logic_vector(67 downto 0);
    updateTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
    updateTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
    updateTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
    updateTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
    getQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
    getQueueElement_call_acks : in   std_logic_vector(0 downto 0);
    getQueueElement_call_data : out  std_logic_vector(67 downto 0);
    getQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
    getQueueElement_return_acks : in   std_logic_vector(0 downto 0);
    getQueueElement_return_data : in   std_logic_vector(31 downto 0);
    getQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
    getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
    getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
    getTotalMessages_call_data : out  std_logic_vector(35 downto 0);
    getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
    getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
    getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
    getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
    getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
    getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
    getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
    getQueueLength_call_data : out  std_logic_vector(35 downto 0);
    getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
    getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
    getQueueLength_return_data : in   std_logic_vector(31 downto 0);
    getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
    getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
    getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
    getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
    getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
    getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
    getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
    getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity popFromQueue;
architecture popFromQueue_arch of popFromQueue is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 37)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 33)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal lock_buffer :  std_logic_vector(0 downto 0);
  signal lock_update_enable: Boolean;
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  -- output port buffer signals
  signal q_r_data_buffer :  std_logic_vector(31 downto 0);
  signal q_r_data_update_enable: Boolean;
  signal status_buffer :  std_logic_vector(0 downto 0);
  signal status_update_enable: Boolean;
  signal popFromQueue_CP_1344_start: Boolean;
  signal popFromQueue_CP_1344_symbol: Boolean;
  -- volatile/operator module components. 
  component releaseLock is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component setQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : in  std_logic_vector(31 downto 0);
      rp : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component acquireLock is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      m_ok : out  std_logic_vector(0 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component updateTotalMessages is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      updated_total_msgs : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getQueueElement is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      read_index : in  std_logic_vector(31 downto 0);
      q_r_data : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getTotalMessages is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      total_msgs : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getQueueLength is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      Queue_Length : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : out  std_logic_vector(31 downto 0);
      rp : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1175_call_req_0 : boolean;
  signal call_stmt_1175_call_ack_0 : boolean;
  signal call_stmt_1175_call_req_1 : boolean;
  signal call_stmt_1175_call_ack_1 : boolean;
  signal call_stmt_1189_call_req_0 : boolean;
  signal call_stmt_1189_call_ack_0 : boolean;
  signal call_stmt_1189_call_req_1 : boolean;
  signal call_stmt_1189_call_ack_1 : boolean;
  signal call_stmt_1194_call_req_0 : boolean;
  signal call_stmt_1194_call_ack_0 : boolean;
  signal call_stmt_1194_call_req_1 : boolean;
  signal call_stmt_1194_call_ack_1 : boolean;
  signal call_stmt_1202_call_req_0 : boolean;
  signal call_stmt_1202_call_ack_0 : boolean;
  signal call_stmt_1202_call_req_1 : boolean;
  signal call_stmt_1202_call_ack_1 : boolean;
  signal call_stmt_1205_call_req_0 : boolean;
  signal call_stmt_1205_call_ack_0 : boolean;
  signal call_stmt_1205_call_req_1 : boolean;
  signal call_stmt_1205_call_ack_1 : boolean;
  signal call_stmt_1225_call_req_0 : boolean;
  signal call_stmt_1225_call_ack_0 : boolean;
  signal call_stmt_1225_call_req_1 : boolean;
  signal call_stmt_1225_call_ack_1 : boolean;
  signal call_stmt_1230_call_req_0 : boolean;
  signal call_stmt_1230_call_ack_0 : boolean;
  signal call_stmt_1230_call_req_1 : boolean;
  signal call_stmt_1230_call_ack_1 : boolean;
  signal call_stmt_1237_call_req_0 : boolean;
  signal call_stmt_1237_call_ack_0 : boolean;
  signal call_stmt_1237_call_req_1 : boolean;
  signal call_stmt_1237_call_ack_1 : boolean;
  signal call_stmt_1248_call_req_0 : boolean;
  signal call_stmt_1248_call_ack_0 : boolean;
  signal call_stmt_1248_call_req_1 : boolean;
  signal call_stmt_1248_call_ack_1 : boolean;
  signal W_status_1249_inst_req_0 : boolean;
  signal W_status_1249_inst_ack_0 : boolean;
  signal W_status_1249_inst_req_1 : boolean;
  signal W_status_1249_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "popFromQueue_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 37) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= lock;
  lock_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(36 downto 1) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(36 downto 1);
  in_buffer_data_in(tag_length + 36 downto 37) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 36 downto 37);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  popFromQueue_CP_1344_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "popFromQueue_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 33) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(31 downto 0) <= q_r_data_buffer;
  q_r_data <= out_buffer_data_out(31 downto 0);
  out_buffer_data_in(32 downto 32) <= status_buffer;
  status <= out_buffer_data_out(32 downto 32);
  out_buffer_data_in(tag_length + 32 downto 33) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 32 downto 33);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= popFromQueue_CP_1344_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= popFromQueue_CP_1344_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= popFromQueue_CP_1344_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  popFromQueue_CP_1344: Block -- control-path 
    signal popFromQueue_CP_1344_elements: BooleanArray(24 downto 0);
    -- 
  begin -- 
    popFromQueue_CP_1344_elements(0) <= popFromQueue_CP_1344_start;
    popFromQueue_CP_1344_symbol <= popFromQueue_CP_1344_elements(24);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_1175_to_call_stmt_1189/$entry
      -- CP-element group 0: 	 call_stmt_1175_to_call_stmt_1189/call_stmt_1175_sample_start_
      -- CP-element group 0: 	 call_stmt_1175_to_call_stmt_1189/call_stmt_1175_update_start_
      -- CP-element group 0: 	 call_stmt_1175_to_call_stmt_1189/call_stmt_1175_Sample/$entry
      -- CP-element group 0: 	 call_stmt_1175_to_call_stmt_1189/call_stmt_1175_Sample/crr
      -- CP-element group 0: 	 call_stmt_1175_to_call_stmt_1189/call_stmt_1175_Update/$entry
      -- CP-element group 0: 	 call_stmt_1175_to_call_stmt_1189/call_stmt_1175_Update/ccr
      -- CP-element group 0: 	 call_stmt_1175_to_call_stmt_1189/call_stmt_1189_update_start_
      -- CP-element group 0: 	 call_stmt_1175_to_call_stmt_1189/call_stmt_1189_Update/$entry
      -- CP-element group 0: 	 call_stmt_1175_to_call_stmt_1189/call_stmt_1189_Update/ccr
      -- 
    crr_1357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1344_elements(0), ack => call_stmt_1175_call_req_0); -- 
    ccr_1362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1344_elements(0), ack => call_stmt_1175_call_req_1); -- 
    ccr_1376_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1376_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1344_elements(0), ack => call_stmt_1189_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_1175_to_call_stmt_1189/call_stmt_1175_sample_completed_
      -- CP-element group 1: 	 call_stmt_1175_to_call_stmt_1189/call_stmt_1175_Sample/$exit
      -- CP-element group 1: 	 call_stmt_1175_to_call_stmt_1189/call_stmt_1175_Sample/cra
      -- 
    cra_1358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1175_call_ack_0, ack => popFromQueue_CP_1344_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 call_stmt_1175_to_call_stmt_1189/call_stmt_1175_update_completed_
      -- CP-element group 2: 	 call_stmt_1175_to_call_stmt_1189/call_stmt_1175_Update/$exit
      -- CP-element group 2: 	 call_stmt_1175_to_call_stmt_1189/call_stmt_1175_Update/cca
      -- CP-element group 2: 	 call_stmt_1175_to_call_stmt_1189/call_stmt_1189_sample_start_
      -- CP-element group 2: 	 call_stmt_1175_to_call_stmt_1189/call_stmt_1189_Sample/$entry
      -- CP-element group 2: 	 call_stmt_1175_to_call_stmt_1189/call_stmt_1189_Sample/crr
      -- 
    cca_1363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1175_call_ack_1, ack => popFromQueue_CP_1344_elements(2)); -- 
    crr_1371_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1371_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1344_elements(2), ack => call_stmt_1189_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 call_stmt_1175_to_call_stmt_1189/call_stmt_1189_sample_completed_
      -- CP-element group 3: 	 call_stmt_1175_to_call_stmt_1189/call_stmt_1189_Sample/$exit
      -- CP-element group 3: 	 call_stmt_1175_to_call_stmt_1189/call_stmt_1189_Sample/cra
      -- 
    cra_1372_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1189_call_ack_0, ack => popFromQueue_CP_1344_elements(3)); -- 
    -- CP-element group 4:  fork  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4: 	6 
    -- CP-element group 4: 	8 
    -- CP-element group 4: 	10 
    -- CP-element group 4: 	13 
    -- CP-element group 4: 	16 
    -- CP-element group 4: 	19 
    -- CP-element group 4:  members (26) 
      -- CP-element group 4: 	 call_stmt_1175_to_call_stmt_1189/$exit
      -- CP-element group 4: 	 call_stmt_1175_to_call_stmt_1189/call_stmt_1189_update_completed_
      -- CP-element group 4: 	 call_stmt_1175_to_call_stmt_1189/call_stmt_1189_Update/$exit
      -- CP-element group 4: 	 call_stmt_1175_to_call_stmt_1189/call_stmt_1189_Update/cca
      -- CP-element group 4: 	 call_stmt_1194_to_call_stmt_1237/$entry
      -- CP-element group 4: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1194_sample_start_
      -- CP-element group 4: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1194_update_start_
      -- CP-element group 4: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1194_Sample/$entry
      -- CP-element group 4: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1194_Sample/crr
      -- CP-element group 4: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1194_Update/$entry
      -- CP-element group 4: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1194_Update/ccr
      -- CP-element group 4: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1202_update_start_
      -- CP-element group 4: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1202_Update/$entry
      -- CP-element group 4: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1202_Update/ccr
      -- CP-element group 4: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1205_update_start_
      -- CP-element group 4: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1205_Update/$entry
      -- CP-element group 4: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1205_Update/ccr
      -- CP-element group 4: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1225_update_start_
      -- CP-element group 4: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1225_Update/$entry
      -- CP-element group 4: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1225_Update/ccr
      -- CP-element group 4: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1230_update_start_
      -- CP-element group 4: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1230_Update/$entry
      -- CP-element group 4: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1230_Update/ccr
      -- CP-element group 4: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1237_update_start_
      -- CP-element group 4: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1237_Update/$entry
      -- CP-element group 4: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1237_Update/ccr
      -- 
    cca_1377_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1189_call_ack_1, ack => popFromQueue_CP_1344_elements(4)); -- 
    crr_1388_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1388_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1344_elements(4), ack => call_stmt_1194_call_req_0); -- 
    ccr_1393_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1393_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1344_elements(4), ack => call_stmt_1194_call_req_1); -- 
    ccr_1407_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1407_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1344_elements(4), ack => call_stmt_1202_call_req_1); -- 
    ccr_1421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1344_elements(4), ack => call_stmt_1205_call_req_1); -- 
    ccr_1435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1344_elements(4), ack => call_stmt_1225_call_req_1); -- 
    ccr_1449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1344_elements(4), ack => call_stmt_1230_call_req_1); -- 
    ccr_1463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1344_elements(4), ack => call_stmt_1237_call_req_1); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1194_sample_completed_
      -- CP-element group 5: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1194_Sample/$exit
      -- CP-element group 5: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1194_Sample/cra
      -- 
    cra_1389_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1194_call_ack_0, ack => popFromQueue_CP_1344_elements(5)); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	4 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	11 
    -- CP-element group 6: 	14 
    -- CP-element group 6: 	17 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1194_update_completed_
      -- CP-element group 6: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1194_Update/$exit
      -- CP-element group 6: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1194_Update/cca
      -- CP-element group 6: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1202_sample_start_
      -- CP-element group 6: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1202_Sample/$entry
      -- CP-element group 6: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1202_Sample/crr
      -- 
    cca_1394_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1194_call_ack_1, ack => popFromQueue_CP_1344_elements(6)); -- 
    crr_1402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1344_elements(6), ack => call_stmt_1202_call_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1202_sample_completed_
      -- CP-element group 7: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1202_Sample/$exit
      -- CP-element group 7: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1202_Sample/cra
      -- 
    cra_1403_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1202_call_ack_0, ack => popFromQueue_CP_1344_elements(7)); -- 
    -- CP-element group 8:  fork  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	4 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8: 	14 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1202_update_completed_
      -- CP-element group 8: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1202_Update/$exit
      -- CP-element group 8: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1202_Update/cca
      -- CP-element group 8: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1205_sample_start_
      -- CP-element group 8: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1205_Sample/$entry
      -- CP-element group 8: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1205_Sample/crr
      -- 
    cca_1408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1202_call_ack_1, ack => popFromQueue_CP_1344_elements(8)); -- 
    crr_1416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1344_elements(8), ack => call_stmt_1205_call_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1205_sample_completed_
      -- CP-element group 9: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1205_Sample/$exit
      -- CP-element group 9: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1205_Sample/cra
      -- 
    cra_1417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1205_call_ack_0, ack => popFromQueue_CP_1344_elements(9)); -- 
    -- CP-element group 10:  fork  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	4 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	17 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1205_update_completed_
      -- CP-element group 10: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1205_Update/$exit
      -- CP-element group 10: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1205_Update/cca
      -- 
    cca_1422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1205_call_ack_1, ack => popFromQueue_CP_1344_elements(10)); -- 
    -- CP-element group 11:  join  transition  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	6 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1225_sample_start_
      -- CP-element group 11: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1225_Sample/$entry
      -- CP-element group 11: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1225_Sample/crr
      -- 
    crr_1430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1344_elements(11), ack => call_stmt_1225_call_req_0); -- 
    popFromQueue_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "popFromQueue_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= popFromQueue_CP_1344_elements(6) & popFromQueue_CP_1344_elements(10);
      gj_popFromQueue_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => popFromQueue_CP_1344_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1225_sample_completed_
      -- CP-element group 12: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1225_Sample/$exit
      -- CP-element group 12: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1225_Sample/cra
      -- 
    cra_1431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1225_call_ack_0, ack => popFromQueue_CP_1344_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	4 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1225_update_completed_
      -- CP-element group 13: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1225_Update/$exit
      -- CP-element group 13: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1225_Update/cca
      -- 
    cca_1436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1225_call_ack_1, ack => popFromQueue_CP_1344_elements(13)); -- 
    -- CP-element group 14:  join  transition  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	6 
    -- CP-element group 14: 	8 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1230_sample_start_
      -- CP-element group 14: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1230_Sample/$entry
      -- CP-element group 14: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1230_Sample/crr
      -- 
    crr_1444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1344_elements(14), ack => call_stmt_1230_call_req_0); -- 
    popFromQueue_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "popFromQueue_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= popFromQueue_CP_1344_elements(6) & popFromQueue_CP_1344_elements(8) & popFromQueue_CP_1344_elements(13);
      gj_popFromQueue_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => popFromQueue_CP_1344_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1230_sample_completed_
      -- CP-element group 15: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1230_Sample/$exit
      -- CP-element group 15: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1230_Sample/cra
      -- 
    cra_1445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1230_call_ack_0, ack => popFromQueue_CP_1344_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	4 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1230_update_completed_
      -- CP-element group 16: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1230_Update/$exit
      -- CP-element group 16: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1230_Update/cca
      -- 
    cca_1450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1230_call_ack_1, ack => popFromQueue_CP_1344_elements(16)); -- 
    -- CP-element group 17:  join  transition  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	6 
    -- CP-element group 17: 	10 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1237_sample_start_
      -- CP-element group 17: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1237_Sample/$entry
      -- CP-element group 17: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1237_Sample/crr
      -- 
    crr_1458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1344_elements(17), ack => call_stmt_1237_call_req_0); -- 
    popFromQueue_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 32) := "popFromQueue_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= popFromQueue_CP_1344_elements(6) & popFromQueue_CP_1344_elements(10) & popFromQueue_CP_1344_elements(16);
      gj_popFromQueue_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => popFromQueue_CP_1344_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1237_sample_completed_
      -- CP-element group 18: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1237_Sample/$exit
      -- CP-element group 18: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1237_Sample/cra
      -- 
    cra_1459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1237_call_ack_0, ack => popFromQueue_CP_1344_elements(18)); -- 
    -- CP-element group 19:  fork  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	4 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19: 	21 
    -- CP-element group 19: 	22 
    -- CP-element group 19: 	23 
    -- CP-element group 19:  members (17) 
      -- CP-element group 19: 	 call_stmt_1194_to_call_stmt_1237/$exit
      -- CP-element group 19: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1237_update_completed_
      -- CP-element group 19: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1237_Update/$exit
      -- CP-element group 19: 	 call_stmt_1194_to_call_stmt_1237/call_stmt_1237_Update/cca
      -- CP-element group 19: 	 call_stmt_1248_to_assign_stmt_1251/$entry
      -- CP-element group 19: 	 call_stmt_1248_to_assign_stmt_1251/call_stmt_1248_sample_start_
      -- CP-element group 19: 	 call_stmt_1248_to_assign_stmt_1251/call_stmt_1248_update_start_
      -- CP-element group 19: 	 call_stmt_1248_to_assign_stmt_1251/call_stmt_1248_Sample/$entry
      -- CP-element group 19: 	 call_stmt_1248_to_assign_stmt_1251/call_stmt_1248_Sample/crr
      -- CP-element group 19: 	 call_stmt_1248_to_assign_stmt_1251/call_stmt_1248_Update/$entry
      -- CP-element group 19: 	 call_stmt_1248_to_assign_stmt_1251/call_stmt_1248_Update/ccr
      -- CP-element group 19: 	 call_stmt_1248_to_assign_stmt_1251/assign_stmt_1251_sample_start_
      -- CP-element group 19: 	 call_stmt_1248_to_assign_stmt_1251/assign_stmt_1251_update_start_
      -- CP-element group 19: 	 call_stmt_1248_to_assign_stmt_1251/assign_stmt_1251_Sample/$entry
      -- CP-element group 19: 	 call_stmt_1248_to_assign_stmt_1251/assign_stmt_1251_Sample/req
      -- CP-element group 19: 	 call_stmt_1248_to_assign_stmt_1251/assign_stmt_1251_Update/$entry
      -- CP-element group 19: 	 call_stmt_1248_to_assign_stmt_1251/assign_stmt_1251_Update/req
      -- 
    cca_1464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1237_call_ack_1, ack => popFromQueue_CP_1344_elements(19)); -- 
    crr_1475_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1475_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1344_elements(19), ack => call_stmt_1248_call_req_0); -- 
    ccr_1480_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1480_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1344_elements(19), ack => call_stmt_1248_call_req_1); -- 
    req_1489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1344_elements(19), ack => W_status_1249_inst_req_0); -- 
    req_1494_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1494_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => popFromQueue_CP_1344_elements(19), ack => W_status_1249_inst_req_1); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 call_stmt_1248_to_assign_stmt_1251/call_stmt_1248_sample_completed_
      -- CP-element group 20: 	 call_stmt_1248_to_assign_stmt_1251/call_stmt_1248_Sample/$exit
      -- CP-element group 20: 	 call_stmt_1248_to_assign_stmt_1251/call_stmt_1248_Sample/cra
      -- 
    cra_1476_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1248_call_ack_0, ack => popFromQueue_CP_1344_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	19 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 call_stmt_1248_to_assign_stmt_1251/call_stmt_1248_update_completed_
      -- CP-element group 21: 	 call_stmt_1248_to_assign_stmt_1251/call_stmt_1248_Update/$exit
      -- CP-element group 21: 	 call_stmt_1248_to_assign_stmt_1251/call_stmt_1248_Update/cca
      -- 
    cca_1481_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1248_call_ack_1, ack => popFromQueue_CP_1344_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 call_stmt_1248_to_assign_stmt_1251/assign_stmt_1251_sample_completed_
      -- CP-element group 22: 	 call_stmt_1248_to_assign_stmt_1251/assign_stmt_1251_Sample/$exit
      -- CP-element group 22: 	 call_stmt_1248_to_assign_stmt_1251/assign_stmt_1251_Sample/ack
      -- 
    ack_1490_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_status_1249_inst_ack_0, ack => popFromQueue_CP_1344_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	19 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 call_stmt_1248_to_assign_stmt_1251/assign_stmt_1251_update_completed_
      -- CP-element group 23: 	 call_stmt_1248_to_assign_stmt_1251/assign_stmt_1251_Update/$exit
      -- CP-element group 23: 	 call_stmt_1248_to_assign_stmt_1251/assign_stmt_1251_Update/ack
      -- 
    ack_1495_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_status_1249_inst_ack_1, ack => popFromQueue_CP_1344_elements(23)); -- 
    -- CP-element group 24:  join  transition  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 $exit
      -- CP-element group 24: 	 call_stmt_1248_to_assign_stmt_1251/$exit
      -- 
    popFromQueue_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "popFromQueue_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= popFromQueue_CP_1344_elements(21) & popFromQueue_CP_1344_elements(23);
      gj_popFromQueue_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => popFromQueue_CP_1344_elements(24), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_1218_wire : std_logic_vector(31 downto 0);
    signal ADD_u36_u36_1171_wire : std_logic_vector(35 downto 0);
    signal NOT_u8_u8_1168_wire_constant : std_logic_vector(7 downto 0);
    signal Queue_Length_1202 : std_logic_vector(31 downto 0);
    signal SUB_u32_u32_1210_wire : std_logic_vector(31 downto 0);
    signal SUB_u32_u32_1236_wire : std_logic_vector(31 downto 0);
    signal ba_and_misc_1175 : std_logic_vector(63 downto 0);
    signal konst_1170_wire_constant : std_logic_vector(35 downto 0);
    signal konst_1209_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1215_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1217_wire_constant : std_logic_vector(31 downto 0);
    signal lock_n_1185 : std_logic_vector(0 downto 0);
    signal m_ok_1189 : std_logic_vector(0 downto 0);
    signal misc_1179 : std_logic_vector(31 downto 0);
    signal next_ri_1220 : std_logic_vector(31 downto 0);
    signal q_empty_1199 : std_logic_vector(0 downto 0);
    signal read_index_1194 : std_logic_vector(31 downto 0);
    signal round_off_1212 : std_logic_vector(0 downto 0);
    signal total_msgs_1205 : std_logic_vector(31 downto 0);
    signal type_cast_1163_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1165_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1173_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1183_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1235_wire_constant : std_logic_vector(31 downto 0);
    signal write_index_1194 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    NOT_u8_u8_1168_wire_constant <= "11111111";
    konst_1170_wire_constant <= "000000000000000000000000000000011000";
    konst_1209_wire_constant <= "00000000000000000000000000000001";
    konst_1215_wire_constant <= "00000000000000000000000000000000";
    konst_1217_wire_constant <= "00000000000000000000000000000001";
    type_cast_1163_wire_constant <= "0";
    type_cast_1165_wire_constant <= "1";
    type_cast_1173_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1183_wire_constant <= "00000000000000000000000000000000";
    type_cast_1235_wire_constant <= "00000000000000000000000000000001";
    -- flow-through select operator MUX_1219_inst
    next_ri_1220 <= konst_1215_wire_constant when (round_off_1212(0) /=  '0') else ADD_u32_u32_1218_wire;
    -- flow-through slice operator slice_1178_inst
    misc_1179 <= ba_and_misc_1175(31 downto 0);
    W_status_1249_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_status_1249_inst_req_0;
      W_status_1249_inst_ack_0<= wack(0);
      rreq(0) <= W_status_1249_inst_req_1;
      W_status_1249_inst_ack_1<= rack(0);
      W_status_1249_inst : InterlockBuffer generic map ( -- 
        name => "W_status_1249_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => q_empty_1199,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => status_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- binary operator ADD_u32_u32_1218_inst
    process(read_index_1194) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(read_index_1194, konst_1217_wire_constant, tmp_var);
      ADD_u32_u32_1218_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u36_u36_1171_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, konst_1170_wire_constant, tmp_var);
      ADD_u36_u36_1171_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1184_inst
    process(misc_1179) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(misc_1179, type_cast_1183_wire_constant, tmp_var);
      lock_n_1185 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1198_inst
    process(write_index_1194, read_index_1194) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(write_index_1194, read_index_1194, tmp_var);
      q_empty_1199 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1211_inst
    process(read_index_1194, SUB_u32_u32_1210_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(read_index_1194, SUB_u32_u32_1210_wire, tmp_var);
      round_off_1212 <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1210_inst
    process(Queue_Length_1202) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(Queue_Length_1202, konst_1209_wire_constant, tmp_var);
      SUB_u32_u32_1210_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1236_inst
    process(total_msgs_1205) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(total_msgs_1205, type_cast_1235_wire_constant, tmp_var);
      SUB_u32_u32_1236_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_1175_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1175_call_req_0;
      call_stmt_1175_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1175_call_req_1;
      call_stmt_1175_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1163_wire_constant & type_cast_1165_wire_constant & NOT_u8_u8_1168_wire_constant & ADD_u36_u36_1171_wire & type_cast_1173_wire_constant;
      ba_and_misc_1175 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1189_call 
    acquireLock_call_group_1: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1189_call_req_0;
      call_stmt_1189_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1189_call_req_1;
      call_stmt_1189_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= lock_n_1185(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      acquireLock_call_group_1_gI: SplitGuardInterface generic map(name => "acquireLock_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      m_ok_1189 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => acquireLock_call_reqs(0),
          ackR => acquireLock_call_acks(0),
          dataR => acquireLock_call_data(35 downto 0),
          tagR => acquireLock_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => acquireLock_return_acks(0), -- cross-over
          ackL => acquireLock_return_reqs(0), -- cross-over
          dataL => acquireLock_return_data(0 downto 0),
          tagL => acquireLock_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1194_call 
    getQueuePointers_call_group_2: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1194_call_req_0;
      call_stmt_1194_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1194_call_req_1;
      call_stmt_1194_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueuePointers_call_group_2_gI: SplitGuardInterface generic map(name => "getQueuePointers_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      write_index_1194 <= data_out(63 downto 32);
      read_index_1194 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueuePointers_call_reqs(0),
          ackR => getQueuePointers_call_acks(0),
          dataR => getQueuePointers_call_data(35 downto 0),
          tagR => getQueuePointers_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueuePointers_return_acks(0), -- cross-over
          ackL => getQueuePointers_return_reqs(0), -- cross-over
          dataL => getQueuePointers_return_data(63 downto 0),
          tagL => getQueuePointers_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_1202_call 
    getQueueLength_call_group_3: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1202_call_req_0;
      call_stmt_1202_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1202_call_req_1;
      call_stmt_1202_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueueLength_call_group_3_gI: SplitGuardInterface generic map(name => "getQueueLength_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      Queue_Length_1202 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueueLength_call_reqs(0),
          ackR => getQueueLength_call_acks(0),
          dataR => getQueueLength_call_data(35 downto 0),
          tagR => getQueueLength_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueueLength_return_acks(0), -- cross-over
          ackL => getQueueLength_return_reqs(0), -- cross-over
          dataL => getQueueLength_return_data(31 downto 0),
          tagL => getQueueLength_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- shared call operator group (4) : call_stmt_1205_call 
    getTotalMessages_call_group_4: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1205_call_req_0;
      call_stmt_1205_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1205_call_req_1;
      call_stmt_1205_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getTotalMessages_call_group_4_gI: SplitGuardInterface generic map(name => "getTotalMessages_call_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      total_msgs_1205 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getTotalMessages_call_reqs(0),
          ackR => getTotalMessages_call_acks(0),
          dataR => getTotalMessages_call_data(35 downto 0),
          tagR => getTotalMessages_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getTotalMessages_return_acks(0), -- cross-over
          ackL => getTotalMessages_return_reqs(0), -- cross-over
          dataL => getTotalMessages_return_data(31 downto 0),
          tagL => getTotalMessages_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 4
    -- shared call operator group (5) : call_stmt_1225_call 
    getQueueElement_call_group_5: Block -- 
      signal data_in: std_logic_vector(67 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1225_call_req_0;
      call_stmt_1225_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1225_call_req_1;
      call_stmt_1225_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_empty_1199(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueueElement_call_group_5_gI: SplitGuardInterface generic map(name => "getQueueElement_call_group_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer & read_index_1194;
      q_r_data_buffer <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 68,
        owidth => 68,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueueElement_call_reqs(0),
          ackR => getQueueElement_call_acks(0),
          dataR => getQueueElement_call_data(67 downto 0),
          tagR => getQueueElement_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueueElement_return_acks(0), -- cross-over
          ackL => getQueueElement_return_reqs(0), -- cross-over
          dataL => getQueueElement_return_data(31 downto 0),
          tagL => getQueueElement_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 5
    -- shared call operator group (6) : call_stmt_1230_call 
    setQueuePointers_call_group_6: Block -- 
      signal data_in: std_logic_vector(99 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1230_call_req_0;
      call_stmt_1230_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1230_call_req_1;
      call_stmt_1230_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_empty_1199(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      setQueuePointers_call_group_6_gI: SplitGuardInterface generic map(name => "setQueuePointers_call_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer & write_index_1194 & next_ri_1220;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 100,
        owidth => 100,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => setQueuePointers_call_reqs(0),
          ackR => setQueuePointers_call_acks(0),
          dataR => setQueuePointers_call_data(99 downto 0),
          tagR => setQueuePointers_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => setQueuePointers_return_acks(0), -- cross-over
          ackL => setQueuePointers_return_reqs(0), -- cross-over
          tagL => setQueuePointers_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 6
    -- shared call operator group (7) : call_stmt_1237_call 
    updateTotalMessages_call_group_7: Block -- 
      signal data_in: std_logic_vector(67 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1237_call_req_0;
      call_stmt_1237_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1237_call_req_1;
      call_stmt_1237_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_empty_1199(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      updateTotalMessages_call_group_7_gI: SplitGuardInterface generic map(name => "updateTotalMessages_call_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer & SUB_u32_u32_1236_wire;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 68,
        owidth => 68,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => updateTotalMessages_call_reqs(0),
          ackR => updateTotalMessages_call_acks(0),
          dataR => updateTotalMessages_call_data(67 downto 0),
          tagR => updateTotalMessages_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => updateTotalMessages_return_acks(0), -- cross-over
          ackL => updateTotalMessages_return_reqs(0), -- cross-over
          tagL => updateTotalMessages_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 7
    -- shared call operator group (8) : call_stmt_1248_call 
    releaseLock_call_group_8: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1248_call_req_0;
      call_stmt_1248_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1248_call_req_1;
      call_stmt_1248_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= lock_n_1185(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      releaseLock_call_group_8_gI: SplitGuardInterface generic map(name => "releaseLock_call_group_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => releaseLock_call_reqs(0),
          ackR => releaseLock_call_acks(0),
          dataR => releaseLock_call_data(35 downto 0),
          tagR => releaseLock_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => releaseLock_return_acks(0), -- cross-over
          ackL => releaseLock_return_reqs(0), -- cross-over
          tagL => releaseLock_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 8
    -- 
  end Block; -- data_path
  -- 
end popFromQueue_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.nic_system_global_package.all;
entity populateRxQueue is -- 
  generic (tag_length : integer); 
  port ( -- 
    rx_buffer_pointer : in  std_logic_vector(35 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX : in std_logic_vector(5 downto 0);
    NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
    LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(5 downto 0);
    AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_call_data : out  std_logic_vector(42 downto 0);
    AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
    AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_return_data : in   std_logic_vector(31 downto 0);
    AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
    pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
    pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity populateRxQueue;
architecture populateRxQueue_arch of populateRxQueue is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rx_buffer_pointer_buffer :  std_logic_vector(35 downto 0);
  signal rx_buffer_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal populateRxQueue_CP_2199_start: Boolean;
  signal populateRxQueue_CP_2199_symbol: Boolean;
  -- volatile/operator module components. 
  component AccessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      register_index : in  std_logic_vector(5 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component pushIntoQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_call_acks : in   std_logic_vector(0 downto 0);
      releaseLock_call_data : out  std_logic_vector(35 downto 0);
      releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_return_acks : in   std_logic_vector(0 downto 0);
      releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_call_acks : in   std_logic_vector(0 downto 0);
      acquireLock_call_data : out  std_logic_vector(35 downto 0);
      acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_return_acks : in   std_logic_vector(0 downto 0);
      acquireLock_return_data : in   std_logic_vector(0 downto 0);
      acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      updateTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_data : out  std_logic_vector(67 downto 0);
      updateTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_call_data : out  std_logic_vector(35 downto 0);
      getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
      getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_call_data : out  std_logic_vector(35 downto 0);
      getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_return_data : in   std_logic_vector(31 downto 0);
      getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_call_data : out  std_logic_vector(99 downto 0);
      setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component delay_time_Operator is -- 
    port ( -- 
      sample_req: in boolean;
      sample_ack: out boolean;
      update_req: in boolean;
      update_ack: out boolean;
      T : in  std_logic_vector(31 downto 0);
      delay_done : out  std_logic_vector(0 downto 0);
      clk, reset: in std_logic
      -- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal n_q_index_1695_1647_buf_req_0 : boolean;
  signal n_q_index_1695_1647_buf_req_1 : boolean;
  signal n_q_index_1695_1647_buf_ack_0 : boolean;
  signal AND_u6_u6_1646_inst_req_1 : boolean;
  signal n_q_index_1695_1647_buf_ack_1 : boolean;
  signal phi_stmt_1637_req_1 : boolean;
  signal AND_u6_u6_1646_inst_ack_1 : boolean;
  signal phi_stmt_1637_ack_0 : boolean;
  signal AND_u6_u6_1646_inst_ack_0 : boolean;
  signal AND_u6_u6_1646_inst_req_0 : boolean;
  signal call_stmt_1668_call_req_0 : boolean;
  signal call_stmt_1668_call_ack_0 : boolean;
  signal call_stmt_1668_call_req_1 : boolean;
  signal call_stmt_1668_call_ack_1 : boolean;
  signal call_stmt_1685_call_req_0 : boolean;
  signal call_stmt_1685_call_ack_0 : boolean;
  signal call_stmt_1685_call_req_1 : boolean;
  signal call_stmt_1685_call_ack_1 : boolean;
  signal if_stmt_1699_branch_req_0 : boolean;
  signal if_stmt_1699_branch_ack_1 : boolean;
  signal if_stmt_1699_branch_ack_0 : boolean;
  signal call_stmt_1704_call_req_0 : boolean;
  signal call_stmt_1704_call_ack_0 : boolean;
  signal call_stmt_1704_call_req_1 : boolean;
  signal call_stmt_1704_call_ack_1 : boolean;
  signal phi_stmt_1637_req_0 : boolean;
  signal if_stmt_1705_branch_req_0 : boolean;
  signal if_stmt_1705_branch_ack_1 : boolean;
  signal if_stmt_1705_branch_ack_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1712_inst_req_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1712_inst_ack_0 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1712_inst_req_1 : boolean;
  signal WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1712_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "populateRxQueue_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= rx_buffer_pointer;
  rx_buffer_pointer_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  populateRxQueue_CP_2199_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "populateRxQueue_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= populateRxQueue_CP_2199_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= populateRxQueue_CP_2199_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= populateRxQueue_CP_2199_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  populateRxQueue_CP_2199: Block -- control-path 
    signal populateRxQueue_CP_2199_elements: BooleanArray(22 downto 0);
    -- 
  begin -- 
    populateRxQueue_CP_2199_elements(0) <= populateRxQueue_CP_2199_start;
    populateRxQueue_CP_2199_symbol <= populateRxQueue_CP_2199_elements(1);
    -- CP-element group 0:  branch  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	14 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1635/$entry
      -- CP-element group 0: 	 branch_block_stmt_1635/branch_block_stmt_1635__entry__
      -- CP-element group 0: 	 branch_block_stmt_1635/merge_stmt_1636__entry__
      -- CP-element group 0: 	 branch_block_stmt_1635/merge_stmt_1636_dead_link/$entry
      -- 
    -- CP-element group 1:  merge  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	11 
    -- CP-element group 1: 	13 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1635/$exit
      -- CP-element group 1: 	 branch_block_stmt_1635/branch_block_stmt_1635__exit__
      -- CP-element group 1: 	 branch_block_stmt_1635/if_stmt_1699__exit__
      -- 
    populateRxQueue_CP_2199_elements(1) <= OrReduce(populateRxQueue_CP_2199_elements(11) & populateRxQueue_CP_2199_elements(13));
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	22 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 branch_block_stmt_1635/assign_stmt_1656_to_assign_stmt_1695/call_stmt_1668_sample_completed_
      -- CP-element group 2: 	 branch_block_stmt_1635/assign_stmt_1656_to_assign_stmt_1695/call_stmt_1668_Sample/$exit
      -- CP-element group 2: 	 branch_block_stmt_1635/assign_stmt_1656_to_assign_stmt_1695/call_stmt_1668_Sample/cra
      -- 
    cra_2224_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1668_call_ack_0, ack => populateRxQueue_CP_2199_elements(2)); -- 
    -- CP-element group 3:  transition  input  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	22 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	4 
    -- CP-element group 3:  members (6) 
      -- CP-element group 3: 	 branch_block_stmt_1635/assign_stmt_1656_to_assign_stmt_1695/call_stmt_1668_update_completed_
      -- CP-element group 3: 	 branch_block_stmt_1635/assign_stmt_1656_to_assign_stmt_1695/call_stmt_1668_Update/$exit
      -- CP-element group 3: 	 branch_block_stmt_1635/assign_stmt_1656_to_assign_stmt_1695/call_stmt_1668_Update/cca
      -- CP-element group 3: 	 branch_block_stmt_1635/assign_stmt_1656_to_assign_stmt_1695/call_stmt_1685_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_1635/assign_stmt_1656_to_assign_stmt_1695/call_stmt_1685_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_1635/assign_stmt_1656_to_assign_stmt_1695/call_stmt_1685_Sample/crr
      -- 
    cca_2229_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1668_call_ack_1, ack => populateRxQueue_CP_2199_elements(3)); -- 
    crr_2237_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2237_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_2199_elements(3), ack => call_stmt_1685_call_req_0); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	3 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (3) 
      -- CP-element group 4: 	 branch_block_stmt_1635/assign_stmt_1656_to_assign_stmt_1695/call_stmt_1685_sample_completed_
      -- CP-element group 4: 	 branch_block_stmt_1635/assign_stmt_1656_to_assign_stmt_1695/call_stmt_1685_Sample/$exit
      -- CP-element group 4: 	 branch_block_stmt_1635/assign_stmt_1656_to_assign_stmt_1695/call_stmt_1685_Sample/cra
      -- 
    cra_2238_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1685_call_ack_0, ack => populateRxQueue_CP_2199_elements(4)); -- 
    -- CP-element group 5:  branch  transition  place  input  output  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	22 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	6 
    -- CP-element group 5: 	7 
    -- CP-element group 5:  members (25) 
      -- CP-element group 5: 	 branch_block_stmt_1635/assign_stmt_1656_to_assign_stmt_1695__exit__
      -- CP-element group 5: 	 branch_block_stmt_1635/if_stmt_1699__entry__
      -- CP-element group 5: 	 branch_block_stmt_1635/assign_stmt_1656_to_assign_stmt_1695/$exit
      -- CP-element group 5: 	 branch_block_stmt_1635/assign_stmt_1656_to_assign_stmt_1695/call_stmt_1685_update_completed_
      -- CP-element group 5: 	 branch_block_stmt_1635/assign_stmt_1656_to_assign_stmt_1695/call_stmt_1685_Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1635/assign_stmt_1656_to_assign_stmt_1695/call_stmt_1685_Update/cca
      -- CP-element group 5: 	 branch_block_stmt_1635/if_stmt_1699_dead_link/$entry
      -- CP-element group 5: 	 branch_block_stmt_1635/if_stmt_1699_eval_test/$entry
      -- CP-element group 5: 	 branch_block_stmt_1635/if_stmt_1699_eval_test/$exit
      -- CP-element group 5: 	 branch_block_stmt_1635/if_stmt_1699_eval_test/NOT_u1_u1_1701/$entry
      -- CP-element group 5: 	 branch_block_stmt_1635/if_stmt_1699_eval_test/NOT_u1_u1_1701/$exit
      -- CP-element group 5: 	 branch_block_stmt_1635/if_stmt_1699_eval_test/NOT_u1_u1_1701/SplitProtocol/$entry
      -- CP-element group 5: 	 branch_block_stmt_1635/if_stmt_1699_eval_test/NOT_u1_u1_1701/SplitProtocol/$exit
      -- CP-element group 5: 	 branch_block_stmt_1635/if_stmt_1699_eval_test/NOT_u1_u1_1701/SplitProtocol/Sample/$entry
      -- CP-element group 5: 	 branch_block_stmt_1635/if_stmt_1699_eval_test/NOT_u1_u1_1701/SplitProtocol/Sample/$exit
      -- CP-element group 5: 	 branch_block_stmt_1635/if_stmt_1699_eval_test/NOT_u1_u1_1701/SplitProtocol/Sample/rr
      -- CP-element group 5: 	 branch_block_stmt_1635/if_stmt_1699_eval_test/NOT_u1_u1_1701/SplitProtocol/Sample/ra
      -- CP-element group 5: 	 branch_block_stmt_1635/if_stmt_1699_eval_test/NOT_u1_u1_1701/SplitProtocol/Update/$entry
      -- CP-element group 5: 	 branch_block_stmt_1635/if_stmt_1699_eval_test/NOT_u1_u1_1701/SplitProtocol/Update/$exit
      -- CP-element group 5: 	 branch_block_stmt_1635/if_stmt_1699_eval_test/NOT_u1_u1_1701/SplitProtocol/Update/cr
      -- CP-element group 5: 	 branch_block_stmt_1635/if_stmt_1699_eval_test/NOT_u1_u1_1701/SplitProtocol/Update/ca
      -- CP-element group 5: 	 branch_block_stmt_1635/if_stmt_1699_eval_test/branch_req
      -- CP-element group 5: 	 branch_block_stmt_1635/NOT_u1_u1_1701_place
      -- CP-element group 5: 	 branch_block_stmt_1635/if_stmt_1699_if_link/$entry
      -- CP-element group 5: 	 branch_block_stmt_1635/if_stmt_1699_else_link/$entry
      -- 
    cca_2243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1685_call_ack_1, ack => populateRxQueue_CP_2199_elements(5)); -- 
    branch_req_2267_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2267_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_2199_elements(5), ack => if_stmt_1699_branch_req_0); -- 
    -- CP-element group 6:  fork  transition  place  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	5 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	8 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (10) 
      -- CP-element group 6: 	 branch_block_stmt_1635/if_stmt_1699_if_link/$exit
      -- CP-element group 6: 	 branch_block_stmt_1635/if_stmt_1699_if_link/if_choice_transition
      -- CP-element group 6: 	 branch_block_stmt_1635/call_stmt_1704__entry__
      -- CP-element group 6: 	 branch_block_stmt_1635/call_stmt_1704/$entry
      -- CP-element group 6: 	 branch_block_stmt_1635/call_stmt_1704/call_stmt_1704_sample_start_
      -- CP-element group 6: 	 branch_block_stmt_1635/call_stmt_1704/call_stmt_1704_update_start_
      -- CP-element group 6: 	 branch_block_stmt_1635/call_stmt_1704/call_stmt_1704_Sample/$entry
      -- CP-element group 6: 	 branch_block_stmt_1635/call_stmt_1704/call_stmt_1704_Sample/crr
      -- CP-element group 6: 	 branch_block_stmt_1635/call_stmt_1704/call_stmt_1704_Update/$entry
      -- CP-element group 6: 	 branch_block_stmt_1635/call_stmt_1704/call_stmt_1704_Update/ccr
      -- 
    if_choice_transition_2272_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1699_branch_ack_1, ack => populateRxQueue_CP_2199_elements(6)); -- 
    crr_2291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_2199_elements(6), ack => call_stmt_1704_call_req_0); -- 
    ccr_2296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_2199_elements(6), ack => call_stmt_1704_call_req_1); -- 
    -- CP-element group 7:  transition  place  input  output  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	5 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	12 
    -- CP-element group 7:  members (7) 
      -- CP-element group 7: 	 branch_block_stmt_1635/if_stmt_1699_else_link/$exit
      -- CP-element group 7: 	 branch_block_stmt_1635/if_stmt_1699_else_link/else_choice_transition
      -- CP-element group 7: 	 branch_block_stmt_1635/assign_stmt_1714__entry__
      -- CP-element group 7: 	 branch_block_stmt_1635/assign_stmt_1714/$entry
      -- CP-element group 7: 	 branch_block_stmt_1635/assign_stmt_1714/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1712_sample_start_
      -- CP-element group 7: 	 branch_block_stmt_1635/assign_stmt_1714/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1712_Sample/$entry
      -- CP-element group 7: 	 branch_block_stmt_1635/assign_stmt_1714/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1712_Sample/req
      -- 
    else_choice_transition_2276_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1699_branch_ack_0, ack => populateRxQueue_CP_2199_elements(7)); -- 
    req_2347_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2347_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_2199_elements(7), ack => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1712_inst_req_0); -- 
    -- CP-element group 8:  transition  input  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	6 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_1635/call_stmt_1704/call_stmt_1704_sample_completed_
      -- CP-element group 8: 	 branch_block_stmt_1635/call_stmt_1704/call_stmt_1704_Sample/$exit
      -- CP-element group 8: 	 branch_block_stmt_1635/call_stmt_1704/call_stmt_1704_Sample/cra
      -- 
    cra_2292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1704_call_ack_0, ack => populateRxQueue_CP_2199_elements(8)); -- 
    -- CP-element group 9:  branch  transition  place  input  output  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	10 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (27) 
      -- CP-element group 9: 	 branch_block_stmt_1635/call_stmt_1704__exit__
      -- CP-element group 9: 	 branch_block_stmt_1635/if_stmt_1705__entry__
      -- CP-element group 9: 	 branch_block_stmt_1635/call_stmt_1704/$exit
      -- CP-element group 9: 	 branch_block_stmt_1635/call_stmt_1704/call_stmt_1704_update_completed_
      -- CP-element group 9: 	 branch_block_stmt_1635/call_stmt_1704/call_stmt_1704_Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_1635/call_stmt_1704/call_stmt_1704_Update/cca
      -- CP-element group 9: 	 branch_block_stmt_1635/if_stmt_1705_dead_link/$entry
      -- CP-element group 9: 	 branch_block_stmt_1635/if_stmt_1705_eval_test/$entry
      -- CP-element group 9: 	 branch_block_stmt_1635/if_stmt_1705_eval_test/$exit
      -- CP-element group 9: 	 branch_block_stmt_1635/if_stmt_1705_eval_test/EQ_u1_u1_1708/$entry
      -- CP-element group 9: 	 branch_block_stmt_1635/if_stmt_1705_eval_test/EQ_u1_u1_1708/$exit
      -- CP-element group 9: 	 branch_block_stmt_1635/if_stmt_1705_eval_test/EQ_u1_u1_1708/EQ_u1_u1_1708_inputs/$entry
      -- CP-element group 9: 	 branch_block_stmt_1635/if_stmt_1705_eval_test/EQ_u1_u1_1708/EQ_u1_u1_1708_inputs/$exit
      -- CP-element group 9: 	 branch_block_stmt_1635/if_stmt_1705_eval_test/EQ_u1_u1_1708/SplitProtocol/$entry
      -- CP-element group 9: 	 branch_block_stmt_1635/if_stmt_1705_eval_test/EQ_u1_u1_1708/SplitProtocol/$exit
      -- CP-element group 9: 	 branch_block_stmt_1635/if_stmt_1705_eval_test/EQ_u1_u1_1708/SplitProtocol/Sample/$entry
      -- CP-element group 9: 	 branch_block_stmt_1635/if_stmt_1705_eval_test/EQ_u1_u1_1708/SplitProtocol/Sample/$exit
      -- CP-element group 9: 	 branch_block_stmt_1635/if_stmt_1705_eval_test/EQ_u1_u1_1708/SplitProtocol/Sample/rr
      -- CP-element group 9: 	 branch_block_stmt_1635/if_stmt_1705_eval_test/EQ_u1_u1_1708/SplitProtocol/Sample/ra
      -- CP-element group 9: 	 branch_block_stmt_1635/if_stmt_1705_eval_test/EQ_u1_u1_1708/SplitProtocol/Update/$entry
      -- CP-element group 9: 	 branch_block_stmt_1635/if_stmt_1705_eval_test/EQ_u1_u1_1708/SplitProtocol/Update/$exit
      -- CP-element group 9: 	 branch_block_stmt_1635/if_stmt_1705_eval_test/EQ_u1_u1_1708/SplitProtocol/Update/cr
      -- CP-element group 9: 	 branch_block_stmt_1635/if_stmt_1705_eval_test/EQ_u1_u1_1708/SplitProtocol/Update/ca
      -- CP-element group 9: 	 branch_block_stmt_1635/if_stmt_1705_eval_test/branch_req
      -- CP-element group 9: 	 branch_block_stmt_1635/EQ_u1_u1_1708_place
      -- CP-element group 9: 	 branch_block_stmt_1635/if_stmt_1705_if_link/$entry
      -- CP-element group 9: 	 branch_block_stmt_1635/if_stmt_1705_else_link/$entry
      -- 
    cca_2297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1704_call_ack_1, ack => populateRxQueue_CP_2199_elements(9)); -- 
    branch_req_2324_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_2324_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_2199_elements(9), ack => if_stmt_1705_branch_req_0); -- 
    -- CP-element group 10:  fork  transition  place  input  output  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	9 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	18 
    -- CP-element group 10: 	19 
    -- CP-element group 10:  members (11) 
      -- CP-element group 10: 	 branch_block_stmt_1635/loopback_PhiReq/phi_stmt_1637/phi_stmt_1637_sources/Interlock/Sample/$entry
      -- CP-element group 10: 	 branch_block_stmt_1635/loopback_PhiReq/phi_stmt_1637/phi_stmt_1637_sources/Interlock/Sample/req
      -- CP-element group 10: 	 branch_block_stmt_1635/loopback_PhiReq/phi_stmt_1637/phi_stmt_1637_sources/Interlock/Update/req
      -- CP-element group 10: 	 branch_block_stmt_1635/loopback_PhiReq/phi_stmt_1637/phi_stmt_1637_sources/Interlock/$entry
      -- CP-element group 10: 	 branch_block_stmt_1635/loopback_PhiReq/phi_stmt_1637/phi_stmt_1637_sources/Interlock/Update/$entry
      -- CP-element group 10: 	 branch_block_stmt_1635/loopback_PhiReq/phi_stmt_1637/phi_stmt_1637_sources/$entry
      -- CP-element group 10: 	 branch_block_stmt_1635/loopback_PhiReq/phi_stmt_1637/$entry
      -- CP-element group 10: 	 branch_block_stmt_1635/loopback_PhiReq/$entry
      -- CP-element group 10: 	 branch_block_stmt_1635/if_stmt_1705_if_link/$exit
      -- CP-element group 10: 	 branch_block_stmt_1635/if_stmt_1705_if_link/if_choice_transition
      -- CP-element group 10: 	 branch_block_stmt_1635/loopback
      -- 
    if_choice_transition_2329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1705_branch_ack_1, ack => populateRxQueue_CP_2199_elements(10)); -- 
    req_2482_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2482_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_2199_elements(10), ack => n_q_index_1695_1647_buf_req_0); -- 
    req_2487_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2487_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_2199_elements(10), ack => n_q_index_1695_1647_buf_req_1); -- 
    -- CP-element group 11:  merge  transition  place  input  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	9 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	1 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 branch_block_stmt_1635/if_stmt_1705__exit__
      -- CP-element group 11: 	 branch_block_stmt_1635/if_stmt_1705_else_link/$exit
      -- CP-element group 11: 	 branch_block_stmt_1635/if_stmt_1705_else_link/else_choice_transition
      -- 
    else_choice_transition_2333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 11_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_1705_branch_ack_0, ack => populateRxQueue_CP_2199_elements(11)); -- 
    -- CP-element group 12:  transition  input  output  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	7 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_1635/assign_stmt_1714/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1712_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1635/assign_stmt_1714/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1712_update_start_
      -- CP-element group 12: 	 branch_block_stmt_1635/assign_stmt_1714/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1712_Sample/$exit
      -- CP-element group 12: 	 branch_block_stmt_1635/assign_stmt_1714/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1712_Sample/ack
      -- CP-element group 12: 	 branch_block_stmt_1635/assign_stmt_1714/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1712_Update/$entry
      -- CP-element group 12: 	 branch_block_stmt_1635/assign_stmt_1714/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1712_Update/req
      -- 
    ack_2348_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1712_inst_ack_0, ack => populateRxQueue_CP_2199_elements(12)); -- 
    req_2352_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2352_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_2199_elements(12), ack => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1712_inst_req_1); -- 
    -- CP-element group 13:  transition  place  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	1 
    -- CP-element group 13:  members (5) 
      -- CP-element group 13: 	 branch_block_stmt_1635/assign_stmt_1714__exit__
      -- CP-element group 13: 	 branch_block_stmt_1635/assign_stmt_1714/$exit
      -- CP-element group 13: 	 branch_block_stmt_1635/assign_stmt_1714/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1712_update_completed_
      -- CP-element group 13: 	 branch_block_stmt_1635/assign_stmt_1714/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1712_Update/$exit
      -- CP-element group 13: 	 branch_block_stmt_1635/assign_stmt_1714/WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1712_Update/ack
      -- 
    ack_2353_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1712_inst_ack_1, ack => populateRxQueue_CP_2199_elements(13)); -- 
    -- CP-element group 14:  join  fork  transition  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	0 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	16 
    -- CP-element group 14:  members (71) 
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/SplitProtocol/$entry
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/SUB_u32_u32_1644/SplitProtocol/Update/ca
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/SplitProtocol/Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/SUB_u32_u32_1644/SplitProtocol/Update/cr
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/SplitProtocol/Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/SUB_u32_u32_1644/SplitProtocol/Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/SUB_u32_u32_1644/SplitProtocol/Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/SplitProtocol/Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/SplitProtocol/$exit
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/SplitProtocol/Update/cr
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/SplitProtocol/Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/SplitProtocol/Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/SplitProtocol/Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/SUB_u32_u32_1644/SplitProtocol/Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/SUB_u32_u32_1644/SplitProtocol/Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/SplitProtocol/Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/SUB_u32_u32_1644/SplitProtocol/Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/SplitProtocol/$entry
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/SplitProtocol/Update/ca
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/SplitProtocol/Update/cr
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/SplitProtocol/Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/SUB_u32_u32_1644/SplitProtocol/Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/SplitProtocol/Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/$entry
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/$entry
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/$entry
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/$entry
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/$entry
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/$exit
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/ADD_u6_u6_1641/$entry
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/ADD_u6_u6_1641/$exit
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/ADD_u6_u6_1641/ADD_u6_u6_1641_inputs/$entry
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/ADD_u6_u6_1641/ADD_u6_u6_1641_inputs/$exit
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/ADD_u6_u6_1641/ADD_u6_u6_1641_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1639/$entry
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/ADD_u6_u6_1641/ADD_u6_u6_1641_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1639/$exit
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/ADD_u6_u6_1641/ADD_u6_u6_1641_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1639/Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/ADD_u6_u6_1641/ADD_u6_u6_1641_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1639/Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/ADD_u6_u6_1641/ADD_u6_u6_1641_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1639/Sample/req
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/ADD_u6_u6_1641/ADD_u6_u6_1641_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1639/Sample/ack
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/ADD_u6_u6_1641/ADD_u6_u6_1641_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1639/Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/ADD_u6_u6_1641/ADD_u6_u6_1641_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1639/Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/ADD_u6_u6_1641/ADD_u6_u6_1641_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1639/Update/req
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/ADD_u6_u6_1641/ADD_u6_u6_1641_inputs/RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1639/Update/ack
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/ADD_u6_u6_1641/SplitProtocol/$entry
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/ADD_u6_u6_1641/SplitProtocol/$exit
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/ADD_u6_u6_1641/SplitProtocol/Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/ADD_u6_u6_1641/SplitProtocol/Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/ADD_u6_u6_1641/SplitProtocol/Sample/rr
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/ADD_u6_u6_1641/SplitProtocol/Sample/ra
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/ADD_u6_u6_1641/SplitProtocol/Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/ADD_u6_u6_1641/SplitProtocol/Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/ADD_u6_u6_1641/SplitProtocol/Update/cr
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/ADD_u6_u6_1641/SplitProtocol/Update/ca
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/$entry
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/$exit
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/SUB_u32_u32_1644/$entry
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/SUB_u32_u32_1644/$exit
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/SUB_u32_u32_1644/SUB_u32_u32_1644_inputs/$entry
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/SUB_u32_u32_1644/SUB_u32_u32_1644_inputs/$exit
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/SUB_u32_u32_1644/SUB_u32_u32_1644_inputs/RPIPE_NUMBER_OF_SERVERS_1642/$entry
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/SUB_u32_u32_1644/SUB_u32_u32_1644_inputs/RPIPE_NUMBER_OF_SERVERS_1642/$exit
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/SUB_u32_u32_1644/SUB_u32_u32_1644_inputs/RPIPE_NUMBER_OF_SERVERS_1642/Sample/$entry
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/SUB_u32_u32_1644/SUB_u32_u32_1644_inputs/RPIPE_NUMBER_OF_SERVERS_1642/Sample/$exit
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/SUB_u32_u32_1644/SUB_u32_u32_1644_inputs/RPIPE_NUMBER_OF_SERVERS_1642/Sample/req
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/SUB_u32_u32_1644/SUB_u32_u32_1644_inputs/RPIPE_NUMBER_OF_SERVERS_1642/Sample/ack
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/SUB_u32_u32_1644/SUB_u32_u32_1644_inputs/RPIPE_NUMBER_OF_SERVERS_1642/Update/$entry
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/SUB_u32_u32_1644/SUB_u32_u32_1644_inputs/RPIPE_NUMBER_OF_SERVERS_1642/Update/$exit
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/SUB_u32_u32_1644/SUB_u32_u32_1644_inputs/RPIPE_NUMBER_OF_SERVERS_1642/Update/req
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/SUB_u32_u32_1644/SUB_u32_u32_1644_inputs/RPIPE_NUMBER_OF_SERVERS_1642/Update/ack
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/SUB_u32_u32_1644/SplitProtocol/$entry
      -- CP-element group 14: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/AND_u6_u6_1646_inputs/type_cast_1645/SUB_u32_u32_1644/SplitProtocol/$exit
      -- 
    rr_2459_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2459_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_2199_elements(14), ack => AND_u6_u6_1646_inst_req_0); -- 
    cr_2464_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2464_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_2199_elements(14), ack => AND_u6_u6_1646_inst_req_1); -- 
    populateRxQueue_CP_2199_elements(14) <= populateRxQueue_CP_2199_elements(0);
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	17 
    -- CP-element group 15:  members (2) 
      -- CP-element group 15: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/SplitProtocol/Sample/ra
      -- CP-element group 15: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/SplitProtocol/Sample/$exit
      -- 
    ra_2460_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u6_u6_1646_inst_ack_0, ack => populateRxQueue_CP_2199_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/SplitProtocol/Update/$exit
      -- CP-element group 16: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/SplitProtocol/Update/ca
      -- 
    ca_2465_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u6_u6_1646_inst_ack_1, ack => populateRxQueue_CP_2199_elements(16)); -- 
    -- CP-element group 17:  join  transition  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	15 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	21 
    -- CP-element group 17:  members (6) 
      -- CP-element group 17: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/SplitProtocol/$exit
      -- CP-element group 17: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_req
      -- CP-element group 17: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/$exit
      -- CP-element group 17: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/$exit
      -- CP-element group 17: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/$exit
      -- CP-element group 17: 	 branch_block_stmt_1635/merge_stmt_1636__entry___PhiReq/phi_stmt_1637/phi_stmt_1637_sources/AND_u6_u6_1646/$exit
      -- 
    phi_stmt_1637_req_2466_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1637_req_2466_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_2199_elements(17), ack => phi_stmt_1637_req_0); -- 
    populateRxQueue_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "populateRxQueue_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= populateRxQueue_CP_2199_elements(15) & populateRxQueue_CP_2199_elements(16);
      gj_populateRxQueue_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => populateRxQueue_CP_2199_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	10 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	20 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1635/loopback_PhiReq/phi_stmt_1637/phi_stmt_1637_sources/Interlock/Sample/$exit
      -- CP-element group 18: 	 branch_block_stmt_1635/loopback_PhiReq/phi_stmt_1637/phi_stmt_1637_sources/Interlock/Sample/ack
      -- 
    ack_2483_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_q_index_1695_1647_buf_ack_0, ack => populateRxQueue_CP_2199_elements(18)); -- 
    -- CP-element group 19:  transition  input  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	10 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_1635/loopback_PhiReq/phi_stmt_1637/phi_stmt_1637_sources/Interlock/Update/$exit
      -- CP-element group 19: 	 branch_block_stmt_1635/loopback_PhiReq/phi_stmt_1637/phi_stmt_1637_sources/Interlock/Update/ack
      -- 
    ack_2488_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_q_index_1695_1647_buf_ack_1, ack => populateRxQueue_CP_2199_elements(19)); -- 
    -- CP-element group 20:  join  transition  output  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	18 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	21 
    -- CP-element group 20:  members (5) 
      -- CP-element group 20: 	 branch_block_stmt_1635/loopback_PhiReq/phi_stmt_1637/phi_stmt_1637_sources/Interlock/$exit
      -- CP-element group 20: 	 branch_block_stmt_1635/loopback_PhiReq/phi_stmt_1637/phi_stmt_1637_req
      -- CP-element group 20: 	 branch_block_stmt_1635/loopback_PhiReq/phi_stmt_1637/phi_stmt_1637_sources/$exit
      -- CP-element group 20: 	 branch_block_stmt_1635/loopback_PhiReq/phi_stmt_1637/$exit
      -- CP-element group 20: 	 branch_block_stmt_1635/loopback_PhiReq/$exit
      -- 
    phi_stmt_1637_req_2489_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1637_req_2489_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_2199_elements(20), ack => phi_stmt_1637_req_1); -- 
    populateRxQueue_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 35) := "populateRxQueue_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= populateRxQueue_CP_2199_elements(18) & populateRxQueue_CP_2199_elements(19);
      gj_populateRxQueue_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => populateRxQueue_CP_2199_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  merge  transition  place  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	17 
    -- CP-element group 21: 	20 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	22 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_1635/merge_stmt_1636_PhiAck/$entry
      -- CP-element group 21: 	 branch_block_stmt_1635/merge_stmt_1636_PhiReqMerge
      -- 
    populateRxQueue_CP_2199_elements(21) <= OrReduce(populateRxQueue_CP_2199_elements(17) & populateRxQueue_CP_2199_elements(20));
    -- CP-element group 22:  merge  fork  transition  place  input  output  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	21 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	2 
    -- CP-element group 22: 	3 
    -- CP-element group 22: 	5 
    -- CP-element group 22:  members (14) 
      -- CP-element group 22: 	 branch_block_stmt_1635/merge_stmt_1636_PhiAck/$exit
      -- CP-element group 22: 	 branch_block_stmt_1635/merge_stmt_1636_PhiAck/phi_stmt_1637_ack
      -- CP-element group 22: 	 branch_block_stmt_1635/merge_stmt_1636__exit__
      -- CP-element group 22: 	 branch_block_stmt_1635/assign_stmt_1656_to_assign_stmt_1695__entry__
      -- CP-element group 22: 	 branch_block_stmt_1635/assign_stmt_1656_to_assign_stmt_1695/$entry
      -- CP-element group 22: 	 branch_block_stmt_1635/assign_stmt_1656_to_assign_stmt_1695/call_stmt_1668_sample_start_
      -- CP-element group 22: 	 branch_block_stmt_1635/assign_stmt_1656_to_assign_stmt_1695/call_stmt_1668_update_start_
      -- CP-element group 22: 	 branch_block_stmt_1635/assign_stmt_1656_to_assign_stmt_1695/call_stmt_1668_Sample/$entry
      -- CP-element group 22: 	 branch_block_stmt_1635/assign_stmt_1656_to_assign_stmt_1695/call_stmt_1668_Sample/crr
      -- CP-element group 22: 	 branch_block_stmt_1635/assign_stmt_1656_to_assign_stmt_1695/call_stmt_1668_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_1635/assign_stmt_1656_to_assign_stmt_1695/call_stmt_1668_Update/ccr
      -- CP-element group 22: 	 branch_block_stmt_1635/assign_stmt_1656_to_assign_stmt_1695/call_stmt_1685_update_start_
      -- CP-element group 22: 	 branch_block_stmt_1635/assign_stmt_1656_to_assign_stmt_1695/call_stmt_1685_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_1635/assign_stmt_1656_to_assign_stmt_1695/call_stmt_1685_Update/ccr
      -- 
    phi_stmt_1637_ack_2494_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1637_ack_0, ack => populateRxQueue_CP_2199_elements(22)); -- 
    crr_2223_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2223_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_2199_elements(22), ack => call_stmt_1668_call_req_0); -- 
    ccr_2228_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2228_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_2199_elements(22), ack => call_stmt_1668_call_req_1); -- 
    ccr_2242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => populateRxQueue_CP_2199_elements(22), ack => call_stmt_1685_call_req_1); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u6_u6_1641_wire : std_logic_vector(5 downto 0);
    signal ADD_u6_u6_1654_wire : std_logic_vector(5 downto 0);
    signal ADD_u6_u6_1689_wire : std_logic_vector(5 downto 0);
    signal AND_u6_u6_1646_wire : std_logic_vector(5 downto 0);
    signal EQ_u1_u1_1708_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1701_wire : std_logic_vector(0 downto 0);
    signal NOT_u4_u4_1663_wire_constant : std_logic_vector(3 downto 0);
    signal RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1639_wire : std_logic_vector(5 downto 0);
    signal RPIPE_NUMBER_OF_SERVERS_1642_wire : std_logic_vector(31 downto 0);
    signal RPIPE_NUMBER_OF_SERVERS_1690_wire : std_logic_vector(31 downto 0);
    signal R_RX_QUEUES_REG_START_OFFSET_1653_wire_constant : std_logic_vector(5 downto 0);
    signal SUB_u32_u32_1644_wire : std_logic_vector(31 downto 0);
    signal SUB_u32_u32_1692_wire : std_logic_vector(31 downto 0);
    signal konst_1640_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1643_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1688_wire_constant : std_logic_vector(5 downto 0);
    signal konst_1691_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1702_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1707_wire_constant : std_logic_vector(0 downto 0);
    signal n_q_index_1695 : std_logic_vector(5 downto 0);
    signal n_q_index_1695_1647_buffered : std_logic_vector(5 downto 0);
    signal push_status_1685 : std_logic_vector(0 downto 0);
    signal q_index_1637 : std_logic_vector(5 downto 0);
    signal register_index_1656 : std_logic_vector(5 downto 0);
    signal rx_queue_pointer_32_1668 : std_logic_vector(31 downto 0);
    signal rx_queue_pointer_36_1674 : std_logic_vector(35 downto 0);
    signal slice_1683_wire : std_logic_vector(31 downto 0);
    signal status_1704 : std_logic_vector(0 downto 0);
    signal type_cast_1645_wire : std_logic_vector(5 downto 0);
    signal type_cast_1660_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1666_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1671_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_1680_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1693_wire : std_logic_vector(5 downto 0);
    -- 
  begin -- 
    NOT_u4_u4_1663_wire_constant <= "1111";
    R_RX_QUEUES_REG_START_OFFSET_1653_wire_constant <= "000010";
    konst_1640_wire_constant <= "000001";
    konst_1643_wire_constant <= "00000000000000000000000000000001";
    konst_1688_wire_constant <= "000001";
    konst_1691_wire_constant <= "00000000000000000000000000000001";
    konst_1702_wire_constant <= "00000000000000000000000000100000";
    konst_1707_wire_constant <= "0";
    type_cast_1660_wire_constant <= "1";
    type_cast_1666_wire_constant <= "00000000000000000000000000000000";
    type_cast_1671_wire_constant <= "0000";
    type_cast_1680_wire_constant <= "1";
    phi_stmt_1637: Block -- phi operator 
      signal idata: std_logic_vector(11 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= AND_u6_u6_1646_wire & n_q_index_1695_1647_buffered;
      req <= phi_stmt_1637_req_0 & phi_stmt_1637_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1637",
          num_reqs => 2,
          bypass_flag => false,
          data_width => 6) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1637_ack_0,
          idata => idata,
          odata => q_index_1637,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1637
    -- flow-through slice operator slice_1683_inst
    slice_1683_wire <= rx_buffer_pointer_buffer(31 downto 0);
    n_q_index_1695_1647_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_q_index_1695_1647_buf_req_0;
      n_q_index_1695_1647_buf_ack_0<= wack(0);
      rreq(0) <= n_q_index_1695_1647_buf_req_1;
      n_q_index_1695_1647_buf_ack_1<= rack(0);
      n_q_index_1695_1647_buf : InterlockBuffer generic map ( -- 
        name => "n_q_index_1695_1647_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 6,
        out_data_width => 6,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_q_index_1695,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_q_index_1695_1647_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_1645_inst
    process(SUB_u32_u32_1644_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := SUB_u32_u32_1644_wire(5 downto 0);
      type_cast_1645_wire <= tmp_var; -- 
    end process;
    -- interlock type_cast_1655_inst
    process(ADD_u6_u6_1654_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := ADD_u6_u6_1654_wire(5 downto 0);
      register_index_1656 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1693_inst
    process(SUB_u32_u32_1692_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := SUB_u32_u32_1692_wire(5 downto 0);
      type_cast_1693_wire <= tmp_var; -- 
    end process;
    if_stmt_1699_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_1701_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1699_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1699_branch_req_0,
          ack0 => if_stmt_1699_branch_ack_0,
          ack1 => if_stmt_1699_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_1705_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= EQ_u1_u1_1708_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_1705_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_1705_branch_req_0,
          ack0 => if_stmt_1705_branch_ack_0,
          ack1 => if_stmt_1705_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u6_u6_1641_inst
    process(RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1639_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1639_wire, konst_1640_wire_constant, tmp_var);
      ADD_u6_u6_1641_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u6_u6_1654_inst
    process(q_index_1637) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_index_1637, R_RX_QUEUES_REG_START_OFFSET_1653_wire_constant, tmp_var);
      ADD_u6_u6_1654_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u6_u6_1689_inst
    process(q_index_1637) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_index_1637, konst_1688_wire_constant, tmp_var);
      ADD_u6_u6_1689_wire <= tmp_var; --
    end process;
    -- shared split operator group (3) : AND_u6_u6_1646_inst 
    ApIntAnd_group_3: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ADD_u6_u6_1641_wire & type_cast_1645_wire;
      AND_u6_u6_1646_wire <= data_out(5 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u6_u6_1646_inst_req_0;
      AND_u6_u6_1646_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u6_u6_1646_inst_req_1;
      AND_u6_u6_1646_inst_ack_1 <= ackR_unguarded(0);
      ApIntAnd_group_3_gI: SplitGuardInterface generic map(name => "ApIntAnd_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 6, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- binary operator AND_u6_u6_1694_inst
    process(ADD_u6_u6_1689_wire, type_cast_1693_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAnd_proc(ADD_u6_u6_1689_wire, type_cast_1693_wire, tmp_var);
      n_q_index_1695 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u4_u36_1673_inst
    process(type_cast_1671_wire_constant, rx_queue_pointer_32_1668) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1671_wire_constant, rx_queue_pointer_32_1668, tmp_var);
      rx_queue_pointer_36_1674 <= tmp_var; --
    end process;
    -- binary operator EQ_u1_u1_1708_inst
    process(status_1704) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(status_1704, konst_1707_wire_constant, tmp_var);
      EQ_u1_u1_1708_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1701_inst
    process(push_status_1685) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", push_status_1685, tmp_var);
      NOT_u1_u1_1701_wire <= tmp_var; -- 
    end process;
    -- binary operator SUB_u32_u32_1644_inst
    process(RPIPE_NUMBER_OF_SERVERS_1642_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(RPIPE_NUMBER_OF_SERVERS_1642_wire, konst_1643_wire_constant, tmp_var);
      SUB_u32_u32_1644_wire <= tmp_var; --
    end process;
    -- binary operator SUB_u32_u32_1692_inst
    process(RPIPE_NUMBER_OF_SERVERS_1690_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(RPIPE_NUMBER_OF_SERVERS_1690_wire, konst_1691_wire_constant, tmp_var);
      SUB_u32_u32_1692_wire <= tmp_var; --
    end process;
    -- read from input-signal LAST_WRITTEN_RX_QUEUE_INDEX
    RPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1639_wire <= LAST_WRITTEN_RX_QUEUE_INDEX;
    -- read from input-signal NUMBER_OF_SERVERS
    RPIPE_NUMBER_OF_SERVERS_1690_wire <= NUMBER_OF_SERVERS;
    RPIPE_NUMBER_OF_SERVERS_1642_wire <= NUMBER_OF_SERVERS;
    -- shared outport operator group (0) : WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1712_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1712_inst_req_0;
      WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1712_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1712_inst_req_1;
      WPIPE_LAST_WRITTEN_RX_QUEUE_INDEX_1712_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= q_index_1637;
      LAST_WRITTEN_RX_QUEUE_INDEX_write_0_gI: SplitGuardInterface generic map(name => "LAST_WRITTEN_RX_QUEUE_INDEX_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      LAST_WRITTEN_RX_QUEUE_INDEX_write_0: OutputPortRevised -- 
        generic map ( name => "LAST_WRITTEN_RX_QUEUE_INDEX", data_width => 6, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req(0),
          oack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack(0),
          odata => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data(5 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared call operator group (0) : call_stmt_1668_call 
    AccessRegister_call_group_0: Block -- 
      signal data_in: std_logic_vector(42 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1668_call_req_0;
      call_stmt_1668_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1668_call_req_1;
      call_stmt_1668_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      AccessRegister_call_group_0_gI: SplitGuardInterface generic map(name => "AccessRegister_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1660_wire_constant & NOT_u4_u4_1663_wire_constant & register_index_1656 & type_cast_1666_wire_constant;
      rx_queue_pointer_32_1668 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 43,
        owidth => 43,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => AccessRegister_call_reqs(0),
          ackR => AccessRegister_call_acks(0),
          dataR => AccessRegister_call_data(42 downto 0),
          tagR => AccessRegister_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => AccessRegister_return_acks(0), -- cross-over
          ackL => AccessRegister_return_reqs(0), -- cross-over
          dataL => AccessRegister_return_data(31 downto 0),
          tagL => AccessRegister_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1685_call 
    pushIntoQueue_call_group_1: Block -- 
      signal data_in: std_logic_vector(68 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1685_call_req_0;
      call_stmt_1685_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1685_call_req_1;
      call_stmt_1685_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      pushIntoQueue_call_group_1_gI: SplitGuardInterface generic map(name => "pushIntoQueue_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1680_wire_constant & rx_queue_pointer_36_1674 & slice_1683_wire;
      push_status_1685 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 69,
        owidth => 69,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => pushIntoQueue_call_reqs(0),
          ackR => pushIntoQueue_call_acks(0),
          dataR => pushIntoQueue_call_data(68 downto 0),
          tagR => pushIntoQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => pushIntoQueue_return_acks(0), -- cross-over
          ackL => pushIntoQueue_return_reqs(0), -- cross-over
          dataL => pushIntoQueue_return_data(0 downto 0),
          tagL => pushIntoQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    operator_delay_time_3871_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_stmt_1704_call_req_0;
      call_stmt_1704_call_ack_0<= sample_ack(0);
      update_req(0) <= call_stmt_1704_call_req_1;
      call_stmt_1704_call_ack_1<= update_ack(0);
      call_stmt_1704_call: delay_time_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        T => konst_1702_wire_constant,
        delay_done => status_1704,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    -- 
  end Block; -- data_path
  -- 
end populateRxQueue_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.nic_system_global_package.all;
entity pushIntoQueue is -- 
  generic (tag_length : integer); 
  port ( -- 
    lock : in  std_logic_vector(0 downto 0);
    q_base_address : in  std_logic_vector(35 downto 0);
    q_w_data : in  std_logic_vector(31 downto 0);
    status : out  std_logic_vector(0 downto 0);
    releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
    releaseLock_call_acks : in   std_logic_vector(0 downto 0);
    releaseLock_call_data : out  std_logic_vector(35 downto 0);
    releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
    releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
    releaseLock_return_acks : in   std_logic_vector(0 downto 0);
    releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
    setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
    setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
    setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
    setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
    setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
    setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
    setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
    acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
    acquireLock_call_acks : in   std_logic_vector(0 downto 0);
    acquireLock_call_data : out  std_logic_vector(35 downto 0);
    acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
    acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
    acquireLock_return_acks : in   std_logic_vector(0 downto 0);
    acquireLock_return_data : in   std_logic_vector(0 downto 0);
    acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    updateTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
    updateTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
    updateTotalMessages_call_data : out  std_logic_vector(67 downto 0);
    updateTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
    updateTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
    updateTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
    updateTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
    getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
    getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
    getTotalMessages_call_data : out  std_logic_vector(35 downto 0);
    getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
    getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
    getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
    getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
    getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
    getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
    getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
    getQueueLength_call_data : out  std_logic_vector(35 downto 0);
    getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
    getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
    getQueueLength_return_data : in   std_logic_vector(31 downto 0);
    getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
    getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
    getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
    getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
    getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
    getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
    getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
    getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
    getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
    setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
    setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
    setQueueElement_call_data : out  std_logic_vector(99 downto 0);
    setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
    setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
    setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
    setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity pushIntoQueue;
architecture pushIntoQueue_arch of pushIntoQueue is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 69)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 1)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal lock_buffer :  std_logic_vector(0 downto 0);
  signal lock_update_enable: Boolean;
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  signal q_w_data_buffer :  std_logic_vector(31 downto 0);
  signal q_w_data_update_enable: Boolean;
  -- output port buffer signals
  signal status_buffer :  std_logic_vector(0 downto 0);
  signal status_update_enable: Boolean;
  signal pushIntoQueue_CP_1948_start: Boolean;
  signal pushIntoQueue_CP_1948_symbol: Boolean;
  -- volatile/operator module components. 
  component releaseLock is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component setQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : in  std_logic_vector(31 downto 0);
      rp : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component acquireLock is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      m_ok : out  std_logic_vector(0 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component updateTotalMessages is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      updated_total_msgs : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getTotalMessages is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      total_msgs : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getQueueLength is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      Queue_Length : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : out  std_logic_vector(31 downto 0);
      rp : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component setQueueElement is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      write_index : in  std_logic_vector(31 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1589_call_req_1 : boolean;
  signal call_stmt_1596_call_ack_1 : boolean;
  signal call_stmt_1596_call_req_0 : boolean;
  signal NOT_u1_u1_1603_inst_req_0 : boolean;
  signal call_stmt_1539_call_req_0 : boolean;
  signal call_stmt_1539_call_req_1 : boolean;
  signal call_stmt_1547_call_req_1 : boolean;
  signal call_stmt_1589_call_ack_0 : boolean;
  signal call_stmt_1539_call_ack_0 : boolean;
  signal call_stmt_1589_call_ack_1 : boolean;
  signal call_stmt_1539_call_ack_1 : boolean;
  signal NOT_u1_u1_1603_inst_ack_0 : boolean;
  signal call_stmt_1547_call_ack_1 : boolean;
  signal call_stmt_1596_call_req_1 : boolean;
  signal call_stmt_1596_call_ack_0 : boolean;
  signal call_stmt_1589_call_req_0 : boolean;
  signal call_stmt_1600_call_ack_1 : boolean;
  signal call_stmt_1600_call_req_1 : boolean;
  signal call_stmt_1525_call_ack_1 : boolean;
  signal call_stmt_1584_call_ack_1 : boolean;
  signal call_stmt_1525_call_req_1 : boolean;
  signal call_stmt_1584_call_req_1 : boolean;
  signal call_stmt_1584_call_ack_0 : boolean;
  signal call_stmt_1550_call_ack_1 : boolean;
  signal call_stmt_1584_call_req_0 : boolean;
  signal call_stmt_1550_call_req_1 : boolean;
  signal call_stmt_1600_call_ack_0 : boolean;
  signal call_stmt_1525_call_ack_0 : boolean;
  signal call_stmt_1525_call_req_0 : boolean;
  signal call_stmt_1550_call_ack_0 : boolean;
  signal call_stmt_1550_call_req_0 : boolean;
  signal call_stmt_1553_call_ack_1 : boolean;
  signal call_stmt_1600_call_req_0 : boolean;
  signal NOT_u1_u1_1603_inst_ack_1 : boolean;
  signal call_stmt_1547_call_ack_0 : boolean;
  signal call_stmt_1553_call_req_1 : boolean;
  signal NOT_u1_u1_1603_inst_req_1 : boolean;
  signal call_stmt_1553_call_ack_0 : boolean;
  signal call_stmt_1553_call_req_0 : boolean;
  signal call_stmt_1547_call_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "pushIntoQueue_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 69) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= lock;
  lock_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(36 downto 1) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(36 downto 1);
  in_buffer_data_in(68 downto 37) <= q_w_data;
  q_w_data_buffer <= in_buffer_data_out(68 downto 37);
  in_buffer_data_in(tag_length + 68 downto 69) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 68 downto 69);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  pushIntoQueue_CP_1948_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "pushIntoQueue_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 1) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(0 downto 0) <= status_buffer;
  status <= out_buffer_data_out(0 downto 0);
  out_buffer_data_in(tag_length + 0 downto 1) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 0 downto 1);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= pushIntoQueue_CP_1948_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= pushIntoQueue_CP_1948_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= pushIntoQueue_CP_1948_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  pushIntoQueue_CP_1948: Block -- control-path 
    signal pushIntoQueue_CP_1948_elements: BooleanArray(24 downto 0);
    -- 
  begin -- 
    pushIntoQueue_CP_1948_elements(0) <= pushIntoQueue_CP_1948_start;
    pushIntoQueue_CP_1948_symbol <= pushIntoQueue_CP_1948_elements(24);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 call_stmt_1525_to_call_stmt_1539/call_stmt_1525_update_start_
      -- CP-element group 0: 	 call_stmt_1525_to_call_stmt_1539/call_stmt_1539_update_start_
      -- CP-element group 0: 	 call_stmt_1525_to_call_stmt_1539/call_stmt_1539_Update/ccr
      -- CP-element group 0: 	 call_stmt_1525_to_call_stmt_1539/call_stmt_1525_sample_start_
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_1525_to_call_stmt_1539/call_stmt_1539_Update/$entry
      -- CP-element group 0: 	 call_stmt_1525_to_call_stmt_1539/$entry
      -- CP-element group 0: 	 call_stmt_1525_to_call_stmt_1539/call_stmt_1525_Update/ccr
      -- CP-element group 0: 	 call_stmt_1525_to_call_stmt_1539/call_stmt_1525_Update/$entry
      -- CP-element group 0: 	 call_stmt_1525_to_call_stmt_1539/call_stmt_1525_Sample/crr
      -- CP-element group 0: 	 call_stmt_1525_to_call_stmt_1539/call_stmt_1525_Sample/$entry
      -- 
    crr_1961_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1961_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1948_elements(0), ack => call_stmt_1525_call_req_0); -- 
    ccr_1966_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1966_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1948_elements(0), ack => call_stmt_1525_call_req_1); -- 
    ccr_1980_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1980_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1948_elements(0), ack => call_stmt_1539_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_1525_to_call_stmt_1539/call_stmt_1525_sample_completed_
      -- CP-element group 1: 	 call_stmt_1525_to_call_stmt_1539/call_stmt_1525_Sample/cra
      -- CP-element group 1: 	 call_stmt_1525_to_call_stmt_1539/call_stmt_1525_Sample/$exit
      -- 
    cra_1962_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1525_call_ack_0, ack => pushIntoQueue_CP_1948_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 call_stmt_1525_to_call_stmt_1539/call_stmt_1539_Sample/$entry
      -- CP-element group 2: 	 call_stmt_1525_to_call_stmt_1539/call_stmt_1539_sample_start_
      -- CP-element group 2: 	 call_stmt_1525_to_call_stmt_1539/call_stmt_1539_Sample/crr
      -- CP-element group 2: 	 call_stmt_1525_to_call_stmt_1539/call_stmt_1525_Update/cca
      -- CP-element group 2: 	 call_stmt_1525_to_call_stmt_1539/call_stmt_1525_Update/$exit
      -- CP-element group 2: 	 call_stmt_1525_to_call_stmt_1539/call_stmt_1525_update_completed_
      -- 
    cca_1967_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1525_call_ack_1, ack => pushIntoQueue_CP_1948_elements(2)); -- 
    crr_1975_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1975_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1948_elements(2), ack => call_stmt_1539_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 call_stmt_1525_to_call_stmt_1539/call_stmt_1539_Sample/$exit
      -- CP-element group 3: 	 call_stmt_1525_to_call_stmt_1539/call_stmt_1539_Sample/cra
      -- CP-element group 3: 	 call_stmt_1525_to_call_stmt_1539/call_stmt_1539_sample_completed_
      -- 
    cra_1976_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1539_call_ack_0, ack => pushIntoQueue_CP_1948_elements(3)); -- 
    -- CP-element group 4:  fork  transition  input  output  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	5 
    -- CP-element group 4: 	6 
    -- CP-element group 4: 	8 
    -- CP-element group 4: 	10 
    -- CP-element group 4: 	13 
    -- CP-element group 4: 	16 
    -- CP-element group 4: 	19 
    -- CP-element group 4:  members (26) 
      -- CP-element group 4: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1589_Update/$entry
      -- CP-element group 4: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1547_sample_start_
      -- CP-element group 4: 	 call_stmt_1547_to_call_stmt_1596/$entry
      -- CP-element group 4: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1589_Update/ccr
      -- CP-element group 4: 	 call_stmt_1525_to_call_stmt_1539/$exit
      -- CP-element group 4: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1553_update_start_
      -- CP-element group 4: 	 call_stmt_1525_to_call_stmt_1539/call_stmt_1539_Update/$exit
      -- CP-element group 4: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1547_Update/ccr
      -- CP-element group 4: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1589_update_start_
      -- CP-element group 4: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1596_Update/$entry
      -- CP-element group 4: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1547_Update/$entry
      -- CP-element group 4: 	 call_stmt_1525_to_call_stmt_1539/call_stmt_1539_update_completed_
      -- CP-element group 4: 	 call_stmt_1525_to_call_stmt_1539/call_stmt_1539_Update/cca
      -- CP-element group 4: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1596_Update/ccr
      -- CP-element group 4: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1547_update_start_
      -- CP-element group 4: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1596_update_start_
      -- CP-element group 4: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1584_Update/ccr
      -- CP-element group 4: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1584_Update/$entry
      -- CP-element group 4: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1584_update_start_
      -- CP-element group 4: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1550_Update/ccr
      -- CP-element group 4: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1550_Update/$entry
      -- CP-element group 4: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1553_Update/ccr
      -- CP-element group 4: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1553_Update/$entry
      -- CP-element group 4: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1547_Sample/crr
      -- CP-element group 4: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1547_Sample/$entry
      -- CP-element group 4: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1550_update_start_
      -- 
    cca_1981_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1539_call_ack_1, ack => pushIntoQueue_CP_1948_elements(4)); -- 
    crr_1992_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1992_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1948_elements(4), ack => call_stmt_1547_call_req_0); -- 
    ccr_1997_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1997_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1948_elements(4), ack => call_stmt_1547_call_req_1); -- 
    ccr_2011_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2011_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1948_elements(4), ack => call_stmt_1550_call_req_1); -- 
    ccr_2025_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2025_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1948_elements(4), ack => call_stmt_1553_call_req_1); -- 
    ccr_2039_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2039_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1948_elements(4), ack => call_stmt_1584_call_req_1); -- 
    ccr_2053_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2053_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1948_elements(4), ack => call_stmt_1589_call_req_1); -- 
    ccr_2067_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2067_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1948_elements(4), ack => call_stmt_1596_call_req_1); -- 
    -- CP-element group 5:  transition  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	4 
    -- CP-element group 5: successors 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1547_sample_completed_
      -- CP-element group 5: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1547_Sample/cra
      -- CP-element group 5: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1547_Sample/$exit
      -- 
    cra_1993_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1547_call_ack_0, ack => pushIntoQueue_CP_1948_elements(5)); -- 
    -- CP-element group 6:  fork  transition  input  output  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	4 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6: 	11 
    -- CP-element group 6: 	14 
    -- CP-element group 6: 	17 
    -- CP-element group 6:  members (6) 
      -- CP-element group 6: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1547_Update/$exit
      -- CP-element group 6: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1547_Update/cca
      -- CP-element group 6: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1550_Sample/crr
      -- CP-element group 6: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1550_Sample/$entry
      -- CP-element group 6: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1547_update_completed_
      -- CP-element group 6: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1550_sample_start_
      -- 
    cca_1998_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1547_call_ack_1, ack => pushIntoQueue_CP_1948_elements(6)); -- 
    crr_2006_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2006_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1948_elements(6), ack => call_stmt_1550_call_req_0); -- 
    -- CP-element group 7:  transition  input  bypass 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1550_Sample/cra
      -- CP-element group 7: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1550_Sample/$exit
      -- CP-element group 7: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1550_sample_completed_
      -- 
    cra_2007_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 7_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1550_call_ack_0, ack => pushIntoQueue_CP_1948_elements(7)); -- 
    -- CP-element group 8:  fork  transition  input  output  bypass 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	4 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8: 	11 
    -- CP-element group 8: 	14 
    -- CP-element group 8: 	17 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1553_Sample/$entry
      -- CP-element group 8: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1553_sample_start_
      -- CP-element group 8: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1550_Update/cca
      -- CP-element group 8: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1550_Update/$exit
      -- CP-element group 8: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1553_Sample/crr
      -- CP-element group 8: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1550_update_completed_
      -- 
    cca_2012_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1550_call_ack_1, ack => pushIntoQueue_CP_1948_elements(8)); -- 
    crr_2020_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2020_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1948_elements(8), ack => call_stmt_1553_call_req_0); -- 
    -- CP-element group 9:  transition  input  bypass 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1553_sample_completed_
      -- CP-element group 9: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1553_Sample/cra
      -- CP-element group 9: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1553_Sample/$exit
      -- 
    cra_2021_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1553_call_ack_0, ack => pushIntoQueue_CP_1948_elements(9)); -- 
    -- CP-element group 10:  fork  transition  input  bypass 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	4 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	11 
    -- CP-element group 10: 	17 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1553_update_completed_
      -- CP-element group 10: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1553_Update/cca
      -- CP-element group 10: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1553_Update/$exit
      -- 
    cca_2026_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 10_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1553_call_ack_1, ack => pushIntoQueue_CP_1948_elements(10)); -- 
    -- CP-element group 11:  join  transition  output  bypass 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	6 
    -- CP-element group 11: 	8 
    -- CP-element group 11: 	10 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	12 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1584_Sample/crr
      -- CP-element group 11: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1584_Sample/$entry
      -- CP-element group 11: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1584_sample_start_
      -- 
    crr_2034_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2034_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1948_elements(11), ack => call_stmt_1584_call_req_0); -- 
    pushIntoQueue_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "pushIntoQueue_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= pushIntoQueue_CP_1948_elements(6) & pushIntoQueue_CP_1948_elements(8) & pushIntoQueue_CP_1948_elements(10);
      gj_pushIntoQueue_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => pushIntoQueue_CP_1948_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  transition  input  bypass 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	11 
    -- CP-element group 12: successors 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1584_Sample/cra
      -- CP-element group 12: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1584_Sample/$exit
      -- CP-element group 12: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1584_sample_completed_
      -- 
    cra_2035_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1584_call_ack_0, ack => pushIntoQueue_CP_1948_elements(12)); -- 
    -- CP-element group 13:  transition  input  bypass 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	4 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1584_Update/cca
      -- CP-element group 13: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1584_Update/$exit
      -- CP-element group 13: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1584_update_completed_
      -- 
    cca_2040_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1584_call_ack_1, ack => pushIntoQueue_CP_1948_elements(13)); -- 
    -- CP-element group 14:  join  transition  output  bypass 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	6 
    -- CP-element group 14: 	8 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1589_Sample/$entry
      -- CP-element group 14: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1589_Sample/crr
      -- CP-element group 14: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1589_sample_start_
      -- 
    crr_2048_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2048_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1948_elements(14), ack => call_stmt_1589_call_req_0); -- 
    pushIntoQueue_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "pushIntoQueue_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= pushIntoQueue_CP_1948_elements(6) & pushIntoQueue_CP_1948_elements(8) & pushIntoQueue_CP_1948_elements(13);
      gj_pushIntoQueue_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => pushIntoQueue_CP_1948_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  transition  input  bypass 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1589_Sample/$exit
      -- CP-element group 15: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1589_Sample/cra
      -- CP-element group 15: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1589_sample_completed_
      -- 
    cra_2049_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 15_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1589_call_ack_0, ack => pushIntoQueue_CP_1948_elements(15)); -- 
    -- CP-element group 16:  transition  input  bypass 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	4 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	17 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1589_Update/$exit
      -- CP-element group 16: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1589_update_completed_
      -- CP-element group 16: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1589_Update/cca
      -- 
    cca_2054_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 16_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1589_call_ack_1, ack => pushIntoQueue_CP_1948_elements(16)); -- 
    -- CP-element group 17:  join  transition  output  bypass 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	6 
    -- CP-element group 17: 	8 
    -- CP-element group 17: 	10 
    -- CP-element group 17: 	16 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	18 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1596_Sample/crr
      -- CP-element group 17: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1596_Sample/$entry
      -- CP-element group 17: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1596_sample_start_
      -- 
    crr_2062_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2062_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1948_elements(17), ack => call_stmt_1596_call_req_0); -- 
    pushIntoQueue_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "pushIntoQueue_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= pushIntoQueue_CP_1948_elements(6) & pushIntoQueue_CP_1948_elements(8) & pushIntoQueue_CP_1948_elements(10) & pushIntoQueue_CP_1948_elements(16);
      gj_pushIntoQueue_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => pushIntoQueue_CP_1948_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  transition  input  bypass 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	17 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1596_Sample/$exit
      -- CP-element group 18: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1596_Sample/cra
      -- CP-element group 18: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1596_sample_completed_
      -- 
    cra_2063_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 18_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1596_call_ack_0, ack => pushIntoQueue_CP_1948_elements(18)); -- 
    -- CP-element group 19:  fork  transition  input  output  bypass 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	4 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	20 
    -- CP-element group 19: 	21 
    -- CP-element group 19: 	22 
    -- CP-element group 19: 	23 
    -- CP-element group 19:  members (17) 
      -- CP-element group 19: 	 call_stmt_1547_to_call_stmt_1596/$exit
      -- CP-element group 19: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1596_Update/cca
      -- CP-element group 19: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1596_Update/$exit
      -- CP-element group 19: 	 call_stmt_1600_to_assign_stmt_1604/NOT_u1_u1_1603_Sample/rr
      -- CP-element group 19: 	 call_stmt_1600_to_assign_stmt_1604/NOT_u1_u1_1603_update_start_
      -- CP-element group 19: 	 call_stmt_1600_to_assign_stmt_1604/NOT_u1_u1_1603_sample_start_
      -- CP-element group 19: 	 call_stmt_1600_to_assign_stmt_1604/NOT_u1_u1_1603_Sample/$entry
      -- CP-element group 19: 	 call_stmt_1547_to_call_stmt_1596/call_stmt_1596_update_completed_
      -- CP-element group 19: 	 call_stmt_1600_to_assign_stmt_1604/call_stmt_1600_Update/ccr
      -- CP-element group 19: 	 call_stmt_1600_to_assign_stmt_1604/call_stmt_1600_Update/$entry
      -- CP-element group 19: 	 call_stmt_1600_to_assign_stmt_1604/call_stmt_1600_sample_start_
      -- CP-element group 19: 	 call_stmt_1600_to_assign_stmt_1604/$entry
      -- CP-element group 19: 	 call_stmt_1600_to_assign_stmt_1604/call_stmt_1600_Sample/crr
      -- CP-element group 19: 	 call_stmt_1600_to_assign_stmt_1604/call_stmt_1600_Sample/$entry
      -- CP-element group 19: 	 call_stmt_1600_to_assign_stmt_1604/NOT_u1_u1_1603_Update/cr
      -- CP-element group 19: 	 call_stmt_1600_to_assign_stmt_1604/call_stmt_1600_update_start_
      -- CP-element group 19: 	 call_stmt_1600_to_assign_stmt_1604/NOT_u1_u1_1603_Update/$entry
      -- 
    cca_2068_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 19_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1596_call_ack_1, ack => pushIntoQueue_CP_1948_elements(19)); -- 
    crr_2079_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2079_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1948_elements(19), ack => call_stmt_1600_call_req_0); -- 
    ccr_2084_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2084_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1948_elements(19), ack => call_stmt_1600_call_req_1); -- 
    rr_2093_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2093_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1948_elements(19), ack => NOT_u1_u1_1603_inst_req_0); -- 
    cr_2098_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2098_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => pushIntoQueue_CP_1948_elements(19), ack => NOT_u1_u1_1603_inst_req_1); -- 
    -- CP-element group 20:  transition  input  bypass 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	19 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (3) 
      -- CP-element group 20: 	 call_stmt_1600_to_assign_stmt_1604/call_stmt_1600_Sample/cra
      -- CP-element group 20: 	 call_stmt_1600_to_assign_stmt_1604/call_stmt_1600_Sample/$exit
      -- CP-element group 20: 	 call_stmt_1600_to_assign_stmt_1604/call_stmt_1600_sample_completed_
      -- 
    cra_2080_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 20_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1600_call_ack_0, ack => pushIntoQueue_CP_1948_elements(20)); -- 
    -- CP-element group 21:  transition  input  bypass 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	19 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	24 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 call_stmt_1600_to_assign_stmt_1604/call_stmt_1600_Update/cca
      -- CP-element group 21: 	 call_stmt_1600_to_assign_stmt_1604/call_stmt_1600_Update/$exit
      -- CP-element group 21: 	 call_stmt_1600_to_assign_stmt_1604/call_stmt_1600_update_completed_
      -- 
    cca_2085_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 21_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1600_call_ack_1, ack => pushIntoQueue_CP_1948_elements(21)); -- 
    -- CP-element group 22:  transition  input  bypass 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	19 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 call_stmt_1600_to_assign_stmt_1604/NOT_u1_u1_1603_sample_completed_
      -- CP-element group 22: 	 call_stmt_1600_to_assign_stmt_1604/NOT_u1_u1_1603_Sample/ra
      -- CP-element group 22: 	 call_stmt_1600_to_assign_stmt_1604/NOT_u1_u1_1603_Sample/$exit
      -- 
    ra_2094_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 22_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1603_inst_ack_0, ack => pushIntoQueue_CP_1948_elements(22)); -- 
    -- CP-element group 23:  transition  input  bypass 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	19 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	24 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 call_stmt_1600_to_assign_stmt_1604/NOT_u1_u1_1603_update_completed_
      -- CP-element group 23: 	 call_stmt_1600_to_assign_stmt_1604/NOT_u1_u1_1603_Update/ca
      -- CP-element group 23: 	 call_stmt_1600_to_assign_stmt_1604/NOT_u1_u1_1603_Update/$exit
      -- 
    ca_2099_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_1603_inst_ack_1, ack => pushIntoQueue_CP_1948_elements(23)); -- 
    -- CP-element group 24:  join  transition  bypass 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	21 
    -- CP-element group 24: 	23 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 $exit
      -- CP-element group 24: 	 call_stmt_1600_to_assign_stmt_1604/$exit
      -- 
    pushIntoQueue_cp_element_group_24: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "pushIntoQueue_cp_element_group_24"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= pushIntoQueue_CP_1948_elements(21) & pushIntoQueue_CP_1948_elements(23);
      gj_pushIntoQueue_cp_element_group_24 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => pushIntoQueue_CP_1948_elements(24), clk => clk, reset => reset); --
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_1566_wire : std_logic_vector(31 downto 0);
    signal ADD_u32_u32_1595_wire : std_logic_vector(31 downto 0);
    signal ADD_u36_u36_1521_wire : std_logic_vector(35 downto 0);
    signal NOT_u8_u8_1518_wire_constant : std_logic_vector(7 downto 0);
    signal Queue_Length_1550 : std_logic_vector(31 downto 0);
    signal SUB_u32_u32_1558_wire : std_logic_vector(31 downto 0);
    signal ba_and_misc_1525 : std_logic_vector(63 downto 0);
    signal konst_1520_wire_constant : std_logic_vector(35 downto 0);
    signal konst_1557_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1563_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1565_wire_constant : std_logic_vector(31 downto 0);
    signal lock_n_1535 : std_logic_vector(0 downto 0);
    signal m_ok_1539 : std_logic_vector(0 downto 0);
    signal misc_1529 : std_logic_vector(31 downto 0);
    signal next_wi_1568 : std_logic_vector(31 downto 0);
    signal q_full_1573 : std_logic_vector(0 downto 0);
    signal read_index_1547 : std_logic_vector(31 downto 0);
    signal round_off_1560 : std_logic_vector(0 downto 0);
    signal total_msgs_1553 : std_logic_vector(31 downto 0);
    signal type_cast_1513_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1515_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1523_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1533_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1594_wire_constant : std_logic_vector(31 downto 0);
    signal write_index_1547 : std_logic_vector(31 downto 0);
    -- 
  begin -- 
    NOT_u8_u8_1518_wire_constant <= "11111111";
    konst_1520_wire_constant <= "000000000000000000000000000000011000";
    konst_1557_wire_constant <= "00000000000000000000000000000001";
    konst_1563_wire_constant <= "00000000000000000000000000000000";
    konst_1565_wire_constant <= "00000000000000000000000000000001";
    type_cast_1513_wire_constant <= "0";
    type_cast_1515_wire_constant <= "1";
    type_cast_1523_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1533_wire_constant <= "00000000000000000000000000000000";
    type_cast_1594_wire_constant <= "00000000000000000000000000000001";
    -- flow-through select operator MUX_1567_inst
    next_wi_1568 <= konst_1563_wire_constant when (round_off_1560(0) /=  '0') else ADD_u32_u32_1566_wire;
    -- flow-through slice operator slice_1528_inst
    misc_1529 <= ba_and_misc_1525(31 downto 0);
    -- binary operator ADD_u32_u32_1566_inst
    process(write_index_1547) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(write_index_1547, konst_1565_wire_constant, tmp_var);
      ADD_u32_u32_1566_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u32_u32_1595_inst
    process(total_msgs_1553) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntAdd_proc(total_msgs_1553, type_cast_1594_wire_constant, tmp_var);
      ADD_u32_u32_1595_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u36_u36_1521_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, konst_1520_wire_constant, tmp_var);
      ADD_u36_u36_1521_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1534_inst
    process(misc_1529) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(misc_1529, type_cast_1533_wire_constant, tmp_var);
      lock_n_1535 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1559_inst
    process(write_index_1547, SUB_u32_u32_1558_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(write_index_1547, SUB_u32_u32_1558_wire, tmp_var);
      round_off_1560 <= tmp_var; --
    end process;
    -- binary operator EQ_u32_u1_1572_inst
    process(next_wi_1568, read_index_1547) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(next_wi_1568, read_index_1547, tmp_var);
      q_full_1573 <= tmp_var; --
    end process;
    -- shared split operator group (6) : NOT_u1_u1_1603_inst 
    ApIntNot_group_6: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= q_full_1573;
      status_buffer <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NOT_u1_u1_1603_inst_req_0;
      NOT_u1_u1_1603_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NOT_u1_u1_1603_inst_req_1;
      NOT_u1_u1_1603_inst_ack_1 <= ackR_unguarded(0);
      ApIntNot_group_6_gI: SplitGuardInterface generic map(name => "ApIntNot_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNot",
          name => "ApIntNot_group_6",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- binary operator SUB_u32_u32_1558_inst
    process(Queue_Length_1550) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(Queue_Length_1550, konst_1557_wire_constant, tmp_var);
      SUB_u32_u32_1558_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_1525_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1525_call_req_0;
      call_stmt_1525_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1525_call_req_1;
      call_stmt_1525_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1513_wire_constant & type_cast_1515_wire_constant & NOT_u8_u8_1518_wire_constant & ADD_u36_u36_1521_wire & type_cast_1523_wire_constant;
      ba_and_misc_1525 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_1539_call 
    acquireLock_call_group_1: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1539_call_req_0;
      call_stmt_1539_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1539_call_req_1;
      call_stmt_1539_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= lock_n_1535(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      acquireLock_call_group_1_gI: SplitGuardInterface generic map(name => "acquireLock_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      m_ok_1539 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => acquireLock_call_reqs(0),
          ackR => acquireLock_call_acks(0),
          dataR => acquireLock_call_data(35 downto 0),
          tagR => acquireLock_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => acquireLock_return_acks(0), -- cross-over
          ackL => acquireLock_return_reqs(0), -- cross-over
          dataL => acquireLock_return_data(0 downto 0),
          tagL => acquireLock_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_1547_call 
    getQueuePointers_call_group_2: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1547_call_req_0;
      call_stmt_1547_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1547_call_req_1;
      call_stmt_1547_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueuePointers_call_group_2_gI: SplitGuardInterface generic map(name => "getQueuePointers_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      write_index_1547 <= data_out(63 downto 32);
      read_index_1547 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueuePointers_call_reqs(0),
          ackR => getQueuePointers_call_acks(0),
          dataR => getQueuePointers_call_data(35 downto 0),
          tagR => getQueuePointers_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueuePointers_return_acks(0), -- cross-over
          ackL => getQueuePointers_return_reqs(0), -- cross-over
          dataL => getQueuePointers_return_data(63 downto 0),
          tagL => getQueuePointers_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_1550_call 
    getQueueLength_call_group_3: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1550_call_req_0;
      call_stmt_1550_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1550_call_req_1;
      call_stmt_1550_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getQueueLength_call_group_3_gI: SplitGuardInterface generic map(name => "getQueueLength_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      Queue_Length_1550 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getQueueLength_call_reqs(0),
          ackR => getQueueLength_call_acks(0),
          dataR => getQueueLength_call_data(35 downto 0),
          tagR => getQueueLength_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getQueueLength_return_acks(0), -- cross-over
          ackL => getQueueLength_return_reqs(0), -- cross-over
          dataL => getQueueLength_return_data(31 downto 0),
          tagL => getQueueLength_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- shared call operator group (4) : call_stmt_1553_call 
    getTotalMessages_call_group_4: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1553_call_req_0;
      call_stmt_1553_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1553_call_req_1;
      call_stmt_1553_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getTotalMessages_call_group_4_gI: SplitGuardInterface generic map(name => "getTotalMessages_call_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      total_msgs_1553 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getTotalMessages_call_reqs(0),
          ackR => getTotalMessages_call_acks(0),
          dataR => getTotalMessages_call_data(35 downto 0),
          tagR => getTotalMessages_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getTotalMessages_return_acks(0), -- cross-over
          ackL => getTotalMessages_return_reqs(0), -- cross-over
          dataL => getTotalMessages_return_data(31 downto 0),
          tagL => getTotalMessages_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 4
    -- shared call operator group (5) : call_stmt_1584_call 
    setQueueElement_call_group_5: Block -- 
      signal data_in: std_logic_vector(99 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1584_call_req_0;
      call_stmt_1584_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1584_call_req_1;
      call_stmt_1584_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_full_1573(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      setQueueElement_call_group_5_gI: SplitGuardInterface generic map(name => "setQueueElement_call_group_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer & write_index_1547 & q_w_data_buffer;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 100,
        owidth => 100,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => setQueueElement_call_reqs(0),
          ackR => setQueueElement_call_acks(0),
          dataR => setQueueElement_call_data(99 downto 0),
          tagR => setQueueElement_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => setQueueElement_return_acks(0), -- cross-over
          ackL => setQueueElement_return_reqs(0), -- cross-over
          tagL => setQueueElement_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 5
    -- shared call operator group (6) : call_stmt_1589_call 
    setQueuePointers_call_group_6: Block -- 
      signal data_in: std_logic_vector(99 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1589_call_req_0;
      call_stmt_1589_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1589_call_req_1;
      call_stmt_1589_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_full_1573(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      setQueuePointers_call_group_6_gI: SplitGuardInterface generic map(name => "setQueuePointers_call_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer & next_wi_1568 & read_index_1547;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 100,
        owidth => 100,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => setQueuePointers_call_reqs(0),
          ackR => setQueuePointers_call_acks(0),
          dataR => setQueuePointers_call_data(99 downto 0),
          tagR => setQueuePointers_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => setQueuePointers_return_acks(0), -- cross-over
          ackL => setQueuePointers_return_reqs(0), -- cross-over
          tagL => setQueuePointers_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 6
    -- shared call operator group (7) : call_stmt_1596_call 
    updateTotalMessages_call_group_7: Block -- 
      signal data_in: std_logic_vector(67 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1596_call_req_0;
      call_stmt_1596_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1596_call_req_1;
      call_stmt_1596_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not q_full_1573(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      updateTotalMessages_call_group_7_gI: SplitGuardInterface generic map(name => "updateTotalMessages_call_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer & ADD_u32_u32_1595_wire;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 68,
        owidth => 68,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => updateTotalMessages_call_reqs(0),
          ackR => updateTotalMessages_call_acks(0),
          dataR => updateTotalMessages_call_data(67 downto 0),
          tagR => updateTotalMessages_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => updateTotalMessages_return_acks(0), -- cross-over
          ackL => updateTotalMessages_return_reqs(0), -- cross-over
          tagL => updateTotalMessages_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 7
    -- shared call operator group (8) : call_stmt_1600_call 
    releaseLock_call_group_8: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1600_call_req_0;
      call_stmt_1600_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1600_call_req_1;
      call_stmt_1600_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= lock_n_1535(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      releaseLock_call_group_8_gI: SplitGuardInterface generic map(name => "releaseLock_call_group_8_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= q_base_address_buffer;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 36,
        owidth => 36,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => releaseLock_call_reqs(0),
          ackR => releaseLock_call_acks(0),
          dataR => releaseLock_call_data(35 downto 0),
          tagR => releaseLock_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => releaseLock_return_acks(0), -- cross-over
          ackL => releaseLock_return_reqs(0), -- cross-over
          tagL => releaseLock_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 8
    -- 
  end Block; -- data_path
  -- 
end pushIntoQueue_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.nic_system_global_package.all;
entity releaseLock is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity releaseLock;
architecture releaseLock_arch of releaseLock is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  -- output port buffer signals
  signal releaseLock_CP_1310_start: Boolean;
  signal releaseLock_CP_1310_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1037_call_ack_0 : boolean;
  signal call_stmt_1155_call_ack_1 : boolean;
  signal call_stmt_1155_call_req_0 : boolean;
  signal call_stmt_1037_call_req_1 : boolean;
  signal call_stmt_1155_call_req_1 : boolean;
  signal call_stmt_1037_call_req_0 : boolean;
  signal call_stmt_1155_call_ack_0 : boolean;
  signal call_stmt_1037_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "releaseLock_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  releaseLock_CP_1310_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "releaseLock_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= releaseLock_CP_1310_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= releaseLock_CP_1310_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= releaseLock_CP_1310_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  releaseLock_CP_1310: Block -- control-path 
    signal releaseLock_CP_1310_elements: BooleanArray(4 downto 0);
    -- 
  begin -- 
    releaseLock_CP_1310_elements(0) <= releaseLock_CP_1310_start;
    releaseLock_CP_1310_symbol <= releaseLock_CP_1310_elements(4);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 assign_stmt_1025_to_call_stmt_1155/call_stmt_1037_Update/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_1025_to_call_stmt_1155/call_stmt_1037_update_start_
      -- CP-element group 0: 	 assign_stmt_1025_to_call_stmt_1155/call_stmt_1037_sample_start_
      -- CP-element group 0: 	 assign_stmt_1025_to_call_stmt_1155/call_stmt_1037_Update/ccr
      -- CP-element group 0: 	 assign_stmt_1025_to_call_stmt_1155/call_stmt_1155_update_start_
      -- CP-element group 0: 	 assign_stmt_1025_to_call_stmt_1155/$entry
      -- CP-element group 0: 	 assign_stmt_1025_to_call_stmt_1155/call_stmt_1155_Update/ccr
      -- CP-element group 0: 	 assign_stmt_1025_to_call_stmt_1155/call_stmt_1155_Update/$entry
      -- CP-element group 0: 	 assign_stmt_1025_to_call_stmt_1155/call_stmt_1037_Sample/crr
      -- CP-element group 0: 	 assign_stmt_1025_to_call_stmt_1155/call_stmt_1037_Sample/$entry
      -- 
    crr_1323_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1323_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => releaseLock_CP_1310_elements(0), ack => call_stmt_1037_call_req_0); -- 
    ccr_1328_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1328_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => releaseLock_CP_1310_elements(0), ack => call_stmt_1037_call_req_1); -- 
    ccr_1342_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1342_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => releaseLock_CP_1310_elements(0), ack => call_stmt_1155_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_1025_to_call_stmt_1155/call_stmt_1037_Sample/cra
      -- CP-element group 1: 	 assign_stmt_1025_to_call_stmt_1155/call_stmt_1037_sample_completed_
      -- CP-element group 1: 	 assign_stmt_1025_to_call_stmt_1155/call_stmt_1037_Sample/$exit
      -- 
    cra_1324_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1037_call_ack_0, ack => releaseLock_CP_1310_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 assign_stmt_1025_to_call_stmt_1155/call_stmt_1155_sample_start_
      -- CP-element group 2: 	 assign_stmt_1025_to_call_stmt_1155/call_stmt_1155_Sample/crr
      -- CP-element group 2: 	 assign_stmt_1025_to_call_stmt_1155/call_stmt_1155_Sample/$entry
      -- CP-element group 2: 	 assign_stmt_1025_to_call_stmt_1155/call_stmt_1037_Update/$exit
      -- CP-element group 2: 	 assign_stmt_1025_to_call_stmt_1155/call_stmt_1037_update_completed_
      -- CP-element group 2: 	 assign_stmt_1025_to_call_stmt_1155/call_stmt_1037_Update/cca
      -- 
    cca_1329_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1037_call_ack_1, ack => releaseLock_CP_1310_elements(2)); -- 
    crr_1337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => releaseLock_CP_1310_elements(2), ack => call_stmt_1155_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 assign_stmt_1025_to_call_stmt_1155/call_stmt_1155_sample_completed_
      -- CP-element group 3: 	 assign_stmt_1025_to_call_stmt_1155/call_stmt_1155_Sample/$exit
      -- CP-element group 3: 	 assign_stmt_1025_to_call_stmt_1155/call_stmt_1155_Sample/cra
      -- 
    cra_1338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1155_call_ack_0, ack => releaseLock_CP_1310_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 $exit
      -- CP-element group 4: 	 assign_stmt_1025_to_call_stmt_1155/call_stmt_1155_Update/cca
      -- CP-element group 4: 	 assign_stmt_1025_to_call_stmt_1155/call_stmt_1155_update_completed_
      -- CP-element group 4: 	 assign_stmt_1025_to_call_stmt_1155/call_stmt_1155_Update/$exit
      -- CP-element group 4: 	 assign_stmt_1025_to_call_stmt_1155/$exit
      -- 
    cca_1343_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1155_call_ack_1, ack => releaseLock_CP_1310_elements(4)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u1_u2_1099_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_1112_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_1126_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_1139_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u2_u4_1113_wire : std_logic_vector(3 downto 0);
    signal CONCAT_u2_u4_1140_wire : std_logic_vector(3 downto 0);
    signal CONCAT_u4_u36_1151_wire : std_logic_vector(35 downto 0);
    signal MUX_1092_wire : std_logic_vector(0 downto 0);
    signal MUX_1098_wire : std_logic_vector(0 downto 0);
    signal MUX_1105_wire : std_logic_vector(0 downto 0);
    signal MUX_1111_wire : std_logic_vector(0 downto 0);
    signal MUX_1119_wire : std_logic_vector(0 downto 0);
    signal MUX_1125_wire : std_logic_vector(0 downto 0);
    signal MUX_1132_wire : std_logic_vector(0 downto 0);
    signal MUX_1138_wire : std_logic_vector(0 downto 0);
    signal NOT_u8_u8_1032_wire_constant : std_logic_vector(7 downto 0);
    signal ignore_1155 : std_logic_vector(63 downto 0);
    signal konst_1048_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1053_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1058_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1063_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1068_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1073_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1078_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1083_wire_constant : std_logic_vector(2 downto 0);
    signal lock_addr_32_1041 : std_logic_vector(31 downto 0);
    signal lock_address_pointer_1025 : std_logic_vector(35 downto 0);
    signal msg_size_plus_lock_1037 : std_logic_vector(63 downto 0);
    signal new_bmask_1142 : std_logic_vector(7 downto 0);
    signal s0_1050 : std_logic_vector(0 downto 0);
    signal s1_1055 : std_logic_vector(0 downto 0);
    signal s2_1060 : std_logic_vector(0 downto 0);
    signal s3_1065 : std_logic_vector(0 downto 0);
    signal s4_1070 : std_logic_vector(0 downto 0);
    signal s5_1075 : std_logic_vector(0 downto 0);
    signal s6_1080 : std_logic_vector(0 downto 0);
    signal s7_1085 : std_logic_vector(0 downto 0);
    signal sel_1045 : std_logic_vector(2 downto 0);
    signal type_cast_1023_wire_constant : std_logic_vector(35 downto 0);
    signal type_cast_1027_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1029_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1035_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_1089_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1091_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1095_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1097_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1102_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1104_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1108_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1110_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1116_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1118_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1122_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1124_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1129_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1131_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1135_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1137_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1144_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1146_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1149_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_1153_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    NOT_u8_u8_1032_wire_constant <= "11111111";
    konst_1048_wire_constant <= "000";
    konst_1053_wire_constant <= "001";
    konst_1058_wire_constant <= "010";
    konst_1063_wire_constant <= "011";
    konst_1068_wire_constant <= "100";
    konst_1073_wire_constant <= "101";
    konst_1078_wire_constant <= "110";
    konst_1083_wire_constant <= "111";
    type_cast_1023_wire_constant <= "000000000000000000000000000000010000";
    type_cast_1027_wire_constant <= "1";
    type_cast_1029_wire_constant <= "1";
    type_cast_1035_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_1089_wire_constant <= "1";
    type_cast_1091_wire_constant <= "0";
    type_cast_1095_wire_constant <= "1";
    type_cast_1097_wire_constant <= "0";
    type_cast_1102_wire_constant <= "1";
    type_cast_1104_wire_constant <= "0";
    type_cast_1108_wire_constant <= "1";
    type_cast_1110_wire_constant <= "0";
    type_cast_1116_wire_constant <= "1";
    type_cast_1118_wire_constant <= "0";
    type_cast_1122_wire_constant <= "1";
    type_cast_1124_wire_constant <= "0";
    type_cast_1129_wire_constant <= "1";
    type_cast_1131_wire_constant <= "0";
    type_cast_1135_wire_constant <= "1";
    type_cast_1137_wire_constant <= "0";
    type_cast_1144_wire_constant <= "0";
    type_cast_1146_wire_constant <= "0";
    type_cast_1149_wire_constant <= "0000";
    type_cast_1153_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    -- flow-through select operator MUX_1092_inst
    MUX_1092_wire <= type_cast_1089_wire_constant when (s0_1050(0) /=  '0') else type_cast_1091_wire_constant;
    -- flow-through select operator MUX_1098_inst
    MUX_1098_wire <= type_cast_1095_wire_constant when (s1_1055(0) /=  '0') else type_cast_1097_wire_constant;
    -- flow-through select operator MUX_1105_inst
    MUX_1105_wire <= type_cast_1102_wire_constant when (s2_1060(0) /=  '0') else type_cast_1104_wire_constant;
    -- flow-through select operator MUX_1111_inst
    MUX_1111_wire <= type_cast_1108_wire_constant when (s3_1065(0) /=  '0') else type_cast_1110_wire_constant;
    -- flow-through select operator MUX_1119_inst
    MUX_1119_wire <= type_cast_1116_wire_constant when (s4_1070(0) /=  '0') else type_cast_1118_wire_constant;
    -- flow-through select operator MUX_1125_inst
    MUX_1125_wire <= type_cast_1122_wire_constant when (s5_1075(0) /=  '0') else type_cast_1124_wire_constant;
    -- flow-through select operator MUX_1132_inst
    MUX_1132_wire <= type_cast_1129_wire_constant when (s6_1080(0) /=  '0') else type_cast_1131_wire_constant;
    -- flow-through select operator MUX_1138_inst
    MUX_1138_wire <= type_cast_1135_wire_constant when (s7_1085(0) /=  '0') else type_cast_1137_wire_constant;
    -- flow-through slice operator slice_1040_inst
    lock_addr_32_1041 <= msg_size_plus_lock_1037(31 downto 0);
    -- flow-through slice operator slice_1044_inst
    sel_1045 <= lock_addr_32_1041(2 downto 0);
    -- binary operator ADD_u36_u36_1024_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, type_cast_1023_wire_constant, tmp_var);
      lock_address_pointer_1025 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_1099_inst
    process(MUX_1092_wire, MUX_1098_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_1092_wire, MUX_1098_wire, tmp_var);
      CONCAT_u1_u2_1099_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_1112_inst
    process(MUX_1105_wire, MUX_1111_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_1105_wire, MUX_1111_wire, tmp_var);
      CONCAT_u1_u2_1112_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_1126_inst
    process(MUX_1119_wire, MUX_1125_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_1119_wire, MUX_1125_wire, tmp_var);
      CONCAT_u1_u2_1126_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_1139_inst
    process(MUX_1132_wire, MUX_1138_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_1132_wire, MUX_1138_wire, tmp_var);
      CONCAT_u1_u2_1139_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u2_u4_1113_inst
    process(CONCAT_u1_u2_1099_wire, CONCAT_u1_u2_1112_wire) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_1099_wire, CONCAT_u1_u2_1112_wire, tmp_var);
      CONCAT_u2_u4_1113_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u2_u4_1140_inst
    process(CONCAT_u1_u2_1126_wire, CONCAT_u1_u2_1139_wire) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_1126_wire, CONCAT_u1_u2_1139_wire, tmp_var);
      CONCAT_u2_u4_1140_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u4_u36_1151_inst
    process(type_cast_1149_wire_constant, lock_addr_32_1041) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1149_wire_constant, lock_addr_32_1041, tmp_var);
      CONCAT_u4_u36_1151_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u4_u8_1141_inst
    process(CONCAT_u2_u4_1113_wire, CONCAT_u2_u4_1140_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u2_u4_1113_wire, CONCAT_u2_u4_1140_wire, tmp_var);
      new_bmask_1142 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1049_inst
    process(sel_1045) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_1045, konst_1048_wire_constant, tmp_var);
      s0_1050 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1054_inst
    process(sel_1045) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_1045, konst_1053_wire_constant, tmp_var);
      s1_1055 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1059_inst
    process(sel_1045) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_1045, konst_1058_wire_constant, tmp_var);
      s2_1060 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1064_inst
    process(sel_1045) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_1045, konst_1063_wire_constant, tmp_var);
      s3_1065 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1069_inst
    process(sel_1045) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_1045, konst_1068_wire_constant, tmp_var);
      s4_1070 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1074_inst
    process(sel_1045) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_1045, konst_1073_wire_constant, tmp_var);
      s5_1075 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1079_inst
    process(sel_1045) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_1045, konst_1078_wire_constant, tmp_var);
      s6_1080 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1084_inst
    process(sel_1045) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(sel_1045, konst_1083_wire_constant, tmp_var);
      s7_1085 <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_1037_call call_stmt_1155_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(219 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_1037_call_req_0;
      reqL_unguarded(0) <= call_stmt_1155_call_req_0;
      call_stmt_1037_call_ack_0 <= ackL_unguarded(1);
      call_stmt_1155_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_1037_call_req_1;
      reqR_unguarded(0) <= call_stmt_1155_call_req_1;
      call_stmt_1037_call_ack_1 <= ackR_unguarded(1);
      call_stmt_1155_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      accessMemory_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1027_wire_constant & type_cast_1029_wire_constant & NOT_u8_u8_1032_wire_constant & lock_address_pointer_1025 & type_cast_1035_wire_constant & type_cast_1144_wire_constant & type_cast_1146_wire_constant & new_bmask_1142 & CONCAT_u4_u36_1151_wire & type_cast_1153_wire_constant;
      msg_size_plus_lock_1037 <= data_out(127 downto 64);
      ignore_1155 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 220,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end releaseLock_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.nic_system_global_package.all;
entity setQueueElement is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    write_index : in  std_logic_vector(31 downto 0);
    q_w_data : in  std_logic_vector(31 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity setQueueElement;
architecture setQueueElement_arch of setQueueElement is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 100)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  signal write_index_buffer :  std_logic_vector(31 downto 0);
  signal write_index_update_enable: Boolean;
  signal q_w_data_buffer :  std_logic_vector(31 downto 0);
  signal q_w_data_update_enable: Boolean;
  -- output port buffer signals
  signal setQueueElement_CP_1928_start: Boolean;
  signal setQueueElement_CP_1928_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1505_call_ack_1 : boolean;
  signal call_stmt_1505_call_req_0 : boolean;
  signal call_stmt_1505_call_req_1 : boolean;
  signal call_stmt_1505_call_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "setQueueElement_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 100) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(67 downto 36) <= write_index;
  write_index_buffer <= in_buffer_data_out(67 downto 36);
  in_buffer_data_in(99 downto 68) <= q_w_data;
  q_w_data_buffer <= in_buffer_data_out(99 downto 68);
  in_buffer_data_in(tag_length + 99 downto 100) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 99 downto 100);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  setQueueElement_CP_1928_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "setQueueElement_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= setQueueElement_CP_1928_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= setQueueElement_CP_1928_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= setQueueElement_CP_1928_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  setQueueElement_CP_1928: Block -- control-path 
    signal setQueueElement_CP_1928_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    setQueueElement_CP_1928_elements(0) <= setQueueElement_CP_1928_start;
    setQueueElement_CP_1928_symbol <= setQueueElement_CP_1928_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 assign_stmt_1449_to_call_stmt_1505/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_1449_to_call_stmt_1505/call_stmt_1505_Update/$entry
      -- CP-element group 0: 	 assign_stmt_1449_to_call_stmt_1505/call_stmt_1505_Sample/crr
      -- CP-element group 0: 	 assign_stmt_1449_to_call_stmt_1505/call_stmt_1505_sample_start_
      -- CP-element group 0: 	 assign_stmt_1449_to_call_stmt_1505/call_stmt_1505_Update/ccr
      -- CP-element group 0: 	 assign_stmt_1449_to_call_stmt_1505/call_stmt_1505_update_start_
      -- CP-element group 0: 	 assign_stmt_1449_to_call_stmt_1505/call_stmt_1505_Sample/$entry
      -- 
    crr_1941_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1941_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueueElement_CP_1928_elements(0), ack => call_stmt_1505_call_req_0); -- 
    ccr_1946_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1946_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueueElement_CP_1928_elements(0), ack => call_stmt_1505_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_1449_to_call_stmt_1505/call_stmt_1505_sample_completed_
      -- CP-element group 1: 	 assign_stmt_1449_to_call_stmt_1505/call_stmt_1505_Sample/cra
      -- CP-element group 1: 	 assign_stmt_1449_to_call_stmt_1505/call_stmt_1505_Sample/$exit
      -- 
    cra_1942_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1505_call_ack_0, ack => setQueueElement_CP_1928_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 assign_stmt_1449_to_call_stmt_1505/call_stmt_1505_Update/cca
      -- CP-element group 2: 	 assign_stmt_1449_to_call_stmt_1505/$exit
      -- CP-element group 2: 	 assign_stmt_1449_to_call_stmt_1505/call_stmt_1505_Update/$exit
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_1449_to_call_stmt_1505/call_stmt_1505_update_completed_
      -- 
    cca_1947_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1505_call_ack_1, ack => setQueueElement_CP_1928_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal BITSEL_u32_u1_1463_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_1481_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u31_u34_1456_wire : std_logic_vector(33 downto 0);
    signal CONCAT_u32_u64_1485_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_1489_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u4_u8_1469_wire_constant : std_logic_vector(7 downto 0);
    signal CONCAT_u4_u8_1475_wire_constant : std_logic_vector(7 downto 0);
    signal bmask_1477 : std_logic_vector(7 downto 0);
    signal buffer_address_1449 : std_logic_vector(35 downto 0);
    signal element_pair_address_1459 : std_logic_vector(35 downto 0);
    signal ignore_1505 : std_logic_vector(63 downto 0);
    signal konst_1462_wire_constant : std_logic_vector(31 downto 0);
    signal konst_1480_wire_constant : std_logic_vector(31 downto 0);
    signal slice_1453_wire : std_logic_vector(30 downto 0);
    signal type_cast_1447_wire_constant : std_logic_vector(35 downto 0);
    signal type_cast_1455_wire_constant : std_logic_vector(2 downto 0);
    signal type_cast_1457_wire : std_logic_vector(35 downto 0);
    signal type_cast_1483_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1488_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_1498_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1500_wire_constant : std_logic_vector(0 downto 0);
    signal wval_1491 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    CONCAT_u4_u8_1469_wire_constant <= "00001111";
    CONCAT_u4_u8_1475_wire_constant <= "11110000";
    konst_1462_wire_constant <= "00000000000000000000000000000000";
    konst_1480_wire_constant <= "00000000000000000000000000000000";
    type_cast_1447_wire_constant <= "000000000000000000000000000000100000";
    type_cast_1455_wire_constant <= "000";
    type_cast_1483_wire_constant <= "00000000000000000000000000000000";
    type_cast_1488_wire_constant <= "00000000000000000000000000000000";
    type_cast_1498_wire_constant <= "0";
    type_cast_1500_wire_constant <= "0";
    -- flow-through select operator MUX_1476_inst
    bmask_1477 <= CONCAT_u4_u8_1469_wire_constant when (BITSEL_u32_u1_1463_wire(0) /=  '0') else CONCAT_u4_u8_1475_wire_constant;
    -- flow-through select operator MUX_1490_inst
    wval_1491 <= CONCAT_u32_u64_1485_wire when (BITSEL_u32_u1_1481_wire(0) /=  '0') else CONCAT_u32_u64_1489_wire;
    -- flow-through slice operator slice_1453_inst
    slice_1453_wire <= write_index_buffer(31 downto 1);
    -- interlock type_cast_1457_inst
    process(CONCAT_u31_u34_1456_wire) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 33 downto 0) := CONCAT_u31_u34_1456_wire(33 downto 0);
      type_cast_1457_wire <= tmp_var; -- 
    end process;
    -- binary operator ADD_u36_u36_1448_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, type_cast_1447_wire_constant, tmp_var);
      buffer_address_1449 <= tmp_var; --
    end process;
    -- binary operator ADD_u36_u36_1458_inst
    process(buffer_address_1449, type_cast_1457_wire) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(buffer_address_1449, type_cast_1457_wire, tmp_var);
      element_pair_address_1459 <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_1463_inst
    process(write_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(write_index_buffer, konst_1462_wire_constant, tmp_var);
      BITSEL_u32_u1_1463_wire <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_1481_inst
    process(write_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(write_index_buffer, konst_1480_wire_constant, tmp_var);
      BITSEL_u32_u1_1481_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u31_u34_1456_inst
    process(slice_1453_wire) -- 
      variable tmp_var : std_logic_vector(33 downto 0); -- 
    begin -- 
      ApConcat_proc(slice_1453_wire, type_cast_1455_wire_constant, tmp_var);
      CONCAT_u31_u34_1456_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u32_u64_1485_inst
    process(type_cast_1483_wire_constant, q_w_data_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_1483_wire_constant, q_w_data_buffer, tmp_var);
      CONCAT_u32_u64_1485_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u32_u64_1489_inst
    process(q_w_data_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(q_w_data_buffer, type_cast_1488_wire_constant, tmp_var);
      CONCAT_u32_u64_1489_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_1505_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1505_call_req_0;
      call_stmt_1505_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1505_call_req_1;
      call_stmt_1505_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1498_wire_constant & type_cast_1500_wire_constant & bmask_1477 & element_pair_address_1459 & wval_1491;
      ignore_1505 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end setQueueElement_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.nic_system_global_package.all;
entity setQueuePointers is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    wp : in  std_logic_vector(31 downto 0);
    rp : in  std_logic_vector(31 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity setQueuePointers;
architecture setQueuePointers_arch of setQueuePointers is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 100)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  signal wp_buffer :  std_logic_vector(31 downto 0);
  signal wp_update_enable: Boolean;
  signal rp_buffer :  std_logic_vector(31 downto 0);
  signal rp_update_enable: Boolean;
  -- output port buffer signals
  signal setQueuePointers_CP_1256_start: Boolean;
  signal setQueuePointers_CP_1256_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_978_call_req_1 : boolean;
  signal call_stmt_978_call_ack_1 : boolean;
  signal call_stmt_996_call_ack_1 : boolean;
  signal call_stmt_996_call_req_1 : boolean;
  signal call_stmt_978_call_req_0 : boolean;
  signal call_stmt_978_call_ack_0 : boolean;
  signal call_stmt_996_call_req_0 : boolean;
  signal call_stmt_996_call_ack_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "setQueuePointers_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 100) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(67 downto 36) <= wp;
  wp_buffer <= in_buffer_data_out(67 downto 36);
  in_buffer_data_in(99 downto 68) <= rp;
  rp_buffer <= in_buffer_data_out(99 downto 68);
  in_buffer_data_in(tag_length + 99 downto 100) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 99 downto 100);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  setQueuePointers_CP_1256_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "setQueuePointers_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= setQueuePointers_CP_1256_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= setQueuePointers_CP_1256_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= setQueuePointers_CP_1256_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  setQueuePointers_CP_1256: Block -- control-path 
    signal setQueuePointers_CP_1256_elements: BooleanArray(4 downto 0);
    -- 
  begin -- 
    setQueuePointers_CP_1256_elements(0) <= setQueuePointers_CP_1256_start;
    setQueuePointers_CP_1256_symbol <= setQueuePointers_CP_1256_elements(4);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	4 
    -- CP-element group 0:  members (11) 
      -- CP-element group 0: 	 call_stmt_978_to_call_stmt_996/$entry
      -- CP-element group 0: 	 call_stmt_978_to_call_stmt_996/call_stmt_978_Update/ccr
      -- CP-element group 0: 	 call_stmt_978_to_call_stmt_996/call_stmt_996_Update/$entry
      -- CP-element group 0: 	 call_stmt_978_to_call_stmt_996/call_stmt_978_Update/$entry
      -- CP-element group 0: 	 call_stmt_978_to_call_stmt_996/call_stmt_996_Update/ccr
      -- CP-element group 0: 	 call_stmt_978_to_call_stmt_996/call_stmt_978_Sample/crr
      -- CP-element group 0: 	 call_stmt_978_to_call_stmt_996/call_stmt_978_update_start_
      -- CP-element group 0: 	 call_stmt_978_to_call_stmt_996/call_stmt_978_sample_start_
      -- CP-element group 0: 	 call_stmt_978_to_call_stmt_996/call_stmt_978_Sample/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_978_to_call_stmt_996/call_stmt_996_update_start_
      -- 
    crr_1269_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1269_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueuePointers_CP_1256_elements(0), ack => call_stmt_978_call_req_0); -- 
    ccr_1274_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1274_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueuePointers_CP_1256_elements(0), ack => call_stmt_978_call_req_1); -- 
    ccr_1288_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1288_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueuePointers_CP_1256_elements(0), ack => call_stmt_996_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_978_to_call_stmt_996/call_stmt_978_sample_completed_
      -- CP-element group 1: 	 call_stmt_978_to_call_stmt_996/call_stmt_978_Sample/$exit
      -- CP-element group 1: 	 call_stmt_978_to_call_stmt_996/call_stmt_978_Sample/cra
      -- 
    cra_1270_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_978_call_ack_0, ack => setQueuePointers_CP_1256_elements(1)); -- 
    -- CP-element group 2:  transition  input  output  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	3 
    -- CP-element group 2:  members (6) 
      -- CP-element group 2: 	 call_stmt_978_to_call_stmt_996/call_stmt_978_Update/cca
      -- CP-element group 2: 	 call_stmt_978_to_call_stmt_996/call_stmt_996_sample_start_
      -- CP-element group 2: 	 call_stmt_978_to_call_stmt_996/call_stmt_978_Update/$exit
      -- CP-element group 2: 	 call_stmt_978_to_call_stmt_996/call_stmt_978_update_completed_
      -- CP-element group 2: 	 call_stmt_978_to_call_stmt_996/call_stmt_996_Sample/crr
      -- CP-element group 2: 	 call_stmt_978_to_call_stmt_996/call_stmt_996_Sample/$entry
      -- 
    cca_1275_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_978_call_ack_1, ack => setQueuePointers_CP_1256_elements(2)); -- 
    crr_1283_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1283_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => setQueuePointers_CP_1256_elements(2), ack => call_stmt_996_call_req_0); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	2 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 call_stmt_978_to_call_stmt_996/call_stmt_996_sample_completed_
      -- CP-element group 3: 	 call_stmt_978_to_call_stmt_996/call_stmt_996_Sample/cra
      -- CP-element group 3: 	 call_stmt_978_to_call_stmt_996/call_stmt_996_Sample/$exit
      -- 
    cra_1284_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_996_call_ack_0, ack => setQueuePointers_CP_1256_elements(3)); -- 
    -- CP-element group 4:  transition  input  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	0 
    -- CP-element group 4: successors 
    -- CP-element group 4:  members (5) 
      -- CP-element group 4: 	 $exit
      -- CP-element group 4: 	 call_stmt_978_to_call_stmt_996/call_stmt_996_Update/cca
      -- CP-element group 4: 	 call_stmt_978_to_call_stmt_996/call_stmt_996_Update/$exit
      -- CP-element group 4: 	 call_stmt_978_to_call_stmt_996/$exit
      -- CP-element group 4: 	 call_stmt_978_to_call_stmt_996/call_stmt_996_update_completed_
      -- 
    cca_1289_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 4_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_996_call_ack_1, ack => setQueuePointers_CP_1256_elements(4)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u36_u36_991_wire : std_logic_vector(35 downto 0);
    signal CONCAT_u32_u64_976_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u32_u64_994_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u4_u8_972_wire_constant : std_logic_vector(7 downto 0);
    signal CONCAT_u4_u8_988_wire_constant : std_logic_vector(7 downto 0);
    signal ignore_1_996 : std_logic_vector(63 downto 0);
    signal ignore_978 : std_logic_vector(63 downto 0);
    signal konst_990_wire_constant : std_logic_vector(35 downto 0);
    signal type_cast_964_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_966_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_980_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_982_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    CONCAT_u4_u8_972_wire_constant <= "00001111";
    CONCAT_u4_u8_988_wire_constant <= "11110000";
    konst_990_wire_constant <= "000000000000000000000000000000001000";
    type_cast_964_wire_constant <= "0";
    type_cast_966_wire_constant <= "0";
    type_cast_980_wire_constant <= "0";
    type_cast_982_wire_constant <= "0";
    -- binary operator ADD_u36_u36_991_inst
    process(q_base_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(q_base_address_buffer, konst_990_wire_constant, tmp_var);
      ADD_u36_u36_991_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u32_u64_976_inst
    process(rp_buffer, rp_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(rp_buffer, rp_buffer, tmp_var);
      CONCAT_u32_u64_976_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u32_u64_994_inst
    process(wp_buffer, wp_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(wp_buffer, wp_buffer, tmp_var);
      CONCAT_u32_u64_994_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_996_call call_stmt_978_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(219 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_996_call_req_0;
      reqL_unguarded(0) <= call_stmt_978_call_req_0;
      call_stmt_996_call_ack_0 <= ackL_unguarded(1);
      call_stmt_978_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_996_call_req_1;
      reqR_unguarded(0) <= call_stmt_978_call_req_1;
      call_stmt_996_call_ack_1 <= ackR_unguarded(1);
      call_stmt_978_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      accessMemory_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_980_wire_constant & type_cast_982_wire_constant & CONCAT_u4_u8_988_wire_constant & ADD_u36_u36_991_wire & CONCAT_u32_u64_994_wire & type_cast_964_wire_constant & type_cast_966_wire_constant & CONCAT_u4_u8_972_wire_constant & q_base_address_buffer & CONCAT_u32_u64_976_wire;
      ignore_1_996 <= data_out(127 downto 64);
      ignore_978 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 220,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end setQueuePointers_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.nic_system_global_package.all;
entity transmitEngineDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    CONTROL_REGISTER : in std_logic_vector(31 downto 0);
    FREE_Q : in std_logic_vector(35 downto 0);
    LAST_READ_TX_QUEUE_INDEX : in std_logic_vector(5 downto 0);
    NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
    LAST_READ_TX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(1 downto 0);
    LAST_READ_TX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(1 downto 0);
    LAST_READ_TX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(11 downto 0);
    AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_call_data : out  std_logic_vector(42 downto 0);
    AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
    AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_return_data : in   std_logic_vector(31 downto 0);
    AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
    pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
    pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
    pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
    pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_call_reqs : out  std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_call_acks : in   std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_call_data : out  std_logic_vector(5 downto 0);
    getTxPacketPointerFromServer_call_tag  :  out  std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_return_reqs : out  std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_return_acks : in   std_logic_vector(0 downto 0);
    getTxPacketPointerFromServer_return_data : in   std_logic_vector(32 downto 0);
    getTxPacketPointerFromServer_return_tag :  in   std_logic_vector(0 downto 0);
    transmitPacket_call_reqs : out  std_logic_vector(0 downto 0);
    transmitPacket_call_acks : in   std_logic_vector(0 downto 0);
    transmitPacket_call_data : out  std_logic_vector(31 downto 0);
    transmitPacket_call_tag  :  out  std_logic_vector(0 downto 0);
    transmitPacket_return_reqs : out  std_logic_vector(0 downto 0);
    transmitPacket_return_acks : in   std_logic_vector(0 downto 0);
    transmitPacket_return_data : in   std_logic_vector(0 downto 0);
    transmitPacket_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity transmitEngineDaemon;
architecture transmitEngineDaemon_arch of transmitEngineDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal transmitEngineDaemon_CP_36381_start: Boolean;
  signal transmitEngineDaemon_CP_36381_symbol: Boolean;
  -- volatile/operator module components. 
  component AccessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      register_index : in  std_logic_vector(5 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component pushIntoQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_call_acks : in   std_logic_vector(0 downto 0);
      releaseLock_call_data : out  std_logic_vector(35 downto 0);
      releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_return_acks : in   std_logic_vector(0 downto 0);
      releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_call_acks : in   std_logic_vector(0 downto 0);
      acquireLock_call_data : out  std_logic_vector(35 downto 0);
      acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_return_acks : in   std_logic_vector(0 downto 0);
      acquireLock_return_data : in   std_logic_vector(0 downto 0);
      acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      updateTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_data : out  std_logic_vector(67 downto 0);
      updateTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_call_data : out  std_logic_vector(35 downto 0);
      getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
      getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_call_data : out  std_logic_vector(35 downto 0);
      getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_return_data : in   std_logic_vector(31 downto 0);
      getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_call_data : out  std_logic_vector(99 downto 0);
      setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getTxPacketPointerFromServer is -- 
    generic (tag_length : integer); 
    port ( -- 
      queue_index : in  std_logic_vector(5 downto 0);
      pkt_pointer : out  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_call_data : out  std_logic_vector(36 downto 0);
      popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_return_data : in   std_logic_vector(32 downto 0);
      popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component transmitPacket is -- 
    generic (tag_length : integer); 
    port ( -- 
      packet_pointer : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_req : out  std_logic_vector(1 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_ack : in   std_logic_vector(1 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_data : out  std_logic_vector(145 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(1 downto 0);
      accessMemory_call_acks : in   std_logic_vector(1 downto 0);
      accessMemory_call_data : out  std_logic_vector(219 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(5 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(1 downto 0);
      accessMemory_return_acks : in   std_logic_vector(1 downto 0);
      accessMemory_return_data : in   std_logic_vector(127 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(5 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_18387_call_req_1 : boolean;
  signal ADD_u32_u32_18391_inst_req_1 : boolean;
  signal call_stmt_18371_call_req_1 : boolean;
  signal do_while_stmt_18315_branch_ack_1 : boolean;
  signal call_stmt_18371_call_ack_1 : boolean;
  signal W_pkt_pointer_17554_delayed_4_0_18362_inst_req_0 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_18404_inst_req_1 : boolean;
  signal call_stmt_18387_call_ack_1 : boolean;
  signal ADD_u32_u32_18391_inst_ack_1 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_18404_inst_ack_1 : boolean;
  signal ADD_u32_u32_18391_inst_ack_0 : boolean;
  signal W_pkt_pointer_17554_delayed_4_0_18362_inst_ack_0 : boolean;
  signal NOT_u1_u1_18352_inst_ack_0 : boolean;
  signal NOT_u1_u1_18352_inst_req_1 : boolean;
  signal NOT_u1_u1_18352_inst_req_0 : boolean;
  signal W_count_17575_delayed_14_0_18393_inst_req_0 : boolean;
  signal ADD_u32_u32_18391_inst_req_0 : boolean;
  signal NOT_u1_u1_18352_inst_ack_1 : boolean;
  signal W_count_17575_delayed_14_0_18393_inst_ack_0 : boolean;
  signal do_while_stmt_18315_branch_ack_0 : boolean;
  signal W_count_17575_delayed_14_0_18393_inst_req_1 : boolean;
  signal call_stmt_18387_call_ack_0 : boolean;
  signal call_stmt_18387_call_req_0 : boolean;
  signal call_stmt_18371_call_ack_0 : boolean;
  signal call_stmt_18371_call_req_0 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_18404_inst_ack_0 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_18404_inst_req_0 : boolean;
  signal W_count_17575_delayed_14_0_18393_inst_ack_1 : boolean;
  signal W_count_17567_delayed_14_0_18375_inst_ack_1 : boolean;
  signal W_count_17567_delayed_14_0_18375_inst_req_1 : boolean;
  signal W_count_17567_delayed_14_0_18375_inst_ack_0 : boolean;
  signal W_pkt_pointer_17554_delayed_4_0_18362_inst_ack_1 : boolean;
  signal W_pkt_pointer_17554_delayed_4_0_18362_inst_req_1 : boolean;
  signal W_count_17567_delayed_14_0_18375_inst_req_0 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_18302_inst_req_0 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_18302_inst_ack_0 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_18302_inst_req_1 : boolean;
  signal WPIPE_LAST_READ_TX_QUEUE_INDEX_18302_inst_ack_1 : boolean;
  signal if_stmt_18307_branch_req_0 : boolean;
  signal if_stmt_18307_branch_ack_1 : boolean;
  signal if_stmt_18307_branch_ack_0 : boolean;
  signal do_while_stmt_18315_branch_req_0 : boolean;
  signal AND_u6_u6_18326_inst_req_0 : boolean;
  signal AND_u6_u6_18326_inst_ack_0 : boolean;
  signal AND_u6_u6_18326_inst_req_1 : boolean;
  signal AND_u6_u6_18326_inst_ack_1 : boolean;
  signal phi_stmt_18327_req_1 : boolean;
  signal phi_stmt_18327_req_0 : boolean;
  signal phi_stmt_18327_ack_0 : boolean;
  signal ncount_18401_18331_buf_req_0 : boolean;
  signal ncount_18401_18331_buf_ack_0 : boolean;
  signal ncount_18401_18331_buf_req_1 : boolean;
  signal ncount_18401_18331_buf_ack_1 : boolean;
  signal call_stmt_18338_call_req_0 : boolean;
  signal call_stmt_18338_call_ack_0 : boolean;
  signal call_stmt_18338_call_req_1 : boolean;
  signal call_stmt_18338_call_ack_1 : boolean;
  signal call_stmt_18342_call_req_0 : boolean;
  signal call_stmt_18342_call_ack_0 : boolean;
  signal call_stmt_18342_call_req_1 : boolean;
  signal call_stmt_18342_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "transmitEngineDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  transmitEngineDaemon_CP_36381_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "transmitEngineDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= transmitEngineDaemon_CP_36381_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= transmitEngineDaemon_CP_36381_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= transmitEngineDaemon_CP_36381_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  transmitEngineDaemon_CP_36381: Block -- control-path 
    signal transmitEngineDaemon_CP_36381_elements: BooleanArray(86 downto 0);
    -- 
  begin -- 
    transmitEngineDaemon_CP_36381_elements(0) <= transmitEngineDaemon_CP_36381_start;
    transmitEngineDaemon_CP_36381_symbol <= transmitEngineDaemon_CP_36381_elements(3);
    -- CP-element group 0:  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_18304/$entry
      -- CP-element group 0: 	 assign_stmt_18304/WPIPE_LAST_READ_TX_QUEUE_INDEX_18302_sample_start_
      -- CP-element group 0: 	 assign_stmt_18304/WPIPE_LAST_READ_TX_QUEUE_INDEX_18302_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_18304/WPIPE_LAST_READ_TX_QUEUE_INDEX_18302_Sample/req
      -- 
    req_36394_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_36394_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_36381_elements(0), ack => WPIPE_LAST_READ_TX_QUEUE_INDEX_18302_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_18304/WPIPE_LAST_READ_TX_QUEUE_INDEX_18302_sample_completed_
      -- CP-element group 1: 	 assign_stmt_18304/WPIPE_LAST_READ_TX_QUEUE_INDEX_18302_update_start_
      -- CP-element group 1: 	 assign_stmt_18304/WPIPE_LAST_READ_TX_QUEUE_INDEX_18302_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_18304/WPIPE_LAST_READ_TX_QUEUE_INDEX_18302_Sample/ack
      -- CP-element group 1: 	 assign_stmt_18304/WPIPE_LAST_READ_TX_QUEUE_INDEX_18302_Update/$entry
      -- CP-element group 1: 	 assign_stmt_18304/WPIPE_LAST_READ_TX_QUEUE_INDEX_18302_Update/req
      -- 
    ack_36395_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_READ_TX_QUEUE_INDEX_18302_inst_ack_0, ack => transmitEngineDaemon_CP_36381_elements(1)); -- 
    req_36399_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_36399_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_36381_elements(1), ack => WPIPE_LAST_READ_TX_QUEUE_INDEX_18302_inst_req_1); -- 
    -- CP-element group 2:  branch  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	86 
    -- CP-element group 2:  members (10) 
      -- CP-element group 2: 	 branch_block_stmt_18305/merge_stmt_18306_dead_link/$entry
      -- CP-element group 2: 	 branch_block_stmt_18305/merge_stmt_18306__entry___PhiReq/$exit
      -- CP-element group 2: 	 branch_block_stmt_18305/merge_stmt_18306__entry___PhiReq/$entry
      -- CP-element group 2: 	 assign_stmt_18304/$exit
      -- CP-element group 2: 	 assign_stmt_18304/WPIPE_LAST_READ_TX_QUEUE_INDEX_18302_update_completed_
      -- CP-element group 2: 	 assign_stmt_18304/WPIPE_LAST_READ_TX_QUEUE_INDEX_18302_Update/$exit
      -- CP-element group 2: 	 assign_stmt_18304/WPIPE_LAST_READ_TX_QUEUE_INDEX_18302_Update/ack
      -- CP-element group 2: 	 branch_block_stmt_18305/$entry
      -- CP-element group 2: 	 branch_block_stmt_18305/branch_block_stmt_18305__entry__
      -- CP-element group 2: 	 branch_block_stmt_18305/merge_stmt_18306__entry__
      -- 
    ack_36400_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_READ_TX_QUEUE_INDEX_18302_inst_ack_1, ack => transmitEngineDaemon_CP_36381_elements(2)); -- 
    -- CP-element group 3:  transition  place  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (3) 
      -- CP-element group 3: 	 $exit
      -- CP-element group 3: 	 branch_block_stmt_18305/$exit
      -- CP-element group 3: 	 branch_block_stmt_18305/branch_block_stmt_18305__exit__
      -- 
    transmitEngineDaemon_CP_36381_elements(3) <= false; 
    -- CP-element group 4:  transition  place  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	85 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	86 
    -- CP-element group 4:  members (4) 
      -- CP-element group 4: 	 branch_block_stmt_18305/disable_loopback_PhiReq/$exit
      -- CP-element group 4: 	 branch_block_stmt_18305/disable_loopback_PhiReq/$entry
      -- CP-element group 4: 	 branch_block_stmt_18305/do_while_stmt_18315__exit__
      -- CP-element group 4: 	 branch_block_stmt_18305/disable_loopback
      -- 
    transmitEngineDaemon_CP_36381_elements(4) <= transmitEngineDaemon_CP_36381_elements(85);
    -- CP-element group 5:  transition  place  input  bypass 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	86 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	86 
    -- CP-element group 5:  members (5) 
      -- CP-element group 5: 	 branch_block_stmt_18305/not_enabled_yet_loopback_PhiReq/$exit
      -- CP-element group 5: 	 branch_block_stmt_18305/not_enabled_yet_loopback_PhiReq/$entry
      -- CP-element group 5: 	 branch_block_stmt_18305/if_stmt_18307_if_link/$exit
      -- CP-element group 5: 	 branch_block_stmt_18305/if_stmt_18307_if_link/if_choice_transition
      -- CP-element group 5: 	 branch_block_stmt_18305/not_enabled_yet_loopback
      -- 
    if_choice_transition_36473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 5_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_18307_branch_ack_1, ack => transmitEngineDaemon_CP_36381_elements(5)); -- 
    -- CP-element group 6:  merge  transition  place  input  bypass 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	86 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	7 
    -- CP-element group 6:  members (4) 
      -- CP-element group 6: 	 branch_block_stmt_18305/if_stmt_18307__exit__
      -- CP-element group 6: 	 branch_block_stmt_18305/do_while_stmt_18315__entry__
      -- CP-element group 6: 	 branch_block_stmt_18305/if_stmt_18307_else_link/$exit
      -- CP-element group 6: 	 branch_block_stmt_18305/if_stmt_18307_else_link/else_choice_transition
      -- 
    else_choice_transition_36477_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 6_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_18307_branch_ack_0, ack => transmitEngineDaemon_CP_36381_elements(6)); -- 
    -- CP-element group 7:  transition  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	6 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	13 
    -- CP-element group 7:  members (2) 
      -- CP-element group 7: 	 branch_block_stmt_18305/do_while_stmt_18315/$entry
      -- CP-element group 7: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315__entry__
      -- 
    transmitEngineDaemon_CP_36381_elements(7) <= transmitEngineDaemon_CP_36381_elements(6);
    -- CP-element group 8:  merge  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	85 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315__exit__
      -- 
    -- Element group transmitEngineDaemon_CP_36381_elements(8) is bound as output of CP function.
    -- CP-element group 9:  merge  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	12 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_18305/do_while_stmt_18315/loop_back
      -- 
    -- Element group transmitEngineDaemon_CP_36381_elements(9) is bound as output of CP function.
    -- CP-element group 10:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	15 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	83 
    -- CP-element group 10: 	84 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 branch_block_stmt_18305/do_while_stmt_18315/loop_exit/$entry
      -- CP-element group 10: 	 branch_block_stmt_18305/do_while_stmt_18315/loop_taken/$entry
      -- CP-element group 10: 	 branch_block_stmt_18305/do_while_stmt_18315/condition_done
      -- 
    transmitEngineDaemon_CP_36381_elements(10) <= transmitEngineDaemon_CP_36381_elements(15);
    -- CP-element group 11:  branch  place  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	82 
    -- CP-element group 11: successors 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_18305/do_while_stmt_18315/loop_body_done
      -- 
    transmitEngineDaemon_CP_36381_elements(11) <= transmitEngineDaemon_CP_36381_elements(82);
    -- CP-element group 12:  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	9 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	29 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/back_edge_to_loop_body
      -- 
    transmitEngineDaemon_CP_36381_elements(12) <= transmitEngineDaemon_CP_36381_elements(9);
    -- CP-element group 13:  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	7 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	31 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/first_time_through_loop_body
      -- 
    transmitEngineDaemon_CP_36381_elements(13) <= transmitEngineDaemon_CP_36381_elements(7);
    -- CP-element group 14:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	81 
    -- CP-element group 14: 	16 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	25 
    -- CP-element group 14: 	26 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/$entry
      -- CP-element group 14: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/loop_body_start
      -- CP-element group 14: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/phi_stmt_18317_sample_start_
      -- 
    -- Element group transmitEngineDaemon_CP_36381_elements(14) is bound as output of CP function.
    -- CP-element group 15:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	81 
    -- CP-element group 15: 	19 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/condition_evaluated
      -- 
    condition_evaluated_36493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_36493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_36381_elements(15), ack => do_while_stmt_18315_branch_req_0); -- 
    transmitEngineDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_36381_elements(81) & transmitEngineDaemon_CP_36381_elements(19);
      gj_transmitEngineDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_36381_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	14 
    -- CP-element group 16: 	25 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	19 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	21 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/aggregated_phi_sample_req
      -- CP-element group 16: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/phi_stmt_18327_sample_start__ps
      -- 
    transmitEngineDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_36381_elements(14) & transmitEngineDaemon_CP_36381_elements(25) & transmitEngineDaemon_CP_36381_elements(19);
      gj_transmitEngineDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_36381_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	23 
    -- CP-element group 17: 	27 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	47 
    -- CP-element group 17: 	51 
    -- CP-element group 17: 	71 
    -- CP-element group 17: 	82 
    -- CP-element group 17: 	75 
    -- CP-element group 17: marked-successors 
    -- CP-element group 17: 	25 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/aggregated_phi_sample_ack
      -- CP-element group 17: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/phi_stmt_18317_sample_completed_
      -- CP-element group 17: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/phi_stmt_18327_sample_completed_
      -- 
    transmitEngineDaemon_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_36381_elements(23) & transmitEngineDaemon_CP_36381_elements(27);
      gj_transmitEngineDaemon_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_36381_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	20 
    -- CP-element group 18: 	26 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	22 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/aggregated_phi_update_req
      -- CP-element group 18: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/phi_stmt_18327_update_start__ps
      -- 
    transmitEngineDaemon_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_36381_elements(20) & transmitEngineDaemon_CP_36381_elements(26);
      gj_transmitEngineDaemon_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_36381_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	24 
    -- CP-element group 19: 	28 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: marked-successors 
    -- CP-element group 19: 	16 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/aggregated_phi_update_ack
      -- 
    transmitEngineDaemon_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_36381_elements(24) & transmitEngineDaemon_CP_36381_elements(28);
      gj_transmitEngineDaemon_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_36381_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	14 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	44 
    -- CP-element group 20: 	79 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	18 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/phi_stmt_18317_update_start_
      -- 
    transmitEngineDaemon_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_36381_elements(14) & transmitEngineDaemon_CP_36381_elements(44) & transmitEngineDaemon_CP_36381_elements(79);
      gj_transmitEngineDaemon_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_36381_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	16 
    -- CP-element group 21: marked-predecessors 
    -- CP-element group 21: 	23 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	23 
    -- CP-element group 21:  members (3) 
      -- CP-element group 21: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/AND_u6_u6_18326_sample_start_
      -- CP-element group 21: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/AND_u6_u6_18326_Sample/$entry
      -- CP-element group 21: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/AND_u6_u6_18326_Sample/rr
      -- 
    rr_36510_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_36510_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_36381_elements(21), ack => AND_u6_u6_18326_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_21: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_21"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_36381_elements(16) & transmitEngineDaemon_CP_36381_elements(23);
      gj_transmitEngineDaemon_cp_element_group_21 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_36381_elements(21), clk => clk, reset => reset); --
    end block;
    -- CP-element group 22:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	18 
    -- CP-element group 22: marked-predecessors 
    -- CP-element group 22: 	24 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	24 
    -- CP-element group 22:  members (3) 
      -- CP-element group 22: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/AND_u6_u6_18326_update_start_
      -- CP-element group 22: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/AND_u6_u6_18326_Update/$entry
      -- CP-element group 22: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/AND_u6_u6_18326_Update/cr
      -- 
    cr_36515_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_36515_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_36381_elements(22), ack => AND_u6_u6_18326_inst_req_1); -- 
    transmitEngineDaemon_cp_element_group_22: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_22"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_36381_elements(18) & transmitEngineDaemon_CP_36381_elements(24);
      gj_transmitEngineDaemon_cp_element_group_22 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_36381_elements(22), clk => clk, reset => reset); --
    end block;
    -- CP-element group 23:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	21 
    -- CP-element group 23: successors 
    -- CP-element group 23: 	17 
    -- CP-element group 23: marked-successors 
    -- CP-element group 23: 	21 
    -- CP-element group 23:  members (3) 
      -- CP-element group 23: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/AND_u6_u6_18326_sample_completed_
      -- CP-element group 23: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/AND_u6_u6_18326_Sample/$exit
      -- CP-element group 23: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/AND_u6_u6_18326_Sample/ra
      -- 
    ra_36511_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u6_u6_18326_inst_ack_0, ack => transmitEngineDaemon_CP_36381_elements(23)); -- 
    -- CP-element group 24:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	22 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	78 
    -- CP-element group 24: 	19 
    -- CP-element group 24: 	42 
    -- CP-element group 24: marked-successors 
    -- CP-element group 24: 	22 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/phi_stmt_18317_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/AND_u6_u6_18326_update_completed_
      -- CP-element group 24: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/AND_u6_u6_18326_Update/$exit
      -- CP-element group 24: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/AND_u6_u6_18326_Update/ca
      -- 
    ca_36516_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u6_u6_18326_inst_ack_1, ack => transmitEngineDaemon_CP_36381_elements(24)); -- 
    -- CP-element group 25:  join  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	14 
    -- CP-element group 25: marked-predecessors 
    -- CP-element group 25: 	53 
    -- CP-element group 25: 	49 
    -- CP-element group 25: 	73 
    -- CP-element group 25: 	77 
    -- CP-element group 25: 	17 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	16 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/phi_stmt_18327_sample_start_
      -- 
    transmitEngineDaemon_cp_element_group_25: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 31,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_25"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_36381_elements(14) & transmitEngineDaemon_CP_36381_elements(53) & transmitEngineDaemon_CP_36381_elements(49) & transmitEngineDaemon_CP_36381_elements(73) & transmitEngineDaemon_CP_36381_elements(77) & transmitEngineDaemon_CP_36381_elements(17);
      gj_transmitEngineDaemon_cp_element_group_25 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_36381_elements(25), clk => clk, reset => reset); --
    end block;
    -- CP-element group 26:  join  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	14 
    -- CP-element group 26: marked-predecessors 
    -- CP-element group 26: 	64 
    -- CP-element group 26: 	72 
    -- CP-element group 26: 	76 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	18 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/phi_stmt_18327_update_start_
      -- 
    transmitEngineDaemon_cp_element_group_26: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_26"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_36381_elements(14) & transmitEngineDaemon_CP_36381_elements(64) & transmitEngineDaemon_CP_36381_elements(72) & transmitEngineDaemon_CP_36381_elements(76);
      gj_transmitEngineDaemon_cp_element_group_26 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_36381_elements(26), clk => clk, reset => reset); --
    end block;
    -- CP-element group 27:  join  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	17 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/phi_stmt_18327_sample_completed__ps
      -- 
    -- Element group transmitEngineDaemon_CP_36381_elements(27) is bound as output of CP function.
    -- CP-element group 28:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	62 
    -- CP-element group 28: 	70 
    -- CP-element group 28: 	74 
    -- CP-element group 28: 	19 
    -- CP-element group 28:  members (2) 
      -- CP-element group 28: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/phi_stmt_18327_update_completed_
      -- CP-element group 28: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/phi_stmt_18327_update_completed__ps
      -- 
    -- Element group transmitEngineDaemon_CP_36381_elements(28) is bound as output of CP function.
    -- CP-element group 29:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	12 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/phi_stmt_18327_loopback_trigger
      -- 
    transmitEngineDaemon_CP_36381_elements(29) <= transmitEngineDaemon_CP_36381_elements(12);
    -- CP-element group 30:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (2) 
      -- CP-element group 30: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/phi_stmt_18327_loopback_sample_req
      -- CP-element group 30: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/phi_stmt_18327_loopback_sample_req_ps
      -- 
    phi_stmt_18327_loopback_sample_req_36526_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_18327_loopback_sample_req_36526_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_36381_elements(30), ack => phi_stmt_18327_req_1); -- 
    -- Element group transmitEngineDaemon_CP_36381_elements(30) is bound as output of CP function.
    -- CP-element group 31:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	13 
    -- CP-element group 31: successors 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/phi_stmt_18327_entry_trigger
      -- 
    transmitEngineDaemon_CP_36381_elements(31) <= transmitEngineDaemon_CP_36381_elements(13);
    -- CP-element group 32:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (2) 
      -- CP-element group 32: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/phi_stmt_18327_entry_sample_req
      -- CP-element group 32: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/phi_stmt_18327_entry_sample_req_ps
      -- 
    phi_stmt_18327_entry_sample_req_36529_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_18327_entry_sample_req_36529_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_36381_elements(32), ack => phi_stmt_18327_req_0); -- 
    -- Element group transmitEngineDaemon_CP_36381_elements(32) is bound as output of CP function.
    -- CP-element group 33:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33:  members (2) 
      -- CP-element group 33: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/phi_stmt_18327_phi_mux_ack
      -- CP-element group 33: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/phi_stmt_18327_phi_mux_ack_ps
      -- 
    phi_stmt_18327_phi_mux_ack_36532_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_18327_ack_0, ack => transmitEngineDaemon_CP_36381_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/type_cast_18330_sample_start__ps
      -- CP-element group 34: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/type_cast_18330_sample_completed__ps
      -- CP-element group 34: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/type_cast_18330_sample_start_
      -- CP-element group 34: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/type_cast_18330_sample_completed_
      -- 
    -- Element group transmitEngineDaemon_CP_36381_elements(34) is bound as output of CP function.
    -- CP-element group 35:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (2) 
      -- CP-element group 35: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/type_cast_18330_update_start__ps
      -- CP-element group 35: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/type_cast_18330_update_start_
      -- 
    -- Element group transmitEngineDaemon_CP_36381_elements(35) is bound as output of CP function.
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	37 
    -- CP-element group 36: successors 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/type_cast_18330_update_completed__ps
      -- 
    transmitEngineDaemon_CP_36381_elements(36) <= transmitEngineDaemon_CP_36381_elements(37);
    -- CP-element group 37:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	36 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/type_cast_18330_update_completed_
      -- 
    -- Element group transmitEngineDaemon_CP_36381_elements(37) is a control-delay.
    cp_element_37_delay: control_delay_element  generic map(name => " 37_delay", delay_value => 1)  port map(req => transmitEngineDaemon_CP_36381_elements(35), ack => transmitEngineDaemon_CP_36381_elements(37), clk => clk, reset =>reset);
    -- CP-element group 38:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	40 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/R_ncount_18331_sample_start__ps
      -- CP-element group 38: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/R_ncount_18331_sample_start_
      -- CP-element group 38: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/R_ncount_18331_Sample/$entry
      -- CP-element group 38: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/R_ncount_18331_Sample/req
      -- 
    req_36553_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_36553_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_36381_elements(38), ack => ncount_18401_18331_buf_req_0); -- 
    -- Element group transmitEngineDaemon_CP_36381_elements(38) is bound as output of CP function.
    -- CP-element group 39:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39:  members (4) 
      -- CP-element group 39: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/R_ncount_18331_update_start__ps
      -- CP-element group 39: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/R_ncount_18331_update_start_
      -- CP-element group 39: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/R_ncount_18331_Update/$entry
      -- CP-element group 39: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/R_ncount_18331_Update/req
      -- 
    req_36558_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_36558_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_36381_elements(39), ack => ncount_18401_18331_buf_req_1); -- 
    -- Element group transmitEngineDaemon_CP_36381_elements(39) is bound as output of CP function.
    -- CP-element group 40:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	38 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (4) 
      -- CP-element group 40: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/R_ncount_18331_sample_completed__ps
      -- CP-element group 40: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/R_ncount_18331_sample_completed_
      -- CP-element group 40: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/R_ncount_18331_Sample/$exit
      -- CP-element group 40: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/R_ncount_18331_Sample/ack
      -- 
    ack_36554_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 40_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ncount_18401_18331_buf_ack_0, ack => transmitEngineDaemon_CP_36381_elements(40)); -- 
    -- CP-element group 41:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (4) 
      -- CP-element group 41: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/R_ncount_18331_update_completed__ps
      -- CP-element group 41: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/R_ncount_18331_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/R_ncount_18331_Update/$exit
      -- CP-element group 41: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/R_ncount_18331_Update/ack
      -- 
    ack_36559_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ncount_18401_18331_buf_ack_1, ack => transmitEngineDaemon_CP_36381_elements(41)); -- 
    -- CP-element group 42:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	24 
    -- CP-element group 42: marked-predecessors 
    -- CP-element group 42: 	61 
    -- CP-element group 42: 	44 
    -- CP-element group 42: 	69 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	44 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18338_sample_start_
      -- CP-element group 42: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18338_Sample/$entry
      -- CP-element group 42: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18338_Sample/crr
      -- 
    crr_36568_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_36568_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_36381_elements(42), ack => call_stmt_18338_call_req_0); -- 
    transmitEngineDaemon_cp_element_group_42: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 1,3 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_42"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_36381_elements(24) & transmitEngineDaemon_CP_36381_elements(61) & transmitEngineDaemon_CP_36381_elements(44) & transmitEngineDaemon_CP_36381_elements(69);
      gj_transmitEngineDaemon_cp_element_group_42 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_36381_elements(42), clk => clk, reset => reset); --
    end block;
    -- CP-element group 43:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: marked-predecessors 
    -- CP-element group 43: 	56 
    -- CP-element group 43: 	61 
    -- CP-element group 43: 	48 
    -- CP-element group 43: 	52 
    -- CP-element group 43: 	69 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	45 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18338_update_start_
      -- CP-element group 43: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18338_Update/$entry
      -- CP-element group 43: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18338_Update/ccr
      -- 
    ccr_36573_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_36573_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_36381_elements(43), ack => call_stmt_18338_call_req_1); -- 
    transmitEngineDaemon_cp_element_group_43: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_43"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_36381_elements(56) & transmitEngineDaemon_CP_36381_elements(61) & transmitEngineDaemon_CP_36381_elements(48) & transmitEngineDaemon_CP_36381_elements(52) & transmitEngineDaemon_CP_36381_elements(69);
      gj_transmitEngineDaemon_cp_element_group_43 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_36381_elements(43), clk => clk, reset => reset); --
    end block;
    -- CP-element group 44:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: successors 
    -- CP-element group 44: marked-successors 
    -- CP-element group 44: 	20 
    -- CP-element group 44: 	42 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18338_sample_completed_
      -- CP-element group 44: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18338_Sample/$exit
      -- CP-element group 44: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18338_Sample/cra
      -- 
    cra_36569_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_18338_call_ack_0, ack => transmitEngineDaemon_CP_36381_elements(44)); -- 
    -- CP-element group 45:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	43 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	54 
    -- CP-element group 45: 	46 
    -- CP-element group 45: 	50 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18338_update_completed_
      -- CP-element group 45: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18338_Update/$exit
      -- CP-element group 45: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18338_Update/cca
      -- 
    cca_36574_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_18338_call_ack_1, ack => transmitEngineDaemon_CP_36381_elements(45)); -- 
    -- CP-element group 46:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	45 
    -- CP-element group 46: marked-predecessors 
    -- CP-element group 46: 	48 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18342_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18342_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18342_Sample/crr
      -- 
    crr_36582_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_36582_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_36381_elements(46), ack => call_stmt_18342_call_req_0); -- 
    transmitEngineDaemon_cp_element_group_46: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_46"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_36381_elements(45) & transmitEngineDaemon_CP_36381_elements(48);
      gj_transmitEngineDaemon_cp_element_group_46 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_36381_elements(46), clk => clk, reset => reset); --
    end block;
    -- CP-element group 47:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	17 
    -- CP-element group 47: marked-predecessors 
    -- CP-element group 47: 	60 
    -- CP-element group 47: 	68 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18342_update_start_
      -- CP-element group 47: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18342_Update/$entry
      -- CP-element group 47: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18342_Update/ccr
      -- 
    ccr_36587_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_36587_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_36381_elements(47), ack => call_stmt_18342_call_req_1); -- 
    transmitEngineDaemon_cp_element_group_47: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_47"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_36381_elements(17) & transmitEngineDaemon_CP_36381_elements(60) & transmitEngineDaemon_CP_36381_elements(68);
      gj_transmitEngineDaemon_cp_element_group_47 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_36381_elements(47), clk => clk, reset => reset); --
    end block;
    -- CP-element group 48:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: marked-successors 
    -- CP-element group 48: 	43 
    -- CP-element group 48: 	46 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18342_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18342_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18342_Sample/cra
      -- 
    cra_36583_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_18342_call_ack_0, ack => transmitEngineDaemon_CP_36381_elements(48)); -- 
    -- CP-element group 49:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	58 
    -- CP-element group 49: 	66 
    -- CP-element group 49: marked-successors 
    -- CP-element group 49: 	25 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18342_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18342_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18342_Update/cca
      -- 
    cca_36588_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_18342_call_ack_1, ack => transmitEngineDaemon_CP_36381_elements(49)); -- 
    -- CP-element group 50:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	45 
    -- CP-element group 50: marked-predecessors 
    -- CP-element group 50: 	52 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/NOT_u1_u1_18352_Sample/$entry
      -- CP-element group 50: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/NOT_u1_u1_18352_Sample/rr
      -- CP-element group 50: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/NOT_u1_u1_18352_sample_start_
      -- 
    rr_36596_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_36596_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_36381_elements(50), ack => NOT_u1_u1_18352_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_36381_elements(45) & transmitEngineDaemon_CP_36381_elements(52);
      gj_transmitEngineDaemon_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_36381_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	17 
    -- CP-element group 51: marked-predecessors 
    -- CP-element group 51: 	60 
    -- CP-element group 51: 	68 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/NOT_u1_u1_18352_Update/$entry
      -- CP-element group 51: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/NOT_u1_u1_18352_Update/cr
      -- CP-element group 51: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/NOT_u1_u1_18352_update_start_
      -- 
    cr_36601_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_36601_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_36381_elements(51), ack => NOT_u1_u1_18352_inst_req_1); -- 
    transmitEngineDaemon_cp_element_group_51: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_51"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_36381_elements(17) & transmitEngineDaemon_CP_36381_elements(60) & transmitEngineDaemon_CP_36381_elements(68);
      gj_transmitEngineDaemon_cp_element_group_51 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_36381_elements(51), clk => clk, reset => reset); --
    end block;
    -- CP-element group 52:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: marked-successors 
    -- CP-element group 52: 	43 
    -- CP-element group 52: 	50 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/NOT_u1_u1_18352_Sample/ra
      -- CP-element group 52: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/NOT_u1_u1_18352_Sample/$exit
      -- CP-element group 52: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/NOT_u1_u1_18352_sample_completed_
      -- 
    ra_36597_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_18352_inst_ack_0, ack => transmitEngineDaemon_CP_36381_elements(52)); -- 
    -- CP-element group 53:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	58 
    -- CP-element group 53: 	66 
    -- CP-element group 53: marked-successors 
    -- CP-element group 53: 	25 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/NOT_u1_u1_18352_update_completed_
      -- CP-element group 53: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/NOT_u1_u1_18352_Update/$exit
      -- CP-element group 53: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/NOT_u1_u1_18352_Update/ca
      -- 
    ca_36602_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => NOT_u1_u1_18352_inst_ack_1, ack => transmitEngineDaemon_CP_36381_elements(53)); -- 
    -- CP-element group 54:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	45 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	56 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18364_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18364_Sample/req
      -- CP-element group 54: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18364_sample_start_
      -- 
    req_36610_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_36610_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_36381_elements(54), ack => W_pkt_pointer_17554_delayed_4_0_18362_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_36381_elements(45) & transmitEngineDaemon_CP_36381_elements(56);
      gj_transmitEngineDaemon_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_36381_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: marked-predecessors 
    -- CP-element group 55: 	60 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18364_Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18364_update_start_
      -- CP-element group 55: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18364_Update/req
      -- 
    req_36615_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_36615_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_36381_elements(55), ack => W_pkt_pointer_17554_delayed_4_0_18362_inst_req_1); -- 
    transmitEngineDaemon_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= transmitEngineDaemon_CP_36381_elements(60);
      gj_transmitEngineDaemon_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_36381_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: marked-successors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: 	43 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18364_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18364_Sample/ack
      -- CP-element group 56: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18364_sample_completed_
      -- 
    ack_36611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_pkt_pointer_17554_delayed_4_0_18362_inst_ack_0, ack => transmitEngineDaemon_CP_36381_elements(56)); -- 
    -- CP-element group 57:  transition  input  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18364_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18364_Update/ack
      -- CP-element group 57: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18364_Update/$exit
      -- 
    ack_36616_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_pkt_pointer_17554_delayed_4_0_18362_inst_ack_1, ack => transmitEngineDaemon_CP_36381_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	53 
    -- CP-element group 58: 	57 
    -- CP-element group 58: 	49 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	60 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18371_Sample/crr
      -- CP-element group 58: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18371_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18371_sample_start_
      -- 
    crr_36624_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_36624_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_36381_elements(58), ack => call_stmt_18371_call_req_0); -- 
    transmitEngineDaemon_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_36381_elements(53) & transmitEngineDaemon_CP_36381_elements(57) & transmitEngineDaemon_CP_36381_elements(49) & transmitEngineDaemon_CP_36381_elements(60);
      gj_transmitEngineDaemon_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_36381_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18371_Update/ccr
      -- CP-element group 59: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18371_Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18371_update_start_
      -- 
    ccr_36629_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_36629_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_36381_elements(59), ack => call_stmt_18371_call_req_1); -- 
    transmitEngineDaemon_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= transmitEngineDaemon_CP_36381_elements(61);
      gj_transmitEngineDaemon_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_36381_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	55 
    -- CP-element group 60: 	58 
    -- CP-element group 60: 	47 
    -- CP-element group 60: 	51 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18371_Sample/cra
      -- CP-element group 60: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18371_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18371_sample_completed_
      -- 
    cra_36625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_18371_call_ack_0, ack => transmitEngineDaemon_CP_36381_elements(60)); -- 
    -- CP-element group 61:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	82 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: 	43 
    -- CP-element group 61: 	42 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18371_Update/cca
      -- CP-element group 61: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18371_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18371_update_completed_
      -- 
    cca_36630_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_18371_call_ack_1, ack => transmitEngineDaemon_CP_36381_elements(61)); -- 
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	28 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	64 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18377_sample_start_
      -- CP-element group 62: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18377_Sample/$entry
      -- CP-element group 62: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18377_Sample/req
      -- 
    req_36638_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_36638_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_36381_elements(62), ack => W_count_17567_delayed_14_0_18375_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_36381_elements(28) & transmitEngineDaemon_CP_36381_elements(64);
      gj_transmitEngineDaemon_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_36381_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: marked-predecessors 
    -- CP-element group 63: 	68 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	65 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18377_update_start_
      -- CP-element group 63: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18377_Update/req
      -- CP-element group 63: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18377_Update/$entry
      -- 
    req_36643_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_36643_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_36381_elements(63), ack => W_count_17567_delayed_14_0_18375_inst_req_1); -- 
    transmitEngineDaemon_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= transmitEngineDaemon_CP_36381_elements(68);
      gj_transmitEngineDaemon_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_36381_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: 	26 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18377_sample_completed_
      -- CP-element group 64: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18377_Sample/$exit
      -- CP-element group 64: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18377_Sample/ack
      -- 
    ack_36639_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_count_17567_delayed_14_0_18375_inst_ack_0, ack => transmitEngineDaemon_CP_36381_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	63 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18377_update_completed_
      -- CP-element group 65: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18377_Update/ack
      -- CP-element group 65: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18377_Update/$exit
      -- 
    ack_36644_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_count_17567_delayed_14_0_18375_inst_ack_1, ack => transmitEngineDaemon_CP_36381_elements(65)); -- 
    -- CP-element group 66:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	53 
    -- CP-element group 66: 	49 
    -- CP-element group 66: 	65 
    -- CP-element group 66: marked-predecessors 
    -- CP-element group 66: 	68 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18387_Sample/crr
      -- CP-element group 66: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18387_Sample/$entry
      -- CP-element group 66: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18387_sample_start_
      -- 
    crr_36652_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_36652_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_36381_elements(66), ack => call_stmt_18387_call_req_0); -- 
    transmitEngineDaemon_cp_element_group_66: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_66"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_36381_elements(53) & transmitEngineDaemon_CP_36381_elements(49) & transmitEngineDaemon_CP_36381_elements(65) & transmitEngineDaemon_CP_36381_elements(68);
      gj_transmitEngineDaemon_cp_element_group_66 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_36381_elements(66), clk => clk, reset => reset); --
    end block;
    -- CP-element group 67:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: marked-predecessors 
    -- CP-element group 67: 	69 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	69 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18387_Update/ccr
      -- CP-element group 67: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18387_Update/$entry
      -- CP-element group 67: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18387_update_start_
      -- 
    ccr_36657_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_36657_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_36381_elements(67), ack => call_stmt_18387_call_req_1); -- 
    transmitEngineDaemon_cp_element_group_67: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_67"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= transmitEngineDaemon_CP_36381_elements(69);
      gj_transmitEngineDaemon_cp_element_group_67 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_36381_elements(67), clk => clk, reset => reset); --
    end block;
    -- CP-element group 68:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68: marked-successors 
    -- CP-element group 68: 	47 
    -- CP-element group 68: 	51 
    -- CP-element group 68: 	63 
    -- CP-element group 68: 	66 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18387_Sample/cra
      -- CP-element group 68: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18387_Sample/$exit
      -- CP-element group 68: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18387_sample_completed_
      -- 
    cra_36653_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_18387_call_ack_0, ack => transmitEngineDaemon_CP_36381_elements(68)); -- 
    -- CP-element group 69:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: 	67 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	82 
    -- CP-element group 69: marked-successors 
    -- CP-element group 69: 	43 
    -- CP-element group 69: 	67 
    -- CP-element group 69: 	42 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18387_Update/$exit
      -- CP-element group 69: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18387_Update/cca
      -- CP-element group 69: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/call_stmt_18387_update_completed_
      -- 
    cca_36658_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 69_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_18387_call_ack_1, ack => transmitEngineDaemon_CP_36381_elements(69)); -- 
    -- CP-element group 70:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	28 
    -- CP-element group 70: marked-predecessors 
    -- CP-element group 70: 	72 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/ADD_u32_u32_18391_sample_start_
      -- CP-element group 70: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/ADD_u32_u32_18391_Sample/$entry
      -- CP-element group 70: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/ADD_u32_u32_18391_Sample/rr
      -- 
    rr_36666_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_36666_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_36381_elements(70), ack => ADD_u32_u32_18391_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_70: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_70"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_36381_elements(28) & transmitEngineDaemon_CP_36381_elements(72);
      gj_transmitEngineDaemon_cp_element_group_70 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_36381_elements(70), clk => clk, reset => reset); --
    end block;
    -- CP-element group 71:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	17 
    -- CP-element group 71: marked-predecessors 
    -- CP-element group 71: 	73 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/ADD_u32_u32_18391_update_start_
      -- CP-element group 71: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/ADD_u32_u32_18391_Update/cr
      -- CP-element group 71: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/ADD_u32_u32_18391_Update/$entry
      -- 
    cr_36671_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_36671_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_36381_elements(71), ack => ADD_u32_u32_18391_inst_req_1); -- 
    transmitEngineDaemon_cp_element_group_71: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_71"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_36381_elements(17) & transmitEngineDaemon_CP_36381_elements(73);
      gj_transmitEngineDaemon_cp_element_group_71 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_36381_elements(71), clk => clk, reset => reset); --
    end block;
    -- CP-element group 72:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: marked-successors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: 	26 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/ADD_u32_u32_18391_sample_completed_
      -- CP-element group 72: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/ADD_u32_u32_18391_Sample/ra
      -- CP-element group 72: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/ADD_u32_u32_18391_Sample/$exit
      -- 
    ra_36667_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 72_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_18391_inst_ack_0, ack => transmitEngineDaemon_CP_36381_elements(72)); -- 
    -- CP-element group 73:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	82 
    -- CP-element group 73: marked-successors 
    -- CP-element group 73: 	71 
    -- CP-element group 73: 	25 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/ADD_u32_u32_18391_update_completed_
      -- CP-element group 73: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/ADD_u32_u32_18391_Update/ca
      -- CP-element group 73: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/ADD_u32_u32_18391_Update/$exit
      -- 
    ca_36672_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 73_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u32_u32_18391_inst_ack_1, ack => transmitEngineDaemon_CP_36381_elements(73)); -- 
    -- CP-element group 74:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	28 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	76 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18395_Sample/$entry
      -- CP-element group 74: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18395_sample_start_
      -- CP-element group 74: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18395_Sample/req
      -- 
    req_36680_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_36680_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_36381_elements(74), ack => W_count_17575_delayed_14_0_18393_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_36381_elements(28) & transmitEngineDaemon_CP_36381_elements(76);
      gj_transmitEngineDaemon_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_36381_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	17 
    -- CP-element group 75: marked-predecessors 
    -- CP-element group 75: 	77 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	77 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18395_Update/$entry
      -- CP-element group 75: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18395_Update/req
      -- CP-element group 75: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18395_update_start_
      -- 
    req_36685_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_36685_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_36381_elements(75), ack => W_count_17575_delayed_14_0_18393_inst_req_1); -- 
    transmitEngineDaemon_cp_element_group_75: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_75"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_36381_elements(17) & transmitEngineDaemon_CP_36381_elements(77);
      gj_transmitEngineDaemon_cp_element_group_75 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_36381_elements(75), clk => clk, reset => reset); --
    end block;
    -- CP-element group 76:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76: marked-successors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: 	26 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18395_Sample/$exit
      -- CP-element group 76: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18395_Sample/ack
      -- CP-element group 76: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18395_sample_completed_
      -- 
    ack_36681_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_count_17575_delayed_14_0_18393_inst_ack_0, ack => transmitEngineDaemon_CP_36381_elements(76)); -- 
    -- CP-element group 77:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	82 
    -- CP-element group 77: marked-successors 
    -- CP-element group 77: 	75 
    -- CP-element group 77: 	25 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18395_update_completed_
      -- CP-element group 77: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18395_Update/$exit
      -- CP-element group 77: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/assign_stmt_18395_Update/ack
      -- 
    ack_36686_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_count_17575_delayed_14_0_18393_inst_ack_1, ack => transmitEngineDaemon_CP_36381_elements(77)); -- 
    -- CP-element group 78:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	24 
    -- CP-element group 78: marked-predecessors 
    -- CP-element group 78: 	80 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_18404_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_18404_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_18404_Sample/req
      -- 
    req_36694_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_36694_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_36381_elements(78), ack => WPIPE_LAST_READ_TX_QUEUE_INDEX_18404_inst_req_0); -- 
    transmitEngineDaemon_cp_element_group_78: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_78"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_36381_elements(24) & transmitEngineDaemon_CP_36381_elements(80);
      gj_transmitEngineDaemon_cp_element_group_78 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_36381_elements(78), clk => clk, reset => reset); --
    end block;
    -- CP-element group 79:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79: marked-successors 
    -- CP-element group 79: 	20 
    -- CP-element group 79:  members (6) 
      -- CP-element group 79: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_18404_Update/req
      -- CP-element group 79: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_18404_update_start_
      -- CP-element group 79: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_18404_sample_completed_
      -- CP-element group 79: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_18404_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_18404_Update/$entry
      -- CP-element group 79: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_18404_Sample/ack
      -- 
    ack_36695_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_READ_TX_QUEUE_INDEX_18404_inst_ack_0, ack => transmitEngineDaemon_CP_36381_elements(79)); -- 
    req_36699_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_36699_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_36381_elements(79), ack => WPIPE_LAST_READ_TX_QUEUE_INDEX_18404_inst_req_1); -- 
    -- CP-element group 80:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	79 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80: marked-successors 
    -- CP-element group 80: 	78 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_18404_Update/ack
      -- CP-element group 80: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_18404_update_completed_
      -- CP-element group 80: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/WPIPE_LAST_READ_TX_QUEUE_INDEX_18404_Update/$exit
      -- 
    ack_36700_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_LAST_READ_TX_QUEUE_INDEX_18404_inst_ack_1, ack => transmitEngineDaemon_CP_36381_elements(80)); -- 
    -- CP-element group 81:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	14 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	15 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group transmitEngineDaemon_CP_36381_elements(81) is a control-delay.
    cp_element_81_delay: control_delay_element  generic map(name => " 81_delay", delay_value => 1)  port map(req => transmitEngineDaemon_CP_36381_elements(14), ack => transmitEngineDaemon_CP_36381_elements(81), clk => clk, reset =>reset);
    -- CP-element group 82:  join  transition  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	61 
    -- CP-element group 82: 	69 
    -- CP-element group 82: 	80 
    -- CP-element group 82: 	73 
    -- CP-element group 82: 	77 
    -- CP-element group 82: 	17 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	11 
    -- CP-element group 82:  members (1) 
      -- CP-element group 82: 	 branch_block_stmt_18305/do_while_stmt_18315/do_while_stmt_18315_loop_body/$exit
      -- 
    transmitEngineDaemon_cp_element_group_82: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 31,1 => 31,2 => 31,3 => 31,4 => 31,5 => 31);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 40) := "transmitEngineDaemon_cp_element_group_82"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= transmitEngineDaemon_CP_36381_elements(61) & transmitEngineDaemon_CP_36381_elements(69) & transmitEngineDaemon_CP_36381_elements(80) & transmitEngineDaemon_CP_36381_elements(73) & transmitEngineDaemon_CP_36381_elements(77) & transmitEngineDaemon_CP_36381_elements(17);
      gj_transmitEngineDaemon_cp_element_group_82 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitEngineDaemon_CP_36381_elements(82), clk => clk, reset => reset); --
    end block;
    -- CP-element group 83:  transition  input  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	10 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_18305/do_while_stmt_18315/loop_exit/$exit
      -- CP-element group 83: 	 branch_block_stmt_18305/do_while_stmt_18315/loop_exit/ack
      -- 
    ack_36705_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_18315_branch_ack_0, ack => transmitEngineDaemon_CP_36381_elements(83)); -- 
    -- CP-element group 84:  transition  input  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	10 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (2) 
      -- CP-element group 84: 	 branch_block_stmt_18305/do_while_stmt_18315/loop_taken/ack
      -- CP-element group 84: 	 branch_block_stmt_18305/do_while_stmt_18315/loop_taken/$exit
      -- 
    ack_36709_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_18315_branch_ack_1, ack => transmitEngineDaemon_CP_36381_elements(84)); -- 
    -- CP-element group 85:  transition  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	8 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	4 
    -- CP-element group 85:  members (1) 
      -- CP-element group 85: 	 branch_block_stmt_18305/do_while_stmt_18315/$exit
      -- 
    transmitEngineDaemon_CP_36381_elements(85) <= transmitEngineDaemon_CP_36381_elements(8);
    -- CP-element group 86:  merge  branch  transition  place  output  bypass 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	2 
    -- CP-element group 86: 	4 
    -- CP-element group 86: 	5 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	5 
    -- CP-element group 86: 	6 
    -- CP-element group 86:  members (49) 
      -- CP-element group 86: 	 branch_block_stmt_18305/merge_stmt_18306_PhiAck/dummy
      -- CP-element group 86: 	 branch_block_stmt_18305/merge_stmt_18306_PhiAck/$exit
      -- CP-element group 86: 	 branch_block_stmt_18305/merge_stmt_18306_PhiAck/$entry
      -- CP-element group 86: 	 branch_block_stmt_18305/merge_stmt_18306_PhiReqMerge
      -- CP-element group 86: 	 branch_block_stmt_18305/merge_stmt_18306__exit__
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307__entry__
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_dead_link/$entry
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/$entry
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/$exit
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/$entry
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/$exit
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/BITSEL_u32_u1_18310/$entry
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/BITSEL_u32_u1_18310/$exit
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/BITSEL_u32_u1_18310/BITSEL_u32_u1_18310_inputs/$entry
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/BITSEL_u32_u1_18310/BITSEL_u32_u1_18310_inputs/$exit
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/BITSEL_u32_u1_18310/BITSEL_u32_u1_18310_inputs/RPIPE_CONTROL_REGISTER_18308/$entry
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/BITSEL_u32_u1_18310/BITSEL_u32_u1_18310_inputs/RPIPE_CONTROL_REGISTER_18308/$exit
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/BITSEL_u32_u1_18310/BITSEL_u32_u1_18310_inputs/RPIPE_CONTROL_REGISTER_18308/Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/BITSEL_u32_u1_18310/BITSEL_u32_u1_18310_inputs/RPIPE_CONTROL_REGISTER_18308/Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/BITSEL_u32_u1_18310/BITSEL_u32_u1_18310_inputs/RPIPE_CONTROL_REGISTER_18308/Sample/req
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/BITSEL_u32_u1_18310/BITSEL_u32_u1_18310_inputs/RPIPE_CONTROL_REGISTER_18308/Sample/ack
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/BITSEL_u32_u1_18310/BITSEL_u32_u1_18310_inputs/RPIPE_CONTROL_REGISTER_18308/Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/BITSEL_u32_u1_18310/BITSEL_u32_u1_18310_inputs/RPIPE_CONTROL_REGISTER_18308/Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/BITSEL_u32_u1_18310/BITSEL_u32_u1_18310_inputs/RPIPE_CONTROL_REGISTER_18308/Update/req
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/BITSEL_u32_u1_18310/BITSEL_u32_u1_18310_inputs/RPIPE_CONTROL_REGISTER_18308/Update/ack
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/BITSEL_u32_u1_18310/SplitProtocol/$entry
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/BITSEL_u32_u1_18310/SplitProtocol/$exit
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/BITSEL_u32_u1_18310/SplitProtocol/Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/BITSEL_u32_u1_18310/SplitProtocol/Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/BITSEL_u32_u1_18310/SplitProtocol/Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/BITSEL_u32_u1_18310/SplitProtocol/Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/BITSEL_u32_u1_18310/SplitProtocol/Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/BITSEL_u32_u1_18310/SplitProtocol/Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/BITSEL_u32_u1_18310/SplitProtocol/Update/cr
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/BITSEL_u32_u1_18310/SplitProtocol/Update/ca
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/SplitProtocol/$entry
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/SplitProtocol/$exit
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/SplitProtocol/Sample/$entry
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/SplitProtocol/Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/SplitProtocol/Sample/rr
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/SplitProtocol/Sample/ra
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/SplitProtocol/Update/$entry
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/SplitProtocol/Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/SplitProtocol/Update/cr
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/NOT_u1_u1_18311/SplitProtocol/Update/ca
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_eval_test/branch_req
      -- CP-element group 86: 	 branch_block_stmt_18305/NOT_u1_u1_18311_place
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_if_link/$entry
      -- CP-element group 86: 	 branch_block_stmt_18305/if_stmt_18307_else_link/$entry
      -- 
    branch_req_36468_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_36468_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitEngineDaemon_CP_36381_elements(86), ack => if_stmt_18307_branch_req_0); -- 
    transmitEngineDaemon_CP_36381_elements(86) <= OrReduce(transmitEngineDaemon_CP_36381_elements(2) & transmitEngineDaemon_CP_36381_elements(4) & transmitEngineDaemon_CP_36381_elements(5));
    transmitEngineDaemon_do_while_stmt_18315_terminator_36710: loop_terminator -- 
      generic map (name => " transmitEngineDaemon_do_while_stmt_18315_terminator_36710", max_iterations_in_flight =>31) 
      port map(loop_body_exit => transmitEngineDaemon_CP_36381_elements(11),loop_continue => transmitEngineDaemon_CP_36381_elements(84),loop_terminate => transmitEngineDaemon_CP_36381_elements(83),loop_back => transmitEngineDaemon_CP_36381_elements(9),loop_exit => transmitEngineDaemon_CP_36381_elements(8),clk => clk, reset => reset); -- 
    phi_stmt_18327_phi_seq_36560_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= transmitEngineDaemon_CP_36381_elements(31);
      transmitEngineDaemon_CP_36381_elements(34)<= src_sample_reqs(0);
      src_sample_acks(0)  <= transmitEngineDaemon_CP_36381_elements(34);
      transmitEngineDaemon_CP_36381_elements(35)<= src_update_reqs(0);
      src_update_acks(0)  <= transmitEngineDaemon_CP_36381_elements(36);
      transmitEngineDaemon_CP_36381_elements(32) <= phi_mux_reqs(0);
      triggers(1)  <= transmitEngineDaemon_CP_36381_elements(29);
      transmitEngineDaemon_CP_36381_elements(38)<= src_sample_reqs(1);
      src_sample_acks(1)  <= transmitEngineDaemon_CP_36381_elements(40);
      transmitEngineDaemon_CP_36381_elements(39)<= src_update_reqs(1);
      src_update_acks(1)  <= transmitEngineDaemon_CP_36381_elements(41);
      transmitEngineDaemon_CP_36381_elements(30) <= phi_mux_reqs(1);
      phi_stmt_18327_phi_seq_36560 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_18327_phi_seq_36560") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => transmitEngineDaemon_CP_36381_elements(16), 
          phi_sample_ack => transmitEngineDaemon_CP_36381_elements(27), 
          phi_update_req => transmitEngineDaemon_CP_36381_elements(18), 
          phi_update_ack => transmitEngineDaemon_CP_36381_elements(28), 
          phi_mux_ack => transmitEngineDaemon_CP_36381_elements(33), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_36494_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= transmitEngineDaemon_CP_36381_elements(12);
        preds(1)  <= transmitEngineDaemon_CP_36381_elements(13);
        entry_tmerge_36494 : transition_merge -- 
          generic map(name => " entry_tmerge_36494")
          port map (preds => preds, symbol_out => transmitEngineDaemon_CP_36381_elements(14));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u32_u32_17574_17574_delayed_14_0_18392 : std_logic_vector(31 downto 0);
    signal ADD_u6_u6_18321_wire : std_logic_vector(5 downto 0);
    signal AND_u6_u6_18326_wire : std_logic_vector(5 downto 0);
    signal BITSEL_u32_u1_18310_wire : std_logic_vector(0 downto 0);
    signal BITSEL_u32_u1_18410_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_17543_17543_delayed_4_0_18353 : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_18311_wire : std_logic_vector(0 downto 0);
    signal NOT_u4_u4_18383_wire_constant : std_logic_vector(3 downto 0);
    signal RPIPE_CONTROL_REGISTER_18308_wire : std_logic_vector(31 downto 0);
    signal RPIPE_CONTROL_REGISTER_18408_wire : std_logic_vector(31 downto 0);
    signal RPIPE_FREE_Q_18368_wire : std_logic_vector(35 downto 0);
    signal RPIPE_LAST_READ_TX_QUEUE_INDEX_18319_wire : std_logic_vector(5 downto 0);
    signal RPIPE_NUMBER_OF_SERVERS_18322_wire : std_logic_vector(31 downto 0);
    signal SUB_u32_u32_18324_wire : std_logic_vector(31 downto 0);
    signal count_17567_delayed_14_0_18377 : std_logic_vector(31 downto 0);
    signal count_17575_delayed_14_0_18395 : std_logic_vector(31 downto 0);
    signal count_18327 : std_logic_vector(31 downto 0);
    signal ignore_resp_18387 : std_logic_vector(31 downto 0);
    signal konst_18303_wire_constant : std_logic_vector(5 downto 0);
    signal konst_18309_wire_constant : std_logic_vector(31 downto 0);
    signal konst_18320_wire_constant : std_logic_vector(5 downto 0);
    signal konst_18323_wire_constant : std_logic_vector(31 downto 0);
    signal konst_18384_wire_constant : std_logic_vector(5 downto 0);
    signal konst_18390_wire_constant : std_logic_vector(31 downto 0);
    signal konst_18409_wire_constant : std_logic_vector(31 downto 0);
    signal ncount_18401 : std_logic_vector(31 downto 0);
    signal ncount_18401_18331_buffered : std_logic_vector(31 downto 0);
    signal pkt_pointer_17554_delayed_4_0_18364 : std_logic_vector(31 downto 0);
    signal pkt_pointer_18338 : std_logic_vector(31 downto 0);
    signal push_pointer_back_to_free_Q_18358 : std_logic_vector(0 downto 0);
    signal push_status_18371 : std_logic_vector(0 downto 0);
    signal transmitted_flag_18342 : std_logic_vector(0 downto 0);
    signal tx_flag_18338 : std_logic_vector(0 downto 0);
    signal tx_q_index_18317 : std_logic_vector(5 downto 0);
    signal type_cast_18325_wire : std_logic_vector(5 downto 0);
    signal type_cast_18330_wire_constant : std_logic_vector(31 downto 0);
    signal type_cast_18367_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_18380_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    NOT_u4_u4_18383_wire_constant <= "1111";
    konst_18303_wire_constant <= "000000";
    konst_18309_wire_constant <= "00000000000000000000000000000000";
    konst_18320_wire_constant <= "000001";
    konst_18323_wire_constant <= "00000000000000000000000000000001";
    konst_18384_wire_constant <= "010101";
    konst_18390_wire_constant <= "00000000000000000000000000000001";
    konst_18409_wire_constant <= "00000000000000000000000000000000";
    type_cast_18330_wire_constant <= "00000000000000000000000000000001";
    type_cast_18367_wire_constant <= "1";
    type_cast_18380_wire_constant <= "0";
    phi_stmt_18327: Block -- phi operator 
      signal idata: std_logic_vector(63 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_18330_wire_constant & ncount_18401_18331_buffered;
      req <= phi_stmt_18327_req_0 & phi_stmt_18327_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_18327",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 32) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_18327_ack_0,
          idata => idata,
          odata => count_18327,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_18327
    -- flow-through select operator MUX_18400_inst
    ncount_18401 <= ADD_u32_u32_17574_17574_delayed_14_0_18392 when (push_pointer_back_to_free_Q_18358(0) /=  '0') else count_17575_delayed_14_0_18395;
    W_count_17567_delayed_14_0_18375_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_count_17567_delayed_14_0_18375_inst_req_0;
      W_count_17567_delayed_14_0_18375_inst_ack_0<= wack(0);
      rreq(0) <= W_count_17567_delayed_14_0_18375_inst_req_1;
      W_count_17567_delayed_14_0_18375_inst_ack_1<= rack(0);
      W_count_17567_delayed_14_0_18375_inst : InterlockBuffer generic map ( -- 
        name => "W_count_17567_delayed_14_0_18375_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_18327,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => count_17567_delayed_14_0_18377,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_count_17575_delayed_14_0_18393_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_count_17575_delayed_14_0_18393_inst_req_0;
      W_count_17575_delayed_14_0_18393_inst_ack_0<= wack(0);
      rreq(0) <= W_count_17575_delayed_14_0_18393_inst_req_1;
      W_count_17575_delayed_14_0_18393_inst_ack_1<= rack(0);
      W_count_17575_delayed_14_0_18393_inst : InterlockBuffer generic map ( -- 
        name => "W_count_17575_delayed_14_0_18393_inst",
        buffer_size => 14,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => count_18327,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => count_17575_delayed_14_0_18395,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_pkt_pointer_17554_delayed_4_0_18362_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_pkt_pointer_17554_delayed_4_0_18362_inst_req_0;
      W_pkt_pointer_17554_delayed_4_0_18362_inst_ack_0<= wack(0);
      rreq(0) <= W_pkt_pointer_17554_delayed_4_0_18362_inst_req_1;
      W_pkt_pointer_17554_delayed_4_0_18362_inst_ack_1<= rack(0);
      W_pkt_pointer_17554_delayed_4_0_18362_inst : InterlockBuffer generic map ( -- 
        name => "W_pkt_pointer_17554_delayed_4_0_18362_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => pkt_pointer_18338,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pkt_pointer_17554_delayed_4_0_18364,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    ncount_18401_18331_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= ncount_18401_18331_buf_req_0;
      ncount_18401_18331_buf_ack_0<= wack(0);
      rreq(0) <= ncount_18401_18331_buf_req_1;
      ncount_18401_18331_buf_ack_1<= rack(0);
      ncount_18401_18331_buf : InterlockBuffer generic map ( -- 
        name => "ncount_18401_18331_buf",
        buffer_size => 2,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 32,
        out_data_width => 32,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ncount_18401,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ncount_18401_18331_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_18317
    process(AND_u6_u6_18326_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := AND_u6_u6_18326_wire(5 downto 0);
      tx_q_index_18317 <= tmp_var; -- 
    end process;
    -- interlock type_cast_18325_inst
    process(SUB_u32_u32_18324_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 5 downto 0) := SUB_u32_u32_18324_wire(5 downto 0);
      type_cast_18325_wire <= tmp_var; -- 
    end process;
    do_while_stmt_18315_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= BITSEL_u32_u1_18410_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_18315_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_18315_branch_req_0,
          ack0 => do_while_stmt_18315_branch_ack_0,
          ack1 => do_while_stmt_18315_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_18307_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_18311_wire;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_18307_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_18307_branch_req_0,
          ack0 => if_stmt_18307_branch_ack_0,
          ack1 => if_stmt_18307_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u32_u32_18391_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 14);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= count_18327;
      ADD_u32_u32_17574_17574_delayed_14_0_18392 <= data_out(31 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u32_u32_18391_inst_req_0;
      ADD_u32_u32_18391_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u32_u32_18391_inst_req_1;
      ADD_u32_u32_18391_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 32,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 32,
          constant_operand => "00000000000000000000000000000001",
          constant_width => 32,
          buffering  => 14,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- binary operator ADD_u6_u6_18321_inst
    process(RPIPE_LAST_READ_TX_QUEUE_INDEX_18319_wire) -- 
      variable tmp_var : std_logic_vector(5 downto 0); -- 
    begin -- 
      ApIntAdd_proc(RPIPE_LAST_READ_TX_QUEUE_INDEX_18319_wire, konst_18320_wire_constant, tmp_var);
      ADD_u6_u6_18321_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_18357_inst
    process(NOT_u1_u1_17543_17543_delayed_4_0_18353, transmitted_flag_18342) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_17543_17543_delayed_4_0_18353, transmitted_flag_18342, tmp_var);
      push_pointer_back_to_free_Q_18358 <= tmp_var; --
    end process;
    -- shared split operator group (3) : AND_u6_u6_18326_inst 
    ApIntAnd_group_3: Block -- 
      signal data_in: std_logic_vector(11 downto 0);
      signal data_out: std_logic_vector(5 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= ADD_u6_u6_18321_wire & type_cast_18325_wire;
      AND_u6_u6_18326_wire <= data_out(5 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u6_u6_18326_inst_req_0;
      AND_u6_u6_18326_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u6_u6_18326_inst_req_1;
      AND_u6_u6_18326_inst_ack_1 <= ackR_unguarded(0);
      ApIntAnd_group_3_gI: SplitGuardInterface generic map(name => "ApIntAnd_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 6,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 6, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 6,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- binary operator BITSEL_u32_u1_18310_inst
    process(RPIPE_CONTROL_REGISTER_18308_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_CONTROL_REGISTER_18308_wire, konst_18309_wire_constant, tmp_var);
      BITSEL_u32_u1_18310_wire <= tmp_var; --
    end process;
    -- binary operator BITSEL_u32_u1_18410_inst
    process(RPIPE_CONTROL_REGISTER_18408_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApBitsel_proc(RPIPE_CONTROL_REGISTER_18408_wire, konst_18409_wire_constant, tmp_var);
      BITSEL_u32_u1_18410_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_18311_inst
    process(BITSEL_u32_u1_18310_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", BITSEL_u32_u1_18310_wire, tmp_var);
      NOT_u1_u1_18311_wire <= tmp_var; -- 
    end process;
    -- shared split operator group (7) : NOT_u1_u1_18352_inst 
    ApIntNot_group_7: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 4);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= tx_flag_18338;
      NOT_u1_u1_17543_17543_delayed_4_0_18353 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= NOT_u1_u1_18352_inst_req_0;
      NOT_u1_u1_18352_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= NOT_u1_u1_18352_inst_req_1;
      NOT_u1_u1_18352_inst_ack_1 <= ackR_unguarded(0);
      ApIntNot_group_7_gI: SplitGuardInterface generic map(name => "ApIntNot_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntNot",
          name => "ApIntNot_group_7",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 4,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- binary operator SUB_u32_u32_18324_inst
    process(RPIPE_NUMBER_OF_SERVERS_18322_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApIntSub_proc(RPIPE_NUMBER_OF_SERVERS_18322_wire, konst_18323_wire_constant, tmp_var);
      SUB_u32_u32_18324_wire <= tmp_var; --
    end process;
    -- read from input-signal CONTROL_REGISTER
    RPIPE_CONTROL_REGISTER_18308_wire <= CONTROL_REGISTER;
    -- read from input-signal CONTROL_REGISTER
    RPIPE_CONTROL_REGISTER_18408_wire <= CONTROL_REGISTER;
    -- read from input-signal FREE_Q
    RPIPE_FREE_Q_18368_wire <= FREE_Q;
    -- read from input-signal LAST_READ_TX_QUEUE_INDEX
    RPIPE_LAST_READ_TX_QUEUE_INDEX_18319_wire <= LAST_READ_TX_QUEUE_INDEX;
    -- read from input-signal NUMBER_OF_SERVERS
    RPIPE_NUMBER_OF_SERVERS_18322_wire <= NUMBER_OF_SERVERS;
    -- shared outport operator group (0) : WPIPE_LAST_READ_TX_QUEUE_INDEX_18302_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_LAST_READ_TX_QUEUE_INDEX_18302_inst_req_0;
      WPIPE_LAST_READ_TX_QUEUE_INDEX_18302_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_LAST_READ_TX_QUEUE_INDEX_18302_inst_req_1;
      WPIPE_LAST_READ_TX_QUEUE_INDEX_18302_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= konst_18303_wire_constant;
      LAST_READ_TX_QUEUE_INDEX_write_0_gI: SplitGuardInterface generic map(name => "LAST_READ_TX_QUEUE_INDEX_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      LAST_READ_TX_QUEUE_INDEX_write_0: OutputPortRevised -- 
        generic map ( name => "LAST_READ_TX_QUEUE_INDEX", data_width => 6, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => LAST_READ_TX_QUEUE_INDEX_pipe_write_req(1),
          oack => LAST_READ_TX_QUEUE_INDEX_pipe_write_ack(1),
          odata => LAST_READ_TX_QUEUE_INDEX_pipe_write_data(11 downto 6),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_LAST_READ_TX_QUEUE_INDEX_18404_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_LAST_READ_TX_QUEUE_INDEX_18404_inst_req_0;
      WPIPE_LAST_READ_TX_QUEUE_INDEX_18404_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_LAST_READ_TX_QUEUE_INDEX_18404_inst_req_1;
      WPIPE_LAST_READ_TX_QUEUE_INDEX_18404_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= tx_q_index_18317;
      LAST_READ_TX_QUEUE_INDEX_write_1_gI: SplitGuardInterface generic map(name => "LAST_READ_TX_QUEUE_INDEX_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      LAST_READ_TX_QUEUE_INDEX_write_1: OutputPortRevised -- 
        generic map ( name => "LAST_READ_TX_QUEUE_INDEX", data_width => 6, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => LAST_READ_TX_QUEUE_INDEX_pipe_write_req(0),
          oack => LAST_READ_TX_QUEUE_INDEX_pipe_write_ack(0),
          odata => LAST_READ_TX_QUEUE_INDEX_pipe_write_data(5 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_18338_call 
    getTxPacketPointerFromServer_call_group_0: Block -- 
      signal data_in: std_logic_vector(5 downto 0);
      signal data_out: std_logic_vector(32 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 10);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_18338_call_req_0;
      call_stmt_18338_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_18338_call_req_1;
      call_stmt_18338_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      getTxPacketPointerFromServer_call_group_0_gI: SplitGuardInterface generic map(name => "getTxPacketPointerFromServer_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= tx_q_index_18317;
      pkt_pointer_18338 <= data_out(32 downto 1);
      tx_flag_18338 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 6,
        owidth => 6,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => getTxPacketPointerFromServer_call_reqs(0),
          ackR => getTxPacketPointerFromServer_call_acks(0),
          dataR => getTxPacketPointerFromServer_call_data(5 downto 0),
          tagR => getTxPacketPointerFromServer_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 33,
          owidth => 33,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => getTxPacketPointerFromServer_return_acks(0), -- cross-over
          ackL => getTxPacketPointerFromServer_return_reqs(0), -- cross-over
          dataL => getTxPacketPointerFromServer_return_data(32 downto 0),
          tagL => getTxPacketPointerFromServer_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_18342_call 
    transmitPacket_call_group_1: Block -- 
      signal data_in: std_logic_vector(31 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_18342_call_req_0;
      call_stmt_18342_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_18342_call_req_1;
      call_stmt_18342_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not tx_flag_18338(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      transmitPacket_call_group_1_gI: SplitGuardInterface generic map(name => "transmitPacket_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= pkt_pointer_18338;
      transmitted_flag_18342 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 32,
        owidth => 32,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => transmitPacket_call_reqs(0),
          ackR => transmitPacket_call_acks(0),
          dataR => transmitPacket_call_data(31 downto 0),
          tagR => transmitPacket_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => transmitPacket_return_acks(0), -- cross-over
          ackL => transmitPacket_return_reqs(0), -- cross-over
          dataL => transmitPacket_return_data(0 downto 0),
          tagL => transmitPacket_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_18371_call 
    pushIntoQueue_call_group_2: Block -- 
      signal data_in: std_logic_vector(68 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_18371_call_req_0;
      call_stmt_18371_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_18371_call_req_1;
      call_stmt_18371_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= push_pointer_back_to_free_Q_18358(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      pushIntoQueue_call_group_2_gI: SplitGuardInterface generic map(name => "pushIntoQueue_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_18367_wire_constant & RPIPE_FREE_Q_18368_wire & pkt_pointer_17554_delayed_4_0_18364;
      push_status_18371 <= data_out(0 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 69,
        owidth => 69,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => pushIntoQueue_call_reqs(0),
          ackR => pushIntoQueue_call_acks(0),
          dataR => pushIntoQueue_call_data(68 downto 0),
          tagR => pushIntoQueue_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 1,
          owidth => 1,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => pushIntoQueue_return_acks(0), -- cross-over
          ackL => pushIntoQueue_return_reqs(0), -- cross-over
          dataL => pushIntoQueue_return_data(0 downto 0),
          tagL => pushIntoQueue_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- shared call operator group (3) : call_stmt_18387_call 
    AccessRegister_call_group_3: Block -- 
      signal data_in: std_logic_vector(42 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_18387_call_req_0;
      call_stmt_18387_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_18387_call_req_1;
      call_stmt_18387_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= push_pointer_back_to_free_Q_18358(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      AccessRegister_call_group_3_gI: SplitGuardInterface generic map(name => "AccessRegister_call_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_18380_wire_constant & NOT_u4_u4_18383_wire_constant & konst_18384_wire_constant & count_17567_delayed_14_0_18377;
      ignore_resp_18387 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 43,
        owidth => 43,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => AccessRegister_call_reqs(0),
          ackR => AccessRegister_call_acks(0),
          dataR => AccessRegister_call_data(42 downto 0),
          tagR => AccessRegister_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => AccessRegister_return_acks(0), -- cross-over
          ackL => AccessRegister_return_reqs(0), -- cross-over
          dataL => AccessRegister_return_data(31 downto 0),
          tagL => AccessRegister_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 3
    -- 
  end Block; -- data_path
  -- 
end transmitEngineDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.nic_system_global_package.all;
entity transmitPacket is -- 
  generic (tag_length : integer); 
  port ( -- 
    packet_pointer : in  std_logic_vector(31 downto 0);
    status : out  std_logic_vector(0 downto 0);
    nic_to_mac_transmit_pipe_pipe_write_req : out  std_logic_vector(1 downto 0);
    nic_to_mac_transmit_pipe_pipe_write_ack : in   std_logic_vector(1 downto 0);
    nic_to_mac_transmit_pipe_pipe_write_data : out  std_logic_vector(145 downto 0);
    AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_call_data : out  std_logic_vector(42 downto 0);
    AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
    AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
    AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
    AccessRegister_return_data : in   std_logic_vector(31 downto 0);
    AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(1 downto 0);
    accessMemory_call_acks : in   std_logic_vector(1 downto 0);
    accessMemory_call_data : out  std_logic_vector(219 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(5 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(1 downto 0);
    accessMemory_return_acks : in   std_logic_vector(1 downto 0);
    accessMemory_return_data : in   std_logic_vector(127 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(5 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity transmitPacket;
architecture transmitPacket_arch of transmitPacket is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 32)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 1)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal packet_pointer_buffer :  std_logic_vector(31 downto 0);
  signal packet_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal status_buffer :  std_logic_vector(0 downto 0);
  signal status_update_enable: Boolean;
  signal transmitPacket_CP_36099_start: Boolean;
  signal transmitPacket_CP_36099_symbol: Boolean;
  -- volatile/operator module components. 
  component AccessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      register_index : in  std_logic_vector(5 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_18227_call_ack_0 : boolean;
  signal SUB_u11_u11_18209_inst_req_1 : boolean;
  signal call_stmt_18245_call_ack_0 : boolean;
  signal do_while_stmt_18203_branch_req_0 : boolean;
  signal call_stmt_18245_call_req_0 : boolean;
  signal call_stmt_18227_call_req_0 : boolean;
  signal do_while_stmt_18203_branch_ack_0 : boolean;
  signal ncount_down_18250_18210_buf_req_1 : boolean;
  signal CONCAT_u65_u73_18234_inst_req_0 : boolean;
  signal phi_stmt_18205_ack_0 : boolean;
  signal CONCAT_u65_u73_18234_inst_ack_1 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_18283_inst_ack_0 : boolean;
  signal phi_stmt_18211_req_1 : boolean;
  signal ncount_down_18250_18210_buf_ack_0 : boolean;
  signal call_stmt_18245_call_ack_1 : boolean;
  signal call_stmt_18245_call_req_1 : boolean;
  signal nmem_addr_18255_18216_buf_ack_1 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_18228_inst_ack_1 : boolean;
  signal ncount_down_18250_18210_buf_req_0 : boolean;
  signal CONCAT_u65_u73_18234_inst_req_1 : boolean;
  signal nmem_addr_18255_18216_buf_req_1 : boolean;
  signal CONCAT_u65_u73_18289_inst_ack_0 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_18283_inst_req_1 : boolean;
  signal EQ_u11_u1_18297_inst_req_0 : boolean;
  signal EQ_u11_u1_18297_inst_ack_0 : boolean;
  signal SUB_u11_u11_18209_inst_ack_0 : boolean;
  signal SUB_u11_u11_18209_inst_req_0 : boolean;
  signal SUB_u11_u11_18209_inst_ack_1 : boolean;
  signal CONCAT_u65_u73_18289_inst_req_0 : boolean;
  signal nmem_addr_18255_18216_buf_ack_0 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_18228_inst_req_1 : boolean;
  signal CONCAT_u65_u73_18234_inst_ack_0 : boolean;
  signal ncount_down_18250_18210_buf_ack_1 : boolean;
  signal phi_stmt_18205_req_1 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_18283_inst_ack_1 : boolean;
  signal do_while_stmt_18203_branch_ack_1 : boolean;
  signal ADD_u36_u36_18215_inst_req_1 : boolean;
  signal CONCAT_u65_u73_18289_inst_req_1 : boolean;
  signal ADD_u36_u36_18215_inst_ack_1 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_18228_inst_req_0 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_18228_inst_ack_0 : boolean;
  signal EQ_u11_u1_18297_inst_req_1 : boolean;
  signal call_stmt_18280_call_ack_1 : boolean;
  signal CONCAT_u65_u73_18289_inst_ack_1 : boolean;
  signal call_stmt_18280_call_ack_0 : boolean;
  signal call_stmt_18280_call_req_1 : boolean;
  signal call_stmt_18280_call_req_0 : boolean;
  signal WPIPE_nic_to_mac_transmit_pipe_18283_inst_req_0 : boolean;
  signal call_stmt_18190_call_req_1 : boolean;
  signal call_stmt_18227_call_req_1 : boolean;
  signal call_stmt_18190_call_ack_1 : boolean;
  signal ADD_u36_u36_18215_inst_req_0 : boolean;
  signal call_stmt_18227_call_ack_1 : boolean;
  signal EQ_u11_u1_18297_inst_ack_1 : boolean;
  signal phi_stmt_18205_req_0 : boolean;
  signal ADD_u36_u36_18215_inst_ack_0 : boolean;
  signal phi_stmt_18211_req_0 : boolean;
  signal call_stmt_18190_call_ack_0 : boolean;
  signal phi_stmt_18211_ack_0 : boolean;
  signal call_stmt_18190_call_req_0 : boolean;
  signal nmem_addr_18255_18216_buf_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "transmitPacket_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 32) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(31 downto 0) <= packet_pointer;
  packet_pointer_buffer <= in_buffer_data_out(31 downto 0);
  in_buffer_data_in(tag_length + 31 downto 32) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 31 downto 32);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  transmitPacket_CP_36099_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "transmitPacket_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 1) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(0 downto 0) <= status_buffer;
  status <= out_buffer_data_out(0 downto 0);
  out_buffer_data_in(tag_length + 0 downto 1) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 0 downto 1);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= transmitPacket_CP_36099_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= transmitPacket_CP_36099_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= transmitPacket_CP_36099_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  transmitPacket_CP_36099: Block -- control-path 
    signal transmitPacket_CP_36099_elements: BooleanArray(85 downto 0);
    -- 
  begin -- 
    transmitPacket_CP_36099_elements(0) <= transmitPacket_CP_36099_start;
    transmitPacket_CP_36099_symbol <= transmitPacket_CP_36099_elements(85);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 assign_stmt_18177_to_assign_stmt_18198/call_stmt_18190_update_start_
      -- CP-element group 0: 	 assign_stmt_18177_to_assign_stmt_18198/call_stmt_18190_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_18177_to_assign_stmt_18198/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_18177_to_assign_stmt_18198/call_stmt_18190_Update/$entry
      -- CP-element group 0: 	 assign_stmt_18177_to_assign_stmt_18198/call_stmt_18190_Update/ccr
      -- CP-element group 0: 	 assign_stmt_18177_to_assign_stmt_18198/call_stmt_18190_sample_start_
      -- CP-element group 0: 	 assign_stmt_18177_to_assign_stmt_18198/call_stmt_18190_Sample/crr
      -- 
    ccr_36117_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_36117_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_36099_elements(0), ack => call_stmt_18190_call_req_1); -- 
    crr_36112_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_36112_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_36099_elements(0), ack => call_stmt_18190_call_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_18177_to_assign_stmt_18198/call_stmt_18190_sample_completed_
      -- CP-element group 1: 	 assign_stmt_18177_to_assign_stmt_18198/call_stmt_18190_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_18177_to_assign_stmt_18198/call_stmt_18190_Sample/cra
      -- 
    cra_36113_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_18190_call_ack_0, ack => transmitPacket_CP_36099_elements(1)); -- 
    -- CP-element group 2:  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	4 
    -- CP-element group 2:  members (7) 
      -- CP-element group 2: 	 assign_stmt_18177_to_assign_stmt_18198/call_stmt_18190_update_completed_
      -- CP-element group 2: 	 assign_stmt_18177_to_assign_stmt_18198/$exit
      -- CP-element group 2: 	 branch_block_stmt_18202/do_while_stmt_18203__entry__
      -- CP-element group 2: 	 assign_stmt_18177_to_assign_stmt_18198/call_stmt_18190_Update/$exit
      -- CP-element group 2: 	 assign_stmt_18177_to_assign_stmt_18198/call_stmt_18190_Update/cca
      -- CP-element group 2: 	 branch_block_stmt_18202/branch_block_stmt_18202__entry__
      -- CP-element group 2: 	 branch_block_stmt_18202/$entry
      -- 
    cca_36118_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_18190_call_ack_1, ack => transmitPacket_CP_36099_elements(2)); -- 
    -- CP-element group 3:  fork  transition  place  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	76 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	77 
    -- CP-element group 3: 	78 
    -- CP-element group 3: 	80 
    -- CP-element group 3: 	83 
    -- CP-element group 3: 	84 
    -- CP-element group 3:  members (18) 
      -- CP-element group 3: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/call_stmt_18280_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/CONCAT_u65_u73_18289_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/EQ_u11_u1_18297_update_start_
      -- CP-element group 3: 	 branch_block_stmt_18202/do_while_stmt_18203__exit__
      -- CP-element group 3: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/EQ_u11_u1_18297_Sample/rr
      -- CP-element group 3: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/call_stmt_18280_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/CONCAT_u65_u73_18289_update_start_
      -- CP-element group 3: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/CONCAT_u65_u73_18289_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/EQ_u11_u1_18297_Update/cr
      -- CP-element group 3: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/EQ_u11_u1_18297_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/EQ_u11_u1_18297_Sample/$entry
      -- CP-element group 3: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/call_stmt_18280_Update/$entry
      -- CP-element group 3: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/call_stmt_18280_Update/ccr
      -- CP-element group 3: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/call_stmt_18280_Sample/crr
      -- CP-element group 3: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/EQ_u11_u1_18297_sample_start_
      -- CP-element group 3: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/$entry
      -- CP-element group 3: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/call_stmt_18280_update_start_
      -- CP-element group 3: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298__entry__
      -- 
    rr_36374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_36374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_36099_elements(3), ack => EQ_u11_u1_18297_inst_req_0); -- 
    cr_36351_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_36351_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_36099_elements(3), ack => CONCAT_u65_u73_18289_inst_req_1); -- 
    cr_36379_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_36379_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_36099_elements(3), ack => EQ_u11_u1_18297_inst_req_1); -- 
    ccr_36337_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_36337_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_36099_elements(3), ack => call_stmt_18280_call_req_1); -- 
    crr_36332_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_36332_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_36099_elements(3), ack => call_stmt_18280_call_req_0); -- 
    transmitPacket_CP_36099_elements(3) <= transmitPacket_CP_36099_elements(76);
    -- CP-element group 4:  transition  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	10 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203__entry__
      -- CP-element group 4: 	 branch_block_stmt_18202/do_while_stmt_18203/$entry
      -- 
    transmitPacket_CP_36099_elements(4) <= transmitPacket_CP_36099_elements(2);
    -- CP-element group 5:  merge  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	76 
    -- CP-element group 5:  members (1) 
      -- CP-element group 5: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203__exit__
      -- 
    -- Element group transmitPacket_CP_36099_elements(5) is bound as output of CP function.
    -- CP-element group 6:  merge  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_18202/do_while_stmt_18203/loop_back
      -- 
    -- Element group transmitPacket_CP_36099_elements(6) is bound as output of CP function.
    -- CP-element group 7:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	12 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	75 
    -- CP-element group 7: 	74 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_18202/do_while_stmt_18203/condition_done
      -- CP-element group 7: 	 branch_block_stmt_18202/do_while_stmt_18203/loop_exit/$entry
      -- CP-element group 7: 	 branch_block_stmt_18202/do_while_stmt_18203/loop_taken/$entry
      -- 
    transmitPacket_CP_36099_elements(7) <= transmitPacket_CP_36099_elements(12);
    -- CP-element group 8:  branch  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	73 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_18202/do_while_stmt_18203/loop_body_done
      -- 
    transmitPacket_CP_36099_elements(8) <= transmitPacket_CP_36099_elements(73);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	21 
    -- CP-element group 9: 	42 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/back_edge_to_loop_body
      -- 
    transmitPacket_CP_36099_elements(9) <= transmitPacket_CP_36099_elements(6);
    -- CP-element group 10:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	4 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	44 
    -- CP-element group 10: 	23 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/first_time_through_loop_body
      -- 
    transmitPacket_CP_36099_elements(10) <= transmitPacket_CP_36099_elements(4);
    -- CP-element group 11:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	17 
    -- CP-element group 11: 	18 
    -- CP-element group 11: 	36 
    -- CP-element group 11: 	37 
    -- CP-element group 11: 	72 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/loop_body_start
      -- CP-element group 11: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/$entry
      -- 
    -- Element group transmitPacket_CP_36099_elements(11) is bound as output of CP function.
    -- CP-element group 12:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	20 
    -- CP-element group 12: 	16 
    -- CP-element group 12: 	72 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	7 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/condition_evaluated
      -- 
    condition_evaluated_36142_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_36142_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_36099_elements(12), ack => do_while_stmt_18203_branch_req_0); -- 
    transmitPacket_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 31,2 => 31);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitPacket_CP_36099_elements(20) & transmitPacket_CP_36099_elements(16) & transmitPacket_CP_36099_elements(72);
      gj_transmitPacket_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_36099_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	17 
    -- CP-element group 13: 	36 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	16 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	38 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/phi_stmt_18205_sample_start__ps
      -- CP-element group 13: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/aggregated_phi_sample_req
      -- 
    transmitPacket_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 31,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitPacket_CP_36099_elements(17) & transmitPacket_CP_36099_elements(36) & transmitPacket_CP_36099_elements(16);
      gj_transmitPacket_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_36099_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	19 
    -- CP-element group 14: 	39 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	73 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	17 
    -- CP-element group 14: 	36 
    -- CP-element group 14:  members (3) 
      -- CP-element group 14: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/aggregated_phi_sample_ack
      -- CP-element group 14: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/phi_stmt_18211_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/phi_stmt_18205_sample_completed_
      -- 
    transmitPacket_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_36099_elements(19) & transmitPacket_CP_36099_elements(39);
      gj_transmitPacket_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_36099_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	18 
    -- CP-element group 15: 	37 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	40 
    -- CP-element group 15:  members (2) 
      -- CP-element group 15: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/aggregated_phi_update_req
      -- CP-element group 15: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/phi_stmt_18205_update_start__ps
      -- 
    transmitPacket_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_36099_elements(18) & transmitPacket_CP_36099_elements(37);
      gj_transmitPacket_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_36099_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	20 
    -- CP-element group 16: 	41 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	12 
    -- CP-element group 16: marked-successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/aggregated_phi_update_ack
      -- 
    transmitPacket_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 31);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_36099_elements(20) & transmitPacket_CP_36099_elements(41);
      gj_transmitPacket_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_36099_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	13 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/phi_stmt_18205_sample_start_
      -- 
    transmitPacket_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_36099_elements(11) & transmitPacket_CP_36099_elements(14);
      gj_transmitPacket_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_36099_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	11 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	20 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	15 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/phi_stmt_18205_update_start_
      -- 
    transmitPacket_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_36099_elements(11) & transmitPacket_CP_36099_elements(20);
      gj_transmitPacket_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_36099_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	14 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/phi_stmt_18205_sample_completed__ps
      -- 
    -- Element group transmitPacket_CP_36099_elements(19) is bound as output of CP function.
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	12 
    -- CP-element group 20: 	16 
    -- CP-element group 20: marked-successors 
    -- CP-element group 20: 	18 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/phi_stmt_18205_update_completed__ps
      -- CP-element group 20: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/phi_stmt_18205_update_completed_
      -- 
    -- Element group transmitPacket_CP_36099_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	9 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/phi_stmt_18205_loopback_trigger
      -- 
    transmitPacket_CP_36099_elements(21) <= transmitPacket_CP_36099_elements(9);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/phi_stmt_18205_loopback_sample_req
      -- CP-element group 22: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/phi_stmt_18205_loopback_sample_req_ps
      -- 
    phi_stmt_18205_loopback_sample_req_36157_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_18205_loopback_sample_req_36157_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_36099_elements(22), ack => phi_stmt_18205_req_1); -- 
    -- Element group transmitPacket_CP_36099_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	10 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/phi_stmt_18205_entry_trigger
      -- 
    transmitPacket_CP_36099_elements(23) <= transmitPacket_CP_36099_elements(10);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/phi_stmt_18205_entry_sample_req_ps
      -- CP-element group 24: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/phi_stmt_18205_entry_sample_req
      -- 
    phi_stmt_18205_entry_sample_req_36160_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_18205_entry_sample_req_36160_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_36099_elements(24), ack => phi_stmt_18205_req_0); -- 
    -- Element group transmitPacket_CP_36099_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/phi_stmt_18205_phi_mux_ack
      -- CP-element group 25: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/phi_stmt_18205_phi_mux_ack_ps
      -- 
    phi_stmt_18205_phi_mux_ack_36163_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_18205_ack_0, ack => transmitPacket_CP_36099_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/SUB_u11_u11_18209_sample_start__ps
      -- 
    -- Element group transmitPacket_CP_36099_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/SUB_u11_u11_18209_update_start__ps
      -- 
    -- Element group transmitPacket_CP_36099_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: marked-predecessors 
    -- CP-element group 28: 	30 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/SUB_u11_u11_18209_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/SUB_u11_u11_18209_Sample/rr
      -- CP-element group 28: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/SUB_u11_u11_18209_sample_start_
      -- 
    rr_36176_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_36176_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_36099_elements(28), ack => SUB_u11_u11_18209_inst_req_0); -- 
    transmitPacket_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_36099_elements(26) & transmitPacket_CP_36099_elements(30);
      gj_transmitPacket_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_36099_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: marked-predecessors 
    -- CP-element group 29: 	31 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/SUB_u11_u11_18209_Update/cr
      -- CP-element group 29: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/SUB_u11_u11_18209_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/SUB_u11_u11_18209_update_start_
      -- 
    cr_36181_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_36181_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_36099_elements(29), ack => SUB_u11_u11_18209_inst_req_1); -- 
    transmitPacket_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_36099_elements(27) & transmitPacket_CP_36099_elements(31);
      gj_transmitPacket_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_36099_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: marked-successors 
    -- CP-element group 30: 	28 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/SUB_u11_u11_18209_sample_completed__ps
      -- CP-element group 30: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/SUB_u11_u11_18209_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/SUB_u11_u11_18209_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/SUB_u11_u11_18209_sample_completed_
      -- 
    ra_36177_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u11_u11_18209_inst_ack_0, ack => transmitPacket_CP_36099_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: marked-successors 
    -- CP-element group 31: 	29 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/SUB_u11_u11_18209_update_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/SUB_u11_u11_18209_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/SUB_u11_u11_18209_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/SUB_u11_u11_18209_update_completed_
      -- 
    ca_36182_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => SUB_u11_u11_18209_inst_ack_1, ack => transmitPacket_CP_36099_elements(31)); -- 
    -- CP-element group 32:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/R_ncount_down_18210_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/R_ncount_down_18210_sample_start__ps
      -- CP-element group 32: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/R_ncount_down_18210_Sample/req
      -- CP-element group 32: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/R_ncount_down_18210_Sample/$entry
      -- 
    req_36194_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_36194_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_36099_elements(32), ack => ncount_down_18250_18210_buf_req_0); -- 
    -- Element group transmitPacket_CP_36099_elements(32) is bound as output of CP function.
    -- CP-element group 33:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/R_ncount_down_18210_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/R_ncount_down_18210_Update/req
      -- CP-element group 33: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/R_ncount_down_18210_update_start_
      -- CP-element group 33: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/R_ncount_down_18210_update_start__ps
      -- 
    req_36199_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_36199_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_36099_elements(33), ack => ncount_down_18250_18210_buf_req_1); -- 
    -- Element group transmitPacket_CP_36099_elements(33) is bound as output of CP function.
    -- CP-element group 34:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/R_ncount_down_18210_sample_completed_
      -- CP-element group 34: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/R_ncount_down_18210_Sample/ack
      -- CP-element group 34: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/R_ncount_down_18210_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/R_ncount_down_18210_sample_completed__ps
      -- 
    ack_36195_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ncount_down_18250_18210_buf_ack_0, ack => transmitPacket_CP_36099_elements(34)); -- 
    -- CP-element group 35:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/R_ncount_down_18210_Update/ack
      -- CP-element group 35: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/R_ncount_down_18210_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/R_ncount_down_18210_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/R_ncount_down_18210_update_completed__ps
      -- 
    ack_36200_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ncount_down_18250_18210_buf_ack_1, ack => transmitPacket_CP_36099_elements(35)); -- 
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	11 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	14 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	13 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/phi_stmt_18211_sample_start_
      -- 
    transmitPacket_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_36099_elements(11) & transmitPacket_CP_36099_elements(14);
      gj_transmitPacket_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_36099_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	11 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	70 
    -- CP-element group 37: 	41 
    -- CP-element group 37: 	59 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	15 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/phi_stmt_18211_update_start_
      -- 
    transmitPacket_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 31,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 1,2 => 1,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= transmitPacket_CP_36099_elements(11) & transmitPacket_CP_36099_elements(70) & transmitPacket_CP_36099_elements(41) & transmitPacket_CP_36099_elements(59);
      gj_transmitPacket_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_36099_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	13 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/phi_stmt_18211_sample_start__ps
      -- 
    transmitPacket_CP_36099_elements(38) <= transmitPacket_CP_36099_elements(13);
    -- CP-element group 39:  join  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	14 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/phi_stmt_18211_sample_completed__ps
      -- 
    -- Element group transmitPacket_CP_36099_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	15 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/phi_stmt_18211_update_start__ps
      -- 
    transmitPacket_CP_36099_elements(40) <= transmitPacket_CP_36099_elements(15);
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	68 
    -- CP-element group 41: 	16 
    -- CP-element group 41: 	57 
    -- CP-element group 41: marked-successors 
    -- CP-element group 41: 	37 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/phi_stmt_18211_update_completed_
      -- CP-element group 41: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/phi_stmt_18211_update_completed__ps
      -- 
    -- Element group transmitPacket_CP_36099_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	9 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/phi_stmt_18211_loopback_trigger
      -- 
    transmitPacket_CP_36099_elements(42) <= transmitPacket_CP_36099_elements(9);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/phi_stmt_18211_loopback_sample_req
      -- CP-element group 43: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/phi_stmt_18211_loopback_sample_req_ps
      -- 
    phi_stmt_18211_loopback_sample_req_36211_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_18211_loopback_sample_req_36211_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_36099_elements(43), ack => phi_stmt_18211_req_1); -- 
    -- Element group transmitPacket_CP_36099_elements(43) is bound as output of CP function.
    -- CP-element group 44:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	10 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/phi_stmt_18211_entry_trigger
      -- 
    transmitPacket_CP_36099_elements(44) <= transmitPacket_CP_36099_elements(10);
    -- CP-element group 45:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/phi_stmt_18211_entry_sample_req_ps
      -- CP-element group 45: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/phi_stmt_18211_entry_sample_req
      -- 
    phi_stmt_18211_entry_sample_req_36214_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_18211_entry_sample_req_36214_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_36099_elements(45), ack => phi_stmt_18211_req_0); -- 
    -- Element group transmitPacket_CP_36099_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/phi_stmt_18211_phi_mux_ack_ps
      -- CP-element group 46: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/phi_stmt_18211_phi_mux_ack
      -- 
    phi_stmt_18211_phi_mux_ack_36217_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_18211_ack_0, ack => transmitPacket_CP_36099_elements(46)); -- 
    -- CP-element group 47:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/ADD_u36_u36_18215_sample_start__ps
      -- 
    -- Element group transmitPacket_CP_36099_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/ADD_u36_u36_18215_update_start__ps
      -- 
    -- Element group transmitPacket_CP_36099_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: marked-predecessors 
    -- CP-element group 49: 	51 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/ADD_u36_u36_18215_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/ADD_u36_u36_18215_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/ADD_u36_u36_18215_Sample/rr
      -- 
    rr_36230_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_36230_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_36099_elements(49), ack => ADD_u36_u36_18215_inst_req_0); -- 
    transmitPacket_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_36099_elements(47) & transmitPacket_CP_36099_elements(51);
      gj_transmitPacket_cp_element_group_49 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_36099_elements(49), clk => clk, reset => reset); --
    end block;
    -- CP-element group 50:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: marked-predecessors 
    -- CP-element group 50: 	52 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/ADD_u36_u36_18215_Update/$entry
      -- CP-element group 50: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/ADD_u36_u36_18215_update_start_
      -- CP-element group 50: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/ADD_u36_u36_18215_Update/cr
      -- 
    cr_36235_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_36235_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_36099_elements(50), ack => ADD_u36_u36_18215_inst_req_1); -- 
    transmitPacket_cp_element_group_50: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_50"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_36099_elements(48) & transmitPacket_CP_36099_elements(52);
      gj_transmitPacket_cp_element_group_50 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_36099_elements(50), clk => clk, reset => reset); --
    end block;
    -- CP-element group 51:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: marked-successors 
    -- CP-element group 51: 	49 
    -- CP-element group 51:  members (4) 
      -- CP-element group 51: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/ADD_u36_u36_18215_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/ADD_u36_u36_18215_sample_completed__ps
      -- CP-element group 51: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/ADD_u36_u36_18215_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/ADD_u36_u36_18215_Sample/ra
      -- 
    ra_36231_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_18215_inst_ack_0, ack => transmitPacket_CP_36099_elements(51)); -- 
    -- CP-element group 52:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52: marked-successors 
    -- CP-element group 52: 	50 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/ADD_u36_u36_18215_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/ADD_u36_u36_18215_update_completed__ps
      -- CP-element group 52: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/ADD_u36_u36_18215_Update/ca
      -- CP-element group 52: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/ADD_u36_u36_18215_Update/$exit
      -- 
    ca_36236_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_18215_inst_ack_1, ack => transmitPacket_CP_36099_elements(52)); -- 
    -- CP-element group 53:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/R_nmem_addr_18216_sample_start_
      -- CP-element group 53: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/R_nmem_addr_18216_sample_start__ps
      -- CP-element group 53: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/R_nmem_addr_18216_Sample/$entry
      -- CP-element group 53: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/R_nmem_addr_18216_Sample/req
      -- 
    req_36248_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_36248_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_36099_elements(53), ack => nmem_addr_18255_18216_buf_req_0); -- 
    -- Element group transmitPacket_CP_36099_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/R_nmem_addr_18216_update_start_
      -- CP-element group 54: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/R_nmem_addr_18216_Update/req
      -- CP-element group 54: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/R_nmem_addr_18216_Update/$entry
      -- CP-element group 54: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/R_nmem_addr_18216_update_start__ps
      -- 
    req_36253_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_36253_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_36099_elements(54), ack => nmem_addr_18255_18216_buf_req_1); -- 
    -- Element group transmitPacket_CP_36099_elements(54) is bound as output of CP function.
    -- CP-element group 55:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55:  members (4) 
      -- CP-element group 55: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/R_nmem_addr_18216_sample_completed_
      -- CP-element group 55: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/R_nmem_addr_18216_sample_completed__ps
      -- CP-element group 55: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/R_nmem_addr_18216_Sample/ack
      -- CP-element group 55: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/R_nmem_addr_18216_Sample/$exit
      -- 
    ack_36249_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmem_addr_18255_18216_buf_ack_0, ack => transmitPacket_CP_36099_elements(55)); -- 
    -- CP-element group 56:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/R_nmem_addr_18216_update_completed__ps
      -- CP-element group 56: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/R_nmem_addr_18216_Update/ack
      -- CP-element group 56: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/R_nmem_addr_18216_Update/$exit
      -- CP-element group 56: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/R_nmem_addr_18216_update_completed_
      -- 
    ack_36254_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nmem_addr_18255_18216_buf_ack_1, ack => transmitPacket_CP_36099_elements(56)); -- 
    -- CP-element group 57:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	41 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	59 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/call_stmt_18227_Sample/crr
      -- CP-element group 57: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/call_stmt_18227_sample_start_
      -- CP-element group 57: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/call_stmt_18227_Sample/$entry
      -- 
    crr_36263_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_36263_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_36099_elements(57), ack => call_stmt_18227_call_req_0); -- 
    transmitPacket_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_36099_elements(41) & transmitPacket_CP_36099_elements(59);
      gj_transmitPacket_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_36099_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	63 
    -- CP-element group 58: 	60 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/call_stmt_18227_update_start_
      -- CP-element group 58: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/call_stmt_18227_Update/$entry
      -- CP-element group 58: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/call_stmt_18227_Update/ccr
      -- 
    ccr_36268_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_36268_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_36099_elements(58), ack => call_stmt_18227_call_req_1); -- 
    transmitPacket_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_36099_elements(63) & transmitPacket_CP_36099_elements(60);
      gj_transmitPacket_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_36099_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: marked-successors 
    -- CP-element group 59: 	37 
    -- CP-element group 59: 	57 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/call_stmt_18227_Sample/cra
      -- CP-element group 59: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/call_stmt_18227_sample_completed_
      -- CP-element group 59: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/call_stmt_18227_Sample/$exit
      -- 
    cra_36264_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_18227_call_ack_0, ack => transmitPacket_CP_36099_elements(59)); -- 
    -- CP-element group 60:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	61 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	58 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/call_stmt_18227_Update/$exit
      -- CP-element group 60: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/call_stmt_18227_update_completed_
      -- CP-element group 60: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/call_stmt_18227_Update/cca
      -- 
    cca_36269_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_18227_call_ack_1, ack => transmitPacket_CP_36099_elements(60)); -- 
    -- CP-element group 61:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	60 
    -- CP-element group 61: marked-predecessors 
    -- CP-element group 61: 	63 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/CONCAT_u65_u73_18234_Sample/rr
      -- CP-element group 61: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/CONCAT_u65_u73_18234_sample_start_
      -- CP-element group 61: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/CONCAT_u65_u73_18234_Sample/$entry
      -- 
    rr_36277_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_36277_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_36099_elements(61), ack => CONCAT_u65_u73_18234_inst_req_0); -- 
    transmitPacket_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_36099_elements(60) & transmitPacket_CP_36099_elements(63);
      gj_transmitPacket_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_36099_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: marked-predecessors 
    -- CP-element group 62: 	64 
    -- CP-element group 62: 	66 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	64 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/CONCAT_u65_u73_18234_update_start_
      -- CP-element group 62: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/CONCAT_u65_u73_18234_Update/cr
      -- CP-element group 62: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/CONCAT_u65_u73_18234_Update/$entry
      -- 
    cr_36282_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_36282_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_36099_elements(62), ack => CONCAT_u65_u73_18234_inst_req_1); -- 
    transmitPacket_cp_element_group_62: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_62"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_36099_elements(64) & transmitPacket_CP_36099_elements(66);
      gj_transmitPacket_cp_element_group_62 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_36099_elements(62), clk => clk, reset => reset); --
    end block;
    -- CP-element group 63:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: marked-successors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: 	58 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/CONCAT_u65_u73_18234_sample_completed_
      -- CP-element group 63: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/CONCAT_u65_u73_18234_Sample/$exit
      -- CP-element group 63: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/CONCAT_u65_u73_18234_Sample/ra
      -- 
    ra_36278_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u65_u73_18234_inst_ack_0, ack => transmitPacket_CP_36099_elements(63)); -- 
    -- CP-element group 64:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	62 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64: marked-successors 
    -- CP-element group 64: 	62 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/CONCAT_u65_u73_18234_update_completed_
      -- CP-element group 64: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/CONCAT_u65_u73_18234_Update/ca
      -- CP-element group 64: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/CONCAT_u65_u73_18234_Update/$exit
      -- 
    ca_36283_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u65_u73_18234_inst_ack_1, ack => transmitPacket_CP_36099_elements(64)); -- 
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	66 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/WPIPE_nic_to_mac_transmit_pipe_18228_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/WPIPE_nic_to_mac_transmit_pipe_18228_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/WPIPE_nic_to_mac_transmit_pipe_18228_Sample/req
      -- 
    req_36291_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_36291_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_36099_elements(65), ack => WPIPE_nic_to_mac_transmit_pipe_18228_inst_req_0); -- 
    transmitPacket_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_36099_elements(64) & transmitPacket_CP_36099_elements(67);
      gj_transmitPacket_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_36099_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	65 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	67 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	62 
    -- CP-element group 66:  members (6) 
      -- CP-element group 66: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/WPIPE_nic_to_mac_transmit_pipe_18228_sample_completed_
      -- CP-element group 66: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/WPIPE_nic_to_mac_transmit_pipe_18228_update_start_
      -- CP-element group 66: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/WPIPE_nic_to_mac_transmit_pipe_18228_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/WPIPE_nic_to_mac_transmit_pipe_18228_Update/req
      -- CP-element group 66: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/WPIPE_nic_to_mac_transmit_pipe_18228_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/WPIPE_nic_to_mac_transmit_pipe_18228_Update/$entry
      -- 
    ack_36292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_to_mac_transmit_pipe_18228_inst_ack_0, ack => transmitPacket_CP_36099_elements(66)); -- 
    req_36296_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_36296_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_36099_elements(66), ack => WPIPE_nic_to_mac_transmit_pipe_18228_inst_req_1); -- 
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	66 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	73 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	65 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/WPIPE_nic_to_mac_transmit_pipe_18228_update_completed_
      -- CP-element group 67: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/WPIPE_nic_to_mac_transmit_pipe_18228_Update/ack
      -- CP-element group 67: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/WPIPE_nic_to_mac_transmit_pipe_18228_Update/$exit
      -- 
    ack_36297_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_to_mac_transmit_pipe_18228_inst_ack_1, ack => transmitPacket_CP_36099_elements(67)); -- 
    -- CP-element group 68:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	41 
    -- CP-element group 68: marked-predecessors 
    -- CP-element group 68: 	70 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/call_stmt_18245_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/call_stmt_18245_Sample/crr
      -- CP-element group 68: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/call_stmt_18245_sample_start_
      -- 
    crr_36305_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_36305_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_36099_elements(68), ack => call_stmt_18245_call_req_0); -- 
    transmitPacket_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 31,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_36099_elements(41) & transmitPacket_CP_36099_elements(70);
      gj_transmitPacket_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_36099_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: marked-predecessors 
    -- CP-element group 69: 	71 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/call_stmt_18245_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/call_stmt_18245_Update/ccr
      -- CP-element group 69: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/call_stmt_18245_update_start_
      -- 
    ccr_36310_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_36310_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_36099_elements(69), ack => call_stmt_18245_call_req_1); -- 
    transmitPacket_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= transmitPacket_CP_36099_elements(71);
      gj_transmitPacket_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_36099_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: marked-successors 
    -- CP-element group 70: 	37 
    -- CP-element group 70: 	68 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/call_stmt_18245_Sample/cra
      -- CP-element group 70: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/call_stmt_18245_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/call_stmt_18245_sample_completed_
      -- 
    cra_36306_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_18245_call_ack_0, ack => transmitPacket_CP_36099_elements(70)); -- 
    -- CP-element group 71:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	73 
    -- CP-element group 71: marked-successors 
    -- CP-element group 71: 	69 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/call_stmt_18245_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/call_stmt_18245_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/call_stmt_18245_Update/cca
      -- 
    cca_36311_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_18245_call_ack_1, ack => transmitPacket_CP_36099_elements(71)); -- 
    -- CP-element group 72:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	11 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	12 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group transmitPacket_CP_36099_elements(72) is a control-delay.
    cp_element_72_delay: control_delay_element  generic map(name => " 72_delay", delay_value => 1)  port map(req => transmitPacket_CP_36099_elements(11), ack => transmitPacket_CP_36099_elements(72), clk => clk, reset =>reset);
    -- CP-element group 73:  join  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	67 
    -- CP-element group 73: 	14 
    -- CP-element group 73: 	71 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	8 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_18202/do_while_stmt_18203/do_while_stmt_18203_loop_body/$exit
      -- 
    transmitPacket_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 31,1 => 31,2 => 31);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= transmitPacket_CP_36099_elements(67) & transmitPacket_CP_36099_elements(14) & transmitPacket_CP_36099_elements(71);
      gj_transmitPacket_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_36099_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	7 
    -- CP-element group 74: successors 
    -- CP-element group 74:  members (2) 
      -- CP-element group 74: 	 branch_block_stmt_18202/do_while_stmt_18203/loop_exit/ack
      -- CP-element group 74: 	 branch_block_stmt_18202/do_while_stmt_18203/loop_exit/$exit
      -- 
    ack_36316_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_18203_branch_ack_0, ack => transmitPacket_CP_36099_elements(74)); -- 
    -- CP-element group 75:  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	7 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (2) 
      -- CP-element group 75: 	 branch_block_stmt_18202/do_while_stmt_18203/loop_taken/ack
      -- CP-element group 75: 	 branch_block_stmt_18202/do_while_stmt_18203/loop_taken/$exit
      -- 
    ack_36320_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_18203_branch_ack_1, ack => transmitPacket_CP_36099_elements(75)); -- 
    -- CP-element group 76:  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	5 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	3 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_18202/do_while_stmt_18203/$exit
      -- 
    transmitPacket_CP_36099_elements(76) <= transmitPacket_CP_36099_elements(5);
    -- CP-element group 77:  transition  input  bypass 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	3 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/call_stmt_18280_Sample/$exit
      -- CP-element group 77: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/call_stmt_18280_Sample/cra
      -- CP-element group 77: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/call_stmt_18280_sample_completed_
      -- 
    cra_36333_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 77_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_18280_call_ack_0, ack => transmitPacket_CP_36099_elements(77)); -- 
    -- CP-element group 78:  transition  input  output  bypass 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	3 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78:  members (6) 
      -- CP-element group 78: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/CONCAT_u65_u73_18289_Sample/$entry
      -- CP-element group 78: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/call_stmt_18280_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/CONCAT_u65_u73_18289_Sample/rr
      -- CP-element group 78: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/call_stmt_18280_Update/cca
      -- CP-element group 78: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/CONCAT_u65_u73_18289_sample_start_
      -- CP-element group 78: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/call_stmt_18280_Update/$exit
      -- 
    cca_36338_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_18280_call_ack_1, ack => transmitPacket_CP_36099_elements(78)); -- 
    rr_36346_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_36346_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_36099_elements(78), ack => CONCAT_u65_u73_18289_inst_req_0); -- 
    -- CP-element group 79:  transition  input  bypass 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/CONCAT_u65_u73_18289_Sample/$exit
      -- CP-element group 79: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/CONCAT_u65_u73_18289_Sample/ra
      -- CP-element group 79: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/CONCAT_u65_u73_18289_sample_completed_
      -- 
    ra_36347_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u65_u73_18289_inst_ack_0, ack => transmitPacket_CP_36099_elements(79)); -- 
    -- CP-element group 80:  transition  input  output  bypass 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	3 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (6) 
      -- CP-element group 80: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/WPIPE_nic_to_mac_transmit_pipe_18283_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/CONCAT_u65_u73_18289_Update/$exit
      -- CP-element group 80: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/WPIPE_nic_to_mac_transmit_pipe_18283_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/CONCAT_u65_u73_18289_Update/ca
      -- CP-element group 80: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/WPIPE_nic_to_mac_transmit_pipe_18283_Sample/req
      -- CP-element group 80: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/CONCAT_u65_u73_18289_update_completed_
      -- 
    ca_36352_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 80_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u65_u73_18289_inst_ack_1, ack => transmitPacket_CP_36099_elements(80)); -- 
    req_36360_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_36360_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_36099_elements(80), ack => WPIPE_nic_to_mac_transmit_pipe_18283_inst_req_0); -- 
    -- CP-element group 81:  transition  input  output  bypass 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81:  members (6) 
      -- CP-element group 81: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/WPIPE_nic_to_mac_transmit_pipe_18283_update_start_
      -- CP-element group 81: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/WPIPE_nic_to_mac_transmit_pipe_18283_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/WPIPE_nic_to_mac_transmit_pipe_18283_Sample/ack
      -- CP-element group 81: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/WPIPE_nic_to_mac_transmit_pipe_18283_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/WPIPE_nic_to_mac_transmit_pipe_18283_Update/req
      -- CP-element group 81: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/WPIPE_nic_to_mac_transmit_pipe_18283_Update/$entry
      -- 
    ack_36361_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_to_mac_transmit_pipe_18283_inst_ack_0, ack => transmitPacket_CP_36099_elements(81)); -- 
    req_36365_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_36365_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => transmitPacket_CP_36099_elements(81), ack => WPIPE_nic_to_mac_transmit_pipe_18283_inst_req_1); -- 
    -- CP-element group 82:  transition  input  bypass 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	85 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/WPIPE_nic_to_mac_transmit_pipe_18283_Update/ack
      -- CP-element group 82: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/WPIPE_nic_to_mac_transmit_pipe_18283_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/WPIPE_nic_to_mac_transmit_pipe_18283_update_completed_
      -- 
    ack_36366_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_nic_to_mac_transmit_pipe_18283_inst_ack_1, ack => transmitPacket_CP_36099_elements(82)); -- 
    -- CP-element group 83:  transition  input  bypass 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	3 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/EQ_u11_u1_18297_sample_completed_
      -- CP-element group 83: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/EQ_u11_u1_18297_Sample/ra
      -- CP-element group 83: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/EQ_u11_u1_18297_Sample/$exit
      -- 
    ra_36375_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u11_u1_18297_inst_ack_0, ack => transmitPacket_CP_36099_elements(83)); -- 
    -- CP-element group 84:  transition  input  bypass 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	3 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	85 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/EQ_u11_u1_18297_Update/$exit
      -- CP-element group 84: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/EQ_u11_u1_18297_update_completed_
      -- CP-element group 84: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/EQ_u11_u1_18297_Update/ca
      -- 
    ca_36380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 84_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => EQ_u11_u1_18297_inst_ack_1, ack => transmitPacket_CP_36099_elements(84)); -- 
    -- CP-element group 85:  join  transition  place  bypass 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	82 
    -- CP-element group 85: 	84 
    -- CP-element group 85: successors 
    -- CP-element group 85:  members (5) 
      -- CP-element group 85: 	 $exit
      -- CP-element group 85: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298__exit__
      -- CP-element group 85: 	 branch_block_stmt_18202/branch_block_stmt_18202__exit__
      -- CP-element group 85: 	 branch_block_stmt_18202/$exit
      -- CP-element group 85: 	 branch_block_stmt_18202/call_stmt_18280_to_assign_stmt_18298/$exit
      -- 
    transmitPacket_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "transmitPacket_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= transmitPacket_CP_36099_elements(82) & transmitPacket_CP_36099_elements(84);
      gj_transmitPacket_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => transmitPacket_CP_36099_elements(85), clk => clk, reset => reset); --
    end block;
    transmitPacket_do_while_stmt_18203_terminator_36321: loop_terminator -- 
      generic map (name => " transmitPacket_do_while_stmt_18203_terminator_36321", max_iterations_in_flight =>31) 
      port map(loop_body_exit => transmitPacket_CP_36099_elements(8),loop_continue => transmitPacket_CP_36099_elements(75),loop_terminate => transmitPacket_CP_36099_elements(74),loop_back => transmitPacket_CP_36099_elements(6),loop_exit => transmitPacket_CP_36099_elements(5),clk => clk, reset => reset); -- 
    phi_stmt_18205_phi_seq_36201_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= transmitPacket_CP_36099_elements(23);
      transmitPacket_CP_36099_elements(26)<= src_sample_reqs(0);
      src_sample_acks(0)  <= transmitPacket_CP_36099_elements(30);
      transmitPacket_CP_36099_elements(27)<= src_update_reqs(0);
      src_update_acks(0)  <= transmitPacket_CP_36099_elements(31);
      transmitPacket_CP_36099_elements(24) <= phi_mux_reqs(0);
      triggers(1)  <= transmitPacket_CP_36099_elements(21);
      transmitPacket_CP_36099_elements(32)<= src_sample_reqs(1);
      src_sample_acks(1)  <= transmitPacket_CP_36099_elements(34);
      transmitPacket_CP_36099_elements(33)<= src_update_reqs(1);
      src_update_acks(1)  <= transmitPacket_CP_36099_elements(35);
      transmitPacket_CP_36099_elements(22) <= phi_mux_reqs(1);
      phi_stmt_18205_phi_seq_36201 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_18205_phi_seq_36201") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => transmitPacket_CP_36099_elements(13), 
          phi_sample_ack => transmitPacket_CP_36099_elements(19), 
          phi_update_req => transmitPacket_CP_36099_elements(15), 
          phi_update_ack => transmitPacket_CP_36099_elements(20), 
          phi_mux_ack => transmitPacket_CP_36099_elements(25), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_18211_phi_seq_36255_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= transmitPacket_CP_36099_elements(44);
      transmitPacket_CP_36099_elements(47)<= src_sample_reqs(0);
      src_sample_acks(0)  <= transmitPacket_CP_36099_elements(51);
      transmitPacket_CP_36099_elements(48)<= src_update_reqs(0);
      src_update_acks(0)  <= transmitPacket_CP_36099_elements(52);
      transmitPacket_CP_36099_elements(45) <= phi_mux_reqs(0);
      triggers(1)  <= transmitPacket_CP_36099_elements(42);
      transmitPacket_CP_36099_elements(53)<= src_sample_reqs(1);
      src_sample_acks(1)  <= transmitPacket_CP_36099_elements(55);
      transmitPacket_CP_36099_elements(54)<= src_update_reqs(1);
      src_update_acks(1)  <= transmitPacket_CP_36099_elements(56);
      transmitPacket_CP_36099_elements(43) <= phi_mux_reqs(1);
      phi_stmt_18211_phi_seq_36255 : phi_sequencer_v2-- 
        generic map (place_capacity => 31, ntriggers => 2, name => "phi_stmt_18211_phi_seq_36255") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => transmitPacket_CP_36099_elements(38), 
          phi_sample_ack => transmitPacket_CP_36099_elements(39), 
          phi_update_req => transmitPacket_CP_36099_elements(40), 
          phi_update_ack => transmitPacket_CP_36099_elements(41), 
          phi_mux_ack => transmitPacket_CP_36099_elements(46), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_36143_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= transmitPacket_CP_36099_elements(9);
        preds(1)  <= transmitPacket_CP_36099_elements(10);
        entry_tmerge_36143 : transition_merge -- 
          generic map(name => " entry_tmerge_36143")
          port map (preds => preds, symbol_out => transmitPacket_CP_36099_elements(11));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u36_u36_18215_wire : std_logic_vector(35 downto 0);
    signal CONCAT_u1_u65_18232_wire : std_logic_vector(64 downto 0);
    signal CONCAT_u1_u65_18287_wire : std_logic_vector(64 downto 0);
    signal CONCAT_u65_u73_18234_wire : std_logic_vector(72 downto 0);
    signal CONCAT_u65_u73_18289_wire : std_logic_vector(72 downto 0);
    signal NOT_u4_u4_18240_wire_constant : std_logic_vector(3 downto 0);
    signal R_FULL_BYTE_MASK_18185_wire_constant : std_logic_vector(7 downto 0);
    signal R_FULL_BYTE_MASK_18222_wire_constant : std_logic_vector(7 downto 0);
    signal R_FULL_BYTE_MASK_18233_wire_constant : std_logic_vector(7 downto 0);
    signal R_FULL_BYTE_MASK_18275_wire_constant : std_logic_vector(7 downto 0);
    signal SUB_u11_u11_18209_wire : std_logic_vector(10 downto 0);
    signal SUB_u36_u36_18295_wire : std_logic_vector(35 downto 0);
    signal control_data_18190 : std_logic_vector(63 downto 0);
    signal control_data_addr_18177 : std_logic_vector(35 downto 0);
    signal count_down_18205 : std_logic_vector(10 downto 0);
    signal data_18227 : std_logic_vector(63 downto 0);
    signal ignore_resp5_18245 : std_logic_vector(31 downto 0);
    signal konst_18208_wire_constant : std_logic_vector(10 downto 0);
    signal konst_18214_wire_constant : std_logic_vector(35 downto 0);
    signal konst_18241_wire_constant : std_logic_vector(5 downto 0);
    signal konst_18248_wire_constant : std_logic_vector(10 downto 0);
    signal konst_18253_wire_constant : std_logic_vector(35 downto 0);
    signal konst_18264_wire_constant : std_logic_vector(10 downto 0);
    signal last_tkeep_18198 : std_logic_vector(7 downto 0);
    signal last_word_18280 : std_logic_vector(63 downto 0);
    signal mem_addr_18211 : std_logic_vector(35 downto 0);
    signal ncount_down_18250 : std_logic_vector(10 downto 0);
    signal ncount_down_18250_18210_buffered : std_logic_vector(10 downto 0);
    signal nmem_addr_18255 : std_logic_vector(35 downto 0);
    signal nmem_addr_18255_18216_buffered : std_logic_vector(35 downto 0);
    signal not_last_word_18266 : std_logic_vector(0 downto 0);
    signal packet_size_18194 : std_logic_vector(10 downto 0);
    signal slice_18243_wire : std_logic_vector(31 downto 0);
    signal type_cast_18182_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_18184_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_18188_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_18219_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_18221_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_18225_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_18230_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_18237_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_18272_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_18274_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_18278_wire_constant : std_logic_vector(63 downto 0);
    signal type_cast_18285_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_18296_wire : std_logic_vector(10 downto 0);
    -- 
  begin -- 
    NOT_u4_u4_18240_wire_constant <= "1111";
    R_FULL_BYTE_MASK_18185_wire_constant <= "11111111";
    R_FULL_BYTE_MASK_18222_wire_constant <= "11111111";
    R_FULL_BYTE_MASK_18233_wire_constant <= "11111111";
    R_FULL_BYTE_MASK_18275_wire_constant <= "11111111";
    konst_18208_wire_constant <= "00000010000";
    konst_18214_wire_constant <= "000000000000000000000000000000011000";
    konst_18241_wire_constant <= "110101";
    konst_18248_wire_constant <= "00000001000";
    konst_18253_wire_constant <= "000000000000000000000000000000001000";
    konst_18264_wire_constant <= "00000001000";
    type_cast_18182_wire_constant <= "0";
    type_cast_18184_wire_constant <= "1";
    type_cast_18188_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_18219_wire_constant <= "0";
    type_cast_18221_wire_constant <= "1";
    type_cast_18225_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_18230_wire_constant <= "0";
    type_cast_18237_wire_constant <= "0";
    type_cast_18272_wire_constant <= "0";
    type_cast_18274_wire_constant <= "1";
    type_cast_18278_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    type_cast_18285_wire_constant <= "1";
    phi_stmt_18205: Block -- phi operator 
      signal idata: std_logic_vector(21 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= SUB_u11_u11_18209_wire & ncount_down_18250_18210_buffered;
      req <= phi_stmt_18205_req_0 & phi_stmt_18205_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_18205",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 11) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_18205_ack_0,
          idata => idata,
          odata => count_down_18205,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_18205
    phi_stmt_18211: Block -- phi operator 
      signal idata: std_logic_vector(71 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= ADD_u36_u36_18215_wire & nmem_addr_18255_18216_buffered;
      req <= phi_stmt_18211_req_0 & phi_stmt_18211_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_18211",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 36) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_18211_ack_0,
          idata => idata,
          odata => mem_addr_18211,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_18211
    -- flow-through slice operator slice_18193_inst
    packet_size_18194 <= control_data_18190(18 downto 8);
    -- flow-through slice operator slice_18197_inst
    last_tkeep_18198 <= control_data_18190(7 downto 0);
    -- flow-through slice operator slice_18243_inst
    slice_18243_wire <= mem_addr_18211(31 downto 0);
    ncount_down_18250_18210_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= ncount_down_18250_18210_buf_req_0;
      ncount_down_18250_18210_buf_ack_0<= wack(0);
      rreq(0) <= ncount_down_18250_18210_buf_req_1;
      ncount_down_18250_18210_buf_ack_1<= rack(0);
      ncount_down_18250_18210_buf : InterlockBuffer generic map ( -- 
        name => "ncount_down_18250_18210_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 11,
        out_data_width => 11,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => ncount_down_18250,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => ncount_down_18250_18210_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nmem_addr_18255_18216_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nmem_addr_18255_18216_buf_req_0;
      nmem_addr_18255_18216_buf_ack_0<= wack(0);
      rreq(0) <= nmem_addr_18255_18216_buf_req_1;
      nmem_addr_18255_18216_buf_ack_1<= rack(0);
      nmem_addr_18255_18216_buf : InterlockBuffer generic map ( -- 
        name => "nmem_addr_18255_18216_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nmem_addr_18255,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nmem_addr_18255_18216_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock type_cast_18176_inst
    process(packet_pointer_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 31 downto 0) := packet_pointer_buffer(31 downto 0);
      control_data_addr_18177 <= tmp_var; -- 
    end process;
    -- interlock type_cast_18296_inst
    process(SUB_u36_u36_18295_wire) -- 
      variable tmp_var : std_logic_vector(10 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 10 downto 0) := SUB_u36_u36_18295_wire(10 downto 0);
      type_cast_18296_wire <= tmp_var; -- 
    end process;
    do_while_stmt_18203_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= not_last_word_18266;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_18203_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_18203_branch_req_0,
          ack0 => do_while_stmt_18203_branch_ack_0,
          ack1 => do_while_stmt_18203_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u36_u36_18215_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= control_data_addr_18177;
      ADD_u36_u36_18215_wire <= data_out(35 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u36_u36_18215_inst_req_0;
      ADD_u36_u36_18215_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u36_u36_18215_inst_req_1;
      ADD_u36_u36_18215_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 36,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 36,
          constant_operand => "000000000000000000000000000000011000",
          constant_width => 36,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- binary operator ADD_u36_u36_18254_inst
    process(mem_addr_18211) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(mem_addr_18211, konst_18253_wire_constant, tmp_var);
      nmem_addr_18255 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u65_18232_inst
    process(type_cast_18230_wire_constant, data_18227) -- 
      variable tmp_var : std_logic_vector(64 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_18230_wire_constant, data_18227, tmp_var);
      CONCAT_u1_u65_18232_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u65_18287_inst
    process(type_cast_18285_wire_constant, last_word_18280) -- 
      variable tmp_var : std_logic_vector(64 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_18285_wire_constant, last_word_18280, tmp_var);
      CONCAT_u1_u65_18287_wire <= tmp_var; --
    end process;
    -- shared split operator group (4) : CONCAT_u65_u73_18234_inst 
    ApConcat_group_4: Block -- 
      signal data_in: std_logic_vector(64 downto 0);
      signal data_out: std_logic_vector(72 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u1_u65_18232_wire;
      CONCAT_u65_u73_18234_wire <= data_out(72 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u65_u73_18234_inst_req_0;
      CONCAT_u65_u73_18234_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u65_u73_18234_inst_req_1;
      CONCAT_u65_u73_18234_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_4_gI: SplitGuardInterface generic map(name => "ApConcat_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_4",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 65,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 73,
          constant_operand => "11111111",
          constant_width => 8,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- shared split operator group (5) : CONCAT_u65_u73_18289_inst 
    ApConcat_group_5: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal data_out: std_logic_vector(72 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u1_u65_18287_wire & last_tkeep_18198;
      CONCAT_u65_u73_18289_wire <= data_out(72 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u65_u73_18289_inst_req_0;
      CONCAT_u65_u73_18289_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u65_u73_18289_inst_req_1;
      CONCAT_u65_u73_18289_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_5_gI: SplitGuardInterface generic map(name => "ApConcat_group_5_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_5",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 65,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 8, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 73,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 5
    -- shared split operator group (6) : EQ_u11_u1_18297_inst 
    ApIntEq_group_6: Block -- 
      signal data_in: std_logic_vector(21 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= packet_size_18194 & type_cast_18296_wire;
      status_buffer <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= EQ_u11_u1_18297_inst_req_0;
      EQ_u11_u1_18297_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= EQ_u11_u1_18297_inst_req_1;
      EQ_u11_u1_18297_inst_ack_1 <= ackR_unguarded(0);
      ApIntEq_group_6_gI: SplitGuardInterface generic map(name => "ApIntEq_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntEq",
          name => "ApIntEq_group_6",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 11, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- shared split operator group (7) : SUB_u11_u11_18209_inst 
    ApIntSub_group_7: Block -- 
      signal data_in: std_logic_vector(10 downto 0);
      signal data_out: std_logic_vector(10 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= packet_size_18194;
      SUB_u11_u11_18209_wire <= data_out(10 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= SUB_u11_u11_18209_inst_req_0;
      SUB_u11_u11_18209_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= SUB_u11_u11_18209_inst_req_1;
      SUB_u11_u11_18209_inst_ack_1 <= ackR_unguarded(0);
      ApIntSub_group_7_gI: SplitGuardInterface generic map(name => "ApIntSub_group_7_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntSub",
          name => "ApIntSub_group_7",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 11,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 11,
          constant_operand => "00000010000",
          constant_width => 11,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 7
    -- binary operator SUB_u11_u11_18249_inst
    process(count_down_18205) -- 
      variable tmp_var : std_logic_vector(10 downto 0); -- 
    begin -- 
      ApIntSub_proc(count_down_18205, konst_18248_wire_constant, tmp_var);
      ncount_down_18250 <= tmp_var; --
    end process;
    -- binary operator SUB_u36_u36_18295_inst
    process(nmem_addr_18255, control_data_addr_18177) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntSub_proc(nmem_addr_18255, control_data_addr_18177, tmp_var);
      SUB_u36_u36_18295_wire <= tmp_var; --
    end process;
    -- binary operator UGT_u11_u1_18265_inst
    process(ncount_down_18250) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUgt_proc(ncount_down_18250, konst_18264_wire_constant, tmp_var);
      not_last_word_18266 <= tmp_var; --
    end process;
    -- shared outport operator group (0) : WPIPE_nic_to_mac_transmit_pipe_18228_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_nic_to_mac_transmit_pipe_18228_inst_req_0;
      WPIPE_nic_to_mac_transmit_pipe_18228_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_nic_to_mac_transmit_pipe_18228_inst_req_1;
      WPIPE_nic_to_mac_transmit_pipe_18228_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= CONCAT_u65_u73_18234_wire;
      nic_to_mac_transmit_pipe_write_0_gI: SplitGuardInterface generic map(name => "nic_to_mac_transmit_pipe_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      nic_to_mac_transmit_pipe_write_0: OutputPortRevised -- 
        generic map ( name => "nic_to_mac_transmit_pipe", data_width => 73, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => nic_to_mac_transmit_pipe_pipe_write_req(1),
          oack => nic_to_mac_transmit_pipe_pipe_write_ack(1),
          odata => nic_to_mac_transmit_pipe_pipe_write_data(145 downto 73),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_nic_to_mac_transmit_pipe_18283_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(72 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_nic_to_mac_transmit_pipe_18283_inst_req_0;
      WPIPE_nic_to_mac_transmit_pipe_18283_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_nic_to_mac_transmit_pipe_18283_inst_req_1;
      WPIPE_nic_to_mac_transmit_pipe_18283_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= CONCAT_u65_u73_18289_wire;
      nic_to_mac_transmit_pipe_write_1_gI: SplitGuardInterface generic map(name => "nic_to_mac_transmit_pipe_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      nic_to_mac_transmit_pipe_write_1: OutputPortRevised -- 
        generic map ( name => "nic_to_mac_transmit_pipe", data_width => 73, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => nic_to_mac_transmit_pipe_pipe_write_req(0),
          oack => nic_to_mac_transmit_pipe_pipe_write_ack(0),
          odata => nic_to_mac_transmit_pipe_pipe_write_data(72 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared call operator group (0) : call_stmt_18190_call call_stmt_18280_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(219 downto 0);
      signal data_out: std_logic_vector(127 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 1 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 1 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 1 downto 0);
      signal guard_vector : std_logic_vector( 1 downto 0);
      constant inBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant outBUFs : IntegerArray(1 downto 0) := (1 => 1, 0 => 1);
      constant guardFlags : BooleanArray(1 downto 0) := (0 => false, 1 => false);
      constant guardBuffering: IntegerArray(1 downto 0)  := (0 => 2, 1 => 2);
      -- 
    begin -- 
      reqL_unguarded(1) <= call_stmt_18190_call_req_0;
      reqL_unguarded(0) <= call_stmt_18280_call_req_0;
      call_stmt_18190_call_ack_0 <= ackL_unguarded(1);
      call_stmt_18280_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(1) <= call_stmt_18190_call_req_1;
      reqR_unguarded(0) <= call_stmt_18280_call_req_1;
      call_stmt_18190_call_ack_1 <= ackR_unguarded(1);
      call_stmt_18280_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      guard_vector(1)  <=  '1';
      accessMemory_call_group_0_accessRegulator_0: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_0", num_slots => 1) -- 
        port map (req => reqL_unregulated(0), -- 
          ack => ackL_unregulated(0),
          regulated_req => reqL(0),
          regulated_ack => ackL(0),
          release_req => reqR(0),
          release_ack => ackR(0),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_accessRegulator_1: access_regulator_base generic map (name => "accessMemory_call_group_0_accessRegulator_1", num_slots => 1) -- 
        port map (req => reqL_unregulated(1), -- 
          ack => ackL_unregulated(1),
          regulated_req => reqL(1),
          regulated_ack => ackL(1),
          release_req => reqR(1),
          release_ack => ackR(1),
          clk => clk, reset => reset); -- 
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 2, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_18182_wire_constant & type_cast_18184_wire_constant & R_FULL_BYTE_MASK_18185_wire_constant & control_data_addr_18177 & type_cast_18188_wire_constant & type_cast_18272_wire_constant & type_cast_18274_wire_constant & R_FULL_BYTE_MASK_18275_wire_constant & nmem_addr_18255 & type_cast_18278_wire_constant;
      control_data_18190 <= data_out(127 downto 64);
      last_word_18280 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 220,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 2,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(1),
          ackR => accessMemory_call_acks(1),
          dataR => accessMemory_call_data(219 downto 110),
          tagR => accessMemory_call_tag(5 downto 3),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 128,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 2) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(1), -- cross-over
          ackL => accessMemory_return_reqs(1), -- cross-over
          dataL => accessMemory_return_data(127 downto 64),
          tagL => accessMemory_return_tag(5 downto 3),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- shared call operator group (1) : call_stmt_18227_call 
    accessMemory_call_group_1: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_18227_call_req_0;
      call_stmt_18227_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_18227_call_req_1;
      call_stmt_18227_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_1_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_18219_wire_constant & type_cast_18221_wire_constant & R_FULL_BYTE_MASK_18222_wire_constant & mem_addr_18211 & type_cast_18225_wire_constant;
      data_18227 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 3,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 1
    -- shared call operator group (2) : call_stmt_18245_call 
    AccessRegister_call_group_2: Block -- 
      signal data_in: std_logic_vector(42 downto 0);
      signal data_out: std_logic_vector(31 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_18245_call_req_0;
      call_stmt_18245_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_18245_call_req_1;
      call_stmt_18245_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      AccessRegister_call_group_2_gI: SplitGuardInterface generic map(name => "AccessRegister_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_18237_wire_constant & NOT_u4_u4_18240_wire_constant & konst_18241_wire_constant & slice_18243_wire;
      ignore_resp5_18245 <= data_out(31 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 43,
        owidth => 43,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 2,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => AccessRegister_call_reqs(0),
          ackR => AccessRegister_call_acks(0),
          dataR => AccessRegister_call_data(42 downto 0),
          tagR => AccessRegister_call_tag(1 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 32,
          owidth => 32,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 2,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => AccessRegister_return_acks(0), -- cross-over
          ackL => AccessRegister_return_reqs(0), -- cross-over
          dataL => AccessRegister_return_data(31 downto 0),
          tagL => AccessRegister_return_tag(1 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end transmitPacket_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.nic_system_global_package.all;
entity updateTotalMessages is -- 
  generic (tag_length : integer); 
  port ( -- 
    q_base_address : in  std_logic_vector(35 downto 0);
    updated_total_msgs : in  std_logic_vector(31 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity updateTotalMessages;
architecture updateTotalMessages_arch of updateTotalMessages is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 68)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal q_base_address_buffer :  std_logic_vector(35 downto 0);
  signal q_base_address_update_enable: Boolean;
  signal updated_total_msgs_buffer :  std_logic_vector(31 downto 0);
  signal updated_total_msgs_update_enable: Boolean;
  -- output port buffer signals
  signal updateTotalMessages_CP_1290_start: Boolean;
  signal updateTotalMessages_CP_1290_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1016_call_req_0 : boolean;
  signal call_stmt_1016_call_ack_0 : boolean;
  signal call_stmt_1016_call_ack_1 : boolean;
  signal call_stmt_1016_call_req_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "updateTotalMessages_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 68) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= q_base_address;
  q_base_address_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(67 downto 36) <= updated_total_msgs;
  updated_total_msgs_buffer <= in_buffer_data_out(67 downto 36);
  in_buffer_data_in(tag_length + 67 downto 68) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 67 downto 68);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  updateTotalMessages_CP_1290_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "updateTotalMessages_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= updateTotalMessages_CP_1290_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= updateTotalMessages_CP_1290_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= updateTotalMessages_CP_1290_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  updateTotalMessages_CP_1290: Block -- control-path 
    signal updateTotalMessages_CP_1290_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    updateTotalMessages_CP_1290_elements(0) <= updateTotalMessages_CP_1290_start;
    updateTotalMessages_CP_1290_symbol <= updateTotalMessages_CP_1290_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 call_stmt_1016/call_stmt_1016_Sample/$entry
      -- CP-element group 0: 	 call_stmt_1016/call_stmt_1016_Sample/crr
      -- CP-element group 0: 	 call_stmt_1016/call_stmt_1016_Update/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 call_stmt_1016/$entry
      -- CP-element group 0: 	 call_stmt_1016/call_stmt_1016_update_start_
      -- CP-element group 0: 	 call_stmt_1016/call_stmt_1016_sample_start_
      -- CP-element group 0: 	 call_stmt_1016/call_stmt_1016_Update/ccr
      -- 
    ccr_1308_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1308_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateTotalMessages_CP_1290_elements(0), ack => call_stmt_1016_call_req_1); -- 
    crr_1303_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1303_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => updateTotalMessages_CP_1290_elements(0), ack => call_stmt_1016_call_req_0); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 call_stmt_1016/call_stmt_1016_Sample/$exit
      -- CP-element group 1: 	 call_stmt_1016/call_stmt_1016_Sample/cra
      -- CP-element group 1: 	 call_stmt_1016/call_stmt_1016_sample_completed_
      -- 
    cra_1304_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1016_call_ack_0, ack => updateTotalMessages_CP_1290_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 call_stmt_1016/call_stmt_1016_update_completed_
      -- CP-element group 2: 	 call_stmt_1016/call_stmt_1016_Update/cca
      -- CP-element group 2: 	 call_stmt_1016/$exit
      -- CP-element group 2: 	 call_stmt_1016/call_stmt_1016_Update/$exit
      -- 
    cca_1309_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1016_call_ack_1, ack => updateTotalMessages_CP_1290_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u32_u64_1014_wire : std_logic_vector(63 downto 0);
    signal CONCAT_u4_u8_1010_wire_constant : std_logic_vector(7 downto 0);
    signal rdata_1016 : std_logic_vector(63 downto 0);
    signal type_cast_1002_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1004_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    CONCAT_u4_u8_1010_wire_constant <= "11110000";
    type_cast_1002_wire_constant <= "0";
    type_cast_1004_wire_constant <= "0";
    -- binary operator CONCAT_u32_u64_1014_inst
    process(updated_total_msgs_buffer, updated_total_msgs_buffer) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(updated_total_msgs_buffer, updated_total_msgs_buffer, tmp_var);
      CONCAT_u32_u64_1014_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_1016_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1016_call_req_0;
      call_stmt_1016_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1016_call_req_1;
      call_stmt_1016_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1002_wire_constant & type_cast_1004_wire_constant & CONCAT_u4_u8_1010_wire_constant & q_base_address_buffer & CONCAT_u32_u64_1014_wire;
      rdata_1016 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end updateTotalMessages_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.nic_system_global_package.all;
entity writeControlInformationToMem is -- 
  generic (tag_length : integer); 
  port ( -- 
    base_buffer_pointer : in  std_logic_vector(35 downto 0);
    packet_size : in  std_logic_vector(10 downto 0);
    last_keep : in  std_logic_vector(7 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity writeControlInformationToMem;
architecture writeControlInformationToMem_arch of writeControlInformationToMem is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 55)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal base_buffer_pointer_buffer :  std_logic_vector(35 downto 0);
  signal base_buffer_pointer_update_enable: Boolean;
  signal packet_size_buffer :  std_logic_vector(10 downto 0);
  signal packet_size_update_enable: Boolean;
  signal last_keep_buffer :  std_logic_vector(7 downto 0);
  signal last_keep_update_enable: Boolean;
  -- output port buffer signals
  signal writeControlInformationToMem_CP_1812_start: Boolean;
  signal writeControlInformationToMem_CP_1812_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal call_stmt_1411_call_req_0 : boolean;
  signal call_stmt_1411_call_ack_0 : boolean;
  signal call_stmt_1411_call_req_1 : boolean;
  signal call_stmt_1411_call_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "writeControlInformationToMem_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 55) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= base_buffer_pointer;
  base_buffer_pointer_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(46 downto 36) <= packet_size;
  packet_size_buffer <= in_buffer_data_out(46 downto 36);
  in_buffer_data_in(54 downto 47) <= last_keep;
  last_keep_buffer <= in_buffer_data_out(54 downto 47);
  in_buffer_data_in(tag_length + 54 downto 55) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 54 downto 55);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  writeControlInformationToMem_CP_1812_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "writeControlInformationToMem_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeControlInformationToMem_CP_1812_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= writeControlInformationToMem_CP_1812_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeControlInformationToMem_CP_1812_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  writeControlInformationToMem_CP_1812: Block -- control-path 
    signal writeControlInformationToMem_CP_1812_elements: BooleanArray(2 downto 0);
    -- 
  begin -- 
    writeControlInformationToMem_CP_1812_elements(0) <= writeControlInformationToMem_CP_1812_start;
    writeControlInformationToMem_CP_1812_symbol <= writeControlInformationToMem_CP_1812_elements(2);
    -- CP-element group 0:  fork  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (8) 
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 assign_stmt_1402_to_call_stmt_1411/$entry
      -- CP-element group 0: 	 assign_stmt_1402_to_call_stmt_1411/call_stmt_1411_sample_start_
      -- CP-element group 0: 	 assign_stmt_1402_to_call_stmt_1411/call_stmt_1411_update_start_
      -- CP-element group 0: 	 assign_stmt_1402_to_call_stmt_1411/call_stmt_1411_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_1402_to_call_stmt_1411/call_stmt_1411_Sample/crr
      -- CP-element group 0: 	 assign_stmt_1402_to_call_stmt_1411/call_stmt_1411_Update/$entry
      -- CP-element group 0: 	 assign_stmt_1402_to_call_stmt_1411/call_stmt_1411_Update/ccr
      -- 
    crr_1825_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1825_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeControlInformationToMem_CP_1812_elements(0), ack => call_stmt_1411_call_req_0); -- 
    ccr_1830_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1830_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeControlInformationToMem_CP_1812_elements(0), ack => call_stmt_1411_call_req_1); -- 
    -- CP-element group 1:  transition  input  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (3) 
      -- CP-element group 1: 	 assign_stmt_1402_to_call_stmt_1411/call_stmt_1411_sample_completed_
      -- CP-element group 1: 	 assign_stmt_1402_to_call_stmt_1411/call_stmt_1411_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_1402_to_call_stmt_1411/call_stmt_1411_Sample/cra
      -- 
    cra_1826_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1411_call_ack_0, ack => writeControlInformationToMem_CP_1812_elements(1)); -- 
    -- CP-element group 2:  transition  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2:  members (5) 
      -- CP-element group 2: 	 $exit
      -- CP-element group 2: 	 assign_stmt_1402_to_call_stmt_1411/$exit
      -- CP-element group 2: 	 assign_stmt_1402_to_call_stmt_1411/call_stmt_1411_update_completed_
      -- CP-element group 2: 	 assign_stmt_1402_to_call_stmt_1411/call_stmt_1411_Update/$exit
      -- CP-element group 2: 	 assign_stmt_1402_to_call_stmt_1411/call_stmt_1411_Update/cca
      -- 
    cca_1831_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1411_call_ack_1, ack => writeControlInformationToMem_CP_1812_elements(2)); -- 
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u11_u19_1400_wire : std_logic_vector(18 downto 0);
    signal R_FULL_BYTE_MASK_1407_wire_constant : std_logic_vector(7 downto 0);
    signal control_data_1402 : std_logic_vector(63 downto 0);
    signal ignore_return_1411 : std_logic_vector(63 downto 0);
    signal type_cast_1404_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1406_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    R_FULL_BYTE_MASK_1407_wire_constant <= "11111111";
    type_cast_1404_wire_constant <= "0";
    type_cast_1406_wire_constant <= "0";
    -- interlock type_cast_1401_inst
    process(CONCAT_u11_u19_1400_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 18 downto 0) := CONCAT_u11_u19_1400_wire(18 downto 0);
      control_data_1402 <= tmp_var; -- 
    end process;
    -- binary operator CONCAT_u11_u19_1400_inst
    process(packet_size_buffer, last_keep_buffer) -- 
      variable tmp_var : std_logic_vector(18 downto 0); -- 
    begin -- 
      ApConcat_proc(packet_size_buffer, last_keep_buffer, tmp_var);
      CONCAT_u11_u19_1400_wire <= tmp_var; --
    end process;
    -- shared call operator group (0) : call_stmt_1411_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1411_call_req_0;
      call_stmt_1411_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1411_call_req_1;
      call_stmt_1411_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1404_wire_constant & type_cast_1406_wire_constant & R_FULL_BYTE_MASK_1407_wire_constant & base_buffer_pointer_buffer & control_data_1402;
      ignore_return_1411 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  false,
        twidth => 3,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => false, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end writeControlInformationToMem_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.nic_system_global_package.all;
entity writeEthernetHeaderToMem is -- 
  generic (tag_length : integer); 
  port ( -- 
    buf_pointer : in  std_logic_vector(35 downto 0);
    buf_position_out : out  std_logic_vector(35 downto 0);
    nic_rx_to_header_pipe_read_req : out  std_logic_vector(0 downto 0);
    nic_rx_to_header_pipe_read_ack : in   std_logic_vector(0 downto 0);
    nic_rx_to_header_pipe_read_data : in   std_logic_vector(72 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity writeEthernetHeaderToMem;
architecture writeEthernetHeaderToMem_arch of writeEthernetHeaderToMem is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 36)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal buf_pointer_buffer :  std_logic_vector(35 downto 0);
  signal buf_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal buf_position_out_buffer :  std_logic_vector(35 downto 0);
  signal buf_position_out_update_enable: Boolean;
  signal writeEthernetHeaderToMem_CP_1496_start: Boolean;
  signal writeEthernetHeaderToMem_CP_1496_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal ADD_u36_u36_1263_inst_req_1 : boolean;
  signal ADD_u36_u36_1263_inst_req_0 : boolean;
  signal ADD_u36_u36_1263_inst_ack_1 : boolean;
  signal nbuf_position_1303_1264_buf_ack_0 : boolean;
  signal nI_1298_1269_buf_req_0 : boolean;
  signal ADD_u36_u36_1263_inst_ack_0 : boolean;
  signal call_stmt_1293_call_req_1 : boolean;
  signal nI_1298_1269_buf_ack_0 : boolean;
  signal nbuf_position_1303_1264_buf_ack_1 : boolean;
  signal nbuf_position_1303_1264_buf_req_1 : boolean;
  signal do_while_stmt_1257_branch_req_0 : boolean;
  signal call_stmt_1293_call_ack_0 : boolean;
  signal call_stmt_1293_call_req_0 : boolean;
  signal do_while_stmt_1257_branch_ack_1 : boolean;
  signal phi_stmt_1259_ack_0 : boolean;
  signal phi_stmt_1259_req_0 : boolean;
  signal do_while_stmt_1257_branch_ack_0 : boolean;
  signal phi_stmt_1259_req_1 : boolean;
  signal RPIPE_nic_rx_to_header_1272_inst_ack_1 : boolean;
  signal RPIPE_nic_rx_to_header_1272_inst_req_1 : boolean;
  signal nbuf_position_1303_1264_buf_req_0 : boolean;
  signal RPIPE_nic_rx_to_header_1272_inst_ack_0 : boolean;
  signal RPIPE_nic_rx_to_header_1272_inst_req_0 : boolean;
  signal phi_stmt_1265_ack_0 : boolean;
  signal call_stmt_1293_call_ack_1 : boolean;
  signal phi_stmt_1265_req_0 : boolean;
  signal W_buf_position_out_1309_inst_ack_1 : boolean;
  signal phi_stmt_1265_req_1 : boolean;
  signal W_buf_position_out_1309_inst_req_1 : boolean;
  signal nI_1298_1269_buf_ack_1 : boolean;
  signal nI_1298_1269_buf_req_1 : boolean;
  signal W_buf_position_out_1309_inst_ack_0 : boolean;
  signal W_buf_position_out_1309_inst_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "writeEthernetHeaderToMem_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 36) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= buf_pointer;
  buf_pointer_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(tag_length + 35 downto 36) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 35 downto 36);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  writeEthernetHeaderToMem_CP_1496_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "writeEthernetHeaderToMem_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 36) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(35 downto 0) <= buf_position_out_buffer;
  buf_position_out <= out_buffer_data_out(35 downto 0);
  out_buffer_data_in(tag_length + 35 downto 36) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 35 downto 36);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeEthernetHeaderToMem_CP_1496_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= writeEthernetHeaderToMem_CP_1496_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeEthernetHeaderToMem_CP_1496_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  writeEthernetHeaderToMem_CP_1496: Block -- control-path 
    signal writeEthernetHeaderToMem_CP_1496_elements: BooleanArray(68 downto 0);
    -- 
  begin -- 
    writeEthernetHeaderToMem_CP_1496_elements(0) <= writeEthernetHeaderToMem_CP_1496_start;
    writeEthernetHeaderToMem_CP_1496_symbol <= writeEthernetHeaderToMem_CP_1496_elements(68);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_1256/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1256/do_while_stmt_1257__entry__
      -- CP-element group 0: 	 branch_block_stmt_1256/branch_block_stmt_1256__entry__
      -- 
    -- CP-element group 1:  fork  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	66 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	67 
    -- CP-element group 1: 	68 
    -- CP-element group 1:  members (10) 
      -- CP-element group 1: 	 assign_stmt_1311/assign_stmt_1311_sample_start_
      -- CP-element group 1: 	 assign_stmt_1311/$entry
      -- CP-element group 1: 	 assign_stmt_1311/assign_stmt_1311_update_start_
      -- CP-element group 1: 	 assign_stmt_1311/assign_stmt_1311_Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_1256/$exit
      -- CP-element group 1: 	 branch_block_stmt_1256/do_while_stmt_1257__exit__
      -- CP-element group 1: 	 assign_stmt_1311/assign_stmt_1311_Update/req
      -- CP-element group 1: 	 assign_stmt_1311/assign_stmt_1311_Update/$entry
      -- CP-element group 1: 	 branch_block_stmt_1256/branch_block_stmt_1256__exit__
      -- CP-element group 1: 	 assign_stmt_1311/assign_stmt_1311_Sample/req
      -- 
    req_1681_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1681_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1496_elements(1), ack => W_buf_position_out_1309_inst_req_1); -- 
    req_1676_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1676_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1496_elements(1), ack => W_buf_position_out_1309_inst_req_0); -- 
    writeEthernetHeaderToMem_CP_1496_elements(1) <= writeEthernetHeaderToMem_CP_1496_elements(66);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1256/do_while_stmt_1257/$entry
      -- CP-element group 2: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257__entry__
      -- 
    writeEthernetHeaderToMem_CP_1496_elements(2) <= writeEthernetHeaderToMem_CP_1496_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	66 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257__exit__
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1496_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1256/do_while_stmt_1257/loop_back
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1496_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	64 
    -- CP-element group 5: 	65 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1256/do_while_stmt_1257/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1256/do_while_stmt_1257/loop_taken/$entry
      -- CP-element group 5: 	 branch_block_stmt_1256/do_while_stmt_1257/loop_exit/$entry
      -- 
    writeEthernetHeaderToMem_CP_1496_elements(5) <= writeEthernetHeaderToMem_CP_1496_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	63 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1256/do_while_stmt_1257/loop_body_done
      -- 
    writeEthernetHeaderToMem_CP_1496_elements(6) <= writeEthernetHeaderToMem_CP_1496_elements(63);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	40 
    -- CP-element group 7: 	21 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/back_edge_to_loop_body
      -- 
    writeEthernetHeaderToMem_CP_1496_elements(7) <= writeEthernetHeaderToMem_CP_1496_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	42 
    -- CP-element group 8: 	23 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/first_time_through_loop_body
      -- 
    writeEthernetHeaderToMem_CP_1496_elements(8) <= writeEthernetHeaderToMem_CP_1496_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	53 
    -- CP-element group 9: 	62 
    -- CP-element group 9: 	36 
    -- CP-element group 9: 	37 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	11 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1270_sample_start_
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1496_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	62 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/condition_evaluated
      -- 
    condition_evaluated_1520_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1520_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1496_elements(10), ack => do_while_stmt_1257_branch_req_0); -- 
    writeEthernetHeaderToMem_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1496_elements(62) & writeEthernetHeaderToMem_CP_1496_elements(14);
      gj_writeEthernetHeaderToMem_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1496_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	36 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	9 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	54 
    -- CP-element group 11: 	17 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/aggregated_phi_sample_req
      -- CP-element group 11: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1265_sample_start__ps
      -- 
    writeEthernetHeaderToMem_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1496_elements(36) & writeEthernetHeaderToMem_CP_1496_elements(15) & writeEthernetHeaderToMem_CP_1496_elements(9) & writeEthernetHeaderToMem_CP_1496_elements(14);
      gj_writeEthernetHeaderToMem_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1496_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	56 
    -- CP-element group 12: 	38 
    -- CP-element group 12: 	18 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	63 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	36 
    -- CP-element group 12: 	15 
    -- CP-element group 12:  members (4) 
      -- CP-element group 12: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1265_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1259_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1270_sample_completed_
      -- 
    writeEthernetHeaderToMem_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1496_elements(56) & writeEthernetHeaderToMem_CP_1496_elements(38) & writeEthernetHeaderToMem_CP_1496_elements(18);
      gj_writeEthernetHeaderToMem_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1496_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	53 
    -- CP-element group 13: 	37 
    -- CP-element group 13: 	16 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	55 
    -- CP-element group 13: 	19 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/aggregated_phi_update_req
      -- CP-element group 13: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1265_update_start__ps
      -- 
    writeEthernetHeaderToMem_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1496_elements(53) & writeEthernetHeaderToMem_CP_1496_elements(37) & writeEthernetHeaderToMem_CP_1496_elements(16);
      gj_writeEthernetHeaderToMem_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1496_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	57 
    -- CP-element group 14: 	39 
    -- CP-element group 14: 	20 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/aggregated_phi_update_ack
      -- 
    writeEthernetHeaderToMem_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1496_elements(57) & writeEthernetHeaderToMem_CP_1496_elements(39) & writeEthernetHeaderToMem_CP_1496_elements(20);
      gj_writeEthernetHeaderToMem_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1496_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1259_sample_start_
      -- 
    writeEthernetHeaderToMem_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1496_elements(9) & writeEthernetHeaderToMem_CP_1496_elements(12);
      gj_writeEthernetHeaderToMem_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1496_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	60 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1259_update_start_
      -- 
    writeEthernetHeaderToMem_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1496_elements(9) & writeEthernetHeaderToMem_CP_1496_elements(60);
      gj_writeEthernetHeaderToMem_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1496_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	11 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1259_sample_start__ps
      -- 
    writeEthernetHeaderToMem_CP_1496_elements(17) <= writeEthernetHeaderToMem_CP_1496_elements(11);
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	12 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1259_sample_completed__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1496_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	13 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1259_update_start__ps
      -- 
    writeEthernetHeaderToMem_CP_1496_elements(19) <= writeEthernetHeaderToMem_CP_1496_elements(13);
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	58 
    -- CP-element group 20: 	14 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1259_update_completed_
      -- CP-element group 20: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1259_update_completed__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1496_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	7 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1259_loopback_trigger
      -- 
    writeEthernetHeaderToMem_CP_1496_elements(21) <= writeEthernetHeaderToMem_CP_1496_elements(7);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1259_loopback_sample_req_ps
      -- CP-element group 22: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1259_loopback_sample_req
      -- 
    phi_stmt_1259_loopback_sample_req_1535_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1259_loopback_sample_req_1535_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1496_elements(22), ack => phi_stmt_1259_req_1); -- 
    -- Element group writeEthernetHeaderToMem_CP_1496_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	8 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1259_entry_trigger
      -- 
    writeEthernetHeaderToMem_CP_1496_elements(23) <= writeEthernetHeaderToMem_CP_1496_elements(8);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1259_entry_sample_req_ps
      -- CP-element group 24: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1259_entry_sample_req
      -- 
    phi_stmt_1259_entry_sample_req_1538_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1259_entry_sample_req_1538_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1496_elements(24), ack => phi_stmt_1259_req_0); -- 
    -- Element group writeEthernetHeaderToMem_CP_1496_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1259_phi_mux_ack_ps
      -- CP-element group 25: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1259_phi_mux_ack
      -- 
    phi_stmt_1259_phi_mux_ack_1541_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 25_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1259_ack_0, ack => writeEthernetHeaderToMem_CP_1496_elements(25)); -- 
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (1) 
      -- CP-element group 26: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/ADD_u36_u36_1263_sample_start__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1496_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27: 	29 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/ADD_u36_u36_1263_update_start__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1496_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: marked-predecessors 
    -- CP-element group 28: 	30 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (3) 
      -- CP-element group 28: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/ADD_u36_u36_1263_Sample/rr
      -- CP-element group 28: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/ADD_u36_u36_1263_Sample/$entry
      -- CP-element group 28: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/ADD_u36_u36_1263_sample_start_
      -- 
    rr_1554_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1554_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1496_elements(28), ack => ADD_u36_u36_1263_inst_req_0); -- 
    writeEthernetHeaderToMem_cp_element_group_28: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_28"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1496_elements(26) & writeEthernetHeaderToMem_CP_1496_elements(30);
      gj_writeEthernetHeaderToMem_cp_element_group_28 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1496_elements(28), clk => clk, reset => reset); --
    end block;
    -- CP-element group 29:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	27 
    -- CP-element group 29: marked-predecessors 
    -- CP-element group 29: 	31 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (3) 
      -- CP-element group 29: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/ADD_u36_u36_1263_Update/cr
      -- CP-element group 29: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/ADD_u36_u36_1263_Update/$entry
      -- CP-element group 29: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/ADD_u36_u36_1263_update_start_
      -- 
    cr_1559_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1559_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1496_elements(29), ack => ADD_u36_u36_1263_inst_req_1); -- 
    writeEthernetHeaderToMem_cp_element_group_29: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_29"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1496_elements(27) & writeEthernetHeaderToMem_CP_1496_elements(31);
      gj_writeEthernetHeaderToMem_cp_element_group_29 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1496_elements(29), clk => clk, reset => reset); --
    end block;
    -- CP-element group 30:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: marked-successors 
    -- CP-element group 30: 	28 
    -- CP-element group 30:  members (4) 
      -- CP-element group 30: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/ADD_u36_u36_1263_Sample/$exit
      -- CP-element group 30: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/ADD_u36_u36_1263_Sample/ra
      -- CP-element group 30: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/ADD_u36_u36_1263_sample_completed_
      -- CP-element group 30: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/ADD_u36_u36_1263_sample_completed__ps
      -- 
    ra_1555_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 30_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_1263_inst_ack_0, ack => writeEthernetHeaderToMem_CP_1496_elements(30)); -- 
    -- CP-element group 31:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: marked-successors 
    -- CP-element group 31: 	29 
    -- CP-element group 31:  members (4) 
      -- CP-element group 31: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/ADD_u36_u36_1263_Update/ca
      -- CP-element group 31: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/ADD_u36_u36_1263_Update/$exit
      -- CP-element group 31: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/ADD_u36_u36_1263_update_completed__ps
      -- CP-element group 31: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/ADD_u36_u36_1263_update_completed_
      -- 
    ca_1560_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 31_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_1263_inst_ack_1, ack => writeEthernetHeaderToMem_CP_1496_elements(31)); -- 
    -- CP-element group 32:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/R_nbuf_position_1264_sample_start_
      -- CP-element group 32: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/R_nbuf_position_1264_sample_start__ps
      -- CP-element group 32: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/R_nbuf_position_1264_Sample/req
      -- CP-element group 32: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/R_nbuf_position_1264_Sample/$entry
      -- 
    req_1572_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1572_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1496_elements(32), ack => nbuf_position_1303_1264_buf_req_0); -- 
    -- Element group writeEthernetHeaderToMem_CP_1496_elements(32) is bound as output of CP function.
    -- CP-element group 33:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/R_nbuf_position_1264_update_start__ps
      -- CP-element group 33: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/R_nbuf_position_1264_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/R_nbuf_position_1264_Update/req
      -- CP-element group 33: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/R_nbuf_position_1264_update_start_
      -- 
    req_1577_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1577_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1496_elements(33), ack => nbuf_position_1303_1264_buf_req_1); -- 
    -- Element group writeEthernetHeaderToMem_CP_1496_elements(33) is bound as output of CP function.
    -- CP-element group 34:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/R_nbuf_position_1264_Sample/ack
      -- CP-element group 34: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/R_nbuf_position_1264_sample_completed__ps
      -- CP-element group 34: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/R_nbuf_position_1264_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/R_nbuf_position_1264_sample_completed_
      -- 
    ack_1573_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nbuf_position_1303_1264_buf_ack_0, ack => writeEthernetHeaderToMem_CP_1496_elements(34)); -- 
    -- CP-element group 35:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/R_nbuf_position_1264_update_completed__ps
      -- CP-element group 35: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/R_nbuf_position_1264_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/R_nbuf_position_1264_Update/ack
      -- CP-element group 35: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/R_nbuf_position_1264_update_completed_
      -- 
    ack_1578_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nbuf_position_1303_1264_buf_ack_1, ack => writeEthernetHeaderToMem_CP_1496_elements(35)); -- 
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	9 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	12 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	11 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1265_sample_start_
      -- 
    writeEthernetHeaderToMem_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1496_elements(9) & writeEthernetHeaderToMem_CP_1496_elements(12);
      gj_writeEthernetHeaderToMem_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1496_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	9 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	39 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	13 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1265_update_start_
      -- 
    writeEthernetHeaderToMem_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1496_elements(9) & writeEthernetHeaderToMem_CP_1496_elements(39);
      gj_writeEthernetHeaderToMem_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1496_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	12 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1265_sample_completed__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1496_elements(38) is bound as output of CP function.
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	14 
    -- CP-element group 39: marked-successors 
    -- CP-element group 39: 	37 
    -- CP-element group 39:  members (2) 
      -- CP-element group 39: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1265_update_completed__ps
      -- CP-element group 39: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1265_update_completed_
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1496_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	7 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1265_loopback_trigger
      -- 
    writeEthernetHeaderToMem_CP_1496_elements(40) <= writeEthernetHeaderToMem_CP_1496_elements(7);
    -- CP-element group 41:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1265_loopback_sample_req_ps
      -- CP-element group 41: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1265_loopback_sample_req
      -- 
    phi_stmt_1265_loopback_sample_req_1589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1265_loopback_sample_req_1589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1496_elements(41), ack => phi_stmt_1265_req_1); -- 
    -- Element group writeEthernetHeaderToMem_CP_1496_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	8 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1265_entry_trigger
      -- 
    writeEthernetHeaderToMem_CP_1496_elements(42) <= writeEthernetHeaderToMem_CP_1496_elements(8);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1265_entry_sample_req_ps
      -- CP-element group 43: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1265_entry_sample_req
      -- 
    phi_stmt_1265_entry_sample_req_1592_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1265_entry_sample_req_1592_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1496_elements(43), ack => phi_stmt_1265_req_0); -- 
    -- Element group writeEthernetHeaderToMem_CP_1496_elements(43) is bound as output of CP function.
    -- CP-element group 44:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1265_phi_mux_ack_ps
      -- CP-element group 44: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1265_phi_mux_ack
      -- 
    phi_stmt_1265_phi_mux_ack_1595_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 44_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1265_ack_0, ack => writeEthernetHeaderToMem_CP_1496_elements(44)); -- 
    -- CP-element group 45:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (4) 
      -- CP-element group 45: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/type_cast_1268_sample_completed_
      -- CP-element group 45: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/type_cast_1268_sample_start_
      -- CP-element group 45: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/type_cast_1268_sample_completed__ps
      -- CP-element group 45: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/type_cast_1268_sample_start__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1496_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/type_cast_1268_update_start_
      -- CP-element group 46: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/type_cast_1268_update_start__ps
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1496_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	48 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/type_cast_1268_update_completed__ps
      -- 
    writeEthernetHeaderToMem_CP_1496_elements(47) <= writeEthernetHeaderToMem_CP_1496_elements(48);
    -- CP-element group 48:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	47 
    -- CP-element group 48:  members (1) 
      -- CP-element group 48: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/type_cast_1268_update_completed_
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1496_elements(48) is a control-delay.
    cp_element_48_delay: control_delay_element  generic map(name => " 48_delay", delay_value => 1)  port map(req => writeEthernetHeaderToMem_CP_1496_elements(46), ack => writeEthernetHeaderToMem_CP_1496_elements(48), clk => clk, reset =>reset);
    -- CP-element group 49:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/R_nI_1269_Sample/req
      -- CP-element group 49: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/R_nI_1269_Sample/$entry
      -- CP-element group 49: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/R_nI_1269_sample_start_
      -- CP-element group 49: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/R_nI_1269_sample_start__ps
      -- 
    req_1616_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1616_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1496_elements(49), ack => nI_1298_1269_buf_req_0); -- 
    -- Element group writeEthernetHeaderToMem_CP_1496_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	52 
    -- CP-element group 50:  members (4) 
      -- CP-element group 50: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/R_nI_1269_update_start_
      -- CP-element group 50: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/R_nI_1269_update_start__ps
      -- CP-element group 50: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/R_nI_1269_Update/req
      -- CP-element group 50: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/R_nI_1269_Update/$entry
      -- 
    req_1621_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1621_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1496_elements(50), ack => nI_1298_1269_buf_req_1); -- 
    -- Element group writeEthernetHeaderToMem_CP_1496_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51:  members (4) 
      -- CP-element group 51: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/R_nI_1269_Sample/$exit
      -- CP-element group 51: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/R_nI_1269_sample_completed_
      -- CP-element group 51: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/R_nI_1269_Sample/ack
      -- CP-element group 51: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/R_nI_1269_sample_completed__ps
      -- 
    ack_1617_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nI_1298_1269_buf_ack_0, ack => writeEthernetHeaderToMem_CP_1496_elements(51)); -- 
    -- CP-element group 52:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	50 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/R_nI_1269_update_completed_
      -- CP-element group 52: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/R_nI_1269_update_completed__ps
      -- CP-element group 52: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/R_nI_1269_Update/ack
      -- CP-element group 52: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/R_nI_1269_Update/$exit
      -- 
    ack_1622_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 52_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nI_1298_1269_buf_ack_1, ack => writeEthernetHeaderToMem_CP_1496_elements(52)); -- 
    -- CP-element group 53:  join  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	9 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	60 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	13 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1270_update_start_
      -- 
    writeEthernetHeaderToMem_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1496_elements(9) & writeEthernetHeaderToMem_CP_1496_elements(60);
      gj_writeEthernetHeaderToMem_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1496_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	11 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	57 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/RPIPE_nic_rx_to_header_1272_Sample/rr
      -- CP-element group 54: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/RPIPE_nic_rx_to_header_1272_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/RPIPE_nic_rx_to_header_1272_sample_start_
      -- 
    rr_1635_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1635_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1496_elements(54), ack => RPIPE_nic_rx_to_header_1272_inst_req_0); -- 
    writeEthernetHeaderToMem_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1496_elements(11) & writeEthernetHeaderToMem_CP_1496_elements(57);
      gj_writeEthernetHeaderToMem_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1496_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	56 
    -- CP-element group 55: 	13 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/RPIPE_nic_rx_to_header_1272_Update/cr
      -- CP-element group 55: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/RPIPE_nic_rx_to_header_1272_Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/RPIPE_nic_rx_to_header_1272_update_start_
      -- 
    cr_1640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1496_elements(55), ack => RPIPE_nic_rx_to_header_1272_inst_req_1); -- 
    writeEthernetHeaderToMem_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1496_elements(56) & writeEthernetHeaderToMem_CP_1496_elements(13);
      gj_writeEthernetHeaderToMem_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1496_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	55 
    -- CP-element group 56: 	12 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/RPIPE_nic_rx_to_header_1272_Sample/ra
      -- CP-element group 56: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/RPIPE_nic_rx_to_header_1272_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/RPIPE_nic_rx_to_header_1272_sample_completed_
      -- 
    ra_1636_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_nic_rx_to_header_1272_inst_ack_0, ack => writeEthernetHeaderToMem_CP_1496_elements(56)); -- 
    -- CP-element group 57:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	58 
    -- CP-element group 57: 	14 
    -- CP-element group 57: marked-successors 
    -- CP-element group 57: 	54 
    -- CP-element group 57:  members (4) 
      -- CP-element group 57: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/RPIPE_nic_rx_to_header_1272_Update/ca
      -- CP-element group 57: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/RPIPE_nic_rx_to_header_1272_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/RPIPE_nic_rx_to_header_1272_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/phi_stmt_1270_update_completed_
      -- 
    ca_1641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_nic_rx_to_header_1272_inst_ack_1, ack => writeEthernetHeaderToMem_CP_1496_elements(57)); -- 
    -- CP-element group 58:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	57 
    -- CP-element group 58: 	20 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	60 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/call_stmt_1293_Sample/$entry
      -- CP-element group 58: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/call_stmt_1293_sample_start_
      -- CP-element group 58: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/call_stmt_1293_Sample/crr
      -- 
    crr_1649_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1649_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1496_elements(58), ack => call_stmt_1293_call_req_0); -- 
    writeEthernetHeaderToMem_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1496_elements(57) & writeEthernetHeaderToMem_CP_1496_elements(20) & writeEthernetHeaderToMem_CP_1496_elements(60);
      gj_writeEthernetHeaderToMem_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1496_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	61 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	61 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/call_stmt_1293_Update/$entry
      -- CP-element group 59: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/call_stmt_1293_Update/ccr
      -- CP-element group 59: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/call_stmt_1293_update_start_
      -- 
    ccr_1654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeEthernetHeaderToMem_CP_1496_elements(59), ack => call_stmt_1293_call_req_1); -- 
    writeEthernetHeaderToMem_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= writeEthernetHeaderToMem_CP_1496_elements(61);
      gj_writeEthernetHeaderToMem_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1496_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: successors 
    -- CP-element group 60: marked-successors 
    -- CP-element group 60: 	53 
    -- CP-element group 60: 	58 
    -- CP-element group 60: 	16 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/call_stmt_1293_Sample/$exit
      -- CP-element group 60: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/call_stmt_1293_sample_completed_
      -- CP-element group 60: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/call_stmt_1293_Sample/cra
      -- 
    cra_1650_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 60_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1293_call_ack_0, ack => writeEthernetHeaderToMem_CP_1496_elements(60)); -- 
    -- CP-element group 61:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	59 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61: marked-successors 
    -- CP-element group 61: 	59 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/call_stmt_1293_Update/$exit
      -- CP-element group 61: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/call_stmt_1293_update_completed_
      -- CP-element group 61: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/call_stmt_1293_Update/cca
      -- 
    cca_1655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1293_call_ack_1, ack => writeEthernetHeaderToMem_CP_1496_elements(61)); -- 
    -- CP-element group 62:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	9 
    -- CP-element group 62: successors 
    -- CP-element group 62: 	10 
    -- CP-element group 62:  members (1) 
      -- CP-element group 62: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group writeEthernetHeaderToMem_CP_1496_elements(62) is a control-delay.
    cp_element_62_delay: control_delay_element  generic map(name => " 62_delay", delay_value => 1)  port map(req => writeEthernetHeaderToMem_CP_1496_elements(9), ack => writeEthernetHeaderToMem_CP_1496_elements(62), clk => clk, reset =>reset);
    -- CP-element group 63:  join  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: 	12 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	6 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_1256/do_while_stmt_1257/do_while_stmt_1257_loop_body/$exit
      -- 
    writeEthernetHeaderToMem_cp_element_group_63: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 44) := "writeEthernetHeaderToMem_cp_element_group_63"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeEthernetHeaderToMem_CP_1496_elements(61) & writeEthernetHeaderToMem_CP_1496_elements(12);
      gj_writeEthernetHeaderToMem_cp_element_group_63 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1496_elements(63), clk => clk, reset => reset); --
    end block;
    -- CP-element group 64:  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	5 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_1256/do_while_stmt_1257/loop_exit/ack
      -- CP-element group 64: 	 branch_block_stmt_1256/do_while_stmt_1257/loop_exit/$exit
      -- 
    ack_1660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1257_branch_ack_0, ack => writeEthernetHeaderToMem_CP_1496_elements(64)); -- 
    -- CP-element group 65:  transition  input  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	5 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_1256/do_while_stmt_1257/loop_taken/ack
      -- CP-element group 65: 	 branch_block_stmt_1256/do_while_stmt_1257/loop_taken/$exit
      -- 
    ack_1664_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1257_branch_ack_1, ack => writeEthernetHeaderToMem_CP_1496_elements(65)); -- 
    -- CP-element group 66:  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	3 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	1 
    -- CP-element group 66:  members (1) 
      -- CP-element group 66: 	 branch_block_stmt_1256/do_while_stmt_1257/$exit
      -- 
    writeEthernetHeaderToMem_CP_1496_elements(66) <= writeEthernetHeaderToMem_CP_1496_elements(3);
    -- CP-element group 67:  transition  input  bypass 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	1 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 assign_stmt_1311/assign_stmt_1311_sample_completed_
      -- CP-element group 67: 	 assign_stmt_1311/assign_stmt_1311_Sample/$exit
      -- CP-element group 67: 	 assign_stmt_1311/assign_stmt_1311_Sample/ack
      -- 
    ack_1677_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_buf_position_out_1309_inst_ack_0, ack => writeEthernetHeaderToMem_CP_1496_elements(67)); -- 
    -- CP-element group 68:  transition  input  bypass 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	1 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (5) 
      -- CP-element group 68: 	 assign_stmt_1311/$exit
      -- CP-element group 68: 	 assign_stmt_1311/assign_stmt_1311_update_completed_
      -- CP-element group 68: 	 $exit
      -- CP-element group 68: 	 assign_stmt_1311/assign_stmt_1311_Update/ack
      -- CP-element group 68: 	 assign_stmt_1311/assign_stmt_1311_Update/$exit
      -- 
    ack_1682_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_buf_position_out_1309_inst_ack_1, ack => writeEthernetHeaderToMem_CP_1496_elements(68)); -- 
    writeEthernetHeaderToMem_do_while_stmt_1257_terminator_1665: loop_terminator -- 
      generic map (name => " writeEthernetHeaderToMem_do_while_stmt_1257_terminator_1665", max_iterations_in_flight =>15) 
      port map(loop_body_exit => writeEthernetHeaderToMem_CP_1496_elements(6),loop_continue => writeEthernetHeaderToMem_CP_1496_elements(65),loop_terminate => writeEthernetHeaderToMem_CP_1496_elements(64),loop_back => writeEthernetHeaderToMem_CP_1496_elements(4),loop_exit => writeEthernetHeaderToMem_CP_1496_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1259_phi_seq_1579_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= writeEthernetHeaderToMem_CP_1496_elements(23);
      writeEthernetHeaderToMem_CP_1496_elements(26)<= src_sample_reqs(0);
      src_sample_acks(0)  <= writeEthernetHeaderToMem_CP_1496_elements(30);
      writeEthernetHeaderToMem_CP_1496_elements(27)<= src_update_reqs(0);
      src_update_acks(0)  <= writeEthernetHeaderToMem_CP_1496_elements(31);
      writeEthernetHeaderToMem_CP_1496_elements(24) <= phi_mux_reqs(0);
      triggers(1)  <= writeEthernetHeaderToMem_CP_1496_elements(21);
      writeEthernetHeaderToMem_CP_1496_elements(32)<= src_sample_reqs(1);
      src_sample_acks(1)  <= writeEthernetHeaderToMem_CP_1496_elements(34);
      writeEthernetHeaderToMem_CP_1496_elements(33)<= src_update_reqs(1);
      src_update_acks(1)  <= writeEthernetHeaderToMem_CP_1496_elements(35);
      writeEthernetHeaderToMem_CP_1496_elements(22) <= phi_mux_reqs(1);
      phi_stmt_1259_phi_seq_1579 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1259_phi_seq_1579") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => writeEthernetHeaderToMem_CP_1496_elements(17), 
          phi_sample_ack => writeEthernetHeaderToMem_CP_1496_elements(18), 
          phi_update_req => writeEthernetHeaderToMem_CP_1496_elements(19), 
          phi_update_ack => writeEthernetHeaderToMem_CP_1496_elements(20), 
          phi_mux_ack => writeEthernetHeaderToMem_CP_1496_elements(25), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_1265_phi_seq_1623_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= writeEthernetHeaderToMem_CP_1496_elements(42);
      writeEthernetHeaderToMem_CP_1496_elements(45)<= src_sample_reqs(0);
      src_sample_acks(0)  <= writeEthernetHeaderToMem_CP_1496_elements(45);
      writeEthernetHeaderToMem_CP_1496_elements(46)<= src_update_reqs(0);
      src_update_acks(0)  <= writeEthernetHeaderToMem_CP_1496_elements(47);
      writeEthernetHeaderToMem_CP_1496_elements(43) <= phi_mux_reqs(0);
      triggers(1)  <= writeEthernetHeaderToMem_CP_1496_elements(40);
      writeEthernetHeaderToMem_CP_1496_elements(49)<= src_sample_reqs(1);
      src_sample_acks(1)  <= writeEthernetHeaderToMem_CP_1496_elements(51);
      writeEthernetHeaderToMem_CP_1496_elements(50)<= src_update_reqs(1);
      src_update_acks(1)  <= writeEthernetHeaderToMem_CP_1496_elements(52);
      writeEthernetHeaderToMem_CP_1496_elements(41) <= phi_mux_reqs(1);
      phi_stmt_1265_phi_seq_1623 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1265_phi_seq_1623") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => writeEthernetHeaderToMem_CP_1496_elements(11), 
          phi_sample_ack => writeEthernetHeaderToMem_CP_1496_elements(38), 
          phi_update_req => writeEthernetHeaderToMem_CP_1496_elements(13), 
          phi_update_ack => writeEthernetHeaderToMem_CP_1496_elements(39), 
          phi_mux_ack => writeEthernetHeaderToMem_CP_1496_elements(44), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1521_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= writeEthernetHeaderToMem_CP_1496_elements(7);
        preds(1)  <= writeEthernetHeaderToMem_CP_1496_elements(8);
        entry_tmerge_1521 : transition_merge -- 
          generic map(name => " entry_tmerge_1521")
          port map (preds => preds, symbol_out => writeEthernetHeaderToMem_CP_1496_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u36_u36_1263_wire : std_logic_vector(35 downto 0);
    signal I_1265 : std_logic_vector(3 downto 0);
    signal RPIPE_nic_rx_to_header_1272_wire : std_logic_vector(72 downto 0);
    signal ULE_u4_u1_1307_wire : std_logic_vector(0 downto 0);
    signal buf_position_1259 : std_logic_vector(35 downto 0);
    signal ethernet_header_1270 : std_logic_vector(72 downto 0);
    signal ignore_return_1293 : std_logic_vector(63 downto 0);
    signal konst_1262_wire_constant : std_logic_vector(35 downto 0);
    signal konst_1296_wire_constant : std_logic_vector(3 downto 0);
    signal konst_1301_wire_constant : std_logic_vector(35 downto 0);
    signal konst_1306_wire_constant : std_logic_vector(3 downto 0);
    signal nI_1298 : std_logic_vector(3 downto 0);
    signal nI_1298_1269_buffered : std_logic_vector(3 downto 0);
    signal nbuf_position_1303 : std_logic_vector(35 downto 0);
    signal nbuf_position_1303_1264_buffered : std_logic_vector(35 downto 0);
    signal type_cast_1268_wire_constant : std_logic_vector(3 downto 0);
    signal type_cast_1286_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1288_wire_constant : std_logic_vector(0 downto 0);
    signal wdata_1280 : std_logic_vector(63 downto 0);
    signal wkeep_1284 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    konst_1262_wire_constant <= "000000000000000000000000000000001000";
    konst_1296_wire_constant <= "0001";
    konst_1301_wire_constant <= "000000000000000000000000000000001000";
    konst_1306_wire_constant <= "0001";
    type_cast_1268_wire_constant <= "0000";
    type_cast_1286_wire_constant <= "0";
    type_cast_1288_wire_constant <= "0";
    phi_stmt_1259: Block -- phi operator 
      signal idata: std_logic_vector(71 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= ADD_u36_u36_1263_wire & nbuf_position_1303_1264_buffered;
      req <= phi_stmt_1259_req_0 & phi_stmt_1259_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1259",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 36) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1259_ack_0,
          idata => idata,
          odata => buf_position_1259,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1259
    phi_stmt_1265: Block -- phi operator 
      signal idata: std_logic_vector(7 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_1268_wire_constant & nI_1298_1269_buffered;
      req <= phi_stmt_1265_req_0 & phi_stmt_1265_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1265",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 4) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1265_ack_0,
          idata => idata,
          odata => I_1265,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1265
    -- flow-through slice operator slice_1279_inst
    wdata_1280 <= ethernet_header_1270(71 downto 8);
    -- flow-through slice operator slice_1283_inst
    wkeep_1284 <= ethernet_header_1270(7 downto 0);
    W_buf_position_out_1309_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_buf_position_out_1309_inst_req_0;
      W_buf_position_out_1309_inst_ack_0<= wack(0);
      rreq(0) <= W_buf_position_out_1309_inst_req_1;
      W_buf_position_out_1309_inst_ack_1<= rack(0);
      W_buf_position_out_1309_inst : InterlockBuffer generic map ( -- 
        name => "W_buf_position_out_1309_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => buf_position_1259,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => buf_position_out_buffer,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nI_1298_1269_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nI_1298_1269_buf_req_0;
      nI_1298_1269_buf_ack_0<= wack(0);
      rreq(0) <= nI_1298_1269_buf_req_1;
      nI_1298_1269_buf_ack_1<= rack(0);
      nI_1298_1269_buf : InterlockBuffer generic map ( -- 
        name => "nI_1298_1269_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 4,
        out_data_width => 4,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nI_1298,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nI_1298_1269_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nbuf_position_1303_1264_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nbuf_position_1303_1264_buf_req_0;
      nbuf_position_1303_1264_buf_ack_0<= wack(0);
      rreq(0) <= nbuf_position_1303_1264_buf_req_1;
      nbuf_position_1303_1264_buf_ack_1<= rack(0);
      nbuf_position_1303_1264_buf : InterlockBuffer generic map ( -- 
        name => "nbuf_position_1303_1264_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nbuf_position_1303,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nbuf_position_1303_1264_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_1270
    process(RPIPE_nic_rx_to_header_1272_wire) -- 
      variable tmp_var : std_logic_vector(72 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 72 downto 0) := RPIPE_nic_rx_to_header_1272_wire(72 downto 0);
      ethernet_header_1270 <= tmp_var; -- 
    end process;
    do_while_stmt_1257_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= ULE_u4_u1_1307_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1257_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1257_branch_req_0,
          ack0 => do_while_stmt_1257_branch_ack_0,
          ack1 => do_while_stmt_1257_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u36_u36_1263_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= buf_pointer_buffer;
      ADD_u36_u36_1263_wire <= data_out(35 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u36_u36_1263_inst_req_0;
      ADD_u36_u36_1263_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u36_u36_1263_inst_req_1;
      ADD_u36_u36_1263_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 36,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 36,
          constant_operand => "000000000000000000000000000000001000",
          constant_width => 36,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- binary operator ADD_u36_u36_1302_inst
    process(buf_position_1259) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(buf_position_1259, konst_1301_wire_constant, tmp_var);
      nbuf_position_1303 <= tmp_var; --
    end process;
    -- binary operator ADD_u4_u4_1297_inst
    process(I_1265) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApIntAdd_proc(I_1265, konst_1296_wire_constant, tmp_var);
      nI_1298 <= tmp_var; --
    end process;
    -- binary operator ULE_u4_u1_1307_inst
    process(nI_1298) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUle_proc(nI_1298, konst_1306_wire_constant, tmp_var);
      ULE_u4_u1_1307_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_nic_rx_to_header_1272_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(72 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_nic_rx_to_header_1272_inst_req_0;
      RPIPE_nic_rx_to_header_1272_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_nic_rx_to_header_1272_inst_req_1;
      RPIPE_nic_rx_to_header_1272_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_nic_rx_to_header_1272_wire <= data_out(72 downto 0);
      nic_rx_to_header_read_0_gI: SplitGuardInterface generic map(name => "nic_rx_to_header_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      nic_rx_to_header_read_0: InputPortRevised -- 
        generic map ( name => "nic_rx_to_header_read_0", data_width => 73,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => nic_rx_to_header_pipe_read_req(0),
          oack => nic_rx_to_header_pipe_read_ack(0),
          odata => nic_rx_to_header_pipe_read_data(72 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared call operator group (0) : call_stmt_1293_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1293_call_req_0;
      call_stmt_1293_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1293_call_req_1;
      call_stmt_1293_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1286_wire_constant & type_cast_1288_wire_constant & wkeep_1284 & buf_position_1259 & wdata_1280;
      ignore_return_1293 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 3,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end writeEthernetHeaderToMem_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.nic_system_global_package.all;
entity writePayloadToMem is -- 
  generic (tag_length : integer); 
  port ( -- 
    base_buf_pointer : in  std_logic_vector(35 downto 0);
    buf_pointer : in  std_logic_vector(35 downto 0);
    packet_size_32 : out  std_logic_vector(10 downto 0);
    bad_packet_identifier : out  std_logic_vector(0 downto 0);
    last_keep : out  std_logic_vector(7 downto 0);
    nic_rx_to_packet_pipe_read_req : out  std_logic_vector(0 downto 0);
    nic_rx_to_packet_pipe_read_ack : in   std_logic_vector(0 downto 0);
    nic_rx_to_packet_pipe_read_data : in   std_logic_vector(72 downto 0);
    accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_call_acks : in   std_logic_vector(0 downto 0);
    accessMemory_call_data : out  std_logic_vector(109 downto 0);
    accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
    accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
    accessMemory_return_acks : in   std_logic_vector(0 downto 0);
    accessMemory_return_data : in   std_logic_vector(63 downto 0);
    accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity writePayloadToMem;
architecture writePayloadToMem_arch of writePayloadToMem is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 72)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 20)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal base_buf_pointer_buffer :  std_logic_vector(35 downto 0);
  signal base_buf_pointer_update_enable: Boolean;
  signal buf_pointer_buffer :  std_logic_vector(35 downto 0);
  signal buf_pointer_update_enable: Boolean;
  -- output port buffer signals
  signal packet_size_32_buffer :  std_logic_vector(10 downto 0);
  signal packet_size_32_update_enable: Boolean;
  signal bad_packet_identifier_buffer :  std_logic_vector(0 downto 0);
  signal bad_packet_identifier_update_enable: Boolean;
  signal last_keep_buffer :  std_logic_vector(7 downto 0);
  signal last_keep_update_enable: Boolean;
  signal writePayloadToMem_CP_1683_start: Boolean;
  signal writePayloadToMem_CP_1683_symbol: Boolean;
  -- volatile/operator module components. 
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal do_while_stmt_1321_branch_req_0 : boolean;
  signal phi_stmt_1323_req_0 : boolean;
  signal phi_stmt_1323_req_1 : boolean;
  signal phi_stmt_1323_ack_0 : boolean;
  signal nbuf_position_1363_1325_buf_req_0 : boolean;
  signal nbuf_position_1363_1325_buf_ack_0 : boolean;
  signal nbuf_position_1363_1325_buf_req_1 : boolean;
  signal nbuf_position_1363_1325_buf_ack_1 : boolean;
  signal ADD_u36_u36_1328_inst_req_0 : boolean;
  signal ADD_u36_u36_1328_inst_ack_0 : boolean;
  signal ADD_u36_u36_1328_inst_req_1 : boolean;
  signal ADD_u36_u36_1328_inst_ack_1 : boolean;
  signal RPIPE_nic_rx_to_packet_1331_inst_req_0 : boolean;
  signal RPIPE_nic_rx_to_packet_1331_inst_ack_0 : boolean;
  signal RPIPE_nic_rx_to_packet_1331_inst_req_1 : boolean;
  signal RPIPE_nic_rx_to_packet_1331_inst_ack_1 : boolean;
  signal call_stmt_1358_call_req_0 : boolean;
  signal call_stmt_1358_call_ack_0 : boolean;
  signal call_stmt_1358_call_req_1 : boolean;
  signal call_stmt_1358_call_ack_1 : boolean;
  signal do_while_stmt_1321_branch_ack_0 : boolean;
  signal do_while_stmt_1321_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "writePayloadToMem_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 72) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(35 downto 0) <= base_buf_pointer;
  base_buf_pointer_buffer <= in_buffer_data_out(35 downto 0);
  in_buffer_data_in(71 downto 36) <= buf_pointer;
  buf_pointer_buffer <= in_buffer_data_out(71 downto 36);
  in_buffer_data_in(tag_length + 71 downto 72) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 71 downto 72);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  writePayloadToMem_CP_1683_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "writePayloadToMem_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 20) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(10 downto 0) <= packet_size_32_buffer;
  packet_size_32 <= out_buffer_data_out(10 downto 0);
  out_buffer_data_in(11 downto 11) <= bad_packet_identifier_buffer;
  bad_packet_identifier <= out_buffer_data_out(11 downto 11);
  out_buffer_data_in(19 downto 12) <= last_keep_buffer;
  last_keep <= out_buffer_data_out(19 downto 12);
  out_buffer_data_in(tag_length + 19 downto 20) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 19 downto 20);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writePayloadToMem_CP_1683_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= writePayloadToMem_CP_1683_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writePayloadToMem_CP_1683_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  writePayloadToMem_CP_1683: Block -- control-path 
    signal writePayloadToMem_CP_1683_elements: BooleanArray(47 downto 0);
    -- 
  begin -- 
    writePayloadToMem_CP_1683_elements(0) <= writePayloadToMem_CP_1683_start;
    writePayloadToMem_CP_1683_symbol <= writePayloadToMem_CP_1683_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_1320/branch_block_stmt_1320__entry__
      -- CP-element group 0: 	 branch_block_stmt_1320/do_while_stmt_1321__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_1320/$entry
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	47 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 $exit
      -- CP-element group 1: 	 branch_block_stmt_1320/branch_block_stmt_1320__exit__
      -- CP-element group 1: 	 branch_block_stmt_1320/do_while_stmt_1321__exit__
      -- CP-element group 1: 	 branch_block_stmt_1320/$exit
      -- CP-element group 1: 	 assign_stmt_1376_to_assign_stmt_1391/$entry
      -- CP-element group 1: 	 assign_stmt_1376_to_assign_stmt_1391/$exit
      -- 
    writePayloadToMem_CP_1683_elements(1) <= writePayloadToMem_CP_1683_elements(47);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_1320/do_while_stmt_1321/$entry
      -- CP-element group 2: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321__entry__
      -- 
    writePayloadToMem_CP_1683_elements(2) <= writePayloadToMem_CP_1683_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	47 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321__exit__
      -- 
    -- Element group writePayloadToMem_CP_1683_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_1320/do_while_stmt_1321/loop_back
      -- 
    -- Element group writePayloadToMem_CP_1683_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	45 
    -- CP-element group 5: 	46 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_1320/do_while_stmt_1321/condition_done
      -- CP-element group 5: 	 branch_block_stmt_1320/do_while_stmt_1321/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_1320/do_while_stmt_1321/loop_taken/$entry
      -- 
    writePayloadToMem_CP_1683_elements(5) <= writePayloadToMem_CP_1683_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	44 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_1320/do_while_stmt_1321/loop_body_done
      -- 
    writePayloadToMem_CP_1683_elements(6) <= writePayloadToMem_CP_1683_elements(44);
    -- CP-element group 7:  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	19 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/back_edge_to_loop_body
      -- 
    writePayloadToMem_CP_1683_elements(7) <= writePayloadToMem_CP_1683_elements(4);
    -- CP-element group 8:  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	21 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/first_time_through_loop_body
      -- 
    writePayloadToMem_CP_1683_elements(8) <= writePayloadToMem_CP_1683_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	43 
    -- CP-element group 9: 	34 
    -- CP-element group 9: 	11 
    -- CP-element group 9: 	15 
    -- CP-element group 9: 	16 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/loop_body_start
      -- CP-element group 9: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1329_sample_start_
      -- 
    -- Element group writePayloadToMem_CP_1683_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	43 
    -- CP-element group 10: 	14 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/condition_evaluated
      -- 
    condition_evaluated_1707_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_1707_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_1683_elements(10), ack => do_while_stmt_1321_branch_req_0); -- 
    writePayloadToMem_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1683_elements(43) & writePayloadToMem_CP_1683_elements(14);
      gj_writePayloadToMem_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1683_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	9 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	14 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	35 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1323_sample_start__ps
      -- CP-element group 11: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/aggregated_phi_sample_req
      -- 
    writePayloadToMem_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1683_elements(15) & writePayloadToMem_CP_1683_elements(9) & writePayloadToMem_CP_1683_elements(14);
      gj_writePayloadToMem_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1683_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	37 
    -- CP-element group 12: 	17 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	44 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	15 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1323_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1329_sample_completed_
      -- 
    writePayloadToMem_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1683_elements(37) & writePayloadToMem_CP_1683_elements(17);
      gj_writePayloadToMem_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1683_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	34 
    -- CP-element group 13: 	16 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	36 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1323_update_start__ps
      -- CP-element group 13: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/aggregated_phi_update_req
      -- 
    writePayloadToMem_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1683_elements(34) & writePayloadToMem_CP_1683_elements(16);
      gj_writePayloadToMem_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1683_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	38 
    -- CP-element group 14: 	18 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	10 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	11 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/aggregated_phi_update_ack
      -- 
    writePayloadToMem_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1683_elements(38) & writePayloadToMem_CP_1683_elements(18);
      gj_writePayloadToMem_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1683_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	9 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	12 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1323_sample_start_
      -- 
    writePayloadToMem_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1683_elements(9) & writePayloadToMem_CP_1683_elements(12);
      gj_writePayloadToMem_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1683_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	41 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1323_update_start_
      -- 
    writePayloadToMem_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1683_elements(9) & writePayloadToMem_CP_1683_elements(41);
      gj_writePayloadToMem_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1683_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1323_sample_completed__ps
      -- 
    -- Element group writePayloadToMem_CP_1683_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: 	39 
    -- CP-element group 18:  members (2) 
      -- CP-element group 18: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1323_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1323_update_completed__ps
      -- 
    -- Element group writePayloadToMem_CP_1683_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	7 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1323_loopback_trigger
      -- 
    writePayloadToMem_CP_1683_elements(19) <= writePayloadToMem_CP_1683_elements(7);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1323_loopback_sample_req
      -- CP-element group 20: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1323_loopback_sample_req_ps
      -- 
    phi_stmt_1323_loopback_sample_req_1722_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1323_loopback_sample_req_1722_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_1683_elements(20), ack => phi_stmt_1323_req_0); -- 
    -- Element group writePayloadToMem_CP_1683_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	8 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1323_entry_trigger
      -- 
    writePayloadToMem_CP_1683_elements(21) <= writePayloadToMem_CP_1683_elements(8);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1323_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1323_entry_sample_req_ps
      -- 
    phi_stmt_1323_entry_sample_req_1725_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_1323_entry_sample_req_1725_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_1683_elements(22), ack => phi_stmt_1323_req_1); -- 
    -- Element group writePayloadToMem_CP_1683_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1323_phi_mux_ack
      -- CP-element group 23: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1323_phi_mux_ack_ps
      -- 
    phi_stmt_1323_phi_mux_ack_1728_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_1323_ack_0, ack => writePayloadToMem_CP_1683_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_nbuf_position_1325_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_nbuf_position_1325_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_nbuf_position_1325_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_nbuf_position_1325_Sample/req
      -- 
    req_1741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_1683_elements(24), ack => nbuf_position_1363_1325_buf_req_0); -- 
    -- Element group writePayloadToMem_CP_1683_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_nbuf_position_1325_update_start__ps
      -- CP-element group 25: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_nbuf_position_1325_update_start_
      -- CP-element group 25: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_nbuf_position_1325_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_nbuf_position_1325_Update/req
      -- 
    req_1746_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_1746_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_1683_elements(25), ack => nbuf_position_1363_1325_buf_req_1); -- 
    -- Element group writePayloadToMem_CP_1683_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_nbuf_position_1325_sample_completed__ps
      -- CP-element group 26: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_nbuf_position_1325_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_nbuf_position_1325_Sample/$exit
      -- CP-element group 26: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_nbuf_position_1325_Sample/ack
      -- 
    ack_1742_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nbuf_position_1363_1325_buf_ack_0, ack => writePayloadToMem_CP_1683_elements(26)); -- 
    -- CP-element group 27:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_nbuf_position_1325_update_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_nbuf_position_1325_update_completed_
      -- CP-element group 27: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_nbuf_position_1325_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/R_nbuf_position_1325_Update/ack
      -- 
    ack_1747_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nbuf_position_1363_1325_buf_ack_1, ack => writePayloadToMem_CP_1683_elements(27)); -- 
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/ADD_u36_u36_1328_sample_start__ps
      -- 
    -- Element group writePayloadToMem_CP_1683_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/ADD_u36_u36_1328_update_start__ps
      -- 
    -- Element group writePayloadToMem_CP_1683_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: marked-predecessors 
    -- CP-element group 30: 	32 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (3) 
      -- CP-element group 30: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/ADD_u36_u36_1328_sample_start_
      -- CP-element group 30: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/ADD_u36_u36_1328_Sample/$entry
      -- CP-element group 30: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/ADD_u36_u36_1328_Sample/rr
      -- 
    rr_1759_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1759_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_1683_elements(30), ack => ADD_u36_u36_1328_inst_req_0); -- 
    writePayloadToMem_cp_element_group_30: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_30"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1683_elements(28) & writePayloadToMem_CP_1683_elements(32);
      gj_writePayloadToMem_cp_element_group_30 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1683_elements(30), clk => clk, reset => reset); --
    end block;
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	33 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/ADD_u36_u36_1328_update_start_
      -- CP-element group 31: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/ADD_u36_u36_1328_Update/$entry
      -- CP-element group 31: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/ADD_u36_u36_1328_Update/cr
      -- 
    cr_1764_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1764_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_1683_elements(31), ack => ADD_u36_u36_1328_inst_req_1); -- 
    writePayloadToMem_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1683_elements(29) & writePayloadToMem_CP_1683_elements(33);
      gj_writePayloadToMem_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1683_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: successors 
    -- CP-element group 32: marked-successors 
    -- CP-element group 32: 	30 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/ADD_u36_u36_1328_sample_completed__ps
      -- CP-element group 32: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/ADD_u36_u36_1328_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/ADD_u36_u36_1328_Sample/$exit
      -- CP-element group 32: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/ADD_u36_u36_1328_Sample/ra
      -- 
    ra_1760_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 32_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_1328_inst_ack_0, ack => writePayloadToMem_CP_1683_elements(32)); -- 
    -- CP-element group 33:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	31 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/ADD_u36_u36_1328_update_completed__ps
      -- CP-element group 33: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/ADD_u36_u36_1328_update_completed_
      -- CP-element group 33: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/ADD_u36_u36_1328_Update/$exit
      -- CP-element group 33: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/ADD_u36_u36_1328_Update/ca
      -- 
    ca_1765_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => ADD_u36_u36_1328_inst_ack_1, ack => writePayloadToMem_CP_1683_elements(33)); -- 
    -- CP-element group 34:  join  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	9 
    -- CP-element group 34: marked-predecessors 
    -- CP-element group 34: 	41 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	13 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1329_update_start_
      -- 
    writePayloadToMem_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1683_elements(9) & writePayloadToMem_CP_1683_elements(41);
      gj_writePayloadToMem_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1683_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	11 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	38 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	37 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_nic_rx_to_packet_1331_sample_start_
      -- CP-element group 35: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_nic_rx_to_packet_1331_Sample/$entry
      -- CP-element group 35: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_nic_rx_to_packet_1331_Sample/rr
      -- 
    rr_1778_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_1778_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_1683_elements(35), ack => RPIPE_nic_rx_to_packet_1331_inst_req_0); -- 
    writePayloadToMem_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1683_elements(11) & writePayloadToMem_CP_1683_elements(38);
      gj_writePayloadToMem_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1683_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	13 
    -- CP-element group 36: 	37 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_nic_rx_to_packet_1331_update_start_
      -- CP-element group 36: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_nic_rx_to_packet_1331_Update/$entry
      -- CP-element group 36: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_nic_rx_to_packet_1331_Update/cr
      -- 
    cr_1783_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_1783_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_1683_elements(36), ack => RPIPE_nic_rx_to_packet_1331_inst_req_1); -- 
    writePayloadToMem_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1683_elements(13) & writePayloadToMem_CP_1683_elements(37);
      gj_writePayloadToMem_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1683_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	35 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	36 
    -- CP-element group 37: 	12 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_nic_rx_to_packet_1331_sample_completed_
      -- CP-element group 37: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_nic_rx_to_packet_1331_Sample/$exit
      -- CP-element group 37: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_nic_rx_to_packet_1331_Sample/ra
      -- 
    ra_1779_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 37_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_nic_rx_to_packet_1331_inst_ack_0, ack => writePayloadToMem_CP_1683_elements(37)); -- 
    -- CP-element group 38:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	14 
    -- CP-element group 38: 	39 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	35 
    -- CP-element group 38:  members (4) 
      -- CP-element group 38: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/phi_stmt_1329_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_nic_rx_to_packet_1331_update_completed_
      -- CP-element group 38: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_nic_rx_to_packet_1331_Update/$exit
      -- CP-element group 38: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/RPIPE_nic_rx_to_packet_1331_Update/ca
      -- 
    ca_1784_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_nic_rx_to_packet_1331_inst_ack_1, ack => writePayloadToMem_CP_1683_elements(38)); -- 
    -- CP-element group 39:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	38 
    -- CP-element group 39: 	18 
    -- CP-element group 39: marked-predecessors 
    -- CP-element group 39: 	41 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	41 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/call_stmt_1358_sample_start_
      -- CP-element group 39: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/call_stmt_1358_Sample/$entry
      -- CP-element group 39: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/call_stmt_1358_Sample/crr
      -- 
    crr_1792_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_1792_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_1683_elements(39), ack => call_stmt_1358_call_req_0); -- 
    writePayloadToMem_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1683_elements(38) & writePayloadToMem_CP_1683_elements(18) & writePayloadToMem_CP_1683_elements(41);
      gj_writePayloadToMem_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1683_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: marked-predecessors 
    -- CP-element group 40: 	42 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	42 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/call_stmt_1358_update_start_
      -- CP-element group 40: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/call_stmt_1358_Update/$entry
      -- CP-element group 40: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/call_stmt_1358_Update/ccr
      -- 
    ccr_1797_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_1797_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writePayloadToMem_CP_1683_elements(40), ack => call_stmt_1358_call_req_1); -- 
    writePayloadToMem_cp_element_group_40: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_40"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= writePayloadToMem_CP_1683_elements(42);
      gj_writePayloadToMem_cp_element_group_40 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1683_elements(40), clk => clk, reset => reset); --
    end block;
    -- CP-element group 41:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	39 
    -- CP-element group 41: successors 
    -- CP-element group 41: marked-successors 
    -- CP-element group 41: 	34 
    -- CP-element group 41: 	16 
    -- CP-element group 41: 	39 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/call_stmt_1358_sample_completed_
      -- CP-element group 41: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/call_stmt_1358_Sample/$exit
      -- CP-element group 41: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/call_stmt_1358_Sample/cra
      -- 
    cra_1793_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 41_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1358_call_ack_0, ack => writePayloadToMem_CP_1683_elements(41)); -- 
    -- CP-element group 42:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	40 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	44 
    -- CP-element group 42: marked-successors 
    -- CP-element group 42: 	40 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/call_stmt_1358_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/call_stmt_1358_Update/$exit
      -- CP-element group 42: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/call_stmt_1358_Update/cca
      -- 
    cca_1798_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_1358_call_ack_1, ack => writePayloadToMem_CP_1683_elements(42)); -- 
    -- CP-element group 43:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	9 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	10 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group writePayloadToMem_CP_1683_elements(43) is a control-delay.
    cp_element_43_delay: control_delay_element  generic map(name => " 43_delay", delay_value => 1)  port map(req => writePayloadToMem_CP_1683_elements(9), ack => writePayloadToMem_CP_1683_elements(43), clk => clk, reset =>reset);
    -- CP-element group 44:  join  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	42 
    -- CP-element group 44: 	12 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	6 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_1320/do_while_stmt_1321/do_while_stmt_1321_loop_body/$exit
      -- 
    writePayloadToMem_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writePayloadToMem_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writePayloadToMem_CP_1683_elements(42) & writePayloadToMem_CP_1683_elements(12);
      gj_writePayloadToMem_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writePayloadToMem_CP_1683_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  transition  input  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	5 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_1320/do_while_stmt_1321/loop_exit/$exit
      -- CP-element group 45: 	 branch_block_stmt_1320/do_while_stmt_1321/loop_exit/ack
      -- 
    ack_1803_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1321_branch_ack_0, ack => writePayloadToMem_CP_1683_elements(45)); -- 
    -- CP-element group 46:  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	5 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_1320/do_while_stmt_1321/loop_taken/$exit
      -- CP-element group 46: 	 branch_block_stmt_1320/do_while_stmt_1321/loop_taken/ack
      -- 
    ack_1807_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_1321_branch_ack_1, ack => writePayloadToMem_CP_1683_elements(46)); -- 
    -- CP-element group 47:  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	3 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	1 
    -- CP-element group 47:  members (1) 
      -- CP-element group 47: 	 branch_block_stmt_1320/do_while_stmt_1321/$exit
      -- 
    writePayloadToMem_CP_1683_elements(47) <= writePayloadToMem_CP_1683_elements(3);
    writePayloadToMem_do_while_stmt_1321_terminator_1808: loop_terminator -- 
      generic map (name => " writePayloadToMem_do_while_stmt_1321_terminator_1808", max_iterations_in_flight =>15) 
      port map(loop_body_exit => writePayloadToMem_CP_1683_elements(6),loop_continue => writePayloadToMem_CP_1683_elements(46),loop_terminate => writePayloadToMem_CP_1683_elements(45),loop_back => writePayloadToMem_CP_1683_elements(4),loop_exit => writePayloadToMem_CP_1683_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_1323_phi_seq_1766_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= writePayloadToMem_CP_1683_elements(19);
      writePayloadToMem_CP_1683_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= writePayloadToMem_CP_1683_elements(26);
      writePayloadToMem_CP_1683_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= writePayloadToMem_CP_1683_elements(27);
      writePayloadToMem_CP_1683_elements(20) <= phi_mux_reqs(0);
      triggers(1)  <= writePayloadToMem_CP_1683_elements(21);
      writePayloadToMem_CP_1683_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= writePayloadToMem_CP_1683_elements(32);
      writePayloadToMem_CP_1683_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= writePayloadToMem_CP_1683_elements(33);
      writePayloadToMem_CP_1683_elements(22) <= phi_mux_reqs(1);
      phi_stmt_1323_phi_seq_1766 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_1323_phi_seq_1766") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => writePayloadToMem_CP_1683_elements(11), 
          phi_sample_ack => writePayloadToMem_CP_1683_elements(17), 
          phi_update_req => writePayloadToMem_CP_1683_elements(13), 
          phi_update_ack => writePayloadToMem_CP_1683_elements(18), 
          phi_mux_ack => writePayloadToMem_CP_1683_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_1708_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= writePayloadToMem_CP_1683_elements(7);
        preds(1)  <= writePayloadToMem_CP_1683_elements(8);
        entry_tmerge_1708 : transition_merge -- 
          generic map(name => " entry_tmerge_1708")
          port map (preds => preds, symbol_out => writePayloadToMem_CP_1683_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u36_u36_1328_wire : std_logic_vector(35 downto 0);
    signal EQ_u64_u1_1371_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_1374_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1366_wire : std_logic_vector(0 downto 0);
    signal RPIPE_nic_rx_to_packet_1331_wire : std_logic_vector(72 downto 0);
    signal R_BAD_PACKET_DATA_1370_wire_constant : std_logic_vector(63 downto 0);
    signal SUB_u36_u36_1380_wire : std_logic_vector(35 downto 0);
    signal buf_position_1323 : std_logic_vector(35 downto 0);
    signal ignore_return_1358 : std_logic_vector(63 downto 0);
    signal konst_1327_wire_constant : std_logic_vector(35 downto 0);
    signal konst_1361_wire_constant : std_logic_vector(35 downto 0);
    signal konst_1373_wire_constant : std_logic_vector(7 downto 0);
    signal last_bit_1336 : std_logic_vector(0 downto 0);
    signal nbuf_position_1363 : std_logic_vector(35 downto 0);
    signal nbuf_position_1363_1325_buffered : std_logic_vector(35 downto 0);
    signal packet_size_11_1382 : std_logic_vector(10 downto 0);
    signal payload_data_1329 : std_logic_vector(72 downto 0);
    signal type_cast_1351_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_1353_wire_constant : std_logic_vector(0 downto 0);
    signal wdata_1340 : std_logic_vector(63 downto 0);
    signal wkeep_1344 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    R_BAD_PACKET_DATA_1370_wire_constant <= "1111111111111111111111111111111111111111111111111111111111111111";
    konst_1327_wire_constant <= "000000000000000000000000000000001000";
    konst_1361_wire_constant <= "000000000000000000000000000000001000";
    konst_1373_wire_constant <= "00000000";
    type_cast_1351_wire_constant <= "0";
    type_cast_1353_wire_constant <= "0";
    phi_stmt_1323: Block -- phi operator 
      signal idata: std_logic_vector(71 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= nbuf_position_1363_1325_buffered & ADD_u36_u36_1328_wire;
      req <= phi_stmt_1323_req_0 & phi_stmt_1323_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_1323",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 36) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_1323_ack_0,
          idata => idata,
          odata => buf_position_1323,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_1323
    -- flow-through slice operator slice_1335_inst
    last_bit_1336 <= payload_data_1329(72 downto 72);
    -- flow-through slice operator slice_1339_inst
    wdata_1340 <= payload_data_1329(71 downto 8);
    -- flow-through slice operator slice_1343_inst
    wkeep_1344 <= payload_data_1329(7 downto 0);
    -- interlock W_last_keep_1389_inst
    process(wkeep_1344) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := wkeep_1344(7 downto 0);
      last_keep_buffer <= tmp_var; -- 
    end process;
    -- interlock W_packet_size_32_1383_inst
    process(packet_size_11_1382) -- 
      variable tmp_var : std_logic_vector(10 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 10 downto 0) := packet_size_11_1382(10 downto 0);
      packet_size_32_buffer <= tmp_var; -- 
    end process;
    nbuf_position_1363_1325_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nbuf_position_1363_1325_buf_req_0;
      nbuf_position_1363_1325_buf_ack_0<= wack(0);
      rreq(0) <= nbuf_position_1363_1325_buf_req_1;
      nbuf_position_1363_1325_buf_ack_1<= rack(0);
      nbuf_position_1363_1325_buf : InterlockBuffer generic map ( -- 
        name => "nbuf_position_1363_1325_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 36,
        out_data_width => 36,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nbuf_position_1363,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nbuf_position_1363_1325_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock ssrc_phi_stmt_1329
    process(RPIPE_nic_rx_to_packet_1331_wire) -- 
      variable tmp_var : std_logic_vector(72 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 72 downto 0) := RPIPE_nic_rx_to_packet_1331_wire(72 downto 0);
      payload_data_1329 <= tmp_var; -- 
    end process;
    -- interlock type_cast_1381_inst
    process(SUB_u36_u36_1380_wire) -- 
      variable tmp_var : std_logic_vector(10 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 10 downto 0) := SUB_u36_u36_1380_wire(10 downto 0);
      packet_size_11_1382 <= tmp_var; -- 
    end process;
    do_while_stmt_1321_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= NOT_u1_u1_1366_wire;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_1321_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_1321_branch_req_0,
          ack0 => do_while_stmt_1321_branch_ack_0,
          ack1 => do_while_stmt_1321_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- shared split operator group (0) : ADD_u36_u36_1328_inst 
    ApIntAdd_group_0: Block -- 
      signal data_in: std_logic_vector(35 downto 0);
      signal data_out: std_logic_vector(35 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= buf_pointer_buffer;
      ADD_u36_u36_1328_wire <= data_out(35 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= ADD_u36_u36_1328_inst_req_0;
      ADD_u36_u36_1328_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= ADD_u36_u36_1328_inst_req_1;
      ADD_u36_u36_1328_inst_ack_1 <= ackR_unguarded(0);
      ApIntAdd_group_0_gI: SplitGuardInterface generic map(name => "ApIntAdd_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAdd",
          name => "ApIntAdd_group_0",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 36,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 0, 
          num_inputs    => 1,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 36,
          constant_operand => "000000000000000000000000000000001000",
          constant_width => 36,
          buffering  => 1,
          flow_through => false,
          full_rate  => true,
          use_constant  => true
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 0
    -- binary operator ADD_u36_u36_1362_inst
    process(buf_position_1323) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntAdd_proc(buf_position_1323, konst_1361_wire_constant, tmp_var);
      nbuf_position_1363 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1375_inst
    process(EQ_u64_u1_1371_wire, EQ_u8_u1_1374_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u64_u1_1371_wire, EQ_u8_u1_1374_wire, tmp_var);
      bad_packet_identifier_buffer <= tmp_var; --
    end process;
    -- binary operator EQ_u64_u1_1371_inst
    process(wdata_1340) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(wdata_1340, R_BAD_PACKET_DATA_1370_wire_constant, tmp_var);
      EQ_u64_u1_1371_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_1374_inst
    process(wkeep_1344) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(wkeep_1344, konst_1373_wire_constant, tmp_var);
      EQ_u8_u1_1374_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1366_inst
    process(last_bit_1336) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", last_bit_1336, tmp_var);
      NOT_u1_u1_1366_wire <= tmp_var; -- 
    end process;
    -- binary operator SUB_u36_u36_1380_inst
    process(buf_position_1323, base_buf_pointer_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApIntSub_proc(buf_position_1323, base_buf_pointer_buffer, tmp_var);
      SUB_u36_u36_1380_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_nic_rx_to_packet_1331_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(72 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_nic_rx_to_packet_1331_inst_req_0;
      RPIPE_nic_rx_to_packet_1331_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_nic_rx_to_packet_1331_inst_req_1;
      RPIPE_nic_rx_to_packet_1331_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_nic_rx_to_packet_1331_wire <= data_out(72 downto 0);
      nic_rx_to_packet_read_0_gI: SplitGuardInterface generic map(name => "nic_rx_to_packet_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      nic_rx_to_packet_read_0: InputPortRevised -- 
        generic map ( name => "nic_rx_to_packet_read_0", data_width => 73,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => nic_rx_to_packet_pipe_read_req(0),
          oack => nic_rx_to_packet_pipe_read_ack(0),
          odata => nic_rx_to_packet_pipe_read_data(72 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared call operator group (0) : call_stmt_1358_call 
    accessMemory_call_group_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_1358_call_req_0;
      call_stmt_1358_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_1358_call_req_1;
      call_stmt_1358_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessMemory_call_group_0_gI: SplitGuardInterface generic map(name => "accessMemory_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_1351_wire_constant & type_cast_1353_wire_constant & wkeep_1344 & buf_position_1323 & wdata_1340;
      ignore_return_1358 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 110,
        owidth => 110,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 3,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessMemory_call_reqs(0),
          ackR => accessMemory_call_acks(0),
          dataR => accessMemory_call_data(109 downto 0),
          tagR => accessMemory_call_tag(2 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 3,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessMemory_return_acks(0), -- cross-over
          ackL => accessMemory_return_reqs(0), -- cross-over
          dataL => accessMemory_return_data(63 downto 0),
          tagL => accessMemory_return_tag(2 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end writePayloadToMem_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
library work;
use work.nic_system_global_package.all;
entity nic_system is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    AFB_NIC_REQUEST_pipe_write_data: in std_logic_vector(73 downto 0);
    AFB_NIC_REQUEST_pipe_write_req : in std_logic_vector(0 downto 0);
    AFB_NIC_REQUEST_pipe_write_ack : out std_logic_vector(0 downto 0);
    AFB_NIC_RESPONSE_pipe_read_data: out std_logic_vector(32 downto 0);
    AFB_NIC_RESPONSE_pipe_read_req : in std_logic_vector(0 downto 0);
    AFB_NIC_RESPONSE_pipe_read_ack : out std_logic_vector(0 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_write_data: in std_logic_vector(64 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_write_req : in std_logic_vector(0 downto 0);
    MEMORY_TO_NIC_RESPONSE_pipe_write_ack : out std_logic_vector(0 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_read_data: out std_logic_vector(109 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_read_req : in std_logic_vector(0 downto 0);
    NIC_TO_MEMORY_REQUEST_pipe_read_ack : out std_logic_vector(0 downto 0);
    enable_mac_pipe_read_data: out std_logic_vector(0 downto 0);
    enable_mac_pipe_read_req : in std_logic_vector(0 downto 0);
    enable_mac_pipe_read_ack : out std_logic_vector(0 downto 0);
    mac_to_nic_data_pipe_write_data: in std_logic_vector(72 downto 0);
    mac_to_nic_data_pipe_write_req : in std_logic_vector(0 downto 0);
    mac_to_nic_data_pipe_write_ack : out std_logic_vector(0 downto 0);
    nic_to_mac_transmit_pipe_pipe_read_data: out std_logic_vector(72 downto 0);
    nic_to_mac_transmit_pipe_pipe_read_req : in std_logic_vector(0 downto 0);
    nic_to_mac_transmit_pipe_pipe_read_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture nic_system_arch  of nic_system is -- system-architecture 
  -- interface signals to connect to memory space memory_space_0
  -- interface signals to connect to memory space memory_space_1
  -- interface signals to connect to memory space memory_space_2
  signal memory_space_2_lr_req :  std_logic_vector(1 downto 0);
  signal memory_space_2_lr_ack : std_logic_vector(1 downto 0);
  signal memory_space_2_lr_addr : std_logic_vector(11 downto 0);
  signal memory_space_2_lr_tag : std_logic_vector(41 downto 0);
  signal memory_space_2_lc_req : std_logic_vector(1 downto 0);
  signal memory_space_2_lc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_2_lc_data : std_logic_vector(63 downto 0);
  signal memory_space_2_lc_tag :  std_logic_vector(5 downto 0);
  signal memory_space_2_sr_req :  std_logic_vector(1 downto 0);
  signal memory_space_2_sr_ack : std_logic_vector(1 downto 0);
  signal memory_space_2_sr_addr : std_logic_vector(11 downto 0);
  signal memory_space_2_sr_data : std_logic_vector(63 downto 0);
  signal memory_space_2_sr_tag : std_logic_vector(41 downto 0);
  signal memory_space_2_sc_req : std_logic_vector(1 downto 0);
  signal memory_space_2_sc_ack :  std_logic_vector(1 downto 0);
  signal memory_space_2_sc_tag :  std_logic_vector(5 downto 0);
  -- declarations related to module AccessRegister
  component AccessRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(3 downto 0);
      register_index : in  std_logic_vector(5 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      rdata : out  std_logic_vector(31 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(32 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(42 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module AccessRegister
  signal AccessRegister_rwbar :  std_logic_vector(0 downto 0);
  signal AccessRegister_bmask :  std_logic_vector(3 downto 0);
  signal AccessRegister_register_index :  std_logic_vector(5 downto 0);
  signal AccessRegister_wdata :  std_logic_vector(31 downto 0);
  signal AccessRegister_rdata :  std_logic_vector(31 downto 0);
  signal AccessRegister_in_args    : std_logic_vector(42 downto 0);
  signal AccessRegister_out_args   : std_logic_vector(31 downto 0);
  signal AccessRegister_tag_in    : std_logic_vector(4 downto 0) := (others => '0');
  signal AccessRegister_tag_out   : std_logic_vector(4 downto 0);
  signal AccessRegister_start_req : std_logic;
  signal AccessRegister_start_ack : std_logic;
  signal AccessRegister_fin_req   : std_logic;
  signal AccessRegister_fin_ack : std_logic;
  -- caller side aggregated signals for module AccessRegister
  signal AccessRegister_call_reqs: std_logic_vector(6 downto 0);
  signal AccessRegister_call_acks: std_logic_vector(6 downto 0);
  signal AccessRegister_return_reqs: std_logic_vector(6 downto 0);
  signal AccessRegister_return_acks: std_logic_vector(6 downto 0);
  signal AccessRegister_call_data: std_logic_vector(300 downto 0);
  signal AccessRegister_call_tag: std_logic_vector(13 downto 0);
  signal AccessRegister_return_data: std_logic_vector(223 downto 0);
  signal AccessRegister_return_tag: std_logic_vector(13 downto 0);
  -- declarations related to module NicRegisterAccessDaemon
  component NicRegisterAccessDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(5 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(5 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(2 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data : in   std_logic_vector(42 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data : out  std_logic_vector(32 downto 0);
      MAC_ENABLE_pipe_write_req : out  std_logic_vector(0 downto 0);
      MAC_ENABLE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      MAC_ENABLE_pipe_write_data : out  std_logic_vector(0 downto 0);
      UpdateRegister_call_reqs : out  std_logic_vector(0 downto 0);
      UpdateRegister_call_acks : in   std_logic_vector(0 downto 0);
      UpdateRegister_call_data : out  std_logic_vector(73 downto 0);
      UpdateRegister_call_tag  :  out  std_logic_vector(0 downto 0);
      UpdateRegister_return_reqs : out  std_logic_vector(0 downto 0);
      UpdateRegister_return_acks : in   std_logic_vector(0 downto 0);
      UpdateRegister_return_data : in   std_logic_vector(31 downto 0);
      UpdateRegister_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module NicRegisterAccessDaemon
  signal NicRegisterAccessDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal NicRegisterAccessDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal NicRegisterAccessDaemon_start_req : std_logic;
  signal NicRegisterAccessDaemon_start_ack : std_logic;
  signal NicRegisterAccessDaemon_fin_req   : std_logic;
  signal NicRegisterAccessDaemon_fin_ack : std_logic;
  -- declarations related to module ReceiveEngineDaemon
  component ReceiveEngineDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      CONTROL_REGISTER : in std_logic_vector(31 downto 0);
      FREE_Q : in std_logic_vector(35 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(5 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_call_data : out  std_logic_vector(36 downto 0);
      popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_return_data : in   std_logic_vector(32 downto 0);
      popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
      pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
      loadBuffer_call_reqs : out  std_logic_vector(0 downto 0);
      loadBuffer_call_acks : in   std_logic_vector(0 downto 0);
      loadBuffer_call_data : out  std_logic_vector(35 downto 0);
      loadBuffer_call_tag  :  out  std_logic_vector(0 downto 0);
      loadBuffer_return_reqs : out  std_logic_vector(0 downto 0);
      loadBuffer_return_acks : in   std_logic_vector(0 downto 0);
      loadBuffer_return_data : in   std_logic_vector(0 downto 0);
      loadBuffer_return_tag :  in   std_logic_vector(0 downto 0);
      populateRxQueue_call_reqs : out  std_logic_vector(0 downto 0);
      populateRxQueue_call_acks : in   std_logic_vector(0 downto 0);
      populateRxQueue_call_data : out  std_logic_vector(35 downto 0);
      populateRxQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      populateRxQueue_return_reqs : out  std_logic_vector(0 downto 0);
      populateRxQueue_return_acks : in   std_logic_vector(0 downto 0);
      populateRxQueue_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module ReceiveEngineDaemon
  signal ReceiveEngineDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal ReceiveEngineDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal ReceiveEngineDaemon_start_req : std_logic;
  signal ReceiveEngineDaemon_start_ack : std_logic;
  signal ReceiveEngineDaemon_fin_req   : std_logic;
  signal ReceiveEngineDaemon_fin_ack : std_logic;
  -- declarations related to module SoftwareRegisterAccessDaemon
  component SoftwareRegisterAccessDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      memory_space_2_lr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lr_addr : out  std_logic_vector(5 downto 0);
      memory_space_2_lr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_lc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_lc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_lc_data : in   std_logic_vector(31 downto 0);
      memory_space_2_lc_tag :  in  std_logic_vector(2 downto 0);
      AFB_NIC_REQUEST_pipe_read_req : out  std_logic_vector(0 downto 0);
      AFB_NIC_REQUEST_pipe_read_ack : in   std_logic_vector(0 downto 0);
      AFB_NIC_REQUEST_pipe_read_data : in   std_logic_vector(73 downto 0);
      MAC_ENABLE : in std_logic_vector(0 downto 0);
      AFB_NIC_RESPONSE_pipe_write_req : out  std_logic_vector(0 downto 0);
      AFB_NIC_RESPONSE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      AFB_NIC_RESPONSE_pipe_write_data : out  std_logic_vector(32 downto 0);
      CONTROL_REGISTER_pipe_write_req : out  std_logic_vector(0 downto 0);
      CONTROL_REGISTER_pipe_write_ack : in   std_logic_vector(0 downto 0);
      CONTROL_REGISTER_pipe_write_data : out  std_logic_vector(31 downto 0);
      FREE_Q_pipe_write_req : out  std_logic_vector(0 downto 0);
      FREE_Q_pipe_write_ack : in   std_logic_vector(0 downto 0);
      FREE_Q_pipe_write_data : out  std_logic_vector(35 downto 0);
      NUMBER_OF_SERVERS_pipe_write_req : out  std_logic_vector(0 downto 0);
      NUMBER_OF_SERVERS_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NUMBER_OF_SERVERS_pipe_write_data : out  std_logic_vector(31 downto 0);
      enable_mac_pipe_write_req : out  std_logic_vector(0 downto 0);
      enable_mac_pipe_write_ack : in   std_logic_vector(0 downto 0);
      enable_mac_pipe_write_data : out  std_logic_vector(0 downto 0);
      UpdateRegister_call_reqs : out  std_logic_vector(0 downto 0);
      UpdateRegister_call_acks : in   std_logic_vector(0 downto 0);
      UpdateRegister_call_data : out  std_logic_vector(73 downto 0);
      UpdateRegister_call_tag  :  out  std_logic_vector(0 downto 0);
      UpdateRegister_return_reqs : out  std_logic_vector(0 downto 0);
      UpdateRegister_return_acks : in   std_logic_vector(0 downto 0);
      UpdateRegister_return_data : in   std_logic_vector(31 downto 0);
      UpdateRegister_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module SoftwareRegisterAccessDaemon
  signal SoftwareRegisterAccessDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal SoftwareRegisterAccessDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal SoftwareRegisterAccessDaemon_start_req : std_logic;
  signal SoftwareRegisterAccessDaemon_start_ack : std_logic;
  signal SoftwareRegisterAccessDaemon_fin_req   : std_logic;
  signal SoftwareRegisterAccessDaemon_fin_ack : std_logic;
  -- declarations related to module UpdateRegister
  component UpdateRegister is -- 
    generic (tag_length : integer); 
    port ( -- 
      bmask : in  std_logic_vector(3 downto 0);
      rval : in  std_logic_vector(31 downto 0);
      wdata : in  std_logic_vector(31 downto 0);
      index : in  std_logic_vector(5 downto 0);
      wval : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sr_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sr_addr : out  std_logic_vector(5 downto 0);
      memory_space_2_sr_data : out  std_logic_vector(31 downto 0);
      memory_space_2_sr_tag :  out  std_logic_vector(20 downto 0);
      memory_space_2_sc_req : out  std_logic_vector(0 downto 0);
      memory_space_2_sc_ack : in   std_logic_vector(0 downto 0);
      memory_space_2_sc_tag :  in  std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module UpdateRegister
  signal UpdateRegister_bmask :  std_logic_vector(3 downto 0);
  signal UpdateRegister_rval :  std_logic_vector(31 downto 0);
  signal UpdateRegister_wdata :  std_logic_vector(31 downto 0);
  signal UpdateRegister_index :  std_logic_vector(5 downto 0);
  signal UpdateRegister_wval :  std_logic_vector(31 downto 0);
  signal UpdateRegister_in_args    : std_logic_vector(73 downto 0);
  signal UpdateRegister_out_args   : std_logic_vector(31 downto 0);
  signal UpdateRegister_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal UpdateRegister_tag_out   : std_logic_vector(2 downto 0);
  signal UpdateRegister_start_req : std_logic;
  signal UpdateRegister_start_ack : std_logic;
  signal UpdateRegister_fin_req   : std_logic;
  signal UpdateRegister_fin_ack : std_logic;
  -- caller side aggregated signals for module UpdateRegister
  signal UpdateRegister_call_reqs: std_logic_vector(1 downto 0);
  signal UpdateRegister_call_acks: std_logic_vector(1 downto 0);
  signal UpdateRegister_return_reqs: std_logic_vector(1 downto 0);
  signal UpdateRegister_return_acks: std_logic_vector(1 downto 0);
  signal UpdateRegister_call_data: std_logic_vector(147 downto 0);
  signal UpdateRegister_call_tag: std_logic_vector(1 downto 0);
  signal UpdateRegister_return_data: std_logic_vector(63 downto 0);
  signal UpdateRegister_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module accessMemory
  component accessMemory is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      bmask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEMORY_TO_NIC_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NIC_TO_MEMORY_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module accessMemory
  signal accessMemory_lock :  std_logic_vector(0 downto 0);
  signal accessMemory_rwbar :  std_logic_vector(0 downto 0);
  signal accessMemory_bmask :  std_logic_vector(7 downto 0);
  signal accessMemory_addr :  std_logic_vector(35 downto 0);
  signal accessMemory_wdata :  std_logic_vector(63 downto 0);
  signal accessMemory_rdata :  std_logic_vector(63 downto 0);
  signal accessMemory_in_args    : std_logic_vector(109 downto 0);
  signal accessMemory_out_args   : std_logic_vector(63 downto 0);
  signal accessMemory_tag_in    : std_logic_vector(7 downto 0) := (others => '0');
  signal accessMemory_tag_out   : std_logic_vector(7 downto 0);
  signal accessMemory_start_req : std_logic;
  signal accessMemory_start_ack : std_logic;
  signal accessMemory_fin_req   : std_logic;
  signal accessMemory_fin_ack : std_logic;
  -- caller side aggregated signals for module accessMemory
  signal accessMemory_call_reqs: std_logic_vector(15 downto 0);
  signal accessMemory_call_acks: std_logic_vector(15 downto 0);
  signal accessMemory_return_reqs: std_logic_vector(15 downto 0);
  signal accessMemory_return_acks: std_logic_vector(15 downto 0);
  signal accessMemory_call_data: std_logic_vector(1759 downto 0);
  signal accessMemory_call_tag: std_logic_vector(47 downto 0);
  signal accessMemory_return_data: std_logic_vector(1023 downto 0);
  signal accessMemory_return_tag: std_logic_vector(47 downto 0);
  -- declarations related to module acquireLock
  component acquireLock is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      m_ok : out  std_logic_vector(0 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module acquireLock
  signal acquireLock_q_base_address :  std_logic_vector(35 downto 0);
  signal acquireLock_m_ok :  std_logic_vector(0 downto 0);
  signal acquireLock_in_args    : std_logic_vector(35 downto 0);
  signal acquireLock_out_args   : std_logic_vector(0 downto 0);
  signal acquireLock_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal acquireLock_tag_out   : std_logic_vector(2 downto 0);
  signal acquireLock_start_req : std_logic;
  signal acquireLock_start_ack : std_logic;
  signal acquireLock_fin_req   : std_logic;
  signal acquireLock_fin_ack : std_logic;
  -- caller side aggregated signals for module acquireLock
  signal acquireLock_call_reqs: std_logic_vector(1 downto 0);
  signal acquireLock_call_acks: std_logic_vector(1 downto 0);
  signal acquireLock_return_reqs: std_logic_vector(1 downto 0);
  signal acquireLock_return_acks: std_logic_vector(1 downto 0);
  signal acquireLock_call_data: std_logic_vector(71 downto 0);
  signal acquireLock_call_tag: std_logic_vector(1 downto 0);
  signal acquireLock_return_data: std_logic_vector(1 downto 0);
  signal acquireLock_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module delay_time
  -- declarations related to module getQueueElement
  component getQueueElement is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      read_index : in  std_logic_vector(31 downto 0);
      q_r_data : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module getQueueElement
  signal getQueueElement_q_base_address :  std_logic_vector(35 downto 0);
  signal getQueueElement_read_index :  std_logic_vector(31 downto 0);
  signal getQueueElement_q_r_data :  std_logic_vector(31 downto 0);
  signal getQueueElement_in_args    : std_logic_vector(67 downto 0);
  signal getQueueElement_out_args   : std_logic_vector(31 downto 0);
  signal getQueueElement_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal getQueueElement_tag_out   : std_logic_vector(1 downto 0);
  signal getQueueElement_start_req : std_logic;
  signal getQueueElement_start_ack : std_logic;
  signal getQueueElement_fin_req   : std_logic;
  signal getQueueElement_fin_ack : std_logic;
  -- caller side aggregated signals for module getQueueElement
  signal getQueueElement_call_reqs: std_logic_vector(0 downto 0);
  signal getQueueElement_call_acks: std_logic_vector(0 downto 0);
  signal getQueueElement_return_reqs: std_logic_vector(0 downto 0);
  signal getQueueElement_return_acks: std_logic_vector(0 downto 0);
  signal getQueueElement_call_data: std_logic_vector(67 downto 0);
  signal getQueueElement_call_tag: std_logic_vector(0 downto 0);
  signal getQueueElement_return_data: std_logic_vector(31 downto 0);
  signal getQueueElement_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module getQueueLength
  component getQueueLength is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      Queue_Length : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module getQueueLength
  signal getQueueLength_q_base_address :  std_logic_vector(35 downto 0);
  signal getQueueLength_Queue_Length :  std_logic_vector(31 downto 0);
  signal getQueueLength_in_args    : std_logic_vector(35 downto 0);
  signal getQueueLength_out_args   : std_logic_vector(31 downto 0);
  signal getQueueLength_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal getQueueLength_tag_out   : std_logic_vector(2 downto 0);
  signal getQueueLength_start_req : std_logic;
  signal getQueueLength_start_ack : std_logic;
  signal getQueueLength_fin_req   : std_logic;
  signal getQueueLength_fin_ack : std_logic;
  -- caller side aggregated signals for module getQueueLength
  signal getQueueLength_call_reqs: std_logic_vector(1 downto 0);
  signal getQueueLength_call_acks: std_logic_vector(1 downto 0);
  signal getQueueLength_return_reqs: std_logic_vector(1 downto 0);
  signal getQueueLength_return_acks: std_logic_vector(1 downto 0);
  signal getQueueLength_call_data: std_logic_vector(71 downto 0);
  signal getQueueLength_call_tag: std_logic_vector(1 downto 0);
  signal getQueueLength_return_data: std_logic_vector(63 downto 0);
  signal getQueueLength_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module getQueuePointers
  component getQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : out  std_logic_vector(31 downto 0);
      rp : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module getQueuePointers
  signal getQueuePointers_q_base_address :  std_logic_vector(35 downto 0);
  signal getQueuePointers_wp :  std_logic_vector(31 downto 0);
  signal getQueuePointers_rp :  std_logic_vector(31 downto 0);
  signal getQueuePointers_in_args    : std_logic_vector(35 downto 0);
  signal getQueuePointers_out_args   : std_logic_vector(63 downto 0);
  signal getQueuePointers_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal getQueuePointers_tag_out   : std_logic_vector(2 downto 0);
  signal getQueuePointers_start_req : std_logic;
  signal getQueuePointers_start_ack : std_logic;
  signal getQueuePointers_fin_req   : std_logic;
  signal getQueuePointers_fin_ack : std_logic;
  -- caller side aggregated signals for module getQueuePointers
  signal getQueuePointers_call_reqs: std_logic_vector(1 downto 0);
  signal getQueuePointers_call_acks: std_logic_vector(1 downto 0);
  signal getQueuePointers_return_reqs: std_logic_vector(1 downto 0);
  signal getQueuePointers_return_acks: std_logic_vector(1 downto 0);
  signal getQueuePointers_call_data: std_logic_vector(71 downto 0);
  signal getQueuePointers_call_tag: std_logic_vector(1 downto 0);
  signal getQueuePointers_return_data: std_logic_vector(127 downto 0);
  signal getQueuePointers_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module getTotalMessages
  component getTotalMessages is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      total_msgs : out  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module getTotalMessages
  signal getTotalMessages_q_base_address :  std_logic_vector(35 downto 0);
  signal getTotalMessages_total_msgs :  std_logic_vector(31 downto 0);
  signal getTotalMessages_in_args    : std_logic_vector(35 downto 0);
  signal getTotalMessages_out_args   : std_logic_vector(31 downto 0);
  signal getTotalMessages_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal getTotalMessages_tag_out   : std_logic_vector(2 downto 0);
  signal getTotalMessages_start_req : std_logic;
  signal getTotalMessages_start_ack : std_logic;
  signal getTotalMessages_fin_req   : std_logic;
  signal getTotalMessages_fin_ack : std_logic;
  -- caller side aggregated signals for module getTotalMessages
  signal getTotalMessages_call_reqs: std_logic_vector(1 downto 0);
  signal getTotalMessages_call_acks: std_logic_vector(1 downto 0);
  signal getTotalMessages_return_reqs: std_logic_vector(1 downto 0);
  signal getTotalMessages_return_acks: std_logic_vector(1 downto 0);
  signal getTotalMessages_call_data: std_logic_vector(71 downto 0);
  signal getTotalMessages_call_tag: std_logic_vector(1 downto 0);
  signal getTotalMessages_return_data: std_logic_vector(63 downto 0);
  signal getTotalMessages_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module getTxPacketPointerFromServer
  component getTxPacketPointerFromServer is -- 
    generic (tag_length : integer); 
    port ( -- 
      queue_index : in  std_logic_vector(5 downto 0);
      pkt_pointer : out  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      popFromQueue_call_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_call_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_call_data : out  std_logic_vector(36 downto 0);
      popFromQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      popFromQueue_return_reqs : out  std_logic_vector(0 downto 0);
      popFromQueue_return_acks : in   std_logic_vector(0 downto 0);
      popFromQueue_return_data : in   std_logic_vector(32 downto 0);
      popFromQueue_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module getTxPacketPointerFromServer
  signal getTxPacketPointerFromServer_queue_index :  std_logic_vector(5 downto 0);
  signal getTxPacketPointerFromServer_pkt_pointer :  std_logic_vector(31 downto 0);
  signal getTxPacketPointerFromServer_status :  std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_in_args    : std_logic_vector(5 downto 0);
  signal getTxPacketPointerFromServer_out_args   : std_logic_vector(32 downto 0);
  signal getTxPacketPointerFromServer_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal getTxPacketPointerFromServer_tag_out   : std_logic_vector(1 downto 0);
  signal getTxPacketPointerFromServer_start_req : std_logic;
  signal getTxPacketPointerFromServer_start_ack : std_logic;
  signal getTxPacketPointerFromServer_fin_req   : std_logic;
  signal getTxPacketPointerFromServer_fin_ack : std_logic;
  -- caller side aggregated signals for module getTxPacketPointerFromServer
  signal getTxPacketPointerFromServer_call_reqs: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_call_acks: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_return_reqs: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_return_acks: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_call_data: std_logic_vector(5 downto 0);
  signal getTxPacketPointerFromServer_call_tag: std_logic_vector(0 downto 0);
  signal getTxPacketPointerFromServer_return_data: std_logic_vector(32 downto 0);
  signal getTxPacketPointerFromServer_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module loadBuffer
  component loadBuffer is -- 
    generic (tag_length : integer); 
    port ( -- 
      rx_buffer_pointer : in  std_logic_vector(35 downto 0);
      bad_packet_identifier : out  std_logic_vector(0 downto 0);
      writePayloadToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writePayloadToMem_call_acks : in   std_logic_vector(0 downto 0);
      writePayloadToMem_call_data : out  std_logic_vector(71 downto 0);
      writePayloadToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writePayloadToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writePayloadToMem_return_acks : in   std_logic_vector(0 downto 0);
      writePayloadToMem_return_data : in   std_logic_vector(19 downto 0);
      writePayloadToMem_return_tag :  in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_acks : in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_call_data : out  std_logic_vector(35 downto 0);
      writeEthernetHeaderToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_acks : in   std_logic_vector(0 downto 0);
      writeEthernetHeaderToMem_return_data : in   std_logic_vector(35 downto 0);
      writeEthernetHeaderToMem_return_tag :  in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_reqs : out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_acks : in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_call_data : out  std_logic_vector(54 downto 0);
      writeControlInformationToMem_call_tag  :  out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_reqs : out  std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_acks : in   std_logic_vector(0 downto 0);
      writeControlInformationToMem_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module loadBuffer
  signal loadBuffer_rx_buffer_pointer :  std_logic_vector(35 downto 0);
  signal loadBuffer_bad_packet_identifier :  std_logic_vector(0 downto 0);
  signal loadBuffer_in_args    : std_logic_vector(35 downto 0);
  signal loadBuffer_out_args   : std_logic_vector(0 downto 0);
  signal loadBuffer_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal loadBuffer_tag_out   : std_logic_vector(1 downto 0);
  signal loadBuffer_start_req : std_logic;
  signal loadBuffer_start_ack : std_logic;
  signal loadBuffer_fin_req   : std_logic;
  signal loadBuffer_fin_ack : std_logic;
  -- caller side aggregated signals for module loadBuffer
  signal loadBuffer_call_reqs: std_logic_vector(0 downto 0);
  signal loadBuffer_call_acks: std_logic_vector(0 downto 0);
  signal loadBuffer_return_reqs: std_logic_vector(0 downto 0);
  signal loadBuffer_return_acks: std_logic_vector(0 downto 0);
  signal loadBuffer_call_data: std_logic_vector(35 downto 0);
  signal loadBuffer_call_tag: std_logic_vector(0 downto 0);
  signal loadBuffer_return_data: std_logic_vector(0 downto 0);
  signal loadBuffer_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module nextLSTATE
  -- declarations related to module nicRxFromMacDaemon
  component nicRxFromMacDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      mac_to_nic_data_pipe_read_req : out  std_logic_vector(0 downto 0);
      mac_to_nic_data_pipe_read_ack : in   std_logic_vector(0 downto 0);
      mac_to_nic_data_pipe_read_data : in   std_logic_vector(72 downto 0);
      CONTROL_REGISTER : in std_logic_vector(31 downto 0);
      nic_rx_to_header_pipe_write_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_write_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_write_data : out  std_logic_vector(72 downto 0);
      nic_rx_to_packet_pipe_write_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_write_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_write_data : out  std_logic_vector(72 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(1 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(1 downto 0);
      AccessRegister_call_data : out  std_logic_vector(85 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(3 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(1 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(1 downto 0);
      AccessRegister_return_data : in   std_logic_vector(63 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(3 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module nicRxFromMacDaemon
  signal nicRxFromMacDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal nicRxFromMacDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal nicRxFromMacDaemon_start_req : std_logic;
  signal nicRxFromMacDaemon_start_ack : std_logic;
  signal nicRxFromMacDaemon_fin_req   : std_logic;
  signal nicRxFromMacDaemon_fin_ack : std_logic;
  -- declarations related to module popFromQueue
  component popFromQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_r_data : out  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_call_acks : in   std_logic_vector(0 downto 0);
      releaseLock_call_data : out  std_logic_vector(35 downto 0);
      releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_return_acks : in   std_logic_vector(0 downto 0);
      releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_call_acks : in   std_logic_vector(0 downto 0);
      acquireLock_call_data : out  std_logic_vector(35 downto 0);
      acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_return_acks : in   std_logic_vector(0 downto 0);
      acquireLock_return_data : in   std_logic_vector(0 downto 0);
      acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      updateTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_data : out  std_logic_vector(67 downto 0);
      updateTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_call_data : out  std_logic_vector(67 downto 0);
      getQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      getQueueElement_return_data : in   std_logic_vector(31 downto 0);
      getQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_call_data : out  std_logic_vector(35 downto 0);
      getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
      getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_call_data : out  std_logic_vector(35 downto 0);
      getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_return_data : in   std_logic_vector(31 downto 0);
      getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module popFromQueue
  signal popFromQueue_lock :  std_logic_vector(0 downto 0);
  signal popFromQueue_q_base_address :  std_logic_vector(35 downto 0);
  signal popFromQueue_q_r_data :  std_logic_vector(31 downto 0);
  signal popFromQueue_status :  std_logic_vector(0 downto 0);
  signal popFromQueue_in_args    : std_logic_vector(36 downto 0);
  signal popFromQueue_out_args   : std_logic_vector(32 downto 0);
  signal popFromQueue_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal popFromQueue_tag_out   : std_logic_vector(2 downto 0);
  signal popFromQueue_start_req : std_logic;
  signal popFromQueue_start_ack : std_logic;
  signal popFromQueue_fin_req   : std_logic;
  signal popFromQueue_fin_ack : std_logic;
  -- caller side aggregated signals for module popFromQueue
  signal popFromQueue_call_reqs: std_logic_vector(1 downto 0);
  signal popFromQueue_call_acks: std_logic_vector(1 downto 0);
  signal popFromQueue_return_reqs: std_logic_vector(1 downto 0);
  signal popFromQueue_return_acks: std_logic_vector(1 downto 0);
  signal popFromQueue_call_data: std_logic_vector(73 downto 0);
  signal popFromQueue_call_tag: std_logic_vector(1 downto 0);
  signal popFromQueue_return_data: std_logic_vector(65 downto 0);
  signal popFromQueue_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module populateRxQueue
  component populateRxQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      rx_buffer_pointer : in  std_logic_vector(35 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX : in std_logic_vector(5 downto 0);
      NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(0 downto 0);
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(5 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
      pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module populateRxQueue
  signal populateRxQueue_rx_buffer_pointer :  std_logic_vector(35 downto 0);
  signal populateRxQueue_in_args    : std_logic_vector(35 downto 0);
  signal populateRxQueue_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal populateRxQueue_tag_out   : std_logic_vector(1 downto 0);
  signal populateRxQueue_start_req : std_logic;
  signal populateRxQueue_start_ack : std_logic;
  signal populateRxQueue_fin_req   : std_logic;
  signal populateRxQueue_fin_ack : std_logic;
  -- caller side aggregated signals for module populateRxQueue
  signal populateRxQueue_call_reqs: std_logic_vector(0 downto 0);
  signal populateRxQueue_call_acks: std_logic_vector(0 downto 0);
  signal populateRxQueue_return_reqs: std_logic_vector(0 downto 0);
  signal populateRxQueue_return_acks: std_logic_vector(0 downto 0);
  signal populateRxQueue_call_data: std_logic_vector(35 downto 0);
  signal populateRxQueue_call_tag: std_logic_vector(0 downto 0);
  signal populateRxQueue_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module pushIntoQueue
  component pushIntoQueue is -- 
    generic (tag_length : integer); 
    port ( -- 
      lock : in  std_logic_vector(0 downto 0);
      q_base_address : in  std_logic_vector(35 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      releaseLock_call_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_call_acks : in   std_logic_vector(0 downto 0);
      releaseLock_call_data : out  std_logic_vector(35 downto 0);
      releaseLock_call_tag  :  out  std_logic_vector(0 downto 0);
      releaseLock_return_reqs : out  std_logic_vector(0 downto 0);
      releaseLock_return_acks : in   std_logic_vector(0 downto 0);
      releaseLock_return_tag :  in   std_logic_vector(0 downto 0);
      setQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_call_data : out  std_logic_vector(99 downto 0);
      setQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      setQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      setQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      acquireLock_call_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_call_acks : in   std_logic_vector(0 downto 0);
      acquireLock_call_data : out  std_logic_vector(35 downto 0);
      acquireLock_call_tag  :  out  std_logic_vector(0 downto 0);
      acquireLock_return_reqs : out  std_logic_vector(0 downto 0);
      acquireLock_return_acks : in   std_logic_vector(0 downto 0);
      acquireLock_return_data : in   std_logic_vector(0 downto 0);
      acquireLock_return_tag :  in   std_logic_vector(0 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      updateTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_call_data : out  std_logic_vector(67 downto 0);
      updateTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      updateTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      updateTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      getTotalMessages_call_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_call_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_call_data : out  std_logic_vector(35 downto 0);
      getTotalMessages_call_tag  :  out  std_logic_vector(0 downto 0);
      getTotalMessages_return_reqs : out  std_logic_vector(0 downto 0);
      getTotalMessages_return_acks : in   std_logic_vector(0 downto 0);
      getTotalMessages_return_data : in   std_logic_vector(31 downto 0);
      getTotalMessages_return_tag :  in   std_logic_vector(0 downto 0);
      getQueueLength_call_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_call_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_call_data : out  std_logic_vector(35 downto 0);
      getQueueLength_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueueLength_return_reqs : out  std_logic_vector(0 downto 0);
      getQueueLength_return_acks : in   std_logic_vector(0 downto 0);
      getQueueLength_return_data : in   std_logic_vector(31 downto 0);
      getQueueLength_return_tag :  in   std_logic_vector(0 downto 0);
      getQueuePointers_call_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_call_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_call_data : out  std_logic_vector(35 downto 0);
      getQueuePointers_call_tag  :  out  std_logic_vector(0 downto 0);
      getQueuePointers_return_reqs : out  std_logic_vector(0 downto 0);
      getQueuePointers_return_acks : in   std_logic_vector(0 downto 0);
      getQueuePointers_return_data : in   std_logic_vector(63 downto 0);
      getQueuePointers_return_tag :  in   std_logic_vector(0 downto 0);
      setQueueElement_call_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_call_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_call_data : out  std_logic_vector(99 downto 0);
      setQueueElement_call_tag  :  out  std_logic_vector(0 downto 0);
      setQueueElement_return_reqs : out  std_logic_vector(0 downto 0);
      setQueueElement_return_acks : in   std_logic_vector(0 downto 0);
      setQueueElement_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module pushIntoQueue
  signal pushIntoQueue_lock :  std_logic_vector(0 downto 0);
  signal pushIntoQueue_q_base_address :  std_logic_vector(35 downto 0);
  signal pushIntoQueue_q_w_data :  std_logic_vector(31 downto 0);
  signal pushIntoQueue_status :  std_logic_vector(0 downto 0);
  signal pushIntoQueue_in_args    : std_logic_vector(68 downto 0);
  signal pushIntoQueue_out_args   : std_logic_vector(0 downto 0);
  signal pushIntoQueue_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal pushIntoQueue_tag_out   : std_logic_vector(2 downto 0);
  signal pushIntoQueue_start_req : std_logic;
  signal pushIntoQueue_start_ack : std_logic;
  signal pushIntoQueue_fin_req   : std_logic;
  signal pushIntoQueue_fin_ack : std_logic;
  -- caller side aggregated signals for module pushIntoQueue
  signal pushIntoQueue_call_reqs: std_logic_vector(2 downto 0);
  signal pushIntoQueue_call_acks: std_logic_vector(2 downto 0);
  signal pushIntoQueue_return_reqs: std_logic_vector(2 downto 0);
  signal pushIntoQueue_return_acks: std_logic_vector(2 downto 0);
  signal pushIntoQueue_call_data: std_logic_vector(206 downto 0);
  signal pushIntoQueue_call_tag: std_logic_vector(2 downto 0);
  signal pushIntoQueue_return_data: std_logic_vector(2 downto 0);
  signal pushIntoQueue_return_tag: std_logic_vector(2 downto 0);
  -- declarations related to module releaseLock
  component releaseLock is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module releaseLock
  signal releaseLock_q_base_address :  std_logic_vector(35 downto 0);
  signal releaseLock_in_args    : std_logic_vector(35 downto 0);
  signal releaseLock_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal releaseLock_tag_out   : std_logic_vector(2 downto 0);
  signal releaseLock_start_req : std_logic;
  signal releaseLock_start_ack : std_logic;
  signal releaseLock_fin_req   : std_logic;
  signal releaseLock_fin_ack : std_logic;
  -- caller side aggregated signals for module releaseLock
  signal releaseLock_call_reqs: std_logic_vector(1 downto 0);
  signal releaseLock_call_acks: std_logic_vector(1 downto 0);
  signal releaseLock_return_reqs: std_logic_vector(1 downto 0);
  signal releaseLock_return_acks: std_logic_vector(1 downto 0);
  signal releaseLock_call_data: std_logic_vector(71 downto 0);
  signal releaseLock_call_tag: std_logic_vector(1 downto 0);
  signal releaseLock_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module setQueueElement
  component setQueueElement is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      write_index : in  std_logic_vector(31 downto 0);
      q_w_data : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module setQueueElement
  signal setQueueElement_q_base_address :  std_logic_vector(35 downto 0);
  signal setQueueElement_write_index :  std_logic_vector(31 downto 0);
  signal setQueueElement_q_w_data :  std_logic_vector(31 downto 0);
  signal setQueueElement_in_args    : std_logic_vector(99 downto 0);
  signal setQueueElement_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal setQueueElement_tag_out   : std_logic_vector(1 downto 0);
  signal setQueueElement_start_req : std_logic;
  signal setQueueElement_start_ack : std_logic;
  signal setQueueElement_fin_req   : std_logic;
  signal setQueueElement_fin_ack : std_logic;
  -- caller side aggregated signals for module setQueueElement
  signal setQueueElement_call_reqs: std_logic_vector(0 downto 0);
  signal setQueueElement_call_acks: std_logic_vector(0 downto 0);
  signal setQueueElement_return_reqs: std_logic_vector(0 downto 0);
  signal setQueueElement_return_acks: std_logic_vector(0 downto 0);
  signal setQueueElement_call_data: std_logic_vector(99 downto 0);
  signal setQueueElement_call_tag: std_logic_vector(0 downto 0);
  signal setQueueElement_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module setQueuePointers
  component setQueuePointers is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      wp : in  std_logic_vector(31 downto 0);
      rp : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module setQueuePointers
  signal setQueuePointers_q_base_address :  std_logic_vector(35 downto 0);
  signal setQueuePointers_wp :  std_logic_vector(31 downto 0);
  signal setQueuePointers_rp :  std_logic_vector(31 downto 0);
  signal setQueuePointers_in_args    : std_logic_vector(99 downto 0);
  signal setQueuePointers_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal setQueuePointers_tag_out   : std_logic_vector(2 downto 0);
  signal setQueuePointers_start_req : std_logic;
  signal setQueuePointers_start_ack : std_logic;
  signal setQueuePointers_fin_req   : std_logic;
  signal setQueuePointers_fin_ack : std_logic;
  -- caller side aggregated signals for module setQueuePointers
  signal setQueuePointers_call_reqs: std_logic_vector(1 downto 0);
  signal setQueuePointers_call_acks: std_logic_vector(1 downto 0);
  signal setQueuePointers_return_reqs: std_logic_vector(1 downto 0);
  signal setQueuePointers_return_acks: std_logic_vector(1 downto 0);
  signal setQueuePointers_call_data: std_logic_vector(199 downto 0);
  signal setQueuePointers_call_tag: std_logic_vector(1 downto 0);
  signal setQueuePointers_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module transmitEngineDaemon
  component transmitEngineDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      CONTROL_REGISTER : in std_logic_vector(31 downto 0);
      FREE_Q : in std_logic_vector(35 downto 0);
      LAST_READ_TX_QUEUE_INDEX : in std_logic_vector(5 downto 0);
      NUMBER_OF_SERVERS : in std_logic_vector(31 downto 0);
      LAST_READ_TX_QUEUE_INDEX_pipe_write_req : out  std_logic_vector(1 downto 0);
      LAST_READ_TX_QUEUE_INDEX_pipe_write_ack : in   std_logic_vector(1 downto 0);
      LAST_READ_TX_QUEUE_INDEX_pipe_write_data : out  std_logic_vector(11 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      pushIntoQueue_call_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_call_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_call_data : out  std_logic_vector(68 downto 0);
      pushIntoQueue_call_tag  :  out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_reqs : out  std_logic_vector(0 downto 0);
      pushIntoQueue_return_acks : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_data : in   std_logic_vector(0 downto 0);
      pushIntoQueue_return_tag :  in   std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_call_reqs : out  std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_call_acks : in   std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_call_data : out  std_logic_vector(5 downto 0);
      getTxPacketPointerFromServer_call_tag  :  out  std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_return_reqs : out  std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_return_acks : in   std_logic_vector(0 downto 0);
      getTxPacketPointerFromServer_return_data : in   std_logic_vector(32 downto 0);
      getTxPacketPointerFromServer_return_tag :  in   std_logic_vector(0 downto 0);
      transmitPacket_call_reqs : out  std_logic_vector(0 downto 0);
      transmitPacket_call_acks : in   std_logic_vector(0 downto 0);
      transmitPacket_call_data : out  std_logic_vector(31 downto 0);
      transmitPacket_call_tag  :  out  std_logic_vector(0 downto 0);
      transmitPacket_return_reqs : out  std_logic_vector(0 downto 0);
      transmitPacket_return_acks : in   std_logic_vector(0 downto 0);
      transmitPacket_return_data : in   std_logic_vector(0 downto 0);
      transmitPacket_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module transmitEngineDaemon
  signal transmitEngineDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal transmitEngineDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal transmitEngineDaemon_start_req : std_logic;
  signal transmitEngineDaemon_start_ack : std_logic;
  signal transmitEngineDaemon_fin_req   : std_logic;
  signal transmitEngineDaemon_fin_ack : std_logic;
  -- declarations related to module transmitPacket
  component transmitPacket is -- 
    generic (tag_length : integer); 
    port ( -- 
      packet_pointer : in  std_logic_vector(31 downto 0);
      status : out  std_logic_vector(0 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_req : out  std_logic_vector(1 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_ack : in   std_logic_vector(1 downto 0);
      nic_to_mac_transmit_pipe_pipe_write_data : out  std_logic_vector(145 downto 0);
      AccessRegister_call_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_call_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_call_data : out  std_logic_vector(42 downto 0);
      AccessRegister_call_tag  :  out  std_logic_vector(1 downto 0);
      AccessRegister_return_reqs : out  std_logic_vector(0 downto 0);
      AccessRegister_return_acks : in   std_logic_vector(0 downto 0);
      AccessRegister_return_data : in   std_logic_vector(31 downto 0);
      AccessRegister_return_tag :  in   std_logic_vector(1 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(1 downto 0);
      accessMemory_call_acks : in   std_logic_vector(1 downto 0);
      accessMemory_call_data : out  std_logic_vector(219 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(5 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(1 downto 0);
      accessMemory_return_acks : in   std_logic_vector(1 downto 0);
      accessMemory_return_data : in   std_logic_vector(127 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(5 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module transmitPacket
  signal transmitPacket_packet_pointer :  std_logic_vector(31 downto 0);
  signal transmitPacket_status :  std_logic_vector(0 downto 0);
  signal transmitPacket_in_args    : std_logic_vector(31 downto 0);
  signal transmitPacket_out_args   : std_logic_vector(0 downto 0);
  signal transmitPacket_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal transmitPacket_tag_out   : std_logic_vector(1 downto 0);
  signal transmitPacket_start_req : std_logic;
  signal transmitPacket_start_ack : std_logic;
  signal transmitPacket_fin_req   : std_logic;
  signal transmitPacket_fin_ack : std_logic;
  -- caller side aggregated signals for module transmitPacket
  signal transmitPacket_call_reqs: std_logic_vector(0 downto 0);
  signal transmitPacket_call_acks: std_logic_vector(0 downto 0);
  signal transmitPacket_return_reqs: std_logic_vector(0 downto 0);
  signal transmitPacket_return_acks: std_logic_vector(0 downto 0);
  signal transmitPacket_call_data: std_logic_vector(31 downto 0);
  signal transmitPacket_call_tag: std_logic_vector(0 downto 0);
  signal transmitPacket_return_data: std_logic_vector(0 downto 0);
  signal transmitPacket_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module updateTotalMessages
  component updateTotalMessages is -- 
    generic (tag_length : integer); 
    port ( -- 
      q_base_address : in  std_logic_vector(35 downto 0);
      updated_total_msgs : in  std_logic_vector(31 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module updateTotalMessages
  signal updateTotalMessages_q_base_address :  std_logic_vector(35 downto 0);
  signal updateTotalMessages_updated_total_msgs :  std_logic_vector(31 downto 0);
  signal updateTotalMessages_in_args    : std_logic_vector(67 downto 0);
  signal updateTotalMessages_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal updateTotalMessages_tag_out   : std_logic_vector(2 downto 0);
  signal updateTotalMessages_start_req : std_logic;
  signal updateTotalMessages_start_ack : std_logic;
  signal updateTotalMessages_fin_req   : std_logic;
  signal updateTotalMessages_fin_ack : std_logic;
  -- caller side aggregated signals for module updateTotalMessages
  signal updateTotalMessages_call_reqs: std_logic_vector(1 downto 0);
  signal updateTotalMessages_call_acks: std_logic_vector(1 downto 0);
  signal updateTotalMessages_return_reqs: std_logic_vector(1 downto 0);
  signal updateTotalMessages_return_acks: std_logic_vector(1 downto 0);
  signal updateTotalMessages_call_data: std_logic_vector(135 downto 0);
  signal updateTotalMessages_call_tag: std_logic_vector(1 downto 0);
  signal updateTotalMessages_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module writeControlInformationToMem
  component writeControlInformationToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      base_buffer_pointer : in  std_logic_vector(35 downto 0);
      packet_size : in  std_logic_vector(10 downto 0);
      last_keep : in  std_logic_vector(7 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module writeControlInformationToMem
  signal writeControlInformationToMem_base_buffer_pointer :  std_logic_vector(35 downto 0);
  signal writeControlInformationToMem_packet_size :  std_logic_vector(10 downto 0);
  signal writeControlInformationToMem_last_keep :  std_logic_vector(7 downto 0);
  signal writeControlInformationToMem_in_args    : std_logic_vector(54 downto 0);
  signal writeControlInformationToMem_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal writeControlInformationToMem_tag_out   : std_logic_vector(1 downto 0);
  signal writeControlInformationToMem_start_req : std_logic;
  signal writeControlInformationToMem_start_ack : std_logic;
  signal writeControlInformationToMem_fin_req   : std_logic;
  signal writeControlInformationToMem_fin_ack : std_logic;
  -- caller side aggregated signals for module writeControlInformationToMem
  signal writeControlInformationToMem_call_reqs: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_call_acks: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_return_reqs: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_return_acks: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_call_data: std_logic_vector(54 downto 0);
  signal writeControlInformationToMem_call_tag: std_logic_vector(0 downto 0);
  signal writeControlInformationToMem_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module writeEthernetHeaderToMem
  component writeEthernetHeaderToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      buf_pointer : in  std_logic_vector(35 downto 0);
      buf_position_out : out  std_logic_vector(35 downto 0);
      nic_rx_to_header_pipe_read_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_read_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_header_pipe_read_data : in   std_logic_vector(72 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module writeEthernetHeaderToMem
  signal writeEthernetHeaderToMem_buf_pointer :  std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_buf_position_out :  std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_in_args    : std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_out_args   : std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal writeEthernetHeaderToMem_tag_out   : std_logic_vector(1 downto 0);
  signal writeEthernetHeaderToMem_start_req : std_logic;
  signal writeEthernetHeaderToMem_start_ack : std_logic;
  signal writeEthernetHeaderToMem_fin_req   : std_logic;
  signal writeEthernetHeaderToMem_fin_ack : std_logic;
  -- caller side aggregated signals for module writeEthernetHeaderToMem
  signal writeEthernetHeaderToMem_call_reqs: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_call_acks: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_return_reqs: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_return_acks: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_call_data: std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_call_tag: std_logic_vector(0 downto 0);
  signal writeEthernetHeaderToMem_return_data: std_logic_vector(35 downto 0);
  signal writeEthernetHeaderToMem_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module writePayloadToMem
  component writePayloadToMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      base_buf_pointer : in  std_logic_vector(35 downto 0);
      buf_pointer : in  std_logic_vector(35 downto 0);
      packet_size_32 : out  std_logic_vector(10 downto 0);
      bad_packet_identifier : out  std_logic_vector(0 downto 0);
      last_keep : out  std_logic_vector(7 downto 0);
      nic_rx_to_packet_pipe_read_req : out  std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_read_ack : in   std_logic_vector(0 downto 0);
      nic_rx_to_packet_pipe_read_data : in   std_logic_vector(72 downto 0);
      accessMemory_call_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_call_acks : in   std_logic_vector(0 downto 0);
      accessMemory_call_data : out  std_logic_vector(109 downto 0);
      accessMemory_call_tag  :  out  std_logic_vector(2 downto 0);
      accessMemory_return_reqs : out  std_logic_vector(0 downto 0);
      accessMemory_return_acks : in   std_logic_vector(0 downto 0);
      accessMemory_return_data : in   std_logic_vector(63 downto 0);
      accessMemory_return_tag :  in   std_logic_vector(2 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module writePayloadToMem
  signal writePayloadToMem_base_buf_pointer :  std_logic_vector(35 downto 0);
  signal writePayloadToMem_buf_pointer :  std_logic_vector(35 downto 0);
  signal writePayloadToMem_packet_size_32 :  std_logic_vector(10 downto 0);
  signal writePayloadToMem_bad_packet_identifier :  std_logic_vector(0 downto 0);
  signal writePayloadToMem_last_keep :  std_logic_vector(7 downto 0);
  signal writePayloadToMem_in_args    : std_logic_vector(71 downto 0);
  signal writePayloadToMem_out_args   : std_logic_vector(19 downto 0);
  signal writePayloadToMem_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal writePayloadToMem_tag_out   : std_logic_vector(1 downto 0);
  signal writePayloadToMem_start_req : std_logic;
  signal writePayloadToMem_start_ack : std_logic;
  signal writePayloadToMem_fin_req   : std_logic;
  signal writePayloadToMem_fin_ack : std_logic;
  -- caller side aggregated signals for module writePayloadToMem
  signal writePayloadToMem_call_reqs: std_logic_vector(0 downto 0);
  signal writePayloadToMem_call_acks: std_logic_vector(0 downto 0);
  signal writePayloadToMem_return_reqs: std_logic_vector(0 downto 0);
  signal writePayloadToMem_return_acks: std_logic_vector(0 downto 0);
  signal writePayloadToMem_call_data: std_logic_vector(71 downto 0);
  signal writePayloadToMem_call_tag: std_logic_vector(0 downto 0);
  signal writePayloadToMem_return_data: std_logic_vector(19 downto 0);
  signal writePayloadToMem_return_tag: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe AFB_NIC_REQUEST
  signal AFB_NIC_REQUEST_pipe_read_data: std_logic_vector(73 downto 0);
  signal AFB_NIC_REQUEST_pipe_read_req: std_logic_vector(0 downto 0);
  signal AFB_NIC_REQUEST_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe AFB_NIC_RESPONSE
  signal AFB_NIC_RESPONSE_pipe_write_data: std_logic_vector(32 downto 0);
  signal AFB_NIC_RESPONSE_pipe_write_req: std_logic_vector(0 downto 0);
  signal AFB_NIC_RESPONSE_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe CONTROL_REGISTER
  signal CONTROL_REGISTER_pipe_write_data: std_logic_vector(31 downto 0);
  signal CONTROL_REGISTER_pipe_write_req: std_logic_vector(0 downto 0);
  signal CONTROL_REGISTER_pipe_write_ack: std_logic_vector(0 downto 0);
  -- signal decl. for read from internal signal pipe CONTROL_REGISTER
  signal CONTROL_REGISTER: std_logic_vector(31 downto 0);
  -- aggregate signals for write to pipe FREE_Q
  signal FREE_Q_pipe_write_data: std_logic_vector(35 downto 0);
  signal FREE_Q_pipe_write_req: std_logic_vector(0 downto 0);
  signal FREE_Q_pipe_write_ack: std_logic_vector(0 downto 0);
  -- signal decl. for read from internal signal pipe FREE_Q
  signal FREE_Q: std_logic_vector(35 downto 0);
  -- aggregate signals for write to pipe LAST_READ_TX_QUEUE_INDEX
  signal LAST_READ_TX_QUEUE_INDEX_pipe_write_data: std_logic_vector(11 downto 0);
  signal LAST_READ_TX_QUEUE_INDEX_pipe_write_req: std_logic_vector(1 downto 0);
  signal LAST_READ_TX_QUEUE_INDEX_pipe_write_ack: std_logic_vector(1 downto 0);
  -- signal decl. for read from internal signal pipe LAST_READ_TX_QUEUE_INDEX
  signal LAST_READ_TX_QUEUE_INDEX: std_logic_vector(5 downto 0);
  -- aggregate signals for write to pipe LAST_WRITTEN_RX_QUEUE_INDEX
  signal LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data: std_logic_vector(11 downto 0);
  signal LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req: std_logic_vector(1 downto 0);
  signal LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack: std_logic_vector(1 downto 0);
  -- signal decl. for read from internal signal pipe LAST_WRITTEN_RX_QUEUE_INDEX
  signal LAST_WRITTEN_RX_QUEUE_INDEX: std_logic_vector(5 downto 0);
  -- aggregate signals for write to pipe MAC_ENABLE
  signal MAC_ENABLE_pipe_write_data: std_logic_vector(0 downto 0);
  signal MAC_ENABLE_pipe_write_req: std_logic_vector(0 downto 0);
  signal MAC_ENABLE_pipe_write_ack: std_logic_vector(0 downto 0);
  -- signal decl. for read from internal signal pipe MAC_ENABLE
  signal MAC_ENABLE: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe MEMORY_TO_NIC_RESPONSE
  signal MEMORY_TO_NIC_RESPONSE_pipe_read_data: std_logic_vector(64 downto 0);
  signal MEMORY_TO_NIC_RESPONSE_pipe_read_req: std_logic_vector(0 downto 0);
  signal MEMORY_TO_NIC_RESPONSE_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe NIC_REQUEST_REGISTER_ACCESS_PIPE
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data: std_logic_vector(42 downto 0);
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req: std_logic_vector(0 downto 0);
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe NIC_REQUEST_REGISTER_ACCESS_PIPE
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data: std_logic_vector(42 downto 0);
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req: std_logic_vector(0 downto 0);
  signal NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe NIC_RESPONSE_REGISTER_ACCESS_PIPE
  signal NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data: std_logic_vector(32 downto 0);
  signal NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req: std_logic_vector(0 downto 0);
  signal NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe NIC_RESPONSE_REGISTER_ACCESS_PIPE
  signal NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data: std_logic_vector(32 downto 0);
  signal NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req: std_logic_vector(0 downto 0);
  signal NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe NIC_TO_MEMORY_REQUEST
  signal NIC_TO_MEMORY_REQUEST_pipe_write_data: std_logic_vector(109 downto 0);
  signal NIC_TO_MEMORY_REQUEST_pipe_write_req: std_logic_vector(0 downto 0);
  signal NIC_TO_MEMORY_REQUEST_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe NUMBER_OF_SERVERS
  signal NUMBER_OF_SERVERS_pipe_write_data: std_logic_vector(31 downto 0);
  signal NUMBER_OF_SERVERS_pipe_write_req: std_logic_vector(0 downto 0);
  signal NUMBER_OF_SERVERS_pipe_write_ack: std_logic_vector(0 downto 0);
  -- signal decl. for read from internal signal pipe NUMBER_OF_SERVERS
  signal NUMBER_OF_SERVERS: std_logic_vector(31 downto 0);
  -- aggregate signals for write to pipe enable_mac
  signal enable_mac_pipe_write_data: std_logic_vector(0 downto 0);
  signal enable_mac_pipe_write_req: std_logic_vector(0 downto 0);
  signal enable_mac_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe mac_to_nic_data
  signal mac_to_nic_data_pipe_read_data: std_logic_vector(72 downto 0);
  signal mac_to_nic_data_pipe_read_req: std_logic_vector(0 downto 0);
  signal mac_to_nic_data_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe nic_rx_to_header
  signal nic_rx_to_header_pipe_write_data: std_logic_vector(72 downto 0);
  signal nic_rx_to_header_pipe_write_req: std_logic_vector(0 downto 0);
  signal nic_rx_to_header_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe nic_rx_to_header
  signal nic_rx_to_header_pipe_read_data: std_logic_vector(72 downto 0);
  signal nic_rx_to_header_pipe_read_req: std_logic_vector(0 downto 0);
  signal nic_rx_to_header_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe nic_rx_to_packet
  signal nic_rx_to_packet_pipe_write_data: std_logic_vector(72 downto 0);
  signal nic_rx_to_packet_pipe_write_req: std_logic_vector(0 downto 0);
  signal nic_rx_to_packet_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe nic_rx_to_packet
  signal nic_rx_to_packet_pipe_read_data: std_logic_vector(72 downto 0);
  signal nic_rx_to_packet_pipe_read_req: std_logic_vector(0 downto 0);
  signal nic_rx_to_packet_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe nic_to_mac_transmit_pipe
  signal nic_to_mac_transmit_pipe_pipe_write_data: std_logic_vector(145 downto 0);
  signal nic_to_mac_transmit_pipe_pipe_write_req: std_logic_vector(1 downto 0);
  signal nic_to_mac_transmit_pipe_pipe_write_ack: std_logic_vector(1 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module AccessRegister
  AccessRegister_rwbar <= AccessRegister_in_args(42 downto 42);
  AccessRegister_bmask <= AccessRegister_in_args(41 downto 38);
  AccessRegister_register_index <= AccessRegister_in_args(37 downto 32);
  AccessRegister_wdata <= AccessRegister_in_args(31 downto 0);
  AccessRegister_out_args <= AccessRegister_rdata ;
  -- call arbiter for module AccessRegister
  AccessRegister_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 7,
      call_data_width => 43,
      return_data_width => 32,
      callee_tag_length => 3,
      caller_tag_length => 2--
    )
    port map(-- 
      call_reqs => AccessRegister_call_reqs,
      call_acks => AccessRegister_call_acks,
      return_reqs => AccessRegister_return_reqs,
      return_acks => AccessRegister_return_acks,
      call_data  => AccessRegister_call_data,
      call_tag  => AccessRegister_call_tag,
      return_tag  => AccessRegister_return_tag,
      call_mtag => AccessRegister_tag_in,
      return_mtag => AccessRegister_tag_out,
      return_data =>AccessRegister_return_data,
      call_mreq => AccessRegister_start_req,
      call_mack => AccessRegister_start_ack,
      return_mreq => AccessRegister_fin_req,
      return_mack => AccessRegister_fin_ack,
      call_mdata => AccessRegister_in_args,
      return_mdata => AccessRegister_out_args,
      clk => clk, 
      reset => reset --
    ); --
  AccessRegister_instance:AccessRegister-- 
    generic map(tag_length => 5)
    port map(-- 
      rwbar => AccessRegister_rwbar,
      bmask => AccessRegister_bmask,
      register_index => AccessRegister_register_index,
      wdata => AccessRegister_wdata,
      rdata => AccessRegister_rdata,
      start_req => AccessRegister_start_req,
      start_ack => AccessRegister_start_ack,
      fin_req => AccessRegister_fin_req,
      fin_ack => AccessRegister_fin_ack,
      clk => clk,
      reset => reset,
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req(0 downto 0),
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack(0 downto 0),
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data(32 downto 0),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req(0 downto 0),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack(0 downto 0),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data(42 downto 0),
      tag_in => AccessRegister_tag_in,
      tag_out => AccessRegister_tag_out-- 
    ); -- 
  -- module NicRegisterAccessDaemon
  NicRegisterAccessDaemon_instance:NicRegisterAccessDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => NicRegisterAccessDaemon_start_req,
      start_ack => NicRegisterAccessDaemon_start_ack,
      fin_req => NicRegisterAccessDaemon_fin_req,
      fin_ack => NicRegisterAccessDaemon_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(1 downto 1),
      memory_space_2_lr_ack => memory_space_2_lr_ack(1 downto 1),
      memory_space_2_lr_addr => memory_space_2_lr_addr(11 downto 6),
      memory_space_2_lr_tag => memory_space_2_lr_tag(41 downto 21),
      memory_space_2_lc_req => memory_space_2_lc_req(1 downto 1),
      memory_space_2_lc_ack => memory_space_2_lc_ack(1 downto 1),
      memory_space_2_lc_data => memory_space_2_lc_data(63 downto 32),
      memory_space_2_lc_tag => memory_space_2_lc_tag(5 downto 3),
      memory_space_2_sr_req => memory_space_2_sr_req(1 downto 1),
      memory_space_2_sr_ack => memory_space_2_sr_ack(1 downto 1),
      memory_space_2_sr_addr => memory_space_2_sr_addr(11 downto 6),
      memory_space_2_sr_data => memory_space_2_sr_data(63 downto 32),
      memory_space_2_sr_tag => memory_space_2_sr_tag(41 downto 21),
      memory_space_2_sc_req => memory_space_2_sc_req(1 downto 1),
      memory_space_2_sc_ack => memory_space_2_sc_ack(1 downto 1),
      memory_space_2_sc_tag => memory_space_2_sc_tag(5 downto 3),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req(0 downto 0),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack(0 downto 0),
      NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data(42 downto 0),
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req(0 downto 0),
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack(0 downto 0),
      NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data(32 downto 0),
      MAC_ENABLE_pipe_write_req => MAC_ENABLE_pipe_write_req(0 downto 0),
      MAC_ENABLE_pipe_write_ack => MAC_ENABLE_pipe_write_ack(0 downto 0),
      MAC_ENABLE_pipe_write_data => MAC_ENABLE_pipe_write_data(0 downto 0),
      UpdateRegister_call_reqs => UpdateRegister_call_reqs(1 downto 1),
      UpdateRegister_call_acks => UpdateRegister_call_acks(1 downto 1),
      UpdateRegister_call_data => UpdateRegister_call_data(147 downto 74),
      UpdateRegister_call_tag => UpdateRegister_call_tag(1 downto 1),
      UpdateRegister_return_reqs => UpdateRegister_return_reqs(1 downto 1),
      UpdateRegister_return_acks => UpdateRegister_return_acks(1 downto 1),
      UpdateRegister_return_data => UpdateRegister_return_data(63 downto 32),
      UpdateRegister_return_tag => UpdateRegister_return_tag(1 downto 1),
      tag_in => NicRegisterAccessDaemon_tag_in,
      tag_out => NicRegisterAccessDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  NicRegisterAccessDaemon_tag_in <= (others => '0');
  NicRegisterAccessDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => NicRegisterAccessDaemon_start_req, start_ack => NicRegisterAccessDaemon_start_ack,  fin_req => NicRegisterAccessDaemon_fin_req,  fin_ack => NicRegisterAccessDaemon_fin_ack);
  -- module ReceiveEngineDaemon
  ReceiveEngineDaemon_instance:ReceiveEngineDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => ReceiveEngineDaemon_start_req,
      start_ack => ReceiveEngineDaemon_start_ack,
      fin_req => ReceiveEngineDaemon_fin_req,
      fin_ack => ReceiveEngineDaemon_fin_ack,
      clk => clk,
      reset => reset,
      CONTROL_REGISTER => CONTROL_REGISTER,
      FREE_Q => FREE_Q,
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req(0 downto 0),
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack(0 downto 0),
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data(5 downto 0),
      AccessRegister_call_reqs => AccessRegister_call_reqs(5 downto 5),
      AccessRegister_call_acks => AccessRegister_call_acks(5 downto 5),
      AccessRegister_call_data => AccessRegister_call_data(257 downto 215),
      AccessRegister_call_tag => AccessRegister_call_tag(11 downto 10),
      AccessRegister_return_reqs => AccessRegister_return_reqs(5 downto 5),
      AccessRegister_return_acks => AccessRegister_return_acks(5 downto 5),
      AccessRegister_return_data => AccessRegister_return_data(191 downto 160),
      AccessRegister_return_tag => AccessRegister_return_tag(11 downto 10),
      popFromQueue_call_reqs => popFromQueue_call_reqs(1 downto 1),
      popFromQueue_call_acks => popFromQueue_call_acks(1 downto 1),
      popFromQueue_call_data => popFromQueue_call_data(73 downto 37),
      popFromQueue_call_tag => popFromQueue_call_tag(1 downto 1),
      popFromQueue_return_reqs => popFromQueue_return_reqs(1 downto 1),
      popFromQueue_return_acks => popFromQueue_return_acks(1 downto 1),
      popFromQueue_return_data => popFromQueue_return_data(65 downto 33),
      popFromQueue_return_tag => popFromQueue_return_tag(1 downto 1),
      loadBuffer_call_reqs => loadBuffer_call_reqs(0 downto 0),
      loadBuffer_call_acks => loadBuffer_call_acks(0 downto 0),
      loadBuffer_call_data => loadBuffer_call_data(35 downto 0),
      loadBuffer_call_tag => loadBuffer_call_tag(0 downto 0),
      loadBuffer_return_reqs => loadBuffer_return_reqs(0 downto 0),
      loadBuffer_return_acks => loadBuffer_return_acks(0 downto 0),
      loadBuffer_return_data => loadBuffer_return_data(0 downto 0),
      loadBuffer_return_tag => loadBuffer_return_tag(0 downto 0),
      pushIntoQueue_call_reqs => pushIntoQueue_call_reqs(1 downto 1),
      pushIntoQueue_call_acks => pushIntoQueue_call_acks(1 downto 1),
      pushIntoQueue_call_data => pushIntoQueue_call_data(137 downto 69),
      pushIntoQueue_call_tag => pushIntoQueue_call_tag(1 downto 1),
      pushIntoQueue_return_reqs => pushIntoQueue_return_reqs(1 downto 1),
      pushIntoQueue_return_acks => pushIntoQueue_return_acks(1 downto 1),
      pushIntoQueue_return_data => pushIntoQueue_return_data(1 downto 1),
      pushIntoQueue_return_tag => pushIntoQueue_return_tag(1 downto 1),
      populateRxQueue_call_reqs => populateRxQueue_call_reqs(0 downto 0),
      populateRxQueue_call_acks => populateRxQueue_call_acks(0 downto 0),
      populateRxQueue_call_data => populateRxQueue_call_data(35 downto 0),
      populateRxQueue_call_tag => populateRxQueue_call_tag(0 downto 0),
      populateRxQueue_return_reqs => populateRxQueue_return_reqs(0 downto 0),
      populateRxQueue_return_acks => populateRxQueue_return_acks(0 downto 0),
      populateRxQueue_return_tag => populateRxQueue_return_tag(0 downto 0),
      tag_in => ReceiveEngineDaemon_tag_in,
      tag_out => ReceiveEngineDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  ReceiveEngineDaemon_tag_in <= (others => '0');
  ReceiveEngineDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => ReceiveEngineDaemon_start_req, start_ack => ReceiveEngineDaemon_start_ack,  fin_req => ReceiveEngineDaemon_fin_req,  fin_ack => ReceiveEngineDaemon_fin_ack);
  -- module SoftwareRegisterAccessDaemon
  SoftwareRegisterAccessDaemon_instance:SoftwareRegisterAccessDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => SoftwareRegisterAccessDaemon_start_req,
      start_ack => SoftwareRegisterAccessDaemon_start_ack,
      fin_req => SoftwareRegisterAccessDaemon_fin_req,
      fin_ack => SoftwareRegisterAccessDaemon_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_lr_req => memory_space_2_lr_req(0 downto 0),
      memory_space_2_lr_ack => memory_space_2_lr_ack(0 downto 0),
      memory_space_2_lr_addr => memory_space_2_lr_addr(5 downto 0),
      memory_space_2_lr_tag => memory_space_2_lr_tag(20 downto 0),
      memory_space_2_lc_req => memory_space_2_lc_req(0 downto 0),
      memory_space_2_lc_ack => memory_space_2_lc_ack(0 downto 0),
      memory_space_2_lc_data => memory_space_2_lc_data(31 downto 0),
      memory_space_2_lc_tag => memory_space_2_lc_tag(2 downto 0),
      AFB_NIC_REQUEST_pipe_read_req => AFB_NIC_REQUEST_pipe_read_req(0 downto 0),
      AFB_NIC_REQUEST_pipe_read_ack => AFB_NIC_REQUEST_pipe_read_ack(0 downto 0),
      AFB_NIC_REQUEST_pipe_read_data => AFB_NIC_REQUEST_pipe_read_data(73 downto 0),
      MAC_ENABLE => MAC_ENABLE,
      AFB_NIC_RESPONSE_pipe_write_req => AFB_NIC_RESPONSE_pipe_write_req(0 downto 0),
      AFB_NIC_RESPONSE_pipe_write_ack => AFB_NIC_RESPONSE_pipe_write_ack(0 downto 0),
      AFB_NIC_RESPONSE_pipe_write_data => AFB_NIC_RESPONSE_pipe_write_data(32 downto 0),
      CONTROL_REGISTER_pipe_write_req => CONTROL_REGISTER_pipe_write_req(0 downto 0),
      CONTROL_REGISTER_pipe_write_ack => CONTROL_REGISTER_pipe_write_ack(0 downto 0),
      CONTROL_REGISTER_pipe_write_data => CONTROL_REGISTER_pipe_write_data(31 downto 0),
      FREE_Q_pipe_write_req => FREE_Q_pipe_write_req(0 downto 0),
      FREE_Q_pipe_write_ack => FREE_Q_pipe_write_ack(0 downto 0),
      FREE_Q_pipe_write_data => FREE_Q_pipe_write_data(35 downto 0),
      NUMBER_OF_SERVERS_pipe_write_req => NUMBER_OF_SERVERS_pipe_write_req(0 downto 0),
      NUMBER_OF_SERVERS_pipe_write_ack => NUMBER_OF_SERVERS_pipe_write_ack(0 downto 0),
      NUMBER_OF_SERVERS_pipe_write_data => NUMBER_OF_SERVERS_pipe_write_data(31 downto 0),
      enable_mac_pipe_write_req => enable_mac_pipe_write_req(0 downto 0),
      enable_mac_pipe_write_ack => enable_mac_pipe_write_ack(0 downto 0),
      enable_mac_pipe_write_data => enable_mac_pipe_write_data(0 downto 0),
      UpdateRegister_call_reqs => UpdateRegister_call_reqs(0 downto 0),
      UpdateRegister_call_acks => UpdateRegister_call_acks(0 downto 0),
      UpdateRegister_call_data => UpdateRegister_call_data(73 downto 0),
      UpdateRegister_call_tag => UpdateRegister_call_tag(0 downto 0),
      UpdateRegister_return_reqs => UpdateRegister_return_reqs(0 downto 0),
      UpdateRegister_return_acks => UpdateRegister_return_acks(0 downto 0),
      UpdateRegister_return_data => UpdateRegister_return_data(31 downto 0),
      UpdateRegister_return_tag => UpdateRegister_return_tag(0 downto 0),
      tag_in => SoftwareRegisterAccessDaemon_tag_in,
      tag_out => SoftwareRegisterAccessDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  SoftwareRegisterAccessDaemon_tag_in <= (others => '0');
  SoftwareRegisterAccessDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => SoftwareRegisterAccessDaemon_start_req, start_ack => SoftwareRegisterAccessDaemon_start_ack,  fin_req => SoftwareRegisterAccessDaemon_fin_req,  fin_ack => SoftwareRegisterAccessDaemon_fin_ack);
  -- module UpdateRegister
  UpdateRegister_bmask <= UpdateRegister_in_args(73 downto 70);
  UpdateRegister_rval <= UpdateRegister_in_args(69 downto 38);
  UpdateRegister_wdata <= UpdateRegister_in_args(37 downto 6);
  UpdateRegister_index <= UpdateRegister_in_args(5 downto 0);
  UpdateRegister_out_args <= UpdateRegister_wval ;
  -- call arbiter for module UpdateRegister
  UpdateRegister_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 74,
      return_data_width => 32,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => UpdateRegister_call_reqs,
      call_acks => UpdateRegister_call_acks,
      return_reqs => UpdateRegister_return_reqs,
      return_acks => UpdateRegister_return_acks,
      call_data  => UpdateRegister_call_data,
      call_tag  => UpdateRegister_call_tag,
      return_tag  => UpdateRegister_return_tag,
      call_mtag => UpdateRegister_tag_in,
      return_mtag => UpdateRegister_tag_out,
      return_data =>UpdateRegister_return_data,
      call_mreq => UpdateRegister_start_req,
      call_mack => UpdateRegister_start_ack,
      return_mreq => UpdateRegister_fin_req,
      return_mack => UpdateRegister_fin_ack,
      call_mdata => UpdateRegister_in_args,
      return_mdata => UpdateRegister_out_args,
      clk => clk, 
      reset => reset --
    ); --
  UpdateRegister_instance:UpdateRegister-- 
    generic map(tag_length => 3)
    port map(-- 
      bmask => UpdateRegister_bmask,
      rval => UpdateRegister_rval,
      wdata => UpdateRegister_wdata,
      index => UpdateRegister_index,
      wval => UpdateRegister_wval,
      start_req => UpdateRegister_start_req,
      start_ack => UpdateRegister_start_ack,
      fin_req => UpdateRegister_fin_req,
      fin_ack => UpdateRegister_fin_ack,
      clk => clk,
      reset => reset,
      memory_space_2_sr_req => memory_space_2_sr_req(0 downto 0),
      memory_space_2_sr_ack => memory_space_2_sr_ack(0 downto 0),
      memory_space_2_sr_addr => memory_space_2_sr_addr(5 downto 0),
      memory_space_2_sr_data => memory_space_2_sr_data(31 downto 0),
      memory_space_2_sr_tag => memory_space_2_sr_tag(20 downto 0),
      memory_space_2_sc_req => memory_space_2_sc_req(0 downto 0),
      memory_space_2_sc_ack => memory_space_2_sc_ack(0 downto 0),
      memory_space_2_sc_tag => memory_space_2_sc_tag(2 downto 0),
      tag_in => UpdateRegister_tag_in,
      tag_out => UpdateRegister_tag_out-- 
    ); -- 
  -- module accessMemory
  accessMemory_lock <= accessMemory_in_args(109 downto 109);
  accessMemory_rwbar <= accessMemory_in_args(108 downto 108);
  accessMemory_bmask <= accessMemory_in_args(107 downto 100);
  accessMemory_addr <= accessMemory_in_args(99 downto 64);
  accessMemory_wdata <= accessMemory_in_args(63 downto 0);
  accessMemory_out_args <= accessMemory_rdata ;
  -- call arbiter for module accessMemory
  accessMemory_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 16,
      call_data_width => 110,
      return_data_width => 64,
      callee_tag_length => 5,
      caller_tag_length => 3--
    )
    port map(-- 
      call_reqs => accessMemory_call_reqs,
      call_acks => accessMemory_call_acks,
      return_reqs => accessMemory_return_reqs,
      return_acks => accessMemory_return_acks,
      call_data  => accessMemory_call_data,
      call_tag  => accessMemory_call_tag,
      return_tag  => accessMemory_return_tag,
      call_mtag => accessMemory_tag_in,
      return_mtag => accessMemory_tag_out,
      return_data =>accessMemory_return_data,
      call_mreq => accessMemory_start_req,
      call_mack => accessMemory_start_ack,
      return_mreq => accessMemory_fin_req,
      return_mack => accessMemory_fin_ack,
      call_mdata => accessMemory_in_args,
      return_mdata => accessMemory_out_args,
      clk => clk, 
      reset => reset --
    ); --
  accessMemory_instance:accessMemory-- 
    generic map(tag_length => 8)
    port map(-- 
      lock => accessMemory_lock,
      rwbar => accessMemory_rwbar,
      bmask => accessMemory_bmask,
      addr => accessMemory_addr,
      wdata => accessMemory_wdata,
      rdata => accessMemory_rdata,
      start_req => accessMemory_start_req,
      start_ack => accessMemory_start_ack,
      fin_req => accessMemory_fin_req,
      fin_ack => accessMemory_fin_ack,
      clk => clk,
      reset => reset,
      MEMORY_TO_NIC_RESPONSE_pipe_read_req => MEMORY_TO_NIC_RESPONSE_pipe_read_req(0 downto 0),
      MEMORY_TO_NIC_RESPONSE_pipe_read_ack => MEMORY_TO_NIC_RESPONSE_pipe_read_ack(0 downto 0),
      MEMORY_TO_NIC_RESPONSE_pipe_read_data => MEMORY_TO_NIC_RESPONSE_pipe_read_data(64 downto 0),
      NIC_TO_MEMORY_REQUEST_pipe_write_req => NIC_TO_MEMORY_REQUEST_pipe_write_req(0 downto 0),
      NIC_TO_MEMORY_REQUEST_pipe_write_ack => NIC_TO_MEMORY_REQUEST_pipe_write_ack(0 downto 0),
      NIC_TO_MEMORY_REQUEST_pipe_write_data => NIC_TO_MEMORY_REQUEST_pipe_write_data(109 downto 0),
      tag_in => accessMemory_tag_in,
      tag_out => accessMemory_tag_out-- 
    ); -- 
  -- module acquireLock
  acquireLock_q_base_address <= acquireLock_in_args(35 downto 0);
  acquireLock_out_args <= acquireLock_m_ok ;
  -- call arbiter for module acquireLock
  acquireLock_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 36,
      return_data_width => 1,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => acquireLock_call_reqs,
      call_acks => acquireLock_call_acks,
      return_reqs => acquireLock_return_reqs,
      return_acks => acquireLock_return_acks,
      call_data  => acquireLock_call_data,
      call_tag  => acquireLock_call_tag,
      return_tag  => acquireLock_return_tag,
      call_mtag => acquireLock_tag_in,
      return_mtag => acquireLock_tag_out,
      return_data =>acquireLock_return_data,
      call_mreq => acquireLock_start_req,
      call_mack => acquireLock_start_ack,
      return_mreq => acquireLock_fin_req,
      return_mack => acquireLock_fin_ack,
      call_mdata => acquireLock_in_args,
      return_mdata => acquireLock_out_args,
      clk => clk, 
      reset => reset --
    ); --
  acquireLock_instance:acquireLock-- 
    generic map(tag_length => 3)
    port map(-- 
      q_base_address => acquireLock_q_base_address,
      m_ok => acquireLock_m_ok,
      start_req => acquireLock_start_req,
      start_ack => acquireLock_start_ack,
      fin_req => acquireLock_fin_req,
      fin_ack => acquireLock_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(13 downto 13),
      accessMemory_call_acks => accessMemory_call_acks(13 downto 13),
      accessMemory_call_data => accessMemory_call_data(1539 downto 1430),
      accessMemory_call_tag => accessMemory_call_tag(41 downto 39),
      accessMemory_return_reqs => accessMemory_return_reqs(13 downto 13),
      accessMemory_return_acks => accessMemory_return_acks(13 downto 13),
      accessMemory_return_data => accessMemory_return_data(895 downto 832),
      accessMemory_return_tag => accessMemory_return_tag(41 downto 39),
      tag_in => acquireLock_tag_in,
      tag_out => acquireLock_tag_out-- 
    ); -- 
  -- module getQueueElement
  getQueueElement_q_base_address <= getQueueElement_in_args(67 downto 32);
  getQueueElement_read_index <= getQueueElement_in_args(31 downto 0);
  getQueueElement_out_args <= getQueueElement_q_r_data ;
  -- call arbiter for module getQueueElement
  getQueueElement_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 68,
      return_data_width => 32,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => getQueueElement_call_reqs,
      call_acks => getQueueElement_call_acks,
      return_reqs => getQueueElement_return_reqs,
      return_acks => getQueueElement_return_acks,
      call_data  => getQueueElement_call_data,
      call_tag  => getQueueElement_call_tag,
      return_tag  => getQueueElement_return_tag,
      call_mtag => getQueueElement_tag_in,
      return_mtag => getQueueElement_tag_out,
      return_data =>getQueueElement_return_data,
      call_mreq => getQueueElement_start_req,
      call_mack => getQueueElement_start_ack,
      return_mreq => getQueueElement_fin_req,
      return_mack => getQueueElement_fin_ack,
      call_mdata => getQueueElement_in_args,
      return_mdata => getQueueElement_out_args,
      clk => clk, 
      reset => reset --
    ); --
  getQueueElement_instance:getQueueElement-- 
    generic map(tag_length => 2)
    port map(-- 
      q_base_address => getQueueElement_q_base_address,
      read_index => getQueueElement_read_index,
      q_r_data => getQueueElement_q_r_data,
      start_req => getQueueElement_start_req,
      start_ack => getQueueElement_start_ack,
      fin_req => getQueueElement_fin_req,
      fin_ack => getQueueElement_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(11 downto 11),
      accessMemory_call_acks => accessMemory_call_acks(11 downto 11),
      accessMemory_call_data => accessMemory_call_data(1319 downto 1210),
      accessMemory_call_tag => accessMemory_call_tag(35 downto 33),
      accessMemory_return_reqs => accessMemory_return_reqs(11 downto 11),
      accessMemory_return_acks => accessMemory_return_acks(11 downto 11),
      accessMemory_return_data => accessMemory_return_data(767 downto 704),
      accessMemory_return_tag => accessMemory_return_tag(35 downto 33),
      tag_in => getQueueElement_tag_in,
      tag_out => getQueueElement_tag_out-- 
    ); -- 
  -- module getQueueLength
  getQueueLength_q_base_address <= getQueueLength_in_args(35 downto 0);
  getQueueLength_out_args <= getQueueLength_Queue_Length ;
  -- call arbiter for module getQueueLength
  getQueueLength_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 36,
      return_data_width => 32,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => getQueueLength_call_reqs,
      call_acks => getQueueLength_call_acks,
      return_reqs => getQueueLength_return_reqs,
      return_acks => getQueueLength_return_acks,
      call_data  => getQueueLength_call_data,
      call_tag  => getQueueLength_call_tag,
      return_tag  => getQueueLength_return_tag,
      call_mtag => getQueueLength_tag_in,
      return_mtag => getQueueLength_tag_out,
      return_data =>getQueueLength_return_data,
      call_mreq => getQueueLength_start_req,
      call_mack => getQueueLength_start_ack,
      return_mreq => getQueueLength_fin_req,
      return_mack => getQueueLength_fin_ack,
      call_mdata => getQueueLength_in_args,
      return_mdata => getQueueLength_out_args,
      clk => clk, 
      reset => reset --
    ); --
  getQueueLength_instance:getQueueLength-- 
    generic map(tag_length => 3)
    port map(-- 
      q_base_address => getQueueLength_q_base_address,
      Queue_Length => getQueueLength_Queue_Length,
      start_req => getQueueLength_start_req,
      start_ack => getQueueLength_start_ack,
      fin_req => getQueueLength_fin_req,
      fin_ack => getQueueLength_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(9 downto 9),
      accessMemory_call_acks => accessMemory_call_acks(9 downto 9),
      accessMemory_call_data => accessMemory_call_data(1099 downto 990),
      accessMemory_call_tag => accessMemory_call_tag(29 downto 27),
      accessMemory_return_reqs => accessMemory_return_reqs(9 downto 9),
      accessMemory_return_acks => accessMemory_return_acks(9 downto 9),
      accessMemory_return_data => accessMemory_return_data(639 downto 576),
      accessMemory_return_tag => accessMemory_return_tag(29 downto 27),
      tag_in => getQueueLength_tag_in,
      tag_out => getQueueLength_tag_out-- 
    ); -- 
  -- module getQueuePointers
  getQueuePointers_q_base_address <= getQueuePointers_in_args(35 downto 0);
  getQueuePointers_out_args <= getQueuePointers_wp & getQueuePointers_rp ;
  -- call arbiter for module getQueuePointers
  getQueuePointers_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 36,
      return_data_width => 64,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => getQueuePointers_call_reqs,
      call_acks => getQueuePointers_call_acks,
      return_reqs => getQueuePointers_return_reqs,
      return_acks => getQueuePointers_return_acks,
      call_data  => getQueuePointers_call_data,
      call_tag  => getQueuePointers_call_tag,
      return_tag  => getQueuePointers_return_tag,
      call_mtag => getQueuePointers_tag_in,
      return_mtag => getQueuePointers_tag_out,
      return_data =>getQueuePointers_return_data,
      call_mreq => getQueuePointers_start_req,
      call_mack => getQueuePointers_start_ack,
      return_mreq => getQueuePointers_fin_req,
      return_mack => getQueuePointers_fin_ack,
      call_mdata => getQueuePointers_in_args,
      return_mdata => getQueuePointers_out_args,
      clk => clk, 
      reset => reset --
    ); --
  getQueuePointers_instance:getQueuePointers-- 
    generic map(tag_length => 3)
    port map(-- 
      q_base_address => getQueuePointers_q_base_address,
      wp => getQueuePointers_wp,
      rp => getQueuePointers_rp,
      start_req => getQueuePointers_start_req,
      start_ack => getQueuePointers_start_ack,
      fin_req => getQueuePointers_fin_req,
      fin_ack => getQueuePointers_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(8 downto 8),
      accessMemory_call_acks => accessMemory_call_acks(8 downto 8),
      accessMemory_call_data => accessMemory_call_data(989 downto 880),
      accessMemory_call_tag => accessMemory_call_tag(26 downto 24),
      accessMemory_return_reqs => accessMemory_return_reqs(8 downto 8),
      accessMemory_return_acks => accessMemory_return_acks(8 downto 8),
      accessMemory_return_data => accessMemory_return_data(575 downto 512),
      accessMemory_return_tag => accessMemory_return_tag(26 downto 24),
      tag_in => getQueuePointers_tag_in,
      tag_out => getQueuePointers_tag_out-- 
    ); -- 
  -- module getTotalMessages
  getTotalMessages_q_base_address <= getTotalMessages_in_args(35 downto 0);
  getTotalMessages_out_args <= getTotalMessages_total_msgs ;
  -- call arbiter for module getTotalMessages
  getTotalMessages_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 36,
      return_data_width => 32,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => getTotalMessages_call_reqs,
      call_acks => getTotalMessages_call_acks,
      return_reqs => getTotalMessages_return_reqs,
      return_acks => getTotalMessages_return_acks,
      call_data  => getTotalMessages_call_data,
      call_tag  => getTotalMessages_call_tag,
      return_tag  => getTotalMessages_return_tag,
      call_mtag => getTotalMessages_tag_in,
      return_mtag => getTotalMessages_tag_out,
      return_data =>getTotalMessages_return_data,
      call_mreq => getTotalMessages_start_req,
      call_mack => getTotalMessages_start_ack,
      return_mreq => getTotalMessages_fin_req,
      return_mack => getTotalMessages_fin_ack,
      call_mdata => getTotalMessages_in_args,
      return_mdata => getTotalMessages_out_args,
      clk => clk, 
      reset => reset --
    ); --
  getTotalMessages_instance:getTotalMessages-- 
    generic map(tag_length => 3)
    port map(-- 
      q_base_address => getTotalMessages_q_base_address,
      total_msgs => getTotalMessages_total_msgs,
      start_req => getTotalMessages_start_req,
      start_ack => getTotalMessages_start_ack,
      fin_req => getTotalMessages_fin_req,
      fin_ack => getTotalMessages_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(10 downto 10),
      accessMemory_call_acks => accessMemory_call_acks(10 downto 10),
      accessMemory_call_data => accessMemory_call_data(1209 downto 1100),
      accessMemory_call_tag => accessMemory_call_tag(32 downto 30),
      accessMemory_return_reqs => accessMemory_return_reqs(10 downto 10),
      accessMemory_return_acks => accessMemory_return_acks(10 downto 10),
      accessMemory_return_data => accessMemory_return_data(703 downto 640),
      accessMemory_return_tag => accessMemory_return_tag(32 downto 30),
      tag_in => getTotalMessages_tag_in,
      tag_out => getTotalMessages_tag_out-- 
    ); -- 
  -- module getTxPacketPointerFromServer
  getTxPacketPointerFromServer_queue_index <= getTxPacketPointerFromServer_in_args(5 downto 0);
  getTxPacketPointerFromServer_out_args <= getTxPacketPointerFromServer_pkt_pointer & getTxPacketPointerFromServer_status ;
  -- call arbiter for module getTxPacketPointerFromServer
  getTxPacketPointerFromServer_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 6,
      return_data_width => 33,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => getTxPacketPointerFromServer_call_reqs,
      call_acks => getTxPacketPointerFromServer_call_acks,
      return_reqs => getTxPacketPointerFromServer_return_reqs,
      return_acks => getTxPacketPointerFromServer_return_acks,
      call_data  => getTxPacketPointerFromServer_call_data,
      call_tag  => getTxPacketPointerFromServer_call_tag,
      return_tag  => getTxPacketPointerFromServer_return_tag,
      call_mtag => getTxPacketPointerFromServer_tag_in,
      return_mtag => getTxPacketPointerFromServer_tag_out,
      return_data =>getTxPacketPointerFromServer_return_data,
      call_mreq => getTxPacketPointerFromServer_start_req,
      call_mack => getTxPacketPointerFromServer_start_ack,
      return_mreq => getTxPacketPointerFromServer_fin_req,
      return_mack => getTxPacketPointerFromServer_fin_ack,
      call_mdata => getTxPacketPointerFromServer_in_args,
      return_mdata => getTxPacketPointerFromServer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  getTxPacketPointerFromServer_instance:getTxPacketPointerFromServer-- 
    generic map(tag_length => 2)
    port map(-- 
      queue_index => getTxPacketPointerFromServer_queue_index,
      pkt_pointer => getTxPacketPointerFromServer_pkt_pointer,
      status => getTxPacketPointerFromServer_status,
      start_req => getTxPacketPointerFromServer_start_req,
      start_ack => getTxPacketPointerFromServer_start_ack,
      fin_req => getTxPacketPointerFromServer_fin_req,
      fin_ack => getTxPacketPointerFromServer_fin_ack,
      clk => clk,
      reset => reset,
      AccessRegister_call_reqs => AccessRegister_call_reqs(4 downto 4),
      AccessRegister_call_acks => AccessRegister_call_acks(4 downto 4),
      AccessRegister_call_data => AccessRegister_call_data(214 downto 172),
      AccessRegister_call_tag => AccessRegister_call_tag(9 downto 8),
      AccessRegister_return_reqs => AccessRegister_return_reqs(4 downto 4),
      AccessRegister_return_acks => AccessRegister_return_acks(4 downto 4),
      AccessRegister_return_data => AccessRegister_return_data(159 downto 128),
      AccessRegister_return_tag => AccessRegister_return_tag(9 downto 8),
      popFromQueue_call_reqs => popFromQueue_call_reqs(0 downto 0),
      popFromQueue_call_acks => popFromQueue_call_acks(0 downto 0),
      popFromQueue_call_data => popFromQueue_call_data(36 downto 0),
      popFromQueue_call_tag => popFromQueue_call_tag(0 downto 0),
      popFromQueue_return_reqs => popFromQueue_return_reqs(0 downto 0),
      popFromQueue_return_acks => popFromQueue_return_acks(0 downto 0),
      popFromQueue_return_data => popFromQueue_return_data(32 downto 0),
      popFromQueue_return_tag => popFromQueue_return_tag(0 downto 0),
      tag_in => getTxPacketPointerFromServer_tag_in,
      tag_out => getTxPacketPointerFromServer_tag_out-- 
    ); -- 
  -- module loadBuffer
  loadBuffer_rx_buffer_pointer <= loadBuffer_in_args(35 downto 0);
  loadBuffer_out_args <= loadBuffer_bad_packet_identifier ;
  -- call arbiter for module loadBuffer
  loadBuffer_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 36,
      return_data_width => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => loadBuffer_call_reqs,
      call_acks => loadBuffer_call_acks,
      return_reqs => loadBuffer_return_reqs,
      return_acks => loadBuffer_return_acks,
      call_data  => loadBuffer_call_data,
      call_tag  => loadBuffer_call_tag,
      return_tag  => loadBuffer_return_tag,
      call_mtag => loadBuffer_tag_in,
      return_mtag => loadBuffer_tag_out,
      return_data =>loadBuffer_return_data,
      call_mreq => loadBuffer_start_req,
      call_mack => loadBuffer_start_ack,
      return_mreq => loadBuffer_fin_req,
      return_mack => loadBuffer_fin_ack,
      call_mdata => loadBuffer_in_args,
      return_mdata => loadBuffer_out_args,
      clk => clk, 
      reset => reset --
    ); --
  loadBuffer_instance:loadBuffer-- 
    generic map(tag_length => 2)
    port map(-- 
      rx_buffer_pointer => loadBuffer_rx_buffer_pointer,
      bad_packet_identifier => loadBuffer_bad_packet_identifier,
      start_req => loadBuffer_start_req,
      start_ack => loadBuffer_start_ack,
      fin_req => loadBuffer_fin_req,
      fin_ack => loadBuffer_fin_ack,
      clk => clk,
      reset => reset,
      writeEthernetHeaderToMem_call_reqs => writeEthernetHeaderToMem_call_reqs(0 downto 0),
      writeEthernetHeaderToMem_call_acks => writeEthernetHeaderToMem_call_acks(0 downto 0),
      writeEthernetHeaderToMem_call_data => writeEthernetHeaderToMem_call_data(35 downto 0),
      writeEthernetHeaderToMem_call_tag => writeEthernetHeaderToMem_call_tag(0 downto 0),
      writeEthernetHeaderToMem_return_reqs => writeEthernetHeaderToMem_return_reqs(0 downto 0),
      writeEthernetHeaderToMem_return_acks => writeEthernetHeaderToMem_return_acks(0 downto 0),
      writeEthernetHeaderToMem_return_data => writeEthernetHeaderToMem_return_data(35 downto 0),
      writeEthernetHeaderToMem_return_tag => writeEthernetHeaderToMem_return_tag(0 downto 0),
      writePayloadToMem_call_reqs => writePayloadToMem_call_reqs(0 downto 0),
      writePayloadToMem_call_acks => writePayloadToMem_call_acks(0 downto 0),
      writePayloadToMem_call_data => writePayloadToMem_call_data(71 downto 0),
      writePayloadToMem_call_tag => writePayloadToMem_call_tag(0 downto 0),
      writePayloadToMem_return_reqs => writePayloadToMem_return_reqs(0 downto 0),
      writePayloadToMem_return_acks => writePayloadToMem_return_acks(0 downto 0),
      writePayloadToMem_return_data => writePayloadToMem_return_data(19 downto 0),
      writePayloadToMem_return_tag => writePayloadToMem_return_tag(0 downto 0),
      writeControlInformationToMem_call_reqs => writeControlInformationToMem_call_reqs(0 downto 0),
      writeControlInformationToMem_call_acks => writeControlInformationToMem_call_acks(0 downto 0),
      writeControlInformationToMem_call_data => writeControlInformationToMem_call_data(54 downto 0),
      writeControlInformationToMem_call_tag => writeControlInformationToMem_call_tag(0 downto 0),
      writeControlInformationToMem_return_reqs => writeControlInformationToMem_return_reqs(0 downto 0),
      writeControlInformationToMem_return_acks => writeControlInformationToMem_return_acks(0 downto 0),
      writeControlInformationToMem_return_tag => writeControlInformationToMem_return_tag(0 downto 0),
      tag_in => loadBuffer_tag_in,
      tag_out => loadBuffer_tag_out-- 
    ); -- 
  -- module nicRxFromMacDaemon
  nicRxFromMacDaemon_instance:nicRxFromMacDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => nicRxFromMacDaemon_start_req,
      start_ack => nicRxFromMacDaemon_start_ack,
      fin_req => nicRxFromMacDaemon_fin_req,
      fin_ack => nicRxFromMacDaemon_fin_ack,
      clk => clk,
      reset => reset,
      CONTROL_REGISTER => CONTROL_REGISTER,
      mac_to_nic_data_pipe_read_req => mac_to_nic_data_pipe_read_req(0 downto 0),
      mac_to_nic_data_pipe_read_ack => mac_to_nic_data_pipe_read_ack(0 downto 0),
      mac_to_nic_data_pipe_read_data => mac_to_nic_data_pipe_read_data(72 downto 0),
      nic_rx_to_header_pipe_write_req => nic_rx_to_header_pipe_write_req(0 downto 0),
      nic_rx_to_header_pipe_write_ack => nic_rx_to_header_pipe_write_ack(0 downto 0),
      nic_rx_to_header_pipe_write_data => nic_rx_to_header_pipe_write_data(72 downto 0),
      nic_rx_to_packet_pipe_write_req => nic_rx_to_packet_pipe_write_req(0 downto 0),
      nic_rx_to_packet_pipe_write_ack => nic_rx_to_packet_pipe_write_ack(0 downto 0),
      nic_rx_to_packet_pipe_write_data => nic_rx_to_packet_pipe_write_data(72 downto 0),
      AccessRegister_call_reqs => AccessRegister_call_reqs(3 downto 2),
      AccessRegister_call_acks => AccessRegister_call_acks(3 downto 2),
      AccessRegister_call_data => AccessRegister_call_data(171 downto 86),
      AccessRegister_call_tag => AccessRegister_call_tag(7 downto 4),
      AccessRegister_return_reqs => AccessRegister_return_reqs(3 downto 2),
      AccessRegister_return_acks => AccessRegister_return_acks(3 downto 2),
      AccessRegister_return_data => AccessRegister_return_data(127 downto 64),
      AccessRegister_return_tag => AccessRegister_return_tag(7 downto 4),
      tag_in => nicRxFromMacDaemon_tag_in,
      tag_out => nicRxFromMacDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  nicRxFromMacDaemon_tag_in <= (others => '0');
  nicRxFromMacDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => nicRxFromMacDaemon_start_req, start_ack => nicRxFromMacDaemon_start_ack,  fin_req => nicRxFromMacDaemon_fin_req,  fin_ack => nicRxFromMacDaemon_fin_ack);
  -- module popFromQueue
  popFromQueue_lock <= popFromQueue_in_args(36 downto 36);
  popFromQueue_q_base_address <= popFromQueue_in_args(35 downto 0);
  popFromQueue_out_args <= popFromQueue_q_r_data & popFromQueue_status ;
  -- call arbiter for module popFromQueue
  popFromQueue_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 37,
      return_data_width => 33,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => popFromQueue_call_reqs,
      call_acks => popFromQueue_call_acks,
      return_reqs => popFromQueue_return_reqs,
      return_acks => popFromQueue_return_acks,
      call_data  => popFromQueue_call_data,
      call_tag  => popFromQueue_call_tag,
      return_tag  => popFromQueue_return_tag,
      call_mtag => popFromQueue_tag_in,
      return_mtag => popFromQueue_tag_out,
      return_data =>popFromQueue_return_data,
      call_mreq => popFromQueue_start_req,
      call_mack => popFromQueue_start_ack,
      return_mreq => popFromQueue_fin_req,
      return_mack => popFromQueue_fin_ack,
      call_mdata => popFromQueue_in_args,
      return_mdata => popFromQueue_out_args,
      clk => clk, 
      reset => reset --
    ); --
  popFromQueue_instance:popFromQueue-- 
    generic map(tag_length => 3)
    port map(-- 
      lock => popFromQueue_lock,
      q_base_address => popFromQueue_q_base_address,
      q_r_data => popFromQueue_q_r_data,
      status => popFromQueue_status,
      start_req => popFromQueue_start_req,
      start_ack => popFromQueue_start_ack,
      fin_req => popFromQueue_fin_req,
      fin_ack => popFromQueue_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(7 downto 7),
      accessMemory_call_acks => accessMemory_call_acks(7 downto 7),
      accessMemory_call_data => accessMemory_call_data(879 downto 770),
      accessMemory_call_tag => accessMemory_call_tag(23 downto 21),
      accessMemory_return_reqs => accessMemory_return_reqs(7 downto 7),
      accessMemory_return_acks => accessMemory_return_acks(7 downto 7),
      accessMemory_return_data => accessMemory_return_data(511 downto 448),
      accessMemory_return_tag => accessMemory_return_tag(23 downto 21),
      acquireLock_call_reqs => acquireLock_call_reqs(1 downto 1),
      acquireLock_call_acks => acquireLock_call_acks(1 downto 1),
      acquireLock_call_data => acquireLock_call_data(71 downto 36),
      acquireLock_call_tag => acquireLock_call_tag(1 downto 1),
      acquireLock_return_reqs => acquireLock_return_reqs(1 downto 1),
      acquireLock_return_acks => acquireLock_return_acks(1 downto 1),
      acquireLock_return_data => acquireLock_return_data(1 downto 1),
      acquireLock_return_tag => acquireLock_return_tag(1 downto 1),
      getQueuePointers_call_reqs => getQueuePointers_call_reqs(1 downto 1),
      getQueuePointers_call_acks => getQueuePointers_call_acks(1 downto 1),
      getQueuePointers_call_data => getQueuePointers_call_data(71 downto 36),
      getQueuePointers_call_tag => getQueuePointers_call_tag(1 downto 1),
      getQueuePointers_return_reqs => getQueuePointers_return_reqs(1 downto 1),
      getQueuePointers_return_acks => getQueuePointers_return_acks(1 downto 1),
      getQueuePointers_return_data => getQueuePointers_return_data(127 downto 64),
      getQueuePointers_return_tag => getQueuePointers_return_tag(1 downto 1),
      getQueueLength_call_reqs => getQueueLength_call_reqs(1 downto 1),
      getQueueLength_call_acks => getQueueLength_call_acks(1 downto 1),
      getQueueLength_call_data => getQueueLength_call_data(71 downto 36),
      getQueueLength_call_tag => getQueueLength_call_tag(1 downto 1),
      getQueueLength_return_reqs => getQueueLength_return_reqs(1 downto 1),
      getQueueLength_return_acks => getQueueLength_return_acks(1 downto 1),
      getQueueLength_return_data => getQueueLength_return_data(63 downto 32),
      getQueueLength_return_tag => getQueueLength_return_tag(1 downto 1),
      getTotalMessages_call_reqs => getTotalMessages_call_reqs(1 downto 1),
      getTotalMessages_call_acks => getTotalMessages_call_acks(1 downto 1),
      getTotalMessages_call_data => getTotalMessages_call_data(71 downto 36),
      getTotalMessages_call_tag => getTotalMessages_call_tag(1 downto 1),
      getTotalMessages_return_reqs => getTotalMessages_return_reqs(1 downto 1),
      getTotalMessages_return_acks => getTotalMessages_return_acks(1 downto 1),
      getTotalMessages_return_data => getTotalMessages_return_data(63 downto 32),
      getTotalMessages_return_tag => getTotalMessages_return_tag(1 downto 1),
      getQueueElement_call_reqs => getQueueElement_call_reqs(0 downto 0),
      getQueueElement_call_acks => getQueueElement_call_acks(0 downto 0),
      getQueueElement_call_data => getQueueElement_call_data(67 downto 0),
      getQueueElement_call_tag => getQueueElement_call_tag(0 downto 0),
      getQueueElement_return_reqs => getQueueElement_return_reqs(0 downto 0),
      getQueueElement_return_acks => getQueueElement_return_acks(0 downto 0),
      getQueueElement_return_data => getQueueElement_return_data(31 downto 0),
      getQueueElement_return_tag => getQueueElement_return_tag(0 downto 0),
      setQueuePointers_call_reqs => setQueuePointers_call_reqs(1 downto 1),
      setQueuePointers_call_acks => setQueuePointers_call_acks(1 downto 1),
      setQueuePointers_call_data => setQueuePointers_call_data(199 downto 100),
      setQueuePointers_call_tag => setQueuePointers_call_tag(1 downto 1),
      setQueuePointers_return_reqs => setQueuePointers_return_reqs(1 downto 1),
      setQueuePointers_return_acks => setQueuePointers_return_acks(1 downto 1),
      setQueuePointers_return_tag => setQueuePointers_return_tag(1 downto 1),
      updateTotalMessages_call_reqs => updateTotalMessages_call_reqs(1 downto 1),
      updateTotalMessages_call_acks => updateTotalMessages_call_acks(1 downto 1),
      updateTotalMessages_call_data => updateTotalMessages_call_data(135 downto 68),
      updateTotalMessages_call_tag => updateTotalMessages_call_tag(1 downto 1),
      updateTotalMessages_return_reqs => updateTotalMessages_return_reqs(1 downto 1),
      updateTotalMessages_return_acks => updateTotalMessages_return_acks(1 downto 1),
      updateTotalMessages_return_tag => updateTotalMessages_return_tag(1 downto 1),
      releaseLock_call_reqs => releaseLock_call_reqs(1 downto 1),
      releaseLock_call_acks => releaseLock_call_acks(1 downto 1),
      releaseLock_call_data => releaseLock_call_data(71 downto 36),
      releaseLock_call_tag => releaseLock_call_tag(1 downto 1),
      releaseLock_return_reqs => releaseLock_return_reqs(1 downto 1),
      releaseLock_return_acks => releaseLock_return_acks(1 downto 1),
      releaseLock_return_tag => releaseLock_return_tag(1 downto 1),
      tag_in => popFromQueue_tag_in,
      tag_out => popFromQueue_tag_out-- 
    ); -- 
  -- module populateRxQueue
  populateRxQueue_rx_buffer_pointer <= populateRxQueue_in_args(35 downto 0);
  -- call arbiter for module populateRxQueue
  populateRxQueue_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 36,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => populateRxQueue_call_reqs,
      call_acks => populateRxQueue_call_acks,
      return_reqs => populateRxQueue_return_reqs,
      return_acks => populateRxQueue_return_acks,
      call_data  => populateRxQueue_call_data,
      call_tag  => populateRxQueue_call_tag,
      return_tag  => populateRxQueue_return_tag,
      call_mtag => populateRxQueue_tag_in,
      return_mtag => populateRxQueue_tag_out,
      call_mreq => populateRxQueue_start_req,
      call_mack => populateRxQueue_start_ack,
      return_mreq => populateRxQueue_fin_req,
      return_mack => populateRxQueue_fin_ack,
      call_mdata => populateRxQueue_in_args,
      clk => clk, 
      reset => reset --
    ); --
  populateRxQueue_instance:populateRxQueue-- 
    generic map(tag_length => 2)
    port map(-- 
      rx_buffer_pointer => populateRxQueue_rx_buffer_pointer,
      start_req => populateRxQueue_start_req,
      start_ack => populateRxQueue_start_ack,
      fin_req => populateRxQueue_fin_req,
      fin_ack => populateRxQueue_fin_ack,
      clk => clk,
      reset => reset,
      LAST_WRITTEN_RX_QUEUE_INDEX => LAST_WRITTEN_RX_QUEUE_INDEX,
      NUMBER_OF_SERVERS => NUMBER_OF_SERVERS,
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req(1 downto 1),
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack(1 downto 1),
      LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data(11 downto 6),
      AccessRegister_call_reqs => AccessRegister_call_reqs(6 downto 6),
      AccessRegister_call_acks => AccessRegister_call_acks(6 downto 6),
      AccessRegister_call_data => AccessRegister_call_data(300 downto 258),
      AccessRegister_call_tag => AccessRegister_call_tag(13 downto 12),
      AccessRegister_return_reqs => AccessRegister_return_reqs(6 downto 6),
      AccessRegister_return_acks => AccessRegister_return_acks(6 downto 6),
      AccessRegister_return_data => AccessRegister_return_data(223 downto 192),
      AccessRegister_return_tag => AccessRegister_return_tag(13 downto 12),
      pushIntoQueue_call_reqs => pushIntoQueue_call_reqs(2 downto 2),
      pushIntoQueue_call_acks => pushIntoQueue_call_acks(2 downto 2),
      pushIntoQueue_call_data => pushIntoQueue_call_data(206 downto 138),
      pushIntoQueue_call_tag => pushIntoQueue_call_tag(2 downto 2),
      pushIntoQueue_return_reqs => pushIntoQueue_return_reqs(2 downto 2),
      pushIntoQueue_return_acks => pushIntoQueue_return_acks(2 downto 2),
      pushIntoQueue_return_data => pushIntoQueue_return_data(2 downto 2),
      pushIntoQueue_return_tag => pushIntoQueue_return_tag(2 downto 2),
      tag_in => populateRxQueue_tag_in,
      tag_out => populateRxQueue_tag_out-- 
    ); -- 
  -- module pushIntoQueue
  pushIntoQueue_lock <= pushIntoQueue_in_args(68 downto 68);
  pushIntoQueue_q_base_address <= pushIntoQueue_in_args(67 downto 32);
  pushIntoQueue_q_w_data <= pushIntoQueue_in_args(31 downto 0);
  pushIntoQueue_out_args <= pushIntoQueue_status ;
  -- call arbiter for module pushIntoQueue
  pushIntoQueue_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 3,
      call_data_width => 69,
      return_data_width => 1,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => pushIntoQueue_call_reqs,
      call_acks => pushIntoQueue_call_acks,
      return_reqs => pushIntoQueue_return_reqs,
      return_acks => pushIntoQueue_return_acks,
      call_data  => pushIntoQueue_call_data,
      call_tag  => pushIntoQueue_call_tag,
      return_tag  => pushIntoQueue_return_tag,
      call_mtag => pushIntoQueue_tag_in,
      return_mtag => pushIntoQueue_tag_out,
      return_data =>pushIntoQueue_return_data,
      call_mreq => pushIntoQueue_start_req,
      call_mack => pushIntoQueue_start_ack,
      return_mreq => pushIntoQueue_fin_req,
      return_mack => pushIntoQueue_fin_ack,
      call_mdata => pushIntoQueue_in_args,
      return_mdata => pushIntoQueue_out_args,
      clk => clk, 
      reset => reset --
    ); --
  pushIntoQueue_instance:pushIntoQueue-- 
    generic map(tag_length => 3)
    port map(-- 
      lock => pushIntoQueue_lock,
      q_base_address => pushIntoQueue_q_base_address,
      q_w_data => pushIntoQueue_q_w_data,
      status => pushIntoQueue_status,
      start_req => pushIntoQueue_start_req,
      start_ack => pushIntoQueue_start_ack,
      fin_req => pushIntoQueue_fin_req,
      fin_ack => pushIntoQueue_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(4 downto 4),
      accessMemory_call_acks => accessMemory_call_acks(4 downto 4),
      accessMemory_call_data => accessMemory_call_data(549 downto 440),
      accessMemory_call_tag => accessMemory_call_tag(14 downto 12),
      accessMemory_return_reqs => accessMemory_return_reqs(4 downto 4),
      accessMemory_return_acks => accessMemory_return_acks(4 downto 4),
      accessMemory_return_data => accessMemory_return_data(319 downto 256),
      accessMemory_return_tag => accessMemory_return_tag(14 downto 12),
      acquireLock_call_reqs => acquireLock_call_reqs(0 downto 0),
      acquireLock_call_acks => acquireLock_call_acks(0 downto 0),
      acquireLock_call_data => acquireLock_call_data(35 downto 0),
      acquireLock_call_tag => acquireLock_call_tag(0 downto 0),
      acquireLock_return_reqs => acquireLock_return_reqs(0 downto 0),
      acquireLock_return_acks => acquireLock_return_acks(0 downto 0),
      acquireLock_return_data => acquireLock_return_data(0 downto 0),
      acquireLock_return_tag => acquireLock_return_tag(0 downto 0),
      getQueuePointers_call_reqs => getQueuePointers_call_reqs(0 downto 0),
      getQueuePointers_call_acks => getQueuePointers_call_acks(0 downto 0),
      getQueuePointers_call_data => getQueuePointers_call_data(35 downto 0),
      getQueuePointers_call_tag => getQueuePointers_call_tag(0 downto 0),
      getQueuePointers_return_reqs => getQueuePointers_return_reqs(0 downto 0),
      getQueuePointers_return_acks => getQueuePointers_return_acks(0 downto 0),
      getQueuePointers_return_data => getQueuePointers_return_data(63 downto 0),
      getQueuePointers_return_tag => getQueuePointers_return_tag(0 downto 0),
      getQueueLength_call_reqs => getQueueLength_call_reqs(0 downto 0),
      getQueueLength_call_acks => getQueueLength_call_acks(0 downto 0),
      getQueueLength_call_data => getQueueLength_call_data(35 downto 0),
      getQueueLength_call_tag => getQueueLength_call_tag(0 downto 0),
      getQueueLength_return_reqs => getQueueLength_return_reqs(0 downto 0),
      getQueueLength_return_acks => getQueueLength_return_acks(0 downto 0),
      getQueueLength_return_data => getQueueLength_return_data(31 downto 0),
      getQueueLength_return_tag => getQueueLength_return_tag(0 downto 0),
      getTotalMessages_call_reqs => getTotalMessages_call_reqs(0 downto 0),
      getTotalMessages_call_acks => getTotalMessages_call_acks(0 downto 0),
      getTotalMessages_call_data => getTotalMessages_call_data(35 downto 0),
      getTotalMessages_call_tag => getTotalMessages_call_tag(0 downto 0),
      getTotalMessages_return_reqs => getTotalMessages_return_reqs(0 downto 0),
      getTotalMessages_return_acks => getTotalMessages_return_acks(0 downto 0),
      getTotalMessages_return_data => getTotalMessages_return_data(31 downto 0),
      getTotalMessages_return_tag => getTotalMessages_return_tag(0 downto 0),
      setQueuePointers_call_reqs => setQueuePointers_call_reqs(0 downto 0),
      setQueuePointers_call_acks => setQueuePointers_call_acks(0 downto 0),
      setQueuePointers_call_data => setQueuePointers_call_data(99 downto 0),
      setQueuePointers_call_tag => setQueuePointers_call_tag(0 downto 0),
      setQueuePointers_return_reqs => setQueuePointers_return_reqs(0 downto 0),
      setQueuePointers_return_acks => setQueuePointers_return_acks(0 downto 0),
      setQueuePointers_return_tag => setQueuePointers_return_tag(0 downto 0),
      updateTotalMessages_call_reqs => updateTotalMessages_call_reqs(0 downto 0),
      updateTotalMessages_call_acks => updateTotalMessages_call_acks(0 downto 0),
      updateTotalMessages_call_data => updateTotalMessages_call_data(67 downto 0),
      updateTotalMessages_call_tag => updateTotalMessages_call_tag(0 downto 0),
      updateTotalMessages_return_reqs => updateTotalMessages_return_reqs(0 downto 0),
      updateTotalMessages_return_acks => updateTotalMessages_return_acks(0 downto 0),
      updateTotalMessages_return_tag => updateTotalMessages_return_tag(0 downto 0),
      releaseLock_call_reqs => releaseLock_call_reqs(0 downto 0),
      releaseLock_call_acks => releaseLock_call_acks(0 downto 0),
      releaseLock_call_data => releaseLock_call_data(35 downto 0),
      releaseLock_call_tag => releaseLock_call_tag(0 downto 0),
      releaseLock_return_reqs => releaseLock_return_reqs(0 downto 0),
      releaseLock_return_acks => releaseLock_return_acks(0 downto 0),
      releaseLock_return_tag => releaseLock_return_tag(0 downto 0),
      setQueueElement_call_reqs => setQueueElement_call_reqs(0 downto 0),
      setQueueElement_call_acks => setQueueElement_call_acks(0 downto 0),
      setQueueElement_call_data => setQueueElement_call_data(99 downto 0),
      setQueueElement_call_tag => setQueueElement_call_tag(0 downto 0),
      setQueueElement_return_reqs => setQueueElement_return_reqs(0 downto 0),
      setQueueElement_return_acks => setQueueElement_return_acks(0 downto 0),
      setQueueElement_return_tag => setQueueElement_return_tag(0 downto 0),
      tag_in => pushIntoQueue_tag_in,
      tag_out => pushIntoQueue_tag_out-- 
    ); -- 
  -- module releaseLock
  releaseLock_q_base_address <= releaseLock_in_args(35 downto 0);
  -- call arbiter for module releaseLock
  releaseLock_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 2,
      call_data_width => 36,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => releaseLock_call_reqs,
      call_acks => releaseLock_call_acks,
      return_reqs => releaseLock_return_reqs,
      return_acks => releaseLock_return_acks,
      call_data  => releaseLock_call_data,
      call_tag  => releaseLock_call_tag,
      return_tag  => releaseLock_return_tag,
      call_mtag => releaseLock_tag_in,
      return_mtag => releaseLock_tag_out,
      call_mreq => releaseLock_start_req,
      call_mack => releaseLock_start_ack,
      return_mreq => releaseLock_fin_req,
      return_mack => releaseLock_fin_ack,
      call_mdata => releaseLock_in_args,
      clk => clk, 
      reset => reset --
    ); --
  releaseLock_instance:releaseLock-- 
    generic map(tag_length => 3)
    port map(-- 
      q_base_address => releaseLock_q_base_address,
      start_req => releaseLock_start_req,
      start_ack => releaseLock_start_ack,
      fin_req => releaseLock_fin_req,
      fin_ack => releaseLock_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(15 downto 15),
      accessMemory_call_acks => accessMemory_call_acks(15 downto 15),
      accessMemory_call_data => accessMemory_call_data(1759 downto 1650),
      accessMemory_call_tag => accessMemory_call_tag(47 downto 45),
      accessMemory_return_reqs => accessMemory_return_reqs(15 downto 15),
      accessMemory_return_acks => accessMemory_return_acks(15 downto 15),
      accessMemory_return_data => accessMemory_return_data(1023 downto 960),
      accessMemory_return_tag => accessMemory_return_tag(47 downto 45),
      tag_in => releaseLock_tag_in,
      tag_out => releaseLock_tag_out-- 
    ); -- 
  -- module setQueueElement
  setQueueElement_q_base_address <= setQueueElement_in_args(99 downto 64);
  setQueueElement_write_index <= setQueueElement_in_args(63 downto 32);
  setQueueElement_q_w_data <= setQueueElement_in_args(31 downto 0);
  -- call arbiter for module setQueueElement
  setQueueElement_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 100,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => setQueueElement_call_reqs,
      call_acks => setQueueElement_call_acks,
      return_reqs => setQueueElement_return_reqs,
      return_acks => setQueueElement_return_acks,
      call_data  => setQueueElement_call_data,
      call_tag  => setQueueElement_call_tag,
      return_tag  => setQueueElement_return_tag,
      call_mtag => setQueueElement_tag_in,
      return_mtag => setQueueElement_tag_out,
      call_mreq => setQueueElement_start_req,
      call_mack => setQueueElement_start_ack,
      return_mreq => setQueueElement_fin_req,
      return_mack => setQueueElement_fin_ack,
      call_mdata => setQueueElement_in_args,
      clk => clk, 
      reset => reset --
    ); --
  setQueueElement_instance:setQueueElement-- 
    generic map(tag_length => 2)
    port map(-- 
      q_base_address => setQueueElement_q_base_address,
      write_index => setQueueElement_write_index,
      q_w_data => setQueueElement_q_w_data,
      start_req => setQueueElement_start_req,
      start_ack => setQueueElement_start_ack,
      fin_req => setQueueElement_fin_req,
      fin_ack => setQueueElement_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(3 downto 3),
      accessMemory_call_acks => accessMemory_call_acks(3 downto 3),
      accessMemory_call_data => accessMemory_call_data(439 downto 330),
      accessMemory_call_tag => accessMemory_call_tag(11 downto 9),
      accessMemory_return_reqs => accessMemory_return_reqs(3 downto 3),
      accessMemory_return_acks => accessMemory_return_acks(3 downto 3),
      accessMemory_return_data => accessMemory_return_data(255 downto 192),
      accessMemory_return_tag => accessMemory_return_tag(11 downto 9),
      tag_in => setQueueElement_tag_in,
      tag_out => setQueueElement_tag_out-- 
    ); -- 
  -- module setQueuePointers
  setQueuePointers_q_base_address <= setQueuePointers_in_args(99 downto 64);
  setQueuePointers_wp <= setQueuePointers_in_args(63 downto 32);
  setQueuePointers_rp <= setQueuePointers_in_args(31 downto 0);
  -- call arbiter for module setQueuePointers
  setQueuePointers_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 2,
      call_data_width => 100,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => setQueuePointers_call_reqs,
      call_acks => setQueuePointers_call_acks,
      return_reqs => setQueuePointers_return_reqs,
      return_acks => setQueuePointers_return_acks,
      call_data  => setQueuePointers_call_data,
      call_tag  => setQueuePointers_call_tag,
      return_tag  => setQueuePointers_return_tag,
      call_mtag => setQueuePointers_tag_in,
      return_mtag => setQueuePointers_tag_out,
      call_mreq => setQueuePointers_start_req,
      call_mack => setQueuePointers_start_ack,
      return_mreq => setQueuePointers_fin_req,
      return_mack => setQueuePointers_fin_ack,
      call_mdata => setQueuePointers_in_args,
      clk => clk, 
      reset => reset --
    ); --
  setQueuePointers_instance:setQueuePointers-- 
    generic map(tag_length => 3)
    port map(-- 
      q_base_address => setQueuePointers_q_base_address,
      wp => setQueuePointers_wp,
      rp => setQueuePointers_rp,
      start_req => setQueuePointers_start_req,
      start_ack => setQueuePointers_start_ack,
      fin_req => setQueuePointers_fin_req,
      fin_ack => setQueuePointers_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(14 downto 14),
      accessMemory_call_acks => accessMemory_call_acks(14 downto 14),
      accessMemory_call_data => accessMemory_call_data(1649 downto 1540),
      accessMemory_call_tag => accessMemory_call_tag(44 downto 42),
      accessMemory_return_reqs => accessMemory_return_reqs(14 downto 14),
      accessMemory_return_acks => accessMemory_return_acks(14 downto 14),
      accessMemory_return_data => accessMemory_return_data(959 downto 896),
      accessMemory_return_tag => accessMemory_return_tag(44 downto 42),
      tag_in => setQueuePointers_tag_in,
      tag_out => setQueuePointers_tag_out-- 
    ); -- 
  -- module transmitEngineDaemon
  transmitEngineDaemon_instance:transmitEngineDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => transmitEngineDaemon_start_req,
      start_ack => transmitEngineDaemon_start_ack,
      fin_req => transmitEngineDaemon_fin_req,
      fin_ack => transmitEngineDaemon_fin_ack,
      clk => clk,
      reset => reset,
      CONTROL_REGISTER => CONTROL_REGISTER,
      FREE_Q => FREE_Q,
      LAST_READ_TX_QUEUE_INDEX => LAST_READ_TX_QUEUE_INDEX,
      NUMBER_OF_SERVERS => NUMBER_OF_SERVERS,
      LAST_READ_TX_QUEUE_INDEX_pipe_write_req => LAST_READ_TX_QUEUE_INDEX_pipe_write_req(1 downto 0),
      LAST_READ_TX_QUEUE_INDEX_pipe_write_ack => LAST_READ_TX_QUEUE_INDEX_pipe_write_ack(1 downto 0),
      LAST_READ_TX_QUEUE_INDEX_pipe_write_data => LAST_READ_TX_QUEUE_INDEX_pipe_write_data(11 downto 0),
      AccessRegister_call_reqs => AccessRegister_call_reqs(0 downto 0),
      AccessRegister_call_acks => AccessRegister_call_acks(0 downto 0),
      AccessRegister_call_data => AccessRegister_call_data(42 downto 0),
      AccessRegister_call_tag => AccessRegister_call_tag(1 downto 0),
      AccessRegister_return_reqs => AccessRegister_return_reqs(0 downto 0),
      AccessRegister_return_acks => AccessRegister_return_acks(0 downto 0),
      AccessRegister_return_data => AccessRegister_return_data(31 downto 0),
      AccessRegister_return_tag => AccessRegister_return_tag(1 downto 0),
      pushIntoQueue_call_reqs => pushIntoQueue_call_reqs(0 downto 0),
      pushIntoQueue_call_acks => pushIntoQueue_call_acks(0 downto 0),
      pushIntoQueue_call_data => pushIntoQueue_call_data(68 downto 0),
      pushIntoQueue_call_tag => pushIntoQueue_call_tag(0 downto 0),
      pushIntoQueue_return_reqs => pushIntoQueue_return_reqs(0 downto 0),
      pushIntoQueue_return_acks => pushIntoQueue_return_acks(0 downto 0),
      pushIntoQueue_return_data => pushIntoQueue_return_data(0 downto 0),
      pushIntoQueue_return_tag => pushIntoQueue_return_tag(0 downto 0),
      getTxPacketPointerFromServer_call_reqs => getTxPacketPointerFromServer_call_reqs(0 downto 0),
      getTxPacketPointerFromServer_call_acks => getTxPacketPointerFromServer_call_acks(0 downto 0),
      getTxPacketPointerFromServer_call_data => getTxPacketPointerFromServer_call_data(5 downto 0),
      getTxPacketPointerFromServer_call_tag => getTxPacketPointerFromServer_call_tag(0 downto 0),
      getTxPacketPointerFromServer_return_reqs => getTxPacketPointerFromServer_return_reqs(0 downto 0),
      getTxPacketPointerFromServer_return_acks => getTxPacketPointerFromServer_return_acks(0 downto 0),
      getTxPacketPointerFromServer_return_data => getTxPacketPointerFromServer_return_data(32 downto 0),
      getTxPacketPointerFromServer_return_tag => getTxPacketPointerFromServer_return_tag(0 downto 0),
      transmitPacket_call_reqs => transmitPacket_call_reqs(0 downto 0),
      transmitPacket_call_acks => transmitPacket_call_acks(0 downto 0),
      transmitPacket_call_data => transmitPacket_call_data(31 downto 0),
      transmitPacket_call_tag => transmitPacket_call_tag(0 downto 0),
      transmitPacket_return_reqs => transmitPacket_return_reqs(0 downto 0),
      transmitPacket_return_acks => transmitPacket_return_acks(0 downto 0),
      transmitPacket_return_data => transmitPacket_return_data(0 downto 0),
      transmitPacket_return_tag => transmitPacket_return_tag(0 downto 0),
      tag_in => transmitEngineDaemon_tag_in,
      tag_out => transmitEngineDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  transmitEngineDaemon_tag_in <= (others => '0');
  transmitEngineDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => transmitEngineDaemon_start_req, start_ack => transmitEngineDaemon_start_ack,  fin_req => transmitEngineDaemon_fin_req,  fin_ack => transmitEngineDaemon_fin_ack);
  -- module transmitPacket
  transmitPacket_packet_pointer <= transmitPacket_in_args(31 downto 0);
  transmitPacket_out_args <= transmitPacket_status ;
  -- call arbiter for module transmitPacket
  transmitPacket_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 32,
      return_data_width => 1,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => transmitPacket_call_reqs,
      call_acks => transmitPacket_call_acks,
      return_reqs => transmitPacket_return_reqs,
      return_acks => transmitPacket_return_acks,
      call_data  => transmitPacket_call_data,
      call_tag  => transmitPacket_call_tag,
      return_tag  => transmitPacket_return_tag,
      call_mtag => transmitPacket_tag_in,
      return_mtag => transmitPacket_tag_out,
      return_data =>transmitPacket_return_data,
      call_mreq => transmitPacket_start_req,
      call_mack => transmitPacket_start_ack,
      return_mreq => transmitPacket_fin_req,
      return_mack => transmitPacket_fin_ack,
      call_mdata => transmitPacket_in_args,
      return_mdata => transmitPacket_out_args,
      clk => clk, 
      reset => reset --
    ); --
  transmitPacket_instance:transmitPacket-- 
    generic map(tag_length => 2)
    port map(-- 
      packet_pointer => transmitPacket_packet_pointer,
      status => transmitPacket_status,
      start_req => transmitPacket_start_req,
      start_ack => transmitPacket_start_ack,
      fin_req => transmitPacket_fin_req,
      fin_ack => transmitPacket_fin_ack,
      clk => clk,
      reset => reset,
      nic_to_mac_transmit_pipe_pipe_write_req => nic_to_mac_transmit_pipe_pipe_write_req(1 downto 0),
      nic_to_mac_transmit_pipe_pipe_write_ack => nic_to_mac_transmit_pipe_pipe_write_ack(1 downto 0),
      nic_to_mac_transmit_pipe_pipe_write_data => nic_to_mac_transmit_pipe_pipe_write_data(145 downto 0),
      AccessRegister_call_reqs => AccessRegister_call_reqs(1 downto 1),
      AccessRegister_call_acks => AccessRegister_call_acks(1 downto 1),
      AccessRegister_call_data => AccessRegister_call_data(85 downto 43),
      AccessRegister_call_tag => AccessRegister_call_tag(3 downto 2),
      AccessRegister_return_reqs => AccessRegister_return_reqs(1 downto 1),
      AccessRegister_return_acks => AccessRegister_return_acks(1 downto 1),
      AccessRegister_return_data => AccessRegister_return_data(63 downto 32),
      AccessRegister_return_tag => AccessRegister_return_tag(3 downto 2),
      accessMemory_call_reqs => accessMemory_call_reqs(1 downto 0),
      accessMemory_call_acks => accessMemory_call_acks(1 downto 0),
      accessMemory_call_data => accessMemory_call_data(219 downto 0),
      accessMemory_call_tag => accessMemory_call_tag(5 downto 0),
      accessMemory_return_reqs => accessMemory_return_reqs(1 downto 0),
      accessMemory_return_acks => accessMemory_return_acks(1 downto 0),
      accessMemory_return_data => accessMemory_return_data(127 downto 0),
      accessMemory_return_tag => accessMemory_return_tag(5 downto 0),
      tag_in => transmitPacket_tag_in,
      tag_out => transmitPacket_tag_out-- 
    ); -- 
  -- module updateTotalMessages
  updateTotalMessages_q_base_address <= updateTotalMessages_in_args(67 downto 32);
  updateTotalMessages_updated_total_msgs <= updateTotalMessages_in_args(31 downto 0);
  -- call arbiter for module updateTotalMessages
  updateTotalMessages_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 2,
      call_data_width => 68,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => updateTotalMessages_call_reqs,
      call_acks => updateTotalMessages_call_acks,
      return_reqs => updateTotalMessages_return_reqs,
      return_acks => updateTotalMessages_return_acks,
      call_data  => updateTotalMessages_call_data,
      call_tag  => updateTotalMessages_call_tag,
      return_tag  => updateTotalMessages_return_tag,
      call_mtag => updateTotalMessages_tag_in,
      return_mtag => updateTotalMessages_tag_out,
      call_mreq => updateTotalMessages_start_req,
      call_mack => updateTotalMessages_start_ack,
      return_mreq => updateTotalMessages_fin_req,
      return_mack => updateTotalMessages_fin_ack,
      call_mdata => updateTotalMessages_in_args,
      clk => clk, 
      reset => reset --
    ); --
  updateTotalMessages_instance:updateTotalMessages-- 
    generic map(tag_length => 3)
    port map(-- 
      q_base_address => updateTotalMessages_q_base_address,
      updated_total_msgs => updateTotalMessages_updated_total_msgs,
      start_req => updateTotalMessages_start_req,
      start_ack => updateTotalMessages_start_ack,
      fin_req => updateTotalMessages_fin_req,
      fin_ack => updateTotalMessages_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(12 downto 12),
      accessMemory_call_acks => accessMemory_call_acks(12 downto 12),
      accessMemory_call_data => accessMemory_call_data(1429 downto 1320),
      accessMemory_call_tag => accessMemory_call_tag(38 downto 36),
      accessMemory_return_reqs => accessMemory_return_reqs(12 downto 12),
      accessMemory_return_acks => accessMemory_return_acks(12 downto 12),
      accessMemory_return_data => accessMemory_return_data(831 downto 768),
      accessMemory_return_tag => accessMemory_return_tag(38 downto 36),
      tag_in => updateTotalMessages_tag_in,
      tag_out => updateTotalMessages_tag_out-- 
    ); -- 
  -- module writeControlInformationToMem
  writeControlInformationToMem_base_buffer_pointer <= writeControlInformationToMem_in_args(54 downto 19);
  writeControlInformationToMem_packet_size <= writeControlInformationToMem_in_args(18 downto 8);
  writeControlInformationToMem_last_keep <= writeControlInformationToMem_in_args(7 downto 0);
  -- call arbiter for module writeControlInformationToMem
  writeControlInformationToMem_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 55,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => writeControlInformationToMem_call_reqs,
      call_acks => writeControlInformationToMem_call_acks,
      return_reqs => writeControlInformationToMem_return_reqs,
      return_acks => writeControlInformationToMem_return_acks,
      call_data  => writeControlInformationToMem_call_data,
      call_tag  => writeControlInformationToMem_call_tag,
      return_tag  => writeControlInformationToMem_return_tag,
      call_mtag => writeControlInformationToMem_tag_in,
      return_mtag => writeControlInformationToMem_tag_out,
      call_mreq => writeControlInformationToMem_start_req,
      call_mack => writeControlInformationToMem_start_ack,
      return_mreq => writeControlInformationToMem_fin_req,
      return_mack => writeControlInformationToMem_fin_ack,
      call_mdata => writeControlInformationToMem_in_args,
      clk => clk, 
      reset => reset --
    ); --
  writeControlInformationToMem_instance:writeControlInformationToMem-- 
    generic map(tag_length => 2)
    port map(-- 
      base_buffer_pointer => writeControlInformationToMem_base_buffer_pointer,
      packet_size => writeControlInformationToMem_packet_size,
      last_keep => writeControlInformationToMem_last_keep,
      start_req => writeControlInformationToMem_start_req,
      start_ack => writeControlInformationToMem_start_ack,
      fin_req => writeControlInformationToMem_fin_req,
      fin_ack => writeControlInformationToMem_fin_ack,
      clk => clk,
      reset => reset,
      accessMemory_call_reqs => accessMemory_call_reqs(2 downto 2),
      accessMemory_call_acks => accessMemory_call_acks(2 downto 2),
      accessMemory_call_data => accessMemory_call_data(329 downto 220),
      accessMemory_call_tag => accessMemory_call_tag(8 downto 6),
      accessMemory_return_reqs => accessMemory_return_reqs(2 downto 2),
      accessMemory_return_acks => accessMemory_return_acks(2 downto 2),
      accessMemory_return_data => accessMemory_return_data(191 downto 128),
      accessMemory_return_tag => accessMemory_return_tag(8 downto 6),
      tag_in => writeControlInformationToMem_tag_in,
      tag_out => writeControlInformationToMem_tag_out-- 
    ); -- 
  -- module writeEthernetHeaderToMem
  writeEthernetHeaderToMem_buf_pointer <= writeEthernetHeaderToMem_in_args(35 downto 0);
  writeEthernetHeaderToMem_out_args <= writeEthernetHeaderToMem_buf_position_out ;
  -- call arbiter for module writeEthernetHeaderToMem
  writeEthernetHeaderToMem_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 36,
      return_data_width => 36,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => writeEthernetHeaderToMem_call_reqs,
      call_acks => writeEthernetHeaderToMem_call_acks,
      return_reqs => writeEthernetHeaderToMem_return_reqs,
      return_acks => writeEthernetHeaderToMem_return_acks,
      call_data  => writeEthernetHeaderToMem_call_data,
      call_tag  => writeEthernetHeaderToMem_call_tag,
      return_tag  => writeEthernetHeaderToMem_return_tag,
      call_mtag => writeEthernetHeaderToMem_tag_in,
      return_mtag => writeEthernetHeaderToMem_tag_out,
      return_data =>writeEthernetHeaderToMem_return_data,
      call_mreq => writeEthernetHeaderToMem_start_req,
      call_mack => writeEthernetHeaderToMem_start_ack,
      return_mreq => writeEthernetHeaderToMem_fin_req,
      return_mack => writeEthernetHeaderToMem_fin_ack,
      call_mdata => writeEthernetHeaderToMem_in_args,
      return_mdata => writeEthernetHeaderToMem_out_args,
      clk => clk, 
      reset => reset --
    ); --
  writeEthernetHeaderToMem_instance:writeEthernetHeaderToMem-- 
    generic map(tag_length => 2)
    port map(-- 
      buf_pointer => writeEthernetHeaderToMem_buf_pointer,
      buf_position_out => writeEthernetHeaderToMem_buf_position_out,
      start_req => writeEthernetHeaderToMem_start_req,
      start_ack => writeEthernetHeaderToMem_start_ack,
      fin_req => writeEthernetHeaderToMem_fin_req,
      fin_ack => writeEthernetHeaderToMem_fin_ack,
      clk => clk,
      reset => reset,
      nic_rx_to_header_pipe_read_req => nic_rx_to_header_pipe_read_req(0 downto 0),
      nic_rx_to_header_pipe_read_ack => nic_rx_to_header_pipe_read_ack(0 downto 0),
      nic_rx_to_header_pipe_read_data => nic_rx_to_header_pipe_read_data(72 downto 0),
      accessMemory_call_reqs => accessMemory_call_reqs(5 downto 5),
      accessMemory_call_acks => accessMemory_call_acks(5 downto 5),
      accessMemory_call_data => accessMemory_call_data(659 downto 550),
      accessMemory_call_tag => accessMemory_call_tag(17 downto 15),
      accessMemory_return_reqs => accessMemory_return_reqs(5 downto 5),
      accessMemory_return_acks => accessMemory_return_acks(5 downto 5),
      accessMemory_return_data => accessMemory_return_data(383 downto 320),
      accessMemory_return_tag => accessMemory_return_tag(17 downto 15),
      tag_in => writeEthernetHeaderToMem_tag_in,
      tag_out => writeEthernetHeaderToMem_tag_out-- 
    ); -- 
  -- module writePayloadToMem
  writePayloadToMem_base_buf_pointer <= writePayloadToMem_in_args(71 downto 36);
  writePayloadToMem_buf_pointer <= writePayloadToMem_in_args(35 downto 0);
  writePayloadToMem_out_args <= writePayloadToMem_packet_size_32 & writePayloadToMem_bad_packet_identifier & writePayloadToMem_last_keep ;
  -- call arbiter for module writePayloadToMem
  writePayloadToMem_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 72,
      return_data_width => 20,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => writePayloadToMem_call_reqs,
      call_acks => writePayloadToMem_call_acks,
      return_reqs => writePayloadToMem_return_reqs,
      return_acks => writePayloadToMem_return_acks,
      call_data  => writePayloadToMem_call_data,
      call_tag  => writePayloadToMem_call_tag,
      return_tag  => writePayloadToMem_return_tag,
      call_mtag => writePayloadToMem_tag_in,
      return_mtag => writePayloadToMem_tag_out,
      return_data =>writePayloadToMem_return_data,
      call_mreq => writePayloadToMem_start_req,
      call_mack => writePayloadToMem_start_ack,
      return_mreq => writePayloadToMem_fin_req,
      return_mack => writePayloadToMem_fin_ack,
      call_mdata => writePayloadToMem_in_args,
      return_mdata => writePayloadToMem_out_args,
      clk => clk, 
      reset => reset --
    ); --
  writePayloadToMem_instance:writePayloadToMem-- 
    generic map(tag_length => 2)
    port map(-- 
      base_buf_pointer => writePayloadToMem_base_buf_pointer,
      buf_pointer => writePayloadToMem_buf_pointer,
      packet_size_32 => writePayloadToMem_packet_size_32,
      bad_packet_identifier => writePayloadToMem_bad_packet_identifier,
      last_keep => writePayloadToMem_last_keep,
      start_req => writePayloadToMem_start_req,
      start_ack => writePayloadToMem_start_ack,
      fin_req => writePayloadToMem_fin_req,
      fin_ack => writePayloadToMem_fin_ack,
      clk => clk,
      reset => reset,
      nic_rx_to_packet_pipe_read_req => nic_rx_to_packet_pipe_read_req(0 downto 0),
      nic_rx_to_packet_pipe_read_ack => nic_rx_to_packet_pipe_read_ack(0 downto 0),
      nic_rx_to_packet_pipe_read_data => nic_rx_to_packet_pipe_read_data(72 downto 0),
      accessMemory_call_reqs => accessMemory_call_reqs(6 downto 6),
      accessMemory_call_acks => accessMemory_call_acks(6 downto 6),
      accessMemory_call_data => accessMemory_call_data(769 downto 660),
      accessMemory_call_tag => accessMemory_call_tag(20 downto 18),
      accessMemory_return_reqs => accessMemory_return_reqs(6 downto 6),
      accessMemory_return_acks => accessMemory_return_acks(6 downto 6),
      accessMemory_return_data => accessMemory_return_data(447 downto 384),
      accessMemory_return_tag => accessMemory_return_tag(20 downto 18),
      tag_in => writePayloadToMem_tag_in,
      tag_out => writePayloadToMem_tag_out-- 
    ); -- 
  AFB_NIC_REQUEST_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe AFB_NIC_REQUEST",
      num_reads => 1,
      num_writes => 1,
      data_width => 74,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => AFB_NIC_REQUEST_pipe_read_req,
      read_ack => AFB_NIC_REQUEST_pipe_read_ack,
      read_data => AFB_NIC_REQUEST_pipe_read_data,
      write_req => AFB_NIC_REQUEST_pipe_write_req,
      write_ack => AFB_NIC_REQUEST_pipe_write_ack,
      write_data => AFB_NIC_REQUEST_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  AFB_NIC_RESPONSE_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe AFB_NIC_RESPONSE",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => AFB_NIC_RESPONSE_pipe_read_req,
      read_ack => AFB_NIC_RESPONSE_pipe_read_ack,
      read_data => AFB_NIC_RESPONSE_pipe_read_data,
      write_req => AFB_NIC_RESPONSE_pipe_write_req,
      write_ack => AFB_NIC_RESPONSE_pipe_write_ack,
      write_data => AFB_NIC_RESPONSE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  CONTROL_REGISTER_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe CONTROL_REGISTER",
      volatile_flag => false,
      num_writes => 1,
      data_width => 32 --
    ) 
    port map( -- 
      read_data => CONTROL_REGISTER,
      write_req => CONTROL_REGISTER_pipe_write_req,
      write_ack => CONTROL_REGISTER_pipe_write_ack,
      write_data => CONTROL_REGISTER_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  FREE_Q_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe FREE_Q",
      volatile_flag => false,
      num_writes => 1,
      data_width => 36 --
    ) 
    port map( -- 
      read_data => FREE_Q,
      write_req => FREE_Q_pipe_write_req,
      write_ack => FREE_Q_pipe_write_ack,
      write_data => FREE_Q_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  LAST_READ_TX_QUEUE_INDEX_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe LAST_READ_TX_QUEUE_INDEX",
      volatile_flag => false,
      num_writes => 2,
      data_width => 6 --
    ) 
    port map( -- 
      read_data => LAST_READ_TX_QUEUE_INDEX,
      write_req => LAST_READ_TX_QUEUE_INDEX_pipe_write_req,
      write_ack => LAST_READ_TX_QUEUE_INDEX_pipe_write_ack,
      write_data => LAST_READ_TX_QUEUE_INDEX_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  LAST_WRITTEN_RX_QUEUE_INDEX_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe LAST_WRITTEN_RX_QUEUE_INDEX",
      volatile_flag => false,
      num_writes => 2,
      data_width => 6 --
    ) 
    port map( -- 
      read_data => LAST_WRITTEN_RX_QUEUE_INDEX,
      write_req => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_req,
      write_ack => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_ack,
      write_data => LAST_WRITTEN_RX_QUEUE_INDEX_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  MAC_ENABLE_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe MAC_ENABLE",
      volatile_flag => false,
      num_writes => 1,
      data_width => 1 --
    ) 
    port map( -- 
      read_data => MAC_ENABLE,
      write_req => MAC_ENABLE_pipe_write_req,
      write_ack => MAC_ENABLE_pipe_write_ack,
      write_data => MAC_ENABLE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  MEMORY_TO_NIC_RESPONSE_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe MEMORY_TO_NIC_RESPONSE",
      num_reads => 1,
      num_writes => 1,
      data_width => 65,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => MEMORY_TO_NIC_RESPONSE_pipe_read_req,
      read_ack => MEMORY_TO_NIC_RESPONSE_pipe_read_ack,
      read_data => MEMORY_TO_NIC_RESPONSE_pipe_read_data,
      write_req => MEMORY_TO_NIC_RESPONSE_pipe_write_req,
      write_ack => MEMORY_TO_NIC_RESPONSE_pipe_write_ack,
      write_data => MEMORY_TO_NIC_RESPONSE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  NIC_REQUEST_REGISTER_ACCESS_PIPE_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe NIC_REQUEST_REGISTER_ACCESS_PIPE",
      num_reads => 1,
      num_writes => 1,
      data_width => 43,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_req,
      read_ack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_ack,
      read_data => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_read_data,
      write_req => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_req,
      write_ack => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_ack,
      write_data => NIC_REQUEST_REGISTER_ACCESS_PIPE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  NIC_RESPONSE_REGISTER_ACCESS_PIPE_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe NIC_RESPONSE_REGISTER_ACCESS_PIPE",
      num_reads => 1,
      num_writes => 1,
      data_width => 33,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_req,
      read_ack => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_ack,
      read_data => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_read_data,
      write_req => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_req,
      write_ack => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_ack,
      write_data => NIC_RESPONSE_REGISTER_ACCESS_PIPE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  NIC_TO_MEMORY_REQUEST_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe NIC_TO_MEMORY_REQUEST",
      num_reads => 1,
      num_writes => 1,
      data_width => 110,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => NIC_TO_MEMORY_REQUEST_pipe_read_req,
      read_ack => NIC_TO_MEMORY_REQUEST_pipe_read_ack,
      read_data => NIC_TO_MEMORY_REQUEST_pipe_read_data,
      write_req => NIC_TO_MEMORY_REQUEST_pipe_write_req,
      write_ack => NIC_TO_MEMORY_REQUEST_pipe_write_ack,
      write_data => NIC_TO_MEMORY_REQUEST_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  NUMBER_OF_SERVERS_Signal: SignalBase -- 
    generic map( -- 
      name => "pipe NUMBER_OF_SERVERS",
      volatile_flag => false,
      num_writes => 1,
      data_width => 32 --
    ) 
    port map( -- 
      read_data => NUMBER_OF_SERVERS,
      write_req => NUMBER_OF_SERVERS_pipe_write_req,
      write_ack => NUMBER_OF_SERVERS_pipe_write_ack,
      write_data => NUMBER_OF_SERVERS_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  enable_mac_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe enable_mac",
      num_reads => 1,
      num_writes => 1,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => enable_mac_pipe_read_req,
      read_ack => enable_mac_pipe_read_ack,
      read_data => enable_mac_pipe_read_data,
      write_req => enable_mac_pipe_write_req,
      write_ack => enable_mac_pipe_write_ack,
      write_data => enable_mac_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  mac_to_nic_data_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe mac_to_nic_data",
      num_reads => 1,
      num_writes => 1,
      data_width => 73,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => mac_to_nic_data_pipe_read_req,
      read_ack => mac_to_nic_data_pipe_read_ack,
      read_data => mac_to_nic_data_pipe_read_data,
      write_req => mac_to_nic_data_pipe_write_req,
      write_ack => mac_to_nic_data_pipe_write_ack,
      write_data => mac_to_nic_data_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  nic_rx_to_header_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe nic_rx_to_header",
      num_reads => 1,
      num_writes => 1,
      data_width => 73,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => nic_rx_to_header_pipe_read_req,
      read_ack => nic_rx_to_header_pipe_read_ack,
      read_data => nic_rx_to_header_pipe_read_data,
      write_req => nic_rx_to_header_pipe_write_req,
      write_ack => nic_rx_to_header_pipe_write_ack,
      write_data => nic_rx_to_header_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  nic_rx_to_packet_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe nic_rx_to_packet",
      num_reads => 1,
      num_writes => 1,
      data_width => 73,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => nic_rx_to_packet_pipe_read_req,
      read_ack => nic_rx_to_packet_pipe_read_ack,
      read_data => nic_rx_to_packet_pipe_read_data,
      write_req => nic_rx_to_packet_pipe_write_req,
      write_ack => nic_rx_to_packet_pipe_write_ack,
      write_data => nic_rx_to_packet_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  nic_to_mac_transmit_pipe_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe nic_to_mac_transmit_pipe",
      num_reads => 1,
      num_writes => 2,
      data_width => 73,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 2 --
    )
    port map( -- 
      read_req => nic_to_mac_transmit_pipe_pipe_read_req,
      read_ack => nic_to_mac_transmit_pipe_pipe_read_ack,
      read_data => nic_to_mac_transmit_pipe_pipe_read_data,
      write_req => nic_to_mac_transmit_pipe_pipe_write_req,
      write_ack => nic_to_mac_transmit_pipe_pipe_write_ack,
      write_data => nic_to_mac_transmit_pipe_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  MemorySpace_memory_space_2: ordered_memory_subsystem -- 
    generic map(-- 
      name => "memory_space_2",
      num_loads => 2,
      num_stores => 2,
      addr_width => 6,
      data_width => 32,
      tag_width => 3,
      time_stamp_width => 18,
      number_of_banks => 1,
      mux_degree => 2,
      demux_degree => 2,
      base_bank_addr_width => 6,
      base_bank_data_width => 32
      ) -- 
    port map(-- 
      lr_addr_in => memory_space_2_lr_addr,
      lr_req_in => memory_space_2_lr_req,
      lr_ack_out => memory_space_2_lr_ack,
      lr_tag_in => memory_space_2_lr_tag,
      lc_req_in => memory_space_2_lc_req,
      lc_ack_out => memory_space_2_lc_ack,
      lc_data_out => memory_space_2_lc_data,
      lc_tag_out => memory_space_2_lc_tag,
      sr_addr_in => memory_space_2_sr_addr,
      sr_data_in => memory_space_2_sr_data,
      sr_req_in => memory_space_2_sr_req,
      sr_ack_out => memory_space_2_sr_ack,
      sr_tag_in => memory_space_2_sr_tag,
      sc_req_in=> memory_space_2_sc_req,
      sc_ack_out => memory_space_2_sc_ack,
      sc_tag_out => memory_space_2_sc_tag,
      clock => clk,
      reset => reset); -- 
  -- 
end nic_system_arch;

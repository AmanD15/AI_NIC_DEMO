

`protect begin_protected
`protect version = 1
`protect encrypt_agent = "XILINX"
`protect encrypt_agent_info = "Xilinx Encryption Tool 2014"
`protect key_keyowner = "Cadence Design Systems.", key_keyname= "cds_rsa_key", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 64)
`protect key_block
hYn4T1Tz8lmB8loeGYuHmgEJp5TdMkRKn5tdK0Pxo3wkkBR/aG2es4RXT0Kx9IkGgy2jVWVPoeKB
usRl+M6Pxw==


`protect key_keyowner = "Mentor Graphics Corporation", key_keyname= "MGC-VERIF-SIM-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
cZOTsELKZdXMGraSgAw9rgqxvSLbW0aT2lTeYBbmmRdIiILVX40Q3XF89sXvrmWq2q7dAJSXvpsX
1JIpxbCUMi40Nuru7hdg9WkNNMs1Q8UJCou9g/GNLxJnh56Wx2JqOiplBqlgeaLjd0T16sGmIYm4
kTNGsNPOASR/dWaldsE=


`protect key_keyowner = "Synopsys", key_keyname= "SNPS-VCS-RSA-1", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 128)
`protect key_block
o6ehD67QiTZFs1auOjL5nkbDEbn3neiXmbyTqqoQKK+v0TaPL6hSxGHE/Fz3NtmR3RIza9+Y9rVH
Je7RNuyq8vsgofAGK5Qpf28P/9kF6eDh0JgLJHOonk7lnG+gufS3pMHIfioCEe/2wyoIxzbwUPNl
TCIJtbzDvWpcCIKBgiQ=


`protect key_keyowner = "Aldec", key_keyname= "ALDEC15_001", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
cASOe3RHelXhU6s/jEEqAnadTjmj4ihjbMuYb8YjKT8lAROht6xaHEt/3WXUlUPXIpDwtJlexClV
csQVUSlNShzZmxBI5epxH/HJqLhQYwkRDFK2BUAagxn++cS1iWJGlow9Gha0EU+PfllVje3OWy4O
LbiqHgQlEG6sIGo0ZCj6KPC87SBAytHtAiVRpovpGAxLS/DLeXSJaavSSwOc7nmWFDaNEi9dJS9i
qixZxDI5QNaDp3uaBFLzKqo9oSPgNj1mYKRZp6XL0ganfqQCHh/snCyymi+o0DC5vSM/+RtCZHXA
A1u3UsiXv/IfegAneXJ/yU2Rpj4P9iaLKgmtjQ==


`protect key_keyowner = "ATRENTA", key_keyname= "ATR-SG-2015-RSA-3", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
kAlIhoAHksCGo5mF85FXcP0dM1NExLuDn6ZkyfgoWH09b5qcw8bLJnQMlkLvdLRrczznUPKBLrRR
nUHSMi9UTzRZ0rrnazgGnHFEV1vyoRgDQDOpkZbrkgl/VynbkoMBhCQXYT59yyHhqjI6WeIYVipR
zyn+NdmUB+/GwlsSYygywX31rotvUxb4RZmCqg+UCemw+N0tS43QuIzJuG1JM+3+SVbU3LuVcClf
rOwWqAFHsOXBSrXNoPX6QeNlYUKy8gcjiaQqPSrbrSJWdgvqshdNnvLWuzkREOLY43TCoAFwM8p5
73h2VUHmwffIqzCELbp3Tee5sQXgMbvJ+Mbfpg==


`protect key_keyowner = "Xilinx", key_keyname= "xilinx_2016_05", key_method = "rsa"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 256)
`protect key_block
CFQ8408huN9E8h2/r246qkePkogHtf4rd5gf8GO4NiUzetOQ2my8cbvxYBjZy3yQSw0/LrN95Drj
cc3uAe9r+wOvBQ3aM7AKnKpRkAvmqyCRt8lkW5NRi37udLv8jQJ5gVByTJ76KIn8s2kfj/iHou8+
VyK641fcvp2Fk/dmC13HALsHzGvO1m9Kg3zHT1aJxtdh2FDGLhOy/TtcAEbSWUhNkclp4pw4r97T
urhhIiarPZZDEkAXG1Ezi9I9ebmvdHMRRa/e9P95Xg7vwS04EHfmVTpFKF7UHncoI46I8za8vjyZ
8MCKLS5zKbgCU1OCJ9lQ6mJX1roD79pJrnKYpw==


`protect data_method = "AES128-CBC"
`protect encoding = (enctype = "BASE64", line_length = 76, bytes = 967856)
`protect data_block
Yb3XkfnvUyyxyVBZ77rD0yReO5JqXnmydY8NMySp3QKRk6SUaUVVSDV7cCUuEJ8RH6x0DT+MeiqV
z6EKaymVN7nRr4VAeH3DiFis5QnvaXV13FL4cyDBPy0sWq/W15Y6WbCdo/uwLGKHPFbNvruOQo7Y
4V/7YTiWceGVi3V64hzDmLCTvFdQM687Rjq7vtS7gFrn0w8qNH/DxECxf0ZJAGgM4ju5gF4g5wFF
CkFY2kR+IvzxSx61sd6Lv4xXPw3VpQ+zMVQe2aW3RWh2xl4rvGcRcMYBt9z1k1L0r+O+mFuF7871
ooENwTw1EWmZnTXOBqDRhzDlF8nbptBUpgdv0YsWu0sAAj/D8GaMqTvoxeV52qDXA1zjldLisNbL
EcV1iOum+t1MpZXTOL0UHPm0oFXbZVoWvhdrkIfcMruSdZMbiV4syN9IxoNolkyYvWgzGSXG7Y0O
U12DIMTsJwzUX24Y6shFQXwaDX+YIoaBE2WIlAE/kgVo4ojdxIrcv/e4hUM4sYQryHPGy47gfFAK
NsW1HbXuE6ZMsbep5NpS7mCb6a5dyyuDQldTQ7cRTBTOnvBL8UDk/eiVXKp6W+0JJygOyUG/KmSB
YheFZaDNlNz2CkYr7I8PAGFNw7DV0iTk/zSROLzQN/GEQcWNaBfzFeh3Ymmi2uPGFoEP+YXQzulB
uYL7dN/XFxig+ZXMx4mYkWsKAFE1z/1M8ODXdzT3R0J/qFfXaYu4Q1Eq4YYVk7aKvyLWZcem7NDe
TFeU7oWd1OnBOKupk+nc9DuLYWu0xutVzYD0vNWTZaFvaNyIdRThIqpIeNT+1YLlOu45Qp1JMgZh
YlaohqlTLTP5jDynZXUjJwRnYH7dOq/WyfhW3XaDaBjtbjbT2wnnzTJoslp6XOrM1EsyckeoVy5Y
GO334ZSok5gn4qi6yaUQV/VoVv20DWCUcz3sABsdy0j8a+8pUJBzhuBPv1TqpNXJFaXsbgc9DHvn
lVp3vcMNjTHqCQimqP9n9SaMHWpxFKh+Uf6RGf0vHd7OwL+8n2A6zFxbWxLVoJ+SMiAUMubKBrwr
tNwqztkFmrPmWbYATODBQL1OOl/2qlZsF6ZqKeTxtOaEVavO/BQ4BjJloTNGFirug90FBaJKdm1C
0YN0Yk+08YgiXitMR51UHE5XFV/j+L6Xw78Cpv+RqemwuiFv9U3p27Kt+/LLqHNrSI7K4ztgeBkM
0xdiXL6wVgweswQCotyJdGUxuAATMD/1DoaDuRiORgOyJ/jxnOPZnnSDMxvd95l0HqvF5wSt/j/+
4+Dad2OkDVM+acZrkvxf0tfvIKzikyZYcFozzkxUgkCSohR9TY3J7p6cqkGxkwRj4BnQtxyAJrKm
hKizb5UIffV7woSBCtN9ZnfOFtz1QcWLsRVGGmc/hvrB9OuTsh+ABXgRpkAhiGV6oKYVg0B8QM/4
k3xm9UtU/givN0i7Ek4VHFe1dMyqhPd+6eOzOGNWzWp+758pKaXtPEWkuEeX/Ec2sUWhI1iSeyxQ
cGclfhZocJIgiGWvcDI5i8DMnWKjOGAG4kihyD066A52wQaWL9X34bSKIS8iL7VQ1g4RcW5KBX8I
zbibIUpD0Hem982RkOVGC9nhcyUmVzOyRn2JjldNhYwJDZkM3zwl2L1Z3WJsBFfWOZp9Isu1Y7jU
6HyAytmDIz82s2pdag5gzeR94ZoglPGl3L99KzKiuQXul7nBpjLrI5mLgKzyt1uSdHFrnGLdFYHX
Wdn/88uI/YTnmVTiFAwiNshrNlqXUG25b6bVDNMiD+vgmZv4sxY9zN4TNPwaywlEnkTziFK2Tbpt
rexrYOPJqY1WlfKBMvsriZ/Aba0KDuTjO4CRdPON+LRmbGPkapgIQIlIh1tVN/6C1ccmHtc/lEw3
qJi/bdCtO2KmtEGJVKm48ZU5Yrkl+rtNsNGZD2NzG+DIgM/BPs/2oPkFsv9qBY5DqfMJK56p9D1u
PNaNwKMWllOgTHlRy0rmLFdskMemXYyC1SpfL2NosJy83JOIvPD1wXtlOen8z6lCBJa+XDjwKy9l
pcJrxpEbXlm60PJE5uWCrmgRDDMUdIv1kwGZRxLsClRFFkZhUrmAntFgbZqu2Dtze7f+VwrCUoQF
wuU+D9m0OSSQekoGfXK4A+euUkcU8pbgjw+HT/CPlB8F8B413CbfKckHACFGBrfsn2hEGC61ZM0i
icZ8QmTwYS4M+hquvUpVnZotSmFiBOlwJIpJtR7VXXc9mWJayV/McJCuZ+/HQcHFP4f1x8ky+i54
FSZ35Rm7ReWdsm+LYUhJUjXFJk4XTbzf8BeGCktHbJyxr+4p+CECjUefSLL+1bYt55bnypm6pPVd
nNcRkM8NRXBVMr4RN4cC+Hom/QbMqNUbZYp5h5GSfqrDLGAbIMfR4HZwWHW/yk3idutwEcLJSI3k
OR0FCJjHjoQUOpcX0MUrNKj3BlSY9Zn7AQBjoqZvFDX4mY/0XMNM0o7gsH+JJRaEAQKW9bLPfaUi
IFKbvsn1U4C6DADGKMQq0KeaPiTUKqpWsQCEhU8eqZ1hcRuwg6hMzP9QqGkifvccm+f/rVW63eaX
cH2ENvXeCllXc7+AHPNBLmXz+OeLyQu48xgfBj0lz1o08Zb6lahGws0RKJDGyjQuqrTmm5Oe0i5E
x28OveTF2xtHwaNsz7J+8YVde8f1qv+w1mI0QnNxtrr9z5lVWNZu8V6pbslz8MnwylUMWkHLOhvo
9rVbessOZihf16gEhetFvE7oRHgSoX7JYLsnWYxsIHiDD3r5aYzGSGe8050fDNxsje4BeMFVC48E
uPH/AtI+WswHrOcrCmjnRDQ3p6Wvbn+axkY7uSKOzWgt++VOAx5VcgsUbX2IF4jboMqrbnQcfLdx
0mHFxfP6uVrKv1GNiAsBaLNX3yv1z4GP/Iu4Cxq5jQn9v5N5O5IhNh2lmxHL2UG21L6MfltPKDzm
vnXR81Hrd/0HICkP33aaBosTp6D/mz8shaMyLxYpd4aaAHcFbK0bDaiwPaDMJEyDmc7yz3KXSTa+
xsW4LEjU4VsHZa/iMp1RV9ObT0zYu04mB14zl1O1CBsN/yMC0ubbAfVoSHkw8vFLfeVDGZvNaZkK
tdM7bZbf3fcc4Cjkd6Pf8+Zxd5xXPA9+97X918fwYirVt14E1DvbHtQulzJ8FRx84T3mIUGnt96D
uGElzi9zmwJGdYGtBvYXRwQd1+56z5RTCocj25KZE/XdtmcrrLTlPKSua/Iyo43BXFH16J6MrOR/
2BdyVkujO3kLw+ZMOlPvIVK4/Cdt0oszoXNJK20EbyQFvieDIB+XiViHLrutpvOGsPc4RP6vdwbh
VRUQBu1B6elcewYO9GFZ1ISbKp0vrYRGK4hTU2tJT9FfX2c4+h3TZx4jmnM3EkweFgEJnYMQEPUw
d5QWtQmYIBYDbGVWPcOfv06wuwnMC/rGBAgi6s+2yEIyk4Q2CSIabtsfjIYRQyqrSBX/X8gWfGit
T1mmDR79G91dTYEfZFrGMpARHhuxzRvY/Tysc6UnxndfpeyTcu/QAYIuyw/R9tvzlqUCTFgFTnxE
lmriTCAs6KWTEopVH4408iFREQ6KESf3jLb1mV7ub0QEOSMa4yrhUzAeWK76OUEcnXkOhS3JjEPp
V591N3U4mkYS8YBjS/QO2m2zT1SkY0c4kX7nU1dH7pArVLAEotvagz4slYGrXRwxL5BAT4I8ZgH1
A1WvA1vqEWPOL6qyA8e0gWf9QX08rM97BNr6tfkK26xmf/diIGhT0N68nRer5ZbBydoegFHWA+af
ODjQtPD2mGrTYTAidbWkvmOUtee4TiyJHIwkFrhrOKxmUZ2gbJ6QRoEpNhWsGHZ3BsApiCnqmI7n
qj5UsQDYsATOsmV0f45FUhSP6DPcH8ZqXW09xZIi0SVEol1YIhG0vCOZD8ifzR429vSXMeGJV+mg
2QBDW59WuxPT4un+TYR8i6S3RVckcZSUNNvXcexiuxXGOft3p+8zQ5NZpE7urMenoyGTHs2S210q
CetEiuJaQ7sxmLNbaddv+Btj5ui76Bzh85aC3CSDAKcLf2Pi/tuJdTdF/dzl1auu2MCmX4DLNHb4
+sL30mX0j7ciawizBVjhyjnOdn6gQsCse+0tpQIbVlbI9RQ8cS8BDDA9KJ1G+JhrspNb2KKGBJMR
7RIppThde73govJwYnj51W/AjH3ogVimNyhQOzEvNei6RU/0w1Xi2fENWdhKSAEJ0PhOhEo+0+HM
Ka4bxa+6NjXCLssIqLwyWsNJBD9cCH9Wfhk9WgwHshpwl0pLE7O0S7GpdbY5WJSyZ5wWg1mVIrwi
6pGTM7aTaKANHhQm7o2HsgugVJWwCGZdxuPuAk3lkWRS+rDIQNQC0IwebcXNs3lFk7M3t3AjavHM
ubUQTQDDQC3EN1tRwDNLQfiv45KkQ2CP8tC4jFTkL7KXRwqfZ+eC9ICHjs9JeO5+8fHxAEUoOsIV
hPGrEQfZrV676CpAW8vjwLj0wZjd5cgiq/V1MbeJ+84QzJZOEk2RErUAMcWOqu89BEbCibaOAjYm
3LXVugGNBMl56dvYsYUngWJ4kSw0+WV7i8ivLtUwqbt4nd5bnOF5hm2wu2SYAGt9zmunUVxYAVal
kUSXUjFlidXzMXCjA2GneLblmFQD13ROehHbPUubs1i7hELmWrhuplMLO/6tl0olLtsjClwQQD/W
0zmRxpd+zj2BAqIKythzEf1mIF3bb8B0DmQYhdYREus0Qxp4PBfAcijITvyeSFdlkqVT7BjJEJNL
Xl618+EwlDL6z5z2X4sjBgL806rMQfedyIjsctXb7mOyR+1yuXjjiUOkli0I4lPfkpD16gEp1ptp
PLyXK2CY87atCLx+WCeviyuJ21RpRh8Htx1W93c0E3PQ8WX30xvil1cQTWeawZuSuyUi8iLCG2KS
Opqnd0p/wnJi7Y0fAtWVdVhnchxGHin/EKdNXe6nOyVHM6bkOm85moLtSTAgPmoOUEzQWpxQE00V
sxuP6eu5QBnwOD3DDIjxst9Gs5BVjgX5OJBdulXdG8BUDwMDWhEAH/Z7s1KdoWh0cY1IEv/MzBFp
HGoASBSx46E4L4Mr7Sz+WXO+9X0b7dT1awphaG8JkoWld+EXrAMO1E2KdQpN3WvkN/NUnBaxkzAU
HPrgl6DT69PbDdTDgnGmXW7pibNpNX+rZzY/bx7xfcciWBq3zzVpxLyT2b5vfh7eaSC4Vz/DVzqy
KTUDuxsCXw/IgTdZb5M7irkH+Pl8b8kFtLW9V1NlFTRtWIs+ssw7KAIXt0LMJ6blYqUqqr7aswAS
t/7fD2bAvWFMSUCLLq8axSV4ySVcr7tXnKPSklKNxsfh2FMADnfBweRoopoE1SATmOCEPwqxc6ej
RmUhW3ca3VCA9MeWDNJP9rEuMKxA1UZkRECv3S/zrPWR5LVvpssNuHIYExLBDaukHOIH1SDRYh6q
8RF7jWKe0xailcrNTKnkdhFAXX1b/DABGmI769zVLuv2bmc+q1WrmZzu93UtuRfL0C9Mdl2nLUgZ
a79JgCa0923xCgW+0UFo26MRIhv4qob5i3XbJiHWeOacO0OSHO85ul/WsDEZk0tx87cbPONFm+Ul
09Imw7ygeoaWG3V1zlS3AzYQu7HPrI4ufN4xTU59e1XZU8iqrF9VdE33D7H1MsXba3Y8RYeoUO/a
kiEcRK2cahl1B01spLevmNJl2O4PKeekozLMiucwMmclZuFGi0/6CvfZaYvw4DvGPuezqEhpAopL
6a/6v/KK7N5AxW7VUDDzixMYHwpye4aQFOHS+fimlh+NzvWgzllzDT4iy74PfovtyhzXVSPcuDgt
jPPVOR14pRfLRc0fOxJ24zFWtuaR8Qmogyk0GMX++UDSizyAE+wROb61mHv8gVvQdL0MhHCHzTgZ
p6f6Ei0rM0qEG9YSBKORnl30jTAKo/SvducbPpdw7GLr+xfJ4WM/kIR/R1Krz723FzuOGUMibmZv
Irkd57jufPHEEpH7R9iN4ESxG+7AJd1IPvt+ZpKTVdQJycTk++hwr3OcEpakGKhti4clxAk4/Pxs
gi2tD1j86Nbo/MgeUh+P+i/0CkZitM+JFPNU+bbFLZIHyIveHg72xqS1rrNlAvkTFttepNsNBx17
fEf6+fiztXBOg5QT0VytU/njzMpPX5kVjl2SEA9693Or+1ky8l81PwsufR9Ev/i5Dfs5amhVvmmT
Et9MPuBCzOdVaxervSFungkN7fjwnTIGK1HAFnfK8exO82ymIwy6sQKItpcJJMjUmrk3OUKNb6Ws
WTbvDBYLqA19GZQT//NVSOhaPelRSFsjPmwJ5HnmSY22qmUyZkqMs9E817JIa4oO/VZlJj5wJ0f2
GdKTPL8F5UTvB7vx+yuowco2DpWzUxKPmQEhrJhQdyaM75RSG4l+qVNvgGMdvuTNW64Oy0DLxnn8
P6irL7Nro9h+R9aP1c4nwPW/khKgjtGz6xRbWq19fSrdMB0+Keg4tpCg9mO69aM/23tl3j0sQrBD
M0pjkQm+N0efFhQILJWfGcjjp/CSMw79okgnc9InOTFiAzTIXKmiP+1q/QiSsVQhf64rP+OA9Fz0
RlmOsYQW+VbtZXb8yOVtQuCJjozY7ZrPMQNl28xOFOn06acqliLHbC9+CxAV2oM3L5LUYHTkEEAe
CrNLWbcMgKGVejS1GbqY5Ll8WWxMLrKTIMLQetT1Rh5MwxYp9SvhtXNILpBCMaAs7z6AUeNXaY71
LxjL0kcTxp7yJklwZJ+SsFtbVUjPwT/QVvg4urjF/A+H1goJ81hmoNlrJ+PkNAw8kBQfPVvwjxKU
MHjETS/UAPdx2/nmcTWKzy7m6uzaie8eNcgGT+Idyq3eemqzPIUxb22d7MzJ0uJD6YwYkqTlOhxC
auEq4bFHmRDxdB2NvYZf+aJfCJEPjU6keAHfdyhu5WBHlYj+PGUNxG7SMksiMWIAPuHrJQAp3Lvx
IieLH6zdxgBrbyWGNPOul2PVaO8CHSqrwOPaJMXn7ZdB5M4X+HpoIpMbtzCLGF04BLazkJ1FQDID
9hL2T6BItuKB1RUdWxCAW7+sCqH4FligoqdYAo9F/eNLPvZUwHmhaMb1jExabHZi6/eC85k1BUXo
3bc71qeOHZvST3gl/uRe9n5ybOkzUqqyJ0fAIWCU4CxFK5phg51ANRkWKv369ze6PfVetR/4E5Y6
GXg4uJhyI0tldeWZT7PIIK7FCFaEJaQy1p1/Ci78wmyuVLp6dZTxKyKyYw6jLoEJIkZjRXRV0dti
GglwbL7ZXBKPwOT+PwxxGWmjjL5V1lM0YKl1S7j30BSrS+ZhlmiSUy0BSSpx3vpLOu9xO8BDa/kX
JDE+RVD115Cn/HTKauPADCoV4qLxJEt+Bj2z4H8hNETm8vZ4hbh28LyK/slRBj7jwBH2Dly08K0I
0eujL02lAUqf/Rs6eCKI8S2iw6/uQbZGXiSzZ1DckwnGdbTkl+PuhecjCU0Bgk2Gh/Dq5AX8LriF
zOKp3wHrJ0la8ZIvaUhfOex0XmYvK2JCJfHyHdmXJ4QCun5k1f6R4UncJO6xB5GwK2SWC12T7oPz
j/FFkAqWHhUvq6+WXBHZZy7o1y3SABB7nY+DEJJuRhjSQJ2fDT1lJcjZPNsUMHUqmnSgJo0hot5s
GTwUkRSSoBf5nwLHrtgSuqdYeTVpP4kUaAnsYjmfoUDf1ej2Tw5k0E7Bcl1Yb8kIM17Q8XeVZg1U
9nJfmTaSNrbOMMiknCDetCNpWXxRKUrw/0J2/IVDv4oypjM7+oMCoGLGAG0PVuQ2IP1C3iUuN+q7
BeeQQcYzszp1K2Ngx5ecVNotGYCjzgRBUlCeGA8ZQzgdgUFHR6ro8lf/CYHpqbcj6cvUpgQrazFs
v/Bv98ZySi44K6+fyHBgvk5EPU/j7V9/zsW1fjOfOcQptWPmPeEngqWRRW/Bf26srSH4uEhcFMZl
E6F6WFqreRcSVCn62TS0Rgzt2wXWhVI7lyTSD7X+57yKDyzLYuI/28zDJTd36C4K7P5IZn0DS26i
sM1qq2kNmqRWOFhblC5peAEQHwt8GDOBaFxAZ3uKS9GZGdLhT+S92AWAoIR0AcbjhRlWvFXxt8dG
mj7344WlkWSJaslM/R/U1BxwiEQs9Eirj98v6+qXLwR/lp77hk+s1ool336NT72lnXTdSyzF8TFn
znuzwsFSY1FvGIGTL6hY/+e8xKm+o2sYq8He7B8aUp4nDtRNlu/rkRS+ZSUINDhbTyMNuJpUzmvj
KVYL2WR+7NLy5LxMzhKr3WPsgEK/M99dUNC+3urNZMd1wML9xmvyXbj1jVvtgA5b6Q+TCySk9XB6
0KyOaCQ/U1BfoTqSeeL7tarJLTqu0VxsaKg9NlgBwAvU2yUNYC3uGhN4WgFE02vqxfaT4mFwa+CK
NnlG4waCalplTfkFIbKuz32SObADJZkrjJ98VpP+CMuNiTkOQCJKZ2OEe1SIjdxZJ/GWhXP8a9Ft
cp+S716hVUYZSN7Sp0akTneSJ5BiOtFTaoKx9Mv/cChVv42aLFZ9EDKrdNxhrS0lnlIgunRD4jXe
K7fQaiVL9MsCI0V9UoXBYiokgkNw8ba9XlbZkfAu3YWZwscdPPyC8FRWnSyUac6rbrFou5Wp77cw
w3Nb2asX5GyUGsO/SAPWN4YSci8v6izg7HSv3zgy+MQCaWZwHCFxwvyiKe2EjThfFUULoo8OaZ88
9I5V0n3RDy3Ya+J/rs3rRawAoiakl/F4VxKWXDgjjFFYgfUAh+UHSFsctAN6NzcOkEDAsVr4tW8Z
HjYCMurvvoN8TF6s3QOtU9e/Bp+n+agGmpPcx3xtmtEk0pdtRYsB5Iehre7OT2dz68ShP+5yXBAF
J9UB7cbp30WZO7wAIJny9Cs35XI9vV9tVhXLFfCpMJvFRNhjk+uFKaRYe/y1O5ajf4VQJGcwXAxO
BmLhyvY5i3xtDJ4PqcX7q1eYCUCKpoMUCG6cR2Jpi+6Q4lsebHCUBTA/h/1Z6bqbRtgUxvtS2L4P
x1GifIDJYCk1O0qQCvdZO0+j+W/arynNLNiomviwNcbv4RpOoiM8oMcOoQWegb4i5NtLFkn1WicF
gMuVkUXvPG7TUvgzsBbMtd8VTYgqhMXWarWcDgubRMWESS9Gm0efp7bvrckVPqQBdaqmHYQ2np8l
AB6bRmfmNisIXOpwtR99yA66nlBdokDpcMPJNMi1Usv9axST2y5GU3cW46YdfkSrYdiqLlZWV3/E
4v11kZKxGD8E8PtVoRAVhx6By8BHLJM91QdZlOwGsMqTB3R/bTuc4WeQN52RGbOsSUUIhXBHO1du
De9eZAfYQfyAxQGUSbt4QCh+Kc4k2rJpJVl4qrcq1WcSgaW+lG+nfMJ8FVeFLyldEet2Q8uI0UXr
9F8jDdHtX0T/qHXkfZ00N1U5oQZHPrsXex2riajJ9sDvT8XCq9M0OaBqM3MlexV/lHZ9dsXeaIX6
Y3tQZBXZ2snvwgM5goahtXvhEYG9eRjLscI3UpBudpXHph1ncGO3Ak5fOvmASGeG7cbOCMQAjJTI
hTOPy60Tj3muMRkUCwqhxNeft5877SVPbR1Y9BsZ1hs2hSe1za5jZrW8G4PK2jMp2xMwqNd6GPW1
WhfAwTrq4AVOW7MLNyXnYbGXpM4b3Oq8spE8HSdOptkpQA6hjp5vd4sR44c5Xe1gGjuBryIy9Hr8
3djeLFV9AUp3HeOX0xphWDW25oiwu0kSf9uu6ISGXRofoIE6WBAPDevEdelhIA9zA1+m66N67pyJ
SHLnFntWbGaSHHXPdWAjp9HCYkDDnSjLxeokU1qBBYRlP4J42Zj1VBUJsiwzUYRiTdLV7b5QHaYr
zMxUAAJp2LBFvl2LmGn4JkDQMhi12cSyjxNf6z3cPpNmxdV8SBx8zal0SYdbJf89O7H5cb20nxq+
KlWJN0UQhhwQZBepPm6PZDC0hbc0AIeUOs70Kp/tuZixkaXlPk6fKZHqzjpfptFUZw5u3kRQ5Hv3
ja9P1W/8V/8KrFQGRo3+NsoHcZreM09iSo3mi4uDYLjgXHEQAUzW+4ScVd1Xw8EAnvIB98KUi1+H
Gd0eG9YeoHOrzvlicsFKihJxEk3vbDNG1Pr0UZHKeu0AevVhTAjYstp/09uNdfNwBPpHd90PbpUg
b7AcZQpx3KpXxNn9B9xZpPgfE+l8EjH6iG8QB0vnQeiYx5WqcMxERCg3excZEbWO+1DWYGe/I3gc
gYrKosdSfauVxBVBCx3Ev8sfr6690NrVDP8lFSL0ZO2C3x6RTV+Ci+oAoje3uGwnhsYpb9Eq4X1D
KAoyEmWRqry6zWEYEttY05HkVjk9VutVh+gSDeHVLNs3DupJFD2m86C6hOZ4jhhlRKE3pu/spv9V
cDkARLHngIv3WxkpotBtU2QRR3bCJac+FJ4HHBrgwI0ZXkb8kaxXxWk58zeZbQXfMy/EfrnSelca
+cL7Qf7YKcKPuKbuUD6MUsjNGUMAHlcUtOqIQc7prQCfDrPfYBUB/+oUvdH4WbEnMuCHNV+lI2an
RTPKxreul0GTcWO7slrFXHzQdcaWB/DoEYWQEfnp5qf/M3E7GKkaT9owBjd4/OQkYZyRQB3txGNa
inAof8mlRN2aiSQRyERfOYSVEQIVBr81Nz49vt7uZYs/zF5gfiIQ5ZmbdRuFzeD/ZYW/BDot4AZ9
OqaaUhksGOhXMcz5bLxkkzVUloAcLCVYBP/eGwxmnXxcI7m+huaZOb+Fl/Ft7zwNtEwqjL3/SBWz
yQ4gu0gVpNpsnhAMTdKq0VeGpLpzeZGUcjwPWQlwoo5rAg28ZGY4DXjJ6VH2OmdaIQZ9LJmS3WPD
Kdcb+WAh8BMkNYwrYYsW6jKldkk7fyPJ4iDt60b5ZTSlqxAWRbNDzXFh7Ox5YQ7YXlatnwNGN8d7
LrGG4dEWbV/2QAl6Csl7PWN6N5Gt5PbHPU054lF/GIJtPi5L1+UPvFcrMdMAY1e8VCQJLZ0s79uR
0BlMlAC+kaTEsNmbKk106EuT/9yb2clfntFZVPvhBupxMSeZDh1hJ0TBaXjiwQgoFFHzGeVuCr69
I2MpPwTAuTV414i1vznTGDA5JoumCe2y9BUOuGkjfAW0pJPgfVN2hsexsBNI0M1oiru6k3lD2awu
UYie5i5FMDvVIPX3s9XrDJVNeZzoP+aLLpRA7nSx4QqFsAX2GwEiY8JHyi4qi2Xzm4zlLQ1Kveki
YK+1Eqw/VJoB/5/3ViKw4qn6BPxgp5YFmWns8DXGm2qckpRai5HDkPWL0gcfQr3e1hZNUbLacFbZ
LbDx1EqVgPYKnWRXjAGvGeKoDXD4ufL8RtvmfSGtwENd6Qi9sXjK1Pt5tkGUZFj+geTpTKn5Ym1c
GcCCiQeDNTCZrvEQsemZ4clIwh5wDxYjRxdiyx6rXEvKT9FkoLZmZ8hzVh/P+jwuA2zlA9PZFxfc
gfcgPW9ami9oeXkfsCzU05By/ZKQcJICTjeqND9htGFub0RwUkdyktNZR4BpHiwu5iSMa6mE/z2i
wj+9oIVffNSN+9VxqdXAwLHypaOuZyiI+2qzDkeGpr1n2rwo5kY/avW/oRGI1yadQJC5R6xrY6HS
/oN3hXcknm08Qj8CMS7DLUARkNMi0d4C53W1AX7Tc4DlWPqKHi6MWmzn/qijfg6Yq1LGVEuNpWmZ
Mu65geZA5KCGRze+YNQoVp8lgHuA6pbD0DBcC9ejqWapAwHmy1R1Krg/3EWGzCuqD5vvqZh01qR6
rgV1uxvkDvGmM977bj3IFBNYt/fuoCFrwNkx8QoIEAKo9hYtaUPHJxi5soT1JDkvay6+mhBqVly4
RvyPJjoslCKBqz0QoyYoXfiQNzNQ8MTIxWApy1UQ1Vsvxve8ODbEYQS/WHIT8Y6IuAK9TJ9NthM7
qCar6+YDs3NcjuAWBZ6EOESx65kl1JPzAMXe1Cx7wVDykGcsbdVEu56F4pslW/wT6VNk8rBnKUWV
TM+/zVH7wV2Ss2GXxcaWfjUqaWt8u8Gi9v1Ij0RsOcdK++CcHfrFvyF3z3CzrvlM578nyuhZvzUt
6yL71vts3p7qKFhmGm9sPdvZRR4r2fRUSaWLPmVCB3CwHpwQDJ/u6hc7QNcMyjWqYohyxiip4sSo
MhpmW3pAgtWuvQKlMQ8S9qVP3RzwhGhcB3V5EQlr5L4Dc/bDoO/eObtuGn0kna56x4RVcdxxWRf6
neggIzR8O9V61BImTBVglse3KKLanwE+Nkbojcb6xnSbREm/SFxRtsXBxj9zGEDAWagIm68jwV6L
ZLaIgQeKZNquZ4W1Z/WHuZdZzhCq++ZxpRnOnjdGfwEvfDj2/z5Pcek6hW1y6h/R3gNU6qeBq2EP
WKWvywCkmljK6NCCKWJYGxV0mzPUZur99VIIBs+Z0QiFBheCTr/j6VS9H8lpoVMAPfAb2tXC95jJ
lUbMSkZKe4ZtLZ+W9T79P4lMYz6lV3S9RYQdB65rh99DdUuy0pFW29B5fRwk/tZj2GNTRQZHOLyv
g5Hfyrlrr7v90bF8U36se9FwDzlBkj+VRTgtm/wNIu0LsiJG4Y2188YHWvC2YPTCge70VbEETF+N
QoFKTcU18VjRvIFY0RCLtKViJgJvovQmAjxSXTi0pdMpudaxiR1LVj+JSAeOrR2dGRqdZOUHVjMI
oXz5D7P/tWVE+iaXv3oOMa01kwJQiV6Ir4s80H4YdUhKhTtxguRoESLBAT5KS1STFNMhRTa0a+hg
zP/KRk0WXrR7jLMj8IQeRJWPmI9Ox62uemR7rE2ZjA9zr4Dv9UnSmYQ2rKCoHOOGz6GsF1jvYsXy
dUYnXrzLW+8tpXq35IzZH0GTrvKvh3qKekYzhGrms3/pz0vcDL+4CeMIe0H4O51eZejtzmXUeizs
orXGOp5Qo8EXwPzXvMrr3bo06qsuWDjY4OjiPy3sYCr/0aCjxReAGg9c74Fd6CzQ+s8B1j+RzJOV
4IbkXjwNn4/lvc0n1adX0VT7PZibUFGMZch/EXNwXoUTyEwu9tCqmVRqrrj1A8WLaDhQ+c26Hv8r
fu5F9fwlUk2OZ79eYgP5/3wy0eVK1s8sDDgLDeTdBVOy8gHpReC7tI+ZI5rZY6UsSQD7ND0pIkQv
XpaQ5Ssa/6c8nI1OGqiVFle4vlY0OUDQTVjzqqY6nUhgAUBcZIC6YoljGNiC4NgujHpVB6TuAvAP
8aI6VsfGW6k8R8cQDu6Kwn5yjW03aCP32MwJ8ZljaVc+vU/Jdrk7dOj5BIoluQeie9pvOHr0Z0WH
kSWthbSN93hkcsNZD9PCWDdgTfl8cueDROQYu68ZXYNNlG1kjkz4qQZT0Bs5CxcOVirevb5e2ml5
HvaCKP8k3OnxVhuBgfBJwUA1GMkkIdL+grmxtPvncsk6iJSl8kfjmXeMNDqpdZbJhGhIEzoiB/D4
TlF4R8JPonPLNWz12foEC9eMGbVmSWAnh7XkExeTdNsQibOzp2MAVGiJPZXIQkj8WpkALVUT25DX
Cqmtnj3AhagI+o6TIzgIKHkHv0zCOXiMPe+T2MkMYrFUACj8NEma1eOU33B7sTQwhESA20s3ocEC
CIMp1CzUE14gFGzVH6MWRx3CiOhom8z711zCsB3X7iGJq0i7gKLWs+9aEzB+FXlqLEuW6ZHsfse6
I3gq0NdVosv1fhmfW3D8J/9m3qIfST/CQTcY6POQpLkfQC9v2bb2vXi6/6tNnzQfCQzynSEpEW9a
L298lwOIZHxeuLwc+TehCz0uGm/eGGWsYmSjYPpK+zouaYxTtWj8ispFektxEsC2vD8/QMuzR7sV
vPjc3qL4GikPO9vNT4Qw7bY8iuHiYzbdZmfnhe0rm6v8d8Xz8Y8sIg/IL9cWzqOGUFpo774QYfRx
FXEKUnRU4PT2Req4x2E+MtKH9rbyn37da5zIkJ/kLr2Ab6zYGo/u4dDmo+iNpHGbMM8omczhdj2p
09WN7GN5b/TmNuZKKhcOvLCeNUWcLt8cNvLxNoHqjLbcn9TRitcHXxZJJtX1Lt14PNJ4x6Ql45Vv
QBwvNqaS/34iJqF+0cXauFMt7dX4yIaWCUy/dDzRZ82bZiJTvk1+D1SEohEk+V+EAUP+Fv0F587E
Bozf/DfYMJ/0KC3r2OPxcE9uduwouKD3+2vEEZjPoDzjhcvlz6o1ugjETGj9GKKFSPJJrxETXtU1
J+FhplMT8M/UqSG6oa8IYT0FYf9KkPeGKjGH1yuceXBN08HPzcTWchRfWbLW06QZr4q2XJZJgOVV
I+QBqz/B56Q87GV0cFtgkXj11POC2mEKr7O6N/cwtzRlLmtsuMw7xhMsN0NJhrxp+jSxnGfpf2va
S9cZy+cxGo81BPCdO9niI1v/G8qOpaqw658jG+AHFnNVC0013p6res1YNlBVD6pp+tq4LIpFXNfK
B5oe6lp+7IE/tQJWm/xV542vMzu7URRyuK4fWEQoHJ3N20j2rhRwz/8SiBNlZER5i+XeOY10RTAE
z2krgU/W44TaxGyd+wygLC2Qffx7RpkMUvAfzFtI4yfeJ3UGvHkQ7UXefdp+fBfG0KqkP3tW2w7E
0Uiyx2k2h/8+JNqYYN0i/UkXMzw5AA89U7D77lxzpNTpqJ3Lg2mHSgQbcpiedPLCFWDllQOa4d0a
YTr5sIY84k3L8elu0fy2Z3tkOd8xrIwEj1DQhkhZJX+1cTphYmYvcbdwcAWDv81E1Oqai6V0L7Rx
mhulfDImmNrpl7A9dc+xwrwKqXOAVhCnPigbgC1reJBZbPKsslvhNZFBKR05EMSJrKBnDwus3pOR
wU/N3BtuwJRoyElUGx2r26+bGVNvCOA0ErAMwjmG0apQrXZYP4WfsMBD4yYi8RwRbtwueaD2yq92
4X7hutAAoBdm1ZL6bMkULrZiDEUDwOCwCxuwA3F+MJKHM9mlwI3lupkrKh2Zi4mem42QCShKO04E
07Z0ltNpI2Axhr4cHNmKwGUJ7MYdZEuHTpGgqZuCZU/yIdP6R7Sx75iVkUo3nCfBm3ovipKo4dSr
WukB+8rLQguKQClcg1qZJKbGBu2KSdH1blQBQDgyRdc8tTdR5sqF0SpXXTqIn/gv8tuXXxtey6Z1
eRsR0T3KT4MdyKPvJfYSIEH1JGpAfJLTdlB1PdozZm4/JH2+UholXgjYAK2WTJR+6b+qA9JHmXZQ
ch96baJGjDfM1F0no/Tspz4FIUvziEKKJMpHfMXHe7ytMHDy+DSpKbRV7pvjgB21tSrniisHZCIK
7xWau+mnfOsR4yB6p6BnSnF3+cGKZ+CkwIVVDEmawz5aumD8NASl1ia9F2hYSkCaG2LLzuJ388Hd
K+hu5GSCks6qEGdKq7+q/DsK9Mst6tqWK3QM9n1YYlMu035jCtrxBtYUbczUIwAQmIW4J+QgdzHR
7CknrThEYbvGuBcFakTMv4V0+O7qLq4K51kKnZ8eZfmEHUcblxxTwxYo7wDQ11NET2KHBtQPOWb+
m59i8wKuaGyCAERXSPG27pdyROhl0YLUg9a+E4teXIyf0q/wZpOzCf9CIf92o3zAyJnJmNbOL3lg
LM5L4im7EtH1uUM5M7x2zLx2+nV4NqM5z3W517V0rqpYt/+KQULyIPRMSioRepA8LplJZSmOJ+rZ
ITCvg4R78l7d9+v8x7KW2lg8KlE9MkchU4A4vY7Vmh6Y95Xf1mSfe/TnoEGkC7jszdAx1Ay821Qb
ImQmlGYjzpCIhmtZoxyRQ03/+j2qyHg+1XbfH69ORg0JEeCs6lE0o3VU54NOL9x3ExyBRKjkc0rT
v6rNiC59wZJaOa9jZ+Q3hnO4Kf7cn3eA9NG12s5TOZI0DMwpz2G97JA1EIMjyjE5QE9h2v8Ipxyp
WU4AhQFjttv3ZGdz2eqBcFN+ohMj6BbOi/P6+5tpTrVEouy4RE72M96lPWq3Xo57M/fwGVBQcvG2
q2JMoqhP0nHu3ryhaPBseOR3QMw8t9OIESCjTg0twXl/0wZFf42OLjTxwoV2PTnVqv5FPcKjbJA5
IJ5EWEf6q77N0ccZsDhEIzaklVxgMIZKWyc6j+yGVQIgFJryGl0oT+zHbJb9JAcsZiK+URJKf3H6
OBn/FpF+yJreZfbg91CLok4ySMlWfqRYU25cJy+quym1BL79J3w5WBTwukDMTCy9hmWb6vhx8rq7
BUAM7az0kzywD1h6M/E7GanESfQ8cT5yLx9dp/L8DSc+9zn+PFeGCd5Kwu2xRd20pOH7L09RpyH2
1cbODtCtv2MjKFXjn8HfjUH33+1KkqjGKY6DqazJLwZiVp5w5/Yd8bZuI2WcwjMRmRS+amRVlah3
jaiwFKo/Wm61wXM7QvhILFjl1QINCO/614l34jwRNKb++8uvlta8NN7yuTDOuf03wHA2Xpclna0s
oGdb1EvnYcjwzjqQ5ivS48GpRPXbkwdxCWHzbyP0yPs6avdxJTltnSLK6RsShDxAlD4fD5Ql2laY
9dceDNTSZJt+1ZN0dl0QGzahRY3K74/AYIZcAwuIS3sBD4e5jHZNWM4Jed83OTh/yxU/z21GieS3
jDd5nxKzpJ+37spkluKrL3bHKpKIg6QqEHnvd1qE/CKqLZryLyJS1dWYblcAt321SuiLbw9wjnUD
kalw9tPcJkyOfY6oYjw4SQsxcUlVaIQv1P/UXhaw3sAqFiLSkILFT+PK0fFvAJ6qdljWEDltwySw
5U6RJAeb014dGlrwlUvR5zLyXC9lObiY2HeuxiGdzHdyTuidkBOr8Avao9RY4OkmBYVpHEu2X4aE
/2dCH88ym6PafhLms70KjTc5wrhJkrPTPY5KP9qHqNnIhWh/PvdiDmAIBdzLh0+N/DuhoS2Rml7U
VxxBhCforBeLNrfFmmNs73XbwJi+a6rjnTafpTy/XJrkzpbLFyIXo/W1dZ5IgjJwCKvJtZs+IjQf
BZPpW46iaP5LUyLohOOYgXZV/395e2gXsIgtOwHAdoBrsimUZrQh43L0qpFELBUQvRhpjTyuerAS
nik4INyDk1cRgcDddqpX92NibKk8/aD9vibSQerIRWNI54ItmRXeav1kNuI5VbMDGP9MwwvO3T6S
1vVxJFG61qs3fnj/ConjxYzOQMc6TNeleHgy9B4ExfQ3vGMixD8JPN1IeIM9i3QeD4W65PltcHls
FHOWL4pPUiJWw2n1o9cPDEoxf90h/RA809R7lecyvv3K97BntccAgpnyYY0tP2H8YUSVcUp29cLg
xmmBNzfZ19C91NrmgBk+8Oz9oHrgMWv8GymxL42pzEZ6O27QFZnfNfY97Tysggd78sHeQgRUdsi8
WrI3vznqZ8PUJM2/7LCsJ2WTTlKDUforCkBKw0xoFshrS9S67TygyBUmsKt7kpWhH1Gi+K5TMiqg
/2s98Dedk6SJsS2+PDS8UKjdZu09nbKSrV3mUzCoVxfYNw4Ycubdv6aH+V7kDDrgHYuJdjqiw9XH
ME89rxn2Q2QYt6C3PloX3PE60beqBFjpi+cCyK2rSpdRgbHuhoIt5eXTSI9E4o0y1PwkLWnp5J8G
7//hEYmRBG9Zdx5BFvs2JD1Kn3ox1FLGS42pQNHGW4Tnn0B76rg9+tZ2bMtevH3l5Qb9bVEUz8G4
xcoN0SbSTnQojG2AqSNHyA5HBdmCd0096EI4fHCGncQRUekzr+ajsdxbHRZDp3HG49e0aCH6u0nu
80OMVwS3KwqNG1gvJ+9pZyr603LFEDoIM84p1dt8TSWowu5ZSeua+0dfwwrhEwnO+WvRgtP/gu1C
ry6y9Yoto+QW3Cwp2cxMm8J+v+Dw3ZC4SSc0gcYl25kyNu/K6RYjl+/apK+GnTQuoGfX27V+86C0
8Wa0pMdAH6f3KvBjZ0mYYe8ZT5G2vryddsMyANztAdu6Ilxc71UeDWGK4CpQXvQ/fAF1n9aWFhB7
sBxizKRHDDzJXUcogYAMfiQAWG+mUumuJDsQPPDm5m0rx4idKtKOgaZlQDJsNl3upl9WpCg7NnJe
TCi44XG7gcwRYl1LvIWNyeylCm/Wq10TqKlpZkT2EUrnZXTS1UT40P8l6VLNWfq0mUIMAvms3n4a
vD7V/2hWncv4g3mlIwZ7LvSzhxiijJCRno5TlDFwKHn7agakT5O306o48YJwnnP99uBinxlYQbLD
5PqZEavodBR30nlzsnGAfthf2XiTm49Iy+ACMVl7MxnO8/f6ZYlU2npKlNx4O7JsamS0qAD8IE/3
t+hhrTKjKhGduy1ItJRJ5TuCnuLwCJ2KVAuszJknm0RA7QcD8C1QKzXV7t/iZX27NzEmH+OxeHmW
E/Ye4TKraZyp0Uocs3MQKCnvd10iA3PeA0uBrfjCfbZoUbqXEM7HMCyFtaiBGQO+1Mf9BgW4SmRU
jQnIXvgIq4RNbuT9HgYqCw/DYSqS9/PMmqghfuw+ILLkSeTtobJd06bNf39CXzxoAM3sJwkszosp
XSJI5SpFJGxxHWCoDFGXnk8fxKJZjOUOzDJpe6hZlQ2L8bA1CMWvvSiuInsIqT2AWyQzJE4haZuS
1QGZVZqD0Xf0er7bw5dNvzq/2lCwmFv2oSxs2hpTM/RwSHgF+8fVztiSGyv8qgQ8EpmTPkYkpv1y
lQxNK0chIYVy7bDv15gmd3XZVfPdSLpwcKpvBbtEY/F7eQNxL9h9NJp8vyra2Yik5Gq7tWSIJ185
KnQUqCFBXTphkSiaP0hjbV5WcZ6uI4Cw9b85zAWNy/d/2Me/FbbfxaMQC8Udtmdo0JL6h2JsgD+S
Htr/Mb1Qm5EFZgL06/DlPrfazdnGvTd1VMN0Ov+zCcKHqB4qKI8qVrPq5Di8GTZuaqwAUOR4khj+
mWKOBxWyb0UNP+XABquGeZ5cpjHmsG4N1DFgjyTz3AsOdcv22nrfQaj31d1j/Ss00Oh/RTP7+BLd
3Ei+Cxia+mInO3ntvSRqQqBQ6lgciRw89TjUyH4jQn/evHGmakdPBUpJYNeOK8L1azGkA2/QOflS
vPnk+nG7dntHtWEn26+0pPYtUgA8xEZKTwaWQ91zxk8w36FZ++EO4+OgL1Ae4hCsY9cxJcwcOzCo
PDf1mqDqkwY72UQN/xWHxLpPykYoZoxfr5FKyJh8eDo5CJe9US6HvG0GnaQ3eYzVINY99CplqXbD
h3uGJQQK8yytYMwGOyTkbFFcFNMsKRNorIb8ih7Pi+0NIUiMYY+g/OmCAE0E9WiY+WCkLe0VSuZ4
4eAy6iV4Iu7pu/gbQQfopFo7gf3U+2TwOavJqoGgSlWy5L5qqpWsXCLqY+wR95pERg+ikaE8PBuO
v6Ht2XozN6fxgjEZ2k+jQB0YGrHL9YPkZItAdiDZpXVREd0IRXkHbNKrnr5imhnkxY8Dk7KqiSiG
FAVNKaDayCRmHTl8q498K7KBwhN2UDGTyoJg92KZJyr4wiGepRfgGgyMA/xCh9n+UCgauoh2kVTN
Z9i6ioAmshpSLSZ4DbPt9CU1x/cvixZ2aEgI2joJcYhHX/mUTA1RXsjw7adJggV0Ep8RStYmbBm/
baTmsHghvBc8EWUl6yKxcFamq0V7uVxHO2l/Cb4BpulxQ0S553AVY8cHgCbr9PznsisdXl1U8IrL
T88VnRAn89V9N7YjQuqc79xYxvqVOps6mk5bfJbnL9nChdUjdjZpR9Ut8MWRLoWk48ognptJ6FJq
B4NHMThW6J3CbhiH+6JAOcr8+nSAOpBZ4tHJIxP70CwEs3kEu5opSDpWGPYgLO5i5mkYgXRtTrtN
HHCHEF+NtkOWKYsaJpPPTUSMs4pB0GaalV99qsezcVNI1/z12pvIbe0F5ccFmjlqCtr9x2O/nmz4
6vaBIwhtJXJK/67WhUkVef4gDvGCAiU66r3G4od4QyVZiSgBdv96mOjaeaHf8pAeucHJcZsSNIr9
7mkh15lAD1kx9c1/CVK/frTbQ1p0hXU0Usnlm2wXwQLRe5gu2XHqGfGV6Qug/l49tySIvULvkxxX
xAS6o803q0//1UzotXgSdwSzEku9gTZeOHUZ/Ibz4ejSG32O7BmAjb0OwMO8sPWmZ7Cy/XR1kp+C
11HWpB0T6Nh/qEPfK/WbkNbaEd7zlgeIPCIERptjzBW5QFrX72vKRibSN4OAnEuStqzlKet494xo
DCvjAv+6vfuq7doWNYyllRmY+1YPAdYqLwfvNcB5EIUJNNT7KChcl7wXL1xkUeuNXSmCmbuHnfm9
qZbFkV9LVRq2dwcUqbxKHXHc5kBMrWhPEwTeHHavpJnh7GN0d8Ph62olxPH4GA2V/owndXv46obE
Sm7pCGueaMF6H5dCRrylw+LbremugD8UJchrvpZLW46+rH+gXinoHIg6FtQCdb22fibtcFw3ttqe
ygQwc7g17HJtbeH4IkEUIXns4uUY/q4cQcTDIcFaYXUvTnX8FfOUFMc1tPXJ87QOn5LLQXDf4Uva
udofAkckeGYuwmnILuFXJEXu7zXp3SqaMnxAEaH8clRJ/tMUa27YKH4rz8c+outj0RdlZfnV4aP+
Yl5gfGLJ8NFtTkP0ZcMCVzMuH2Qfk7JA+hb8kIMa3Io83aoJej6ody+nXrddHZLg9dwwgmHbdcdu
kDuGcONToTW26wDGj/mT8DNh3ta93k4TMEBdbXJwbbiZJqleJ+/6SmeGZ5rS7h+vNXmH8qhvNCwl
78LZWiWpx4XDrCqr6nB558rVc5MSyDQ8qK9UWUD3gPUTk9rFTKld12eKxcq61BndjbgbeCGXwDhO
C/FBbbS8dfv3pPNdPZPuIr5H2NZMzIDGCpAH6F5Ro5F6e34ou4fJw9NdJIKboT4W6y9XrkZsXz80
oMFBniZpa9hPjVE3TBDiMo+s8mCLV6Lz9fjJh8G7lkQDx+Fa2o5gSB64cM7usLuyQ2adNbwSg2n5
iAV5xeB3LeFDMOCCI+496dT1sup2qAf3n6zKu6rfQbWRIQcsMGTigIlFFSvOS3b948ip1pr0VekR
Xyl3FS/q68z3Uul+rCH2U5DweldAdFz+cJFnGheCxKyRc8SNEnwyKyIiNGeprgm4CLMNZAsoV6oD
E2G/VzT1LtQmHn6BoXINP/sw/FFMtTXMWi+c3qVx0crPn8n0Jvwfw9181qgYdsZKNlvb4Fyjp1jK
sVB6E1tDKzaxpy+tHe5n86a6q0eWYD591e9js2LmvAvbraqZdkteX4lRKetTtH7RgGDqoeh0rtOa
se5lcAww7HOMt2KhZRjWpRIyRilmPe8Jamc2UWot7+98YibLzzB/tactulYUQssSBgBzY0chO29u
TLM0wyzoCVBGJJ/kmY5BWSxzpYOLx9oH4bqoZOL7HMkYwBTSJ62YlPUXloHMPQ1dUxVw6LYWpv/B
uBXT6dIQTXYEHW87y8MarzicjdodX4hS/yaeSWAaCzAmMTfyTSkdl2qugNPuyXlgnoS06iEPKx55
EiwFtJvf/Afr7RrPDqZ/ZXahUGndTU4l9m9yxQwCWFjFb2JvKNLVD1hGnTpxgqs+O/MmphXeT9kh
bIsGMEmX+MeXg7Pow8deoEwa+uE95Pjjh6jeQWQbQYrbsSJbjbwI/cgL7lC5YZNAuU1QIFwIBKji
M239NKAbqap4GiUNHqvw3xthiLRwcHk5R+FWXgx/VfBAamSFHaAFthrEouE2mgEzz/43Lez7jJPI
pOxj1W9HbHJ2nKnDzhJdtaivUpikdueyePNQdZVyGpgrKWhUP09bTZjxwh/8+eRA9Lq9RPNQpXqo
ipfqIFoGcIEVYb2yI6lIqY2TKPec0F8/CM2ftPbBn2CZpVYiG/mVdxNa7JCcrN/AQ/jHQErLmT7d
iAicrocrwUflmk72voCDsc872VR95Mr3Z72naVivmHZI3wBFBYofKSJRIYEbFWxDxG3ge5zq5ZVf
RBSFyIHvV16Ci1iW6vOoBuAYs0ppLKrdG3fD63YGxJmZeq5YMOE42fErWnG6F+gCOKKk1ybsgwfA
v7Sz+UYo4Bv2e6anQyWKmjGo4D3mTKMUbyY9CO2p4NBEHsZhx67p6JlKjBiQqnTGLCQs4JFYklav
zMHmSqybnSe1wLbPKSBE5Hqb6S+NDqYXo4dy/HoRAYY4quuzZr1qhbN0QkDeKSmzByaiUkV2Cb2x
/YWQy1fVTna9pfr8eRu/NN3R6tmyPU2tvsT/rnm1BIbEzEwEim8HbL3bhgoRwwry5PYmdwDh6CP0
RgOqf/3oRF3frFHxkR8nSRj1Tgc0Pv5c30Vj5XpCADhH++z1v48CE2GEA+nlsSM9NYTLFKIWl6H1
Yyabl1mfy9fS9v45Io71z8WROf166/MRx/HT+NhvsZ9idRqQNget2eTv9bvQ2lNRyUkcu6pa+pg3
DUKh6VDgFjhbluUxXFXx5ERLt+UMn6X2jOZmD81bpjKBmtX4esJBdQ7BPfQTTEk/HvSC2OOyEeHp
D+j+UaTwsQ4E9W01UfuZrEdUxzZZIOUlxRWOZcfHTyhnSc8Pf3cZ/S6I3a5AEuih1EBJHAaXCswV
KJHn3fcRZQPVIqfxxXzpgS3SO4ZyGxYHOeVXQgyVq4ivU8sMA960+Tlf5NhVh00EdwRvUfuk9iZM
d0Bk1Vt20WwQN2zxHxXwC6ojwSswvK2gpsc8yz3OKCgr7tqMme00WMNXu6hHLRMS6vk9AfiQgdqW
iul2sRHNk3Cu3Kdg+N3YDglbcBoZ9JoNENlRdmKKtZzaAJSMi4Vl/kc+gPw2UYA72eYrcmnuGHQG
Yq1LejxLEezoXSOOMsMT6+cWvQREHiRJJnQL5nN01vCOp7EvFrFiM/1BFscsZv4mvsRBZ0hUuJK6
MHrPopmUoo52RxpAZYFvVWGRX3bmmyZjDT8dF1EcNc1QkJjLVnC9aoF3YGjhRYlclXJnzTLdW0z1
mmp4CrgGoX+psbR3Nz1WFQ2DYvdYnbguHqcn1uu6u3diTsB1G1juGGWJtEJwgCJgsfjnrcSmoyyV
9Go5CVstUR2/JnPK1wvGrFv3VLUeSP0oOhn0MRrtaazzwhOzo0zfqAzBMLblwiggYtoVDGex/QsK
0XU78Gzhwx3iB5TjKggUm/QLMUBuKMLBhywkfe4k+80rKbV1Ov0R4BvgLm21q/8+4GSqXQwn7Xfo
7LPTQNp8tCFi06O6UKej+JeC4kbW48qbVpzRgPD+/VuTd3nYjU8KC3jj3F+A7u5CUnVMZRdNjtj1
ibcLqMiR5bWUkc0jKbA1N2mmmcxLgt/c95N1aWT2+IlNqTO/zYXNBkIjglMEfnFK5yoev+iAsYZM
yo0+ciiTskjKizXTw5YqRAKjOG3tIdDUUf49xjean6H+9brSWS7JmgBaCIVl9WPic0fJri076dFs
G/XMQarIduXRC0gzngfa8+D81YWTBm6YDpafm6zbkbz7pQxPkwvu8wVpl6kNkx7HkZ6BlBr7uIY+
+FKbA2xYa1AzKFXehsDo8gZEkND+bzwGrZU8v1Xl1zkikuWzhoZgifPqLS1s6WvJPE5mRC/4jZtq
ZbMqZMCZyheG89qHW/AyRGus+tgXxjWM1mvl90QmTUM3qKLCsoioDs2egMUcx+/HAaIgA0BGR08h
GFYT4J+nKajl2bNYenaIzFd666QLE0qljEJ7ZRU5EskGhpPqNXGRu111JtfCOOrzHjAKbdY7W0yW
XMCEPizAbxHPejV10V2V3c/wCQoyZMpOLtXvSw5/AQm7Z8fGxETTrUbw1dkXO73a+KnhHNjZsoeQ
n68yKrZqmQhlVgYC4YLYk6WxfIxsfWlqar7Kr8hSUTsAEVAldM1oMCbFFZujwx5LGIbJLpL6TdyG
SV1TkJcwSwdE3LDfYYfzorL71e/F2ua74F80Utq6BTsdPjmfhZFsythnUvqeOMu+aToHNlNEIPCm
oiSt9kkvfoWe5AZzc6VC3cHmdh+y5vuM6Q99yXwkbaXJLbmzmRvSvEy9DFgEr1ON1SymRoipNz+1
7ZMgfrSQ70o+G24TBBs3eFy9P1zPTFs9ZIqy8YG7lqtIU9FBuN1iYB6fUxSNxWctlr44Ynd2vQWq
a2WZNSB24sQ14JIoCO7BWkpse+zybUQnB6HolRJ5fHWAmiyhApPhlyzUGiXwkSNMi/hoiJ62wpAi
3ndAm2Si1WauiQAaTWita/Ohr7zs8/5OolS0yEw9pVufIPKgUaYxDuyDL4btGNStCDolrsi7PcIM
NqI4KrkNZ3hVevcAlVXn+1MkCQm1cDzk77G2/aMNcGidWAOLc8NpiRVWckhjOLPKKGSaSOcSv5vr
WKKnBNDSCzMfRTn+i3ESPCnsLY+d3amS016HU1NZsFh4uyJ60c0qQMuSkQenN6qeGWMc+Nir+1YC
RtuIfIXqViz54lDjONVr8pgwyIWikkEg7S2EyK6UOZ+8gRtJE+0zsUotuXY5h0J1XyUU3kWhe/hg
oRBSV7Zf2rcuWurbTaIxHco+4KMzJl3eMOU0oP4tipEg9marquZ9vEe6Lm4L4Ko/b58o8AEFKjni
PZ/PN7K2ikzV0Slxyb1xz9ZWTSTNuFgltTjxYW7lv+Il2yIf5VK+1nvDV1A2HLVWW8wKAbUq/dt9
SGuxYA2ymLe/BUydKitDQ0/NhXQkn4/lIjIFAMyKa8nut+zHCTIB4Dnc8FGmKhNy9mumGTQ+VCwk
lJMi0jBqirJd7svvb0Y5tHDJ3iD/zwbapu2oNn9OQCwgMObVis/PeCF5RgefnR9FkVXy5B1mnkBm
slP04KWRU/eMh/30aG+68ddWh84VNYELXNNWjiShRBYrP63dkuf/262vvGs5McFrxzpydxGn/f64
b2uLvpwE8fkbfSwbe8q5+UQgTdkIGXIk2sKhkW+OrLw9xjAEFhkKC1TV9xGpmndw3/BjJO2Z/wBN
+RVNtPaV+p6RymhbhK86R2O3k8ExvJfQUztli6Pzm0UXZ6jl53hX7XN+15DzcTTlLwGCCEqLKBh+
mLiYFvlbjUqXnI/wE+wTS2O35WT0ShqiuG6zeNbvHVfwQCBDci/SNUl1/6q/kQU25HiQtjunQmW5
jyECwX825i3Hcmr9GCmS7RHEgXUaakwwv7cIwdeR2guCinnjV8GBhwcxMxDie4hsZWIW6L9oYiFB
tN0ctd5dDqQe/SVvyCsywIjosnghiqBepYPctLRbBgZU2BB/HpZ/qL/0N3RacHgfvrkHsziCeAig
G8OkVPdHXLs6M3jUHA4ZbfIr7lwAtxzEkX5Bq93u3yJ9lDPBFKK5U7c4Wuw05MWyL1lsrWJh6mvK
djpeDVei/ajdy6Ol02mi0+UgnGv/l5OIPgN023w5HebA49SZVKvABf/j72j2F+wHUdnLbGoJwtcn
TQoax9c62al3z3alxdE7wjXpqWKqMe382RWzWVo6Vp+iYSAhGhcXhfbKKwlVcRSTjqTY1FQDfCaW
AVwIoESepFBZYjr7Hm5EkwpeEgvQLHSw4VxIS7jviM6FXA5RPILp7EXJ1iS/xW0ywJulzhnjm8fp
YL0bHwpOvCMOzrhUP1pvLzqUCcVxjINhLN5MEIKa4FueKTEht3cNeL9tGWCyO0VpjPcimYtQIva3
9L11cHXF95MHY0cb6g+OnpFZSlDcuvmy5AgpjdgWfLa+iU99xdNDjcWVX8v2zytZpP9oed64FnJv
Zw6fdifdDjmqJE9Xz2OxNmBnHqjYzIykEPcmpof+egsJliFrHeso+fkKQ2QxF/92IaK+LJ5w1y6U
PIHns6koHnOAAJ0FaEIKankLqT+RZTwe1qP2o/z5bFlzO+nNLRVQl8MKdWKhAPl17FfEV/8bjMkQ
FFFTFz6Qu/vfeAPLRejEM6zP5XVtwO5ME2e9fjWAKFGrgT+kWIYF5W0RK2N7mI935Qu+saAVy1sK
RkUeoIdKjo2dxzySFM2e7ErSXS+Sfl2wCZm5fihsAPQVP9LAUfFm64dtTKpAPXrA4W1+hw/bZbUD
114g+Ik21uHzyamGKa2XWwcAekJaV4BxQObX/ZI7mK7cQnHN+6XWnm6K+3kAyqCJYAntSwaSvo7q
+iDG+N5oVmow+3mEUEB1XGmedTZS8tY77kEqFQk4mZPwnXVMl/3OL5HEMyoFsT6MxTD8Wh4HomsP
herZkSM9AXh5xZRYHwZ6v3ChSkrNU7DMfhaYhnIuU32zq8zoPMXQ9uFyXBCgXL5sd6P100WDHoPe
qz67nUqmU4R6LbbV6X4tUGO4DBL++9D1/oxIGAOa4RYw2psojHtqJsOUd5jOPj39zuP2gbW6aNd+
t+N/H0g6abX1yvuNwWNV4hd164/jlOk9Ppgfzcm+79+B09huUL/7RryQV9q8EXy0soPkHxcZIAEQ
TDA2c8j0CYy/9CBgy1Dd8XLZfslM4/dbc/W2HzzydX00i00YcxDmKmjcLcPwsmnc4lLrAcmAY4aa
UJvmObtP93LC6M+W1ct6ViNzACQReXVuKVS4pTAMa9neVsaRxnKX2MbSK5zxQv7UlUPmaTNAcUpG
3uRdShIK1hPFKUXmsnDzMazFYBOvIP+BYbBcpG2+WrRDLevqAQtWKpl020nmrA0vb01jXhmu8IlV
VVRWfxLyGgdzYNP6fNds9sM8WnFZitrM1ZS9JdYif+JBnFLayj7ihkfpb1AIZahTPWsjegGG3/Ml
Lfpqu5PF8Cz3KnqSbS2YnGBj0EnI7zqBcz8pJiCBZD2LKjdIJS0EjHXA61NEAzAWGNjlk0d0stED
lCVMfb+0+MGLmuE/FjH4z2fXVXJRF0W9GPfGKpnDLvWNHaSw5oSb3aLfHkx3QpsgtOsbytK8PbQ0
sOAC3jDLIpCwDKma/1Vs2YdSYMSmNdseizZ867sz4MQ86xCN9WAPd5OSpeu6QHKm20nDLyjaAtoi
OfCvP4YpFciYNWCq3OU8Oy75JE9gfpXLbaEORVx6rCmZHCYnrts9e3wSND0m2r38PJIDKDEXKeOh
hiejQmcr0ZGkk35bOmkCmtMoJsyxe6IAiBm8jAuycA4LN2wBw5LbxIzpGxATXFDqsGP5ePVZXBYP
ZAh6tPn1poZbUtytvZ8QFN0mPjMUslS3xDTcoDEDejPVGT+lduwSkl0TSEQ/gekVM76yJNFcoTXz
kacLlp1EtURJ2ss5XJgFhmQCCqZdrdjyzODEjx84AvGUJMgdKlWggK9P8IKFI0hAIpzsAcOIJnAF
UpkmSMHi4wBZyxt9Fm08NfGxYMDKDk3LzCoPz2KR9YNtmOrWXCvp87flnrPpD8xcGlRi2KRBMfAZ
eypUaxNwgeBmfwV0s2jqHfqJrGXkNYq0HQuMUYSKhchgtqDIdZHwKn+Xn8uQfBv4eWlelBZHIvjA
pqpOKGfBxNR6zKirc+IZ7mbo+gU0TFe8hJHciikooI8q49RFYQNB3tNBUSmuduNfH3gWj8FzbDoR
0hX8Wv5g82y0dRiVMCmjLvytwNTT8V3FvyNB9dLB/yU7b1BIIeFIl3dIFa6R2e4Sh7i0jXEOq9Ag
CaLm1XlBDjnUHGqTGqfCE2aT42i4hZOhKjbtOHoGsQeUmgH4DqOBNHxlbU9B+E8BV50rTT4UZRYS
CAlgBYuuI4uLvgcLf77r7YDbPjsRw36P6WH+H6QalD6AWJZFHS2vfIImiAmhrIYo/wfVkI3CqEYI
3+yHgI0CZx/8D8xtv489efZklPZTYjABKLXS39Hffmd9WuvqMr1YOsQlolju1i/UMc/FDEZKSjOq
VsgNYxmFVICCRsMae2/ll3uzBCHGtcMlZnGtKs0aawKFBoqyYW8/o5vDX/FF9cZ73CFikEtsznCx
n/NNEGjkEJLIetp6MZ5sBoHV1Me7LAiw0ifH1fD8gBEzDDMX5C2LSl7LretOjxsEXUJIfpddZXsb
4BY+5yjnRy/SH4ceML79fn5jHciixf/xpbVGfY88Z4a7DS5r8PIfAwXVlL9FF/D29w66+3BuM7of
GCWUygC1jgTu+ua7GIr2NrTwstjfMwGNrBl8UvtLO1fq+gWEMhQ4fijwM+kDMkoXG323F+I64+zs
WJmIGADsbYbL+WIM9vqNhT5Ze1kPYr5ym7cvyMdpacjQgjOb03DvwSxTAi1b8ZnnNWD/6npmkfiu
5FYhqFXK+LTxk1bqrCDokvKIONXZcwq9ts8kdcUBT1gGGfF1pM/F9NJH1H2AHhIbQfw29yk2oE0d
xP3F2+UzqxxyNTtdbQS3Fxc94xKp55mQcdO6auvAv95Wa4X1g9r37ELxM524YoCPN03gm1ewlHDg
CeOYG0jtEz5/uVCcBSNizEnAsZyl5stpTue+Z4lbUZgRUeExmCiUUgQPFJ9UYZcyCrMVXSSzqwRs
wmHuK2+5uUHytAGG/gRJRmUzGFigek72cVxUW2oPudRKF5wgjnemEVXeI0AefJL4nehvtmKTZ1xL
XaT9WxI1L4l2kZ86megnbJOiqa2mga/EgcFPjsfULMjVW5yCGKSEwA+gCI365IGUyawkftnKCvml
i9bUdYvKpxl2kpbUXTKzUyiGxgExe7uHkvfDaE7EipWD3xUF515vKGoMy/swsg1F0QlnBudz56Di
i102hgXbuRsGaqIbGMZwatk2SBCnM99ypAdTKnrmjcZ2kZzdTKTw6FxGo1hZaZBj1tk47hMiC6lT
YELxwQ+y0PFLFfP4nqv+QYG8wHEi2n1uqp2qcIhfXo5OQgHSD6EYAxLfKKb9GYn1xWCQTnXgxQSe
dJc/Fg76aIMmR8PUPwBRssUCDYeKY0EoH0Mnpqd44Uf247j/lTKZ1kokForfPgPV9OCkz9yXK2pf
kHNRvJ4hQXpUreXC0JhiHOWkUJPNdng7plWolnsx+soJmQSsXbTEzpo+SxIWZg400pzc13OgOemC
lskXUnWGqCwONDcxtqAVYLffe7vFCV2StTls0fb9EkLI/ffPklUPyq2dJ1Piivt4tm0/cixyN4o2
X1CBQRSzjvhRCGBgg1SdPPNhU4k9EzPjmpcfpbrauYdnFeqvPRDeDsSddwk2DKoWDgwVnrKKnmkV
XkGsOeIMZAmJj00kQmzet4vMhnbghFdlVpHJSnmwJ8WujDAZVSfg/afS8L1xL8yXUzEUEnhWqwcg
Hm+Z2wGITDWUbnzn+4uQnC+5rkAxdxYI4egPVsF6ZSN8r/+2nKhjT9VcaYSe4QD1ynMqc2813T4c
tNRQZSxOZqBSKO8eqw43qj0Tv9mgOhEsOUfhXgpa7c9GFEu/oDhsbacvfh6zDqUZBe2rWvv5EBV7
JJJ8l89k2SHwQM0+EgymO23o3RtVHSIRtTyO2UJ4mPF0cvvSdN1mOyKzWQvjgf5NS+L4R7iCsVWz
szJhqShjsUL3K/hu6Mpp9SFFK4QoeDkIxTlHiRRnCoiAXL1YELCtc0vRJMVuzXdI/5iGn2qNTQP+
pJywmj6j2MXgHijqTqq7qV0voRu9ipqy95u0f6j6qEp0OJgXnKNJcSN3n0AejNp5a+T+3b4OhL2A
akWNaQYa0aK2rHrK5pY+tMtMykgJ87yysVXBqywAvmASBJBD+iJABw3g18tVcVwOMHsURF2TE4Wu
hhk+dOcCRRqTXFuO1ONcdv0HG1lr4o+zxs+GPhfd4eR0jqvGWB9l+re5YqLvQHVIsYr8U4XidLJJ
Q4aLrWK3JxyDKMDWAQXfXq8ZMAkxwBi6lEqaGUtapxaJfsuWbDfDi8a2enQBSjfgxZ/APDQUb72Z
X/rRHnws7tnTJTeAgUq0DOAkDE2eeCxp1fu23qEM9A9i1FeLExPSJvclwKWwDLhWG6mpJWEU/h14
ZnbWtaQvm1P0SB0d/NkKrs4h2SpOvTbit6UkeLeLwOMzyibviDsTL8XDXSSbUgMDHku9EbTlAmuw
+i7GjZIXfaQLct9sDkmeLqhuGqK84xsx6K6IjNu3Ltdw0pPx/Guw7IVGxLmze2vZqRxfjF2WC3Ci
53QK/rA17uWCPzGpn3lHwx2WpqH5maf+CvyLs1fcttSR+JRSUsFseoidILql8m4l3VJtvY9CqJPN
du4H9bhUdlX8gyg4l7TyFq+xP1iRAJMKxgP+f4sngBWgUe5CXzRuiCRYhZdf1BH27MQqncHXrC1h
1aKBWA81iPFRgZ0z6jBt0gymtMWS3P9ntuYnABOL2PgIKblH2GRNYIgZjue7IpOgh54PD0rrF/k2
0ac8kxv/g/2JYM/I+bnYhBUupFFkU2ZyG05HSjKHW77uhJVC4tswI2gzT3qgcxbTtgfSBi4oFtZR
pmiNbYjYgzUQzP4//2gNW6J7b49kVcY6+43wo1Im6aLkChLk4FaMfy3ovSB7iN/+Q9bVL4rt7H3x
dtBxbz5ap2vfi88ZUEV2ytNF2UDZI7NMyBMFaHyIskgcd/QEdpGlLc9vstqiQb7Wcx5d7zPWy9pv
kWfS0bv8insAr2vnW9dYlBPsO4MDRRssFOhi7zdeUenN3ecs53zDyEoCupR5jMRKYFYjqf05gTUi
kv3oA63JXg8RXgUrvMSB/09Q8koys8SsG3DQPPymf+CyhBGkTkHWfCFF5ncVICXwUvZBMq32lpZZ
Gc2kW2d7sxU9Bk9axq4tSzFrS/IV5j78cDaiIEYTeJAL7RnNZTgM1zDtECEDWW18faMBu+mjuaAA
ZU6e5s91kRteVWEnDuAAVk7MGj8UEDnuxCBOGyVj7hVejQTQgOdY9gkyou1rqfF8C6Nx1GFeS2YM
U3CSB/DsywzoLRSsUuES0wcWCpfB2DoUDaZ6iPoJ0FuWzv61ZslEHRjnXIXbjX0vZQM8AUQeGRl2
I/7UbvSl6sMA4JcrsK64aES8NTM6UYPR/w9DUVMbrWimggiC4xWY9yklXPWqGc+w22Pv7vgOg3oC
ucUb35kR4rX0pepVbMxT9oF5PePMnSD4tYJ2BIJ33r3689RBEa5oQ/PYHYn81fhJ5/EK5MuQEm8G
zq81EmCpLh72PIyTLaz4z8oaQiDqo6YGhP5tniiNfDAwrXAzPZAYMRXRAPyN5+gIKXZ6bT1J7IM7
MEYYhr8+dym54Nm5MBDvu/YBCuXdB0omxKuZ/I7cSxj7h4WbBykbl6cEaAYzuMl83vs6Nle61z/3
kPji3vR7dOyPXP9QBdAFwXQx/il3FsZa94HXeKE8NCYpSrCT0bhI/sAvWoDnRfeVJIr5EyK+1Iwb
OQ72Nv/URNePwnWReX4bM7BMmD5iymAXnU+L9g3dZDJxxuQ395T6ZmJWT1okIsfs3Conj9F6NICb
ugax0OZy/2mGvsT50tN609FmiJAhgyzwdgpMYlaWmdh0uVTGKYY/zPPz1vy5xZshZSqOtir5Bqsx
C3ptLMVpzatrLInbbS73lO+RiCtmOG3zNnoaNlTpFMWyuF0MUGx8w7GOisZGYCXEIt/ZxkukylaD
y4/0Ny0llvz+EE6zavZ/qcaMm5roLE/C2fYFJzFxofbnyS7X4rsqqC4FY9bGBZ0RiMA4soHhBzeW
ThQFvbz/BZ5UyjdZjsz1pY8lNaLeXU3sKKQYjtg9XAwYhxsekRgVBvjP9DWh0oIj9Z76N+hInxfe
2KCWrf4HVaehXRQRd41DNvtm+7iLnie7pSrO2FhyUvah5c5/Hj5ZRnRMIZKv/5Q2RpfWN8R+6cyd
kEAHD8faTfSHUHjaBDfi1+QHdmIEvJ7qAruv9QzqD247iQ0TY4pt1eKhrPHCBFI3MLSz1EdJdUVm
I9zrzVpHEVGN2hE7C2QwtZy0FThcFzW4eUF4CTmqribDImjmvoD4HCF9MRSMUHCMRBGuQ55V26x7
ROqoHoxM23BIxqoOvtqvWehNQeqngBimxeLHchO/sj35FLqtY3yw0D4mS74pNDUneKczOTRdC7VY
ReYfDi5mlv2GTDyIpo35FExI182HqgY6Vvc3nwf/Id4wH1Ls4BQqBQ+frMAYYDenoXYanurnNynC
Q2X5KBSgqFesyGqENhMXd5kGb/f/5h+gHwG8dGBFXuanfz4c0YZL09Bl0MlltDv/EK3VcL/RnKXC
w9g5dFLQjGboVhyTyOA1dUC0g8vIaxD8/UnXy7pQvbKvm93Vtc4vj2oOW3c94WpEEb033LcREyN0
Ome2UA0XIFFU1fX1X6rFU62fW7kMJdpqyU9Jd7WwuCgpjIq/OGzPggO6uF/gIDLVn2xs/FuA2kwz
GrOU2FkXd506N+et1W3AluIf9k5QqnxGo70ukpyeEm5Q37N+MpD+DbEaYdLvyxNpIeiAe1cjQaMF
0e0mp5S8SmccN2cBcQaGcVQpvRhXEwfpAfwh7cn0lm/fruftitsuV044OcADH6oYfpJ56+L9uInJ
qCShmNeC3p0vkVrH/5m6GZcTbIvYsUi0DmoBzZZaQEsqk72WyfZwUnp1hd7hLU4Sqc9FBNeXKhjP
ZJZYQ6+CMfKZg3AgbvvISKLU4ZAHE5TJeWqE2GVg41xpv6SNhTQniCqlAeGL5q1PXQGJutzDtJKj
uy58WVgh6pvVl/06ev73IL7lfdPHjF85CC/yX3FsItQqTp4SADolsBet0i4LmGogI1pvKqAuvesH
aBvA0ZNJK3JlGOuVvevg9YcQeq9Vxd/zshntTm9OZ2a99LkzfAdRW6FiDRKRMp8GxWe3DU/Vr88w
VP62rnq29Kcd8N1inFL7V1Egbn1LK28cSa+5DE77yto1eI0Snfw8m/uH3aPgRv9JYyna2e6yjoJd
L0Lpikx5lG/OqN6ceC12brzg+t/voKinzhfcZg46nMpr1OrrHxfpaqzaFePRMEZurJzj0zrnxosv
bil9cr44l7f/NkamYgDE7SZiSvjfFeiUDxXq5lsmfb8o6bjpKLoPda124wC04BiaekhLr+Vtui7t
h4+6ODxu6sFZB9XjBzp6Aqd89vVWNvGPbhcOLpXhE36cDOeWykry8cA6Rkb6wvji4N4z7sYc4ah9
MoS1J2exrFGnqMk2iv9s3xwlCaTf4cfRhmzjmUiv/OprtuvPTT+aeNkkQsnSXQrFHjU2LBd5x2de
H1mvOZD2G01BdwIdKvncIV67oD8sQXRXfxub8o1Lup/YLvcnuvzIYfd32znENse+9Nbfi1orHe74
q+0AqGBV7KY3tNwkQcCu7p5LbZgXMRnTE85VvfzlHkqWaiSo2HNgPto843ZUEdblj5oA1TAetFWc
aTeEOlvtmuVsUHjDqL4z7lkWLcoBCF9M04JSpkOwTUa7SCYVqbnb/ABaddJQdybKso9m66MrZaaq
3J0a1QTGrz3gL9eVaVDZFiuOf3i5ZgTYpmMzNSNJ3i4xL2EOmT7jApJbaLI4wI8ed0sygM5f39oN
MKpoDzIM8uil9L5L4TNhmkqECFvRM/t+iX+uqAI5+ILB/Rgby+KAduQBqJa1QVX1Go9BCVV1hi2o
mPBhXxvtpCdkaerZoYgqX5W70xmD0FMrvD83N2Qgt4s1DHrV4QQmnKfuF7K4Ir1E4KzP0AIfgqIK
xAyyHehnJof7gCKT0qZRYpNClP8cIEubZhIfR7ckgq8Y1Ga08cP4sGQr+t8ihppnqjO9MNd4qca1
SdANzdsL4azT6saqjMqERXXYxBZTjutvLmd8tWo2sc2tursKPLDQo4AA2vR93ub9AKligA+DaLHk
7VHI3QoibOFYn0lDC3hkVPpfAkXCiTyOaf70r70UQtSs51+snlNukW8RQJcz9fl81ENsxzFtCRTf
E9SNm3LlNO4gcoGFWUhxzmjTeX4JWcPdvpaZYL8I0BdfB2RfdK8E/2whtYgCSOsJ2taj0VpEegRX
MiZMaeIjukGkGFyu9mSJghOZfs4TialdKCsq56bTu2lp/Nm4jcGJrXDgjlZRJjoMPkGKLhCFm0w8
bfGEIiV0sRopso5hLspIY3EWmUmZDWzbchUL91wloq4XTnFyIEo4k7bU5Epp4esg/oPyT19DxmHA
r9OXY8ojQWygYDB6jVs8yiKzmJKz3721b7SM9quU0nrEWeA5JQbPx7eEVJU3Mt0eKfnfEg4I+H8m
+hKCaSV+Zf2yfGyhYErHRsDPtfsKBy3nY3aZZkz1t3OZ864JnZasTG7M86QD0VBeRw0ALSzdBSIj
A+AB7IdgiTQEcavDbTUE59BV1oSJyApcMdXjiegB0uG1Md7xML9H9b5ghLclbNdcrD2gTIO13j0R
g9npfpIk9NVWqVGpptNCCNSCDt9HYTRe2GV7gIljZllyamUpMymCBh1IVfCQxNl8TKz3REDE32pZ
YiTqektrkj+st4S1gnveRqIfX+oGIiaHDFaxQabMRKzCfC6M3wEvyXFLJG6GCYOZEzP29ZvsB4If
GH2kaSIChejD9k+UQFmFRKDumzosiaAoUDsKCGjz7bhOWSpQFuTQm4cusDOmrBHqZndqL7zHJuGr
tMYPLpQyF25/O3nB40kapStauIUoDK/XmvxIbQRH+ulS2I3d+qxCxcuv3qMVBXaO7h/nph0WySVx
uCShf9at8ievaUBKDup4Pm6ePPMjpQXlX/V6wOF6faM52m07Kd1pHyyXhiVq/KUOvJg06v1oOJ+/
ePzPZqUBYO0s4h+q+i+xAn3Mi2yj0Qj/fSReyvW11iHsDV0xqOC7lMvQeNUYSI/6lIzhTqkXP4fy
IxOZ5/vDQobQ9raJ/8x8wdCxadvL3hCUI9WGnBYXVV5dwuQBAve1/7QPpn6aX+UBAVJx5/IxpRGC
5dJ6uRDHuWaulAgonIS6AkGYKjVeYd9aUWQkIMaPtGTnn8BEJKK6NIoqeY9V50XYWhjkO9B70rUG
ztFD2n2bLxKXaN9/T7EwdOkfcTmklGZaS5FdFdwLsdRSQYuCreTsUdVIxR0PBoJxERFXAUp7i7N+
ucNttPT4z5nw7F+9CLjp/SLLsNxG3H2TKw3Cd4cu18ITZpvdR2zgpenAKaOvyBL5OMJv2mTdNmrh
1w4xH7W/MOjZGUymyRcEa28QYYm4SHtsXj8Qxr+96AFN06fXYbMWeP/oIPTobnRUo44ycUTh/FwJ
HUwkDVBQNMx5zhiKyueXfEC+sY+lWm3rHsNL85RpE85QhHOPoC/92mKZU4bp+3USSCmLRSEfGUcs
TsZ73j0hpXhjZxicf2lODaT4tmBCSCMsp80tIU3R+8myTZqmgVxHMz8qRDYmnoLC2Rfx7blrV2xk
gSkFf8tNoXi8RJ9BiLxtzPKem4pWzuguHJFsV4cjrldRJ1zbyxfo+5pCmD6lMZM3KLxGlCvYyKQ+
bfGMZZ33n7wO+6OcSfb6tEY5/gsCt6jAvPo+h3IfTHnOmtBAO/sJNIG5av1ExeRlgBgjkQje890G
fv5qRqL5sOu2h3KjII+zLAb5EQ/geMCNdIvHfATpf8r7Pvp5IWhXsiyMfAoj7QVtPqUeP++zevFD
AylahfyvgB41msMHTbTxnoK+tzq3VPjb72wAw/AT15R6FArTThvk5KJpFv7ZgFXaGhGDmv0aABmq
7JO28S9ZTi8L2JcvI1eFzzpKl4HUP8a0bcmGbOwMDKd2gAlldon19wCLe36/JSUaEL/hfGtxKKiE
qrmYm7Z6KNjMuNvSBGJq0DCKH5nAxn93OWJcGsnHPpQzyJv+XZUZMsqPYrYRNTTYaYpFnmNnY115
rCuh6eCFLZFYDmFdGCSznjscC2O5ir9LemDosjH5O8xHPBmpYcW9k893V1psXCmIiqQimryItdyD
dKjABkov+x/ysVKI1Q9kfJI4/oI2EpDXeACJ+JRV6LcF1QLpiFVR5HG92HBcc2I8WW70mpT0EgqP
sTO9uxua3qbqu4IYEO0QGa0FO10R9iPDh8Rs61o96rxIVKIjCogTiStBdId4lMNZEL101G2FQdkV
zLZCCIzWJUo5ysJAwtqxu6HVCgGaQ4PUrl+CfLV4mEkQXRO9gqvn8bRfNGF48NW0u5R5z+I2NfD6
cPdSd2K2NlcSpdXkGJhMwAWSOzbLiC2iKcOfyhecn9o1YJxWhqz3q/E2mV0ZJnqhQj5BnSGxtGJT
ha/GtulmIa5AmK680QcI2G8idJDMoWgJfYkjs9KnZrhTV6ezVp8xV3ZgTd3xjYbMd+wYHU8V4Q6O
qUQHuZDrTYNzyks1rISCxlq0pmn6T99rr687EWN/rX8KvGTO2qI2H3v/skXDkydGwyi8tZ+KHoiE
GCZddgulmZJ/OW1kCsr0QlakxkOWTV2W13Ed8hxUgs4/gJ22tvkFO14rV79MrpST86W676nYoXyc
fr2r8BIcG+cwITQ+HV6+UqVUkIL5uL+bPZHqa0pSPXrcAKAEyIHfEEuBYlAbj/DJh526TifNpX8q
NMowGafA1SSUR/jVtB9O7X371QRgjU+FsGvS2v/cjbjodIGljziyCQo2IW82mN1I59Kt3gvw56Vv
RIQu1ZRvzcz6B2i4F5EPLFwNII6u6CL8AbbyccUhdl6vqrtRdEuCcIt4yjkrqL214SqtGJHlnC9M
wlt4y5+cRPGOkASc1sgA3zDWNwc7X7iRm56RaR4yOWXNfSx/BbWoymMVDQ1s84JJ83mC81CELWAk
LvAgwbsnE9dEVXaZfQGo4nptEzBApTP2Bw7JHjvIlRGnuAwlB9x8RhwiHpCNSnA3RqEib9WKYg6j
rArfLgyS4xNUMrdnWNcvJAy0pwqI6VNXo/Hjm0yvHDuhip/CXyJUF9We0Yb+orjqIAv62DyQh7Zp
cdUpvZQqXIXD1ZBJe34HnPsjdF58bWaMFDkyu3zw7UiMh6bhdfrGWwe4MGPVrNrmT0kGbUA1gr6g
5jeXBPGo3Vf6aHSLTRFXmLEgc6Vd8+GG57PJlEj4wlxIPC+EkCNHSaIYLsjgcEbBlwf1+inVnrbu
Ag2EYs+rQv6hwDpKoyhI5YKAvJ1WudcKi5xrQyUEO5fNYpAmSE03lv6NlsqIa2INyn6y+q8ugdF6
jfdNVtuLczihrlTt53zKL89j05SRswc6q2XL7Rbl47Obfv+ibhQVD+2RqWooQTdtraJRMz9sSND1
+4PSYKsE0cy+QE6U8V/InJpb/K03CelAJRWqKenEADywkK387YOk9QFag1QnH9vEjfgQ5EfuP79X
jdm/huN1YaatbfPzGlcxMZtl9WU9bFm/K1ujrUhQZX3lqMM9D+AUq7Sk/RmQ/eDAOAvRJygq+LoZ
OKw7F8w6tSbn0k6CauCZx0HM8/DvwoZ851prXlGx+5KXUjmHFjoUl0z14LfB2kxy9/B+jVRrJb5M
G/UbOOIYLnB4/5d3cEIeY6WnIum804NsGEyiuCMxIeusE7I1toUVkdMlRIKxfa1OqvYjBcFaNGD3
px7G2SQa61Bm/rVX8LgxA+XdcAFYILU1oDc6s3Wg13V2506waAu6bV6kQo7cQrNDthr/KN+MkQV/
QczWcghB4XNwzEgH64r1A3lSi+juEH1crd1beNLWA4sLVfIBmUBtBk+fgvNh16/morDlHoTbrxhh
YeYQh2TUfQ/QiPlNefje6sfmJnWurH25XXcngLft7f60u8RLW/8F1lUDu/VJsgTH/8DlEgjnafGx
uHGpuRWJ3QigKphjFf3N1V/dQsFzJbiENnmvj7VWK+EuDNIYd28wtlpQWT9aa76pIFnyZSKaLTvB
sDHiOn2gkCuEZotEYUPMqk5Gu1+GgmN/tHmhFrhEWA+7Ciy1V0MO0BKbl3BuUJxQ1G9b5Y9NW/99
ussJ12525bWivw91yXOMM+0zeLTDWV9C6Gz0xopBTsU0ZkwmmeRZWMno8cEIE4FXAstYY4xjkPkK
t4GqIikwzHQagjPA1BCZdU3VA1VxCm4HjUhMs8fIYhX53wK6Ro1iSN1H6YvlWDpWDMsshoaVY2sE
OepfyCg0DABCXBalW67WhJ5FnKAYMRz2ulZmfy7KhZsqoA85zyuEK19xrTK7stXMeUeOBoA8YnLE
2Axn7i3lZCmeIQmt7sPsM407rmUCz2dpuvlLysNE5IXmAK7T0PMQQRfYXg69wdk4vP0WUt4tBYDE
AafWSlNpBdHlRXc1wEXtuJ0G7HGaLGVBpAR9JP7S6EvcIugUUTIneiydRwWRa9hhKk9dxZaqtYYd
3pKmHocUmw1SP1RqDqfa3J8LuZahDh632DWA59hfqU/8Oup9SnozIBAvITD2VHlBYKlQtkVrBDd8
9lesdZRwzeafvEcPHxONTqodFbbE4r3y30LOtFGLG31JhAN9H2MO1McUzyYZou8o9tzSYbQ/tte5
3PfKEoOh3512lWznG/lA6GVuJXGWa8eodLyGqAJgfTTf/BYh7Vz7E5HxQyBS8oLh8Mtjd3buP7GE
trbjPcjf2AaooifprQ/6+Y2s6PtZu7Pq7uih9kFx/OJ9ESuYFhxZ5BVZlDEIKtTCjRslR56y3QQx
224hmIoescLyx1QK8pKWAv4JRAWqmaldCFMAHe+uEiTil3IINng3l5btEtBATcsVWGbSGtGpnVTB
X6F6Kq3NAZNhEgEhYInpzEB5/VxZQxS4HBRp/JyyyzrTP0ZPTDr5SGcQKIfHADB17kKWCQeY6Aog
o25hQ1AmXS9Psmqpw6hcQQO62wfcAXV/dN4Hg6qjsO7zY15cmxBM3GtroURNFmzDLJVaQuHPW4Cc
0Y2E8r1YhrxMXZdVSrsOQhwEevdvbutJ7E6tnYLqiIJ4noVFiwFwLbRIvIjMkXZzyxNFnAMlwszP
iVAPcE9Xl/vT+veEo1JUBsgICoeC9/ORZyVQURhYuMUWoH8wk9bzvujcE6zFnUBDBUqifvuIH23n
zNoz8Qpv3mrOO2taR2hGQ4J7itfNSSv/cYdoKCz0fWx0g9pZUTw96jluWzuLIrvYG7fbORO3ZCih
EN1LPbEpsRo7Z6ZcCVMDbOGOHui8HoTfTMJ593B3IK0DgYruAPs18m+qo6AiNoZWGFy/zf69U9qr
gCl/6DV30/T4MnzSYzD+wwPwrGck4IJuaUpsTt3Xowsc1oHkmd3LfAWudGVedbP/jRRrBiefCjBA
K7Gq4pwg5fy5DKaqeqQiVeDovmFj/yqt4ugQ4/AAIyaKKJI6EevjyLbZkkglQuNntW5djTgR4jCQ
lAkye/auTpDFmM7OdNxYBLCIoksQ+DAHV9xglgDR1op6nn9o7Gp05LbAKCsEIW+MJoBs5ITvF8AQ
eq4uEpHB+eh9AvegNU4j2RoTeoxO+/p/bGRE1S5vg/oRMx0/ijh/zvLWLU4uhNfgfyF+NbQdxE2z
QgC30cuL7scgJdf5u8PiD4zd/gi5RQsY3Fwgxq29gL64xCIf3PSDQKn6jSxZ7z4yKWgG72hoxBI/
yaqBd7Dw/YNoQLAVzlUO7YK4FOlOsbhPugoARtV0Tv9Wc0xYrdDzEZZN1rDW8od3Ls4MFDha36x/
sbKJQ94+khKAEiQaNNdvAwjVq1tNQDI3j/Z/6Jzy9LbJGjXoTIwnP1AlXe68gAJQC6EQ3YUXDk1Q
8M6aJpjPHfbPky0NmkoVo5YiIzdi/nTn5Y2jz5ZJ++WUozPopKI/N4Yu94zfMEdluuY9CJhy0aMx
8+ZqAn9syeTwpbgb0uRtBagD++ND5s02776Cx9n4vZ/vBCqpqop3FnYn61MYJA4EtXixgimcPeMG
qMlT7d5Kh32x3pRfBrPLSfucSlU7Z0cohzAyB0kkWktcrsEKWWi3sOFGe3O/wtif4taQVqMWEvIH
jp8qx5WWywB3aOqwMbGz5APXu1MqbYDyTP0t/H0MykWdoF6lkHlBsjzQoMCqN4e6Xq4n9Spc069I
qb7Vm53jxqw1F8O+DbWaa3FHX8ijlib+Uz6FWrNKOSBQx1FICAM2wOJBeGZK2CIr6f984Sg5w44G
w/8uaQgdakjSWXWBLq2ZX3feWlUhgCA19mOtUlk8wJFVAfzMyb+xH42GqCCaj9rlWzpyRK3aKggt
J2rb4chavWFiB4Yx64RP4uuCYb7i2oGGAVIzrfFyAJ0wNtC2SRfswHRct/kjk72JdrLmbHOKO6XV
W1xGnMKvHI4jE6vq+9zvUTum4gL9+6BjkL+nr/Z+pMXIgxBrNB7vEvm2lZd6QfXM4nhe6OeLo5M4
wcAAZ5/DXnlIRKgR3cMknyEbP3oW6r6eMLSkw86vJWD0xQJQ480S1OBkivg7aGgop0stdpXwj7Wp
stOoO9OS7G4Gei6HuxJu05sWw0L8XYZNsb5i+bHrX+nZH5+Dsmo9p9idd7VVQwz1pfr280grCjGR
beFTgYIw2D1gtuEkMx7FtLYGwmA7eCxcpwR/hfls5d9186dlnOI7pTO1HAVVyuMSoQsAB+tTwpt/
Naizwzhfy/3RqMGwaK3fAgWI6bnEYwqVcU4Bod2bTpPDCwIlBBU1USR57FXJ2qIg2g1zypsWzEu7
uFG1AD0b2W43ImKu6cGaiVhGuFsPxHyppYGk0vaJpUJPzp5DK4s+W8rFkYPWxGqqGafcGbFmIkZ1
AgWABIb4Ibzi6vDAxonflKP3I+1KkqfnZDj2gs6KGW+pBs3BpY3BC5qoLBb2vJuuE2bb0VbGC7kG
iHY6a4uWzkD9qeNnV0mUfZFT6mTu4ntPju101S29ZhOnGOxchMcAQLMgHYrlDQa310fI8dHpvRW2
e5J5IhrizDNGC5vFh7pnGF3+pikcK2G13y/xc9WczRB7gkESISUU6oejKEmW9ttFjgMa3I784G0r
5u5p5mbc+IW8IFBXIc7H/XiqvbHdPQklfHfWVCRiECwToodaYcMLg+fzv2bFpQ+dgFhJFypBCm9S
hYnOw9gLwUXffIHkJIEpuHI1OBX59+paUUM4Cx1zQ6ck8zKn8BcndlmTNkO4Ive8F/IUY/IONiwu
vVI4u1oN+fjAXp72euy9Cs/6H2qws/11TGZBDUV725rkh6olHSfEu/MnZX/lD2ZPGXh/BDC5A7dR
PqAaBYoaY3Xf+0bgJ3FRLYmZ+IEKPui0Yz2J/wdc4B57yYqpasclRX8wyJ9zDHtgmV8QtrCk1JnQ
Hbg5zojoqhJnuOvsu+PSRiY1wcjcZkAQ6zeuMCnZ8lYmxDaihv5+gQLb1+6SndGkR/loSxDQQmJu
I+sLYUfTs2HZbOyqhqg1yM+bS69Qa9Al5CL7JKge9UrUcLyulpG1DNRU2Y2cAnj5N2ydpAFNdlvR
txDIix+ljG0owBKVRsXJDJ9SAUQFUHm5uEC8JBMiRaGVNpX/bayIW7tctUZ3CbpMxvylIJYsqwOQ
M7YAHDLWsvDjZTs50Epu6lpSPmck/O/Yi5al6CK6W1Lx9DyFYwdD0HnauxU9USaS2bmwJz00D7sp
HVfD/3aZFZh0SHl6htF7kjsLKOS+E/wevc6WLuxfq3UugP9GoV7JuAY7WEspsYeLuJ9haLmNlTrN
eC5RRrk8zyTGIQozOTJ2jWQoYix33FuzqWtfPAV9YytxCkDfL84c7rCPWw+U7UE+hn0kqqGvGkcr
/6HoSA2Vq2fEwS3e47EdpJxYaiWetOdRkXoq5UguyvNnIZyunW5bQ35wQv/T1G74Bdh51afWGmBK
cqTyv6K7D2O9QodKQlY5TT+Oel9HZiQoVrm2muIAG2SYD+DXDgPy+XguS9+V/mMmjTSjkz62AjQF
+KhULA6qQ73YY/hwBA/sP1lGvgYMtqTNrU6vAJ/KPehDR/Td2v2CFej2S88rbaTlZ0Tja43fQjQR
Gym26BnVV9QtgaN0rCctC6aC+17KkfaWRfsy4TMN4Uu1Jhhq2ROw21qlZG1xQugcpghdARBmgUF6
08+PiddvQOxj9O3L6E6dvbG2NRPI+XqhBwVUS02BsBMROOqHKL/mRaGqBeC7k2lUPdjmd3MFMtQy
9HfD+/X/exEToClHGakE/GI6H6p6vc9rkwGwiflb3fwtAoe4Zb5UUh9A2YtqkPjk9Yyfd+D/hIEt
2N+VWoF193FWRbOwp7cpTeQz4aAX+qKVe2I6iSai/1o8OwlNGOMdH/T2f6m8EqHYe0PnLJJiwWHf
hcF4GBEc0vlEbRFfZmDD7J+8xLD/qyjw740ei7bL9KaBgwHm+j/lved/kx1da7jXX950lANuoRHu
82DacINwPKpuPIH8+KQePtCL27xWwa9waTbk1a26y6Oq+VAqRO8aCs8wKzVIvFoFk8WSbF4S5YPw
b8eUcgiug65RGWPXqjTKNM1hXQaK4jHTlZWEXXmYN7jkJt2xazg8twnmtZRzibiZxGrK2dVMLkqZ
KemS1b9IRMsbbWKX6VpCB7je534GdWy/cmB015hL1FJHhjQ87HTXNchJcGmd3B9cGca8CKhIB2c2
BhNcP92lQLhznbLMEn5YWMnAHBB/V3XALlAJLJ7yYuaX7GLootWCeBGpyMCMFJU8QDDdfu60YzPb
UIT+hEePH9/o8R18Ew5hd3wLbLgJJ1G364raVs9IIv0x0vOehGLt2ECjz/CN7tlt8puzV1RMa8AB
mwOdsQ7c/q8eBdNyNoA3tbgBUgjSIMluJe6GzND602hBMrRgZ7fH855L5EQ0nGB++mp5Drypj4Dt
XUvHGJPqzv/CijWLsb6rn9/KAIV+hah4mWwyHYlDl4SwN1M5Jv+b5qmoQpjni84hoOTiqq7fwvYI
tC45/s+/K/5+ns+SpT+oWwZkl1cCEq1Hka5Oq5Ghue9yGHt1Ssk8K3LLrrSYtW6qvxspztlf0SKT
FBgnKaTMpz3gKZdd+edVJtCv+msMgYo6ywRsedla+7pcntGjYzQub5ZH7mFdy3LajXZKQdj1c6a8
FTCH62jucx2Udu7iqvpfzP4BSxVIhyWBsuFsL7xvEeeomL+o6DRk6RARIg2FEVTTqI60tMqcihlc
lFQ6xS24k0PcwxGgwzrvMrz//Xm70gW7PGL2LlnRTHKu6Cm+a004u4vi6At5Za1YdzgHMyskgrKK
RvQ4pF4/mKqkaeXHXsEQb39WPj+6EZlj8mdv+DQDiDcv4JhacxMfbtCiPP7/IMvizje+bZy3i2A8
alOsvawm73Q5f4FEiA+nfyuHNLPv/F0JMnijJt3a/u84MzraZ8xIuA6FbUom1kpfVwSODgCml83l
suCSuB6MWjVzH8s4FakEbGBKSLHA6nBwSvnqZg6BkLX9btH2sv2pjxm/WzJ5bkU1yND2MD+qy5lF
lpOPNhO182qKhjX/xDoISAwuolmT73BpobT7W9kW2V77Dp4C/Vjjioa45b8YIcN2TQxy6A1GjXGR
PdWbUFf+lM1nkCjHPjAL/Tr++0lhfcTwCcEJYxO2+Mf+4Z1uCqSKrqCe3hDDxHc85ywph/OZ38sr
7NPswZ3ODE1WtA1p3T13npit9AoxASpyir9Z9V1cyzcErt9AzfCrr0VdH2yFibcmk00PYp8uWdxB
RyDkcb2RS0slNcfhVPk0CxjiONex6gZCk43fmXyHVthk4EWR+fKyYcuGI2gYNgzNp/LxjV5vlUcB
tyghuAt5qxEF59tlJyOGA6Tq9Qs6IA7TUWJmWKBUHNnAv8r2YPZ9a50F2bp+qmjsaF0j8gk65AMD
vCs+lp7PPUUaK8ovGM7c4zMGMUtjvj7M/uhgGocfpO0p61GOQq2N2U/CAVg2CCUPgKRA/rIWah0a
VgkI+dJUVnF8Tb2NpexujceZyEkgV4UilYFJLp9LC8u8a5HwTMnTTZN41az+XiBSojvuJ4JG7WPo
2auC+yx3RKv9rfjicqvp3wz0MM1T4MZvDnlExyClmsvbwiPEX94bDSF+dEGeaWLrP71xLGKkHp0V
co+Riio0Zmw9GwAzzo4n6U9AYMu4U2t7xzQbgUfYLIV4apXS6PfvTgMi6LlTlfwKiAmTgS1vHwa4
/SULFkNJ/vsVDNPYeQsmbc7wY2eAuSPKyDqb/RehJG01eLGKBCDZHbf6IL0Zwyvv4bWZTIpapkh7
5dBfRyYX9MorMceH22MbJUHon0fEMKFnz//8LID1RobBHeMBgsSEzcUbFvzZ1L6nOQE3rW8Joq+8
+xe1O8kOH9j79B41claXmKDHG7plLFKOh7emGRXRUNJ9VOt3czzNAvgyuJ1Txq1jqD0ft0m877kR
ZNl9i4RId2AtyVhwwTh8TOASqbORlLwGvSmbdH5qwl2aYbJI7Z15K0j1d0DuvcUaDyxJlnzPlm78
CUAW0KEV2akg9BrZ4kAmCQgB/tWkhOlols16nolUfpRzEtIzdrSf5yVcK0iuMGsZ4RlMsjkOsjj2
bNzJNtQE72rXwV3aa9H5vILHSV/sj67waeOFflbm0iSgc6aszfB8CVxrzcmEC+BVxyBhE8iv/qSK
5gYaV62ReSSaOTqZhndMtLXT4y2PQcOTRbaQSJrFMoFLbW6CEsqqlkI/XHxwz59pz49R+/7k83AB
sk/p4nL0NEGXvFVsJGPQWvOmtW00OP9FGZIJzeqnm8KUXtWW/vN4taB8xBDIf3uDjL1XHQ+h3Gyc
SaNx+Yvtk6UoHLpU6p0geh3pbNroXGrfNvy7acbNaZoCpaK4vptPjCLbEQBDqtCrZw9RIAb8aeGQ
rna3+1M3SqtfPULVLJIIDnX7OX/FypQreLgsgvn9/eN5oGYS6NXRzT2bVFQqzQ/i2bKe842dy0su
6zsGS4gp8qhuIcLds1l0noGhwoGS1FqTS58muwXKbykzOdlFbuzufRrbuvPW3TzL02Pv2g+fILV0
+OcZ7BFroZgUxQ/VniKck3PG0hSzBR2iSqB4Sdf610d5sjX8qZS681nTtk6THDy4/evcHllYMu7K
RQCdi3ImaD0SgzJac77bWIWbXjEEwuj6tHvE14yieUW/P/a4JKDypEHtStetqY6DeLTO466gTzs/
y4M4UaKtFycPb3GtQNghk8cBQuFa/Pycq5wPF9QKtrfnTXsuI+/nPq4Hf8Fj8cfrgirqhYgWzloa
/fuEG/VHJbMwOodBv6L60nOFnGzyYt+/yI2nWCQu2HH+rxdRhMsxyQyO7rgnfePCru7G13mdy0F9
mYGJM2i51wXNkqhLjTuZXr1AO+/XIHMf9n4r5y451LgVziL7thkXWjr2qnX/dQhOspk9iPX2Zx+Z
LD6A/6hN0oKRMl9htpK1iDGXDMPA1YM2u8APqjQn2EDZL94be/JBSj3fHKXJ0DF/pYFc9zxa4hhQ
VoXB9HhxxwNH6R7LUPtFT7jO6F2+x0+nwvHSpvrs9mO6pRnlrR2G/Akj/HuL7k7oOvA/n4tM3GsK
Yyq9AEUy7AP9H14lJIcVuOrojihi9hvJb9SSmMznbh2SAy1jU8SIhTsz32nlGHLCXPWsAQBvnLq8
UVBmoNT2MzfWG0EUJln3/CF/PGqQBYgqqcmB5eoBa9RqXiwlzWz6U1qcAB+TdV5UIaVB2IjabmPi
9/dbE5dCE/4UpH1Y/FgRu3Yr/oI25Ssb9edvD4aN9qazu5Lwbo0fSYV3i0SudkNJcbDzyAVjSeoZ
duBvGAIEWKisSEPlkpmb+IljtmH7Z/H+SpSw115hWGClbAbpX8721gucV6Odjm5JoQZMFonKngYw
mbffS2kWLm/Oi5tfjZ1OFPu3KCZCmCwymHwL6M4aulfvAvrWw4ftmHNW1Zy3Mc+Z7RIRPeppTzjZ
QIPGx9EzjRIETReKxWuKdDIedZ0un+MuLchrrOmrUaodn7ZpMex84OE4agOTvFZfBhQBzs/9TqPj
XIkZ8sNcHI2twmkupjpKpeffhInMlBZm63AlhiJ1KlM7xCd1ZMGu2q8v08AUc1cZH1q+RyAog2jx
eAUUroErWQt1aURhbYR+/zjayuWa7g79gb1ZZF9EECLMqCtLfCaT7otvqmhl22t5coojYeBk426H
OJd5zhDTLbJkWXvD9ccxh/lEbpQklJCUbEbqST+oXkWELZ7f9XpwSqMwCPewPUJknU5PxF3oiUZZ
/lmML5mo2ifVNxXYSt4AHYNZaQpzCktWHELQeMSj4wbibRhqPqNEAz0WiMZMALoavkid2LtG3dju
ItYTfG9QQlIOnbCE8F9QuvIdIMqEpDxFVzhaVD0hMwbnhnp25R9BatcNjI6Xjl5N0KxBMB6hVeP2
iZEWFhvNxO/Kccs2QgX/KLF0et6Ik2W4alpKCIZX3ON5qG0D2qeoGwbT37kfXwzBoLhPO6Ve2HRy
UUJbSI9DdBWTCg+FtU5eH+Z2qTPlE9XWoPxKDW2l4V3dGZS1cZJcS4bwwbUotmI4N8FDHDSz38YY
56FAlARDZg3oOAZwwz+80kqALwYEek94gogSjscamODr+rLOvGW0i70Koid+bhlF49Bmfp3VvA9x
4d4Lo7ozae0kq6Oj+x/IopmioRtW4ueILmyVduOsLTKWUzgqYOKjwWWo9FgyghhZbzyvmJmPT91/
LjrUjAtN8+F1tU042J85P6qMOTXXWoVzm96T5XtdXrTekO7ctFj2RLvXF2LmBi4wLAbB0hOW3vN3
JSIGgbJh0NgE6bbzH1e5mSDpkxFnv0sJFwXjQQjw6JoW0D9xJMbbzOOhGHSKQ+3PDVPtIcnEThJm
FkS56m2HK1ym0T//q2vz9JhxAPuK0rlTkLMYO0f0VcAE/J4/nD49sWZuJ/htbHKQmsqNr67coysb
fWc8OdB6jLLM+1Lqo28IUK6RFvdjSb0yXAUZFk79mWrhyTbg2HsAZJyB/FO3ESeZKk4k7exqlujz
5VSXKHVWSyfOVpsBDOqz5TPWLEJ8psFq9Wu25kzgYbG6KEC/BXrOFE79P1Q1H2scnyxDM4VtYMiK
lQhq/g9DyinRI33Pr618fVLpX73gVxijsyHfdoj0q3KzBRtZvU7V1+45rTanvrh9N3AQdpDRJBTQ
xMQj/K21Bmt3+NLxxNkrAT3Bs2Bahk0S1rSUCjrS2v4ZWcBbfzLbE+RhnJxkX4Kpoc1/EgKK4+Oh
yCDtnQ73FsebCpT+1rEjaVfgZOUHy2rr96hkxqL82N2hCgbDgKlrG187LWdR6FGEkeBubBD75E9z
hlk/g98mxapzmHdfqeLgleIh0ZrHUOa9vlmPBBEg3CQHH1JM0jJqS11RgItopMJQEAGWIe7AG6PR
2iIKWbC6LhR4zuEJBYacfSK+avuUPWSZwaxWkMcwVTcnIkSMNrwAdGDMJUuPUBG9HhvdE8wru4QL
HZXkEauesNYiq3RzgWPArOcZdUM5GmhV/Z94LYSXFtVSwJuK2dEISn9IAVTkUtYnuD7nBVD3uYzu
P30e+3kZokuutEzaAZAORgvpW5Y3+Yy5pC+qYWNuWg13kt+OxI22fBTLcJr9TCaPcvysBInNAYTf
WXx1MEgEwOArClYTgQgOd075YUsOa8hmhrUSAghxBUR+CDNm/ktVAkznoVZVo+q8UrWdih6VBz2K
J82FUFWdhaBIWeYNayXhViQu+ioaQ05NGjZMVxryPY4IOf05ndsIjSKbbMqGZZW4jTbXuTytfoXx
2Ncr1Dn0ipKG6N8yvOVcDAsYfsayXIHikB8nsetL+m9jpFqDzffiYtESObK3fDqh3pDSOb9yrss1
Fn7IHuALzsx2+fbuZKltauZP1wbCtWZRk4op/tYkMT3ig10uqPJNC7r29bdDfk/yGwsk6WOT29S7
+rYHBleQXHYwvEcmfKhdUHMLCi88hQBxaCVdEhcToY3cR+N/XpW2e27nmOWZXgLd42DqVYVPNd5F
LUQTcWUdsuldlftpOYZD8yUtitP/8IppvXGLWKtXRAQG+DHPo+cL/gEPdH0jX48oqzR3sZeYJ0tT
uh0xzppXDHuKKrEWP5wnoaZ/Eqn9Spl3WLVVk0KZujVvphuTI9p4CB1h3e0QOHDHEgwDAEbJ7Fnm
3sqazeIYdwKuEqXzGMFKCmiQv4phXgJlxvmBYMtISb939xlMmaSgG4EBB8SaVzftZaC74xfwlvvO
g9kzZwiH/RTjUsL6dCqIiWS5bxyXkhnsmCgS4HoymLTf+mGtDuIkA0o+kT2ppLX8WPTs3Iv88TM/
BzhQwR8R34QpEkQnAga/RFgS3JqQXuMdyyttnNg79eKvNTrTIPXjK32dm+0kcLOclZ+9vaVt28IE
egSd/Pnkt57y0v+fEhUixKH3OUHD+CngtwqAdAPapmIFj568x2LrnydED9pqV2PqNH9Plkgrs7gd
Pe7sGwbb33p0N2reof4lSlYMgU4Ds+cGnSUDg1FPuUvct6TCFWgsCcrl+YYD54dXZBVNtmN8zSrj
1wHgO5Tm7KuCbH9jMXfyfMfmbifRmafe1dzOCN1IzAhkbqC9SFp9rsYjZ4R49An2rpNKy1IOvkVy
eimNfi72QXdKaYv1ysEBazD/DjkH32fnXOXiQ3s9dKpKoxmmZ2VCJRhawtQXDNILfWPH3bpuht3C
fHDruulHBDH2O6f4AyHsw2tFA6s/MeuRgiTOQ923SAWJsa2jnfOItbXs144+vzdomGSeR40zndUf
rZmCnr0po5DTA4AkfxtVdm4YhQh7W3CTzrIPwdW7SSaEmsXxG6iMozGUIHpJNuKp1nZxDwUAw5pI
Et2iR8CmhWGKV9j1ZqGSyEVNHcT0y+5meWlnt3Y0R5hhb+BoNPiqlc1OPDjmdBszBzFYo9fqotLE
1EihdiRleaEhHDF3EvNNrq1g/XJnVZJjyU2n4x0s/smhLnLcuMK8lPgJWV9fkLkmLwImbQfyxtLI
6SuB/VOXao8/JbCta5NH0Kj8XDOqLzkJEmBKrrzfthYZNDrEmsZvd5cBRHY2tagv032lwgvVG5ih
Bj3AiQ6bErmZFVL10pIHCJEc+fZmqNYzRiccv0ZYGhEtYtyoiyLAkK2hjjoPMlGW0WppDy8lP5C9
ncfYMqLbijdqcllqb5B73PuSpD9fcKBHw9yvlnoBAicZWulzsKZBhypdFJNYFbjc0dQv5a8Y3vW5
LSwYTRSKsNzHEHyGLl2/iZJjeH+YnS8uQnoZKyDPgk+PN1UeIX/QWI8wdD1LQGfH/VyVV3QktcDN
57xCor3Kp2FlTXVVsGwlggQS/1GaMbwSdsyATvt5zn8iDzmfkIPUUIr3zN5Lrt+K7hsUR0IFr+Pv
+bkjw8ueIO/4CckGdsTY3z08oB+H4BZRqXlmtWOKDgjvf3MvjkYMjs8Y7j0GQRs6vm9ylHmNwE5J
3rCTVC1a4lIMLA8Vr3ckifgTdxgYD74r6io8d1jNkKekcG9zPMCuBgAHFLX5YubawW9kUbvCA32y
sGP/Vy34AzOsRkHEHPkTai+Z21LeDsKo8Enr3ufS8pba1fmYzgI1/+OSZKjSd4fRfhiR2+21U+ZK
XUxBKklMdZ9ro4f5xtzUdNq73PwZMJD5ORQ2ojb7H+CmM8egT/ZCX8+9eKFupzJtKGCI9ty1w7nM
2FoSvMlTmr/SOKacBUxzz98eA46qGhiIJ3wr/zcorFLEODV/TWaacLdl1gyrNZw8kcj2whjA2p5c
KtR0eRjSGnsWjPH8TxLWJQKR9RBXNJGIzT5BtmB+3mse0+4PuKSEijwvg1IhlxMuvctkH/I7NiQy
vm7lXD1NztP0+ZtFBvD0FqSUM82xxx/IbPPUn2fySWbP1PAku+OI9f4aLFqfnhhM4aitkv8Cc40x
r9aGaX6Mqg86CL6kZcgaDpOAFCS92OoTEOWBu5r79vosYlghChqzUeWr0Rq3MweERmTqt+gxa0aL
T/GaCcrauG5+qGfa0lmU+W0eClRmexFL4G2VRLlDfUn2ZaugV4/7F9QS37sbvUKVle0aA5ks/0AK
RlO3250x3ad1QIDreVneAS5q+xUwJ9quUUXSlKjPgrREcsNDSmu/Fa20zLzYt+XIygw0JL0kcqRy
raOJ8EwVm8GRAaiGUptqspGeGokSiDglJ3NREJ6xFrA0nqw3y2btZwqgKNLRmRcB0B81tCPM/UDg
0qFjHfYr1sPVWUote+HGXFzjmj+4q42YP++aPi27pR7oAzUQwDhCkP6+9MNsABf8pKQR4gATI8Xo
F6qru+bk6blllUFIoX/4zyCP3yRdiDp8azAzdXtuFF6kqN8bfxWBEP5QYlDZxNsT5ZEVEuEblRvf
HJ5lGoktg8zwR/tuytvxA5fkuVQNdj6dwCOxfTHajPE07tzHpgi8WIrztlpgK3jIGUiX9YEd65Ye
4SUufQG20we6L3rtQ20EE5BHZPh//rOZZ+4PxTXN/crqiv9lsIQIQErDXMD+iNj4d3Bc7QQm6UVy
Bt3vdm7U/Qeq3CmKtEpzikeNKrCccOMRHhTS6v0apEZi6sSAYDaUqgu0hpgQDAUXNOr409Z9QI/m
cCfAvYqC+LUQcMKJ9CEje2sRzjpCXcVABz+iG6esiUvXzL8xhUwm1NNtTGo8BIKaU3ck3ydaIYfG
4LdBO6m/2N3j+hMLoVGFOsUDYYqxiWE2hIoBSx8iNxT7W3dXVMJFeZJL5wNW0NgZKQR7bKBXwvl5
hmzBn/cDGCQgraw6dORUq7h5N9q4UFIxphlWu4qFAm14g8IuIuyHvXhM3yiWuuDtWmnaKNo2rdJy
yDGDEv1ZCsKSQgS33uWdxXpNIBvF3hRzOt799o074099w+S+smRHF+y5+o2i7JtvMbExMicS6Ljq
rFo97ci/YCLz29xQtHTk45fZVO1xKX42uOgKEXivC4KcZAlfJ7Oj/Dp1h/eYMQw8wIg0+csdSZXc
3Hr3VtI61mu77FEr5Xxebs6FWTfpucar2VZj/tqsLhgvnwaZKmDPh6oWsRqQnUBBOgcGXMRaRvxE
q7azaZhiClz9uefneadw2eNXrvNzqZBEGWpWS1fZXqcYTKsR9UADGwYyRUoWZB9OeCwZLNKz60Br
FZLjpSI8a0wu5l5RBlKbQdj8K3iG++3y2qUTShjb4+EZkxe9O/AVMdJGwAq/d/Skbe1muRfl0R2W
hdB7xQ5So/Qd5aJKyp9O7ge3tF60qG6sbJpev200pJ3KtwwAWRcyaolvNYyZjkGZ8ZTlAbhLvKbL
vPfmN2kqnbR1QsUnuxAtZo2FS7Xdu/tfnEXM6xjom9muQ/5gZHHR7XXRwB1QzckFwzCx/2lIyFG2
zlz8dyRIL/KEtIyTKNEOjcynt1VJuHwQLCfYjbek1AzPqANv8BkxZ6OzjPEbG2VOLeJ7s32/606z
OdPCY4GFEz6dCzgyu2NW+RuhJhFbEa0clcYGkk9CYvR/zVtiYMXs/XQiQ4jIg9GzwCYRKWJgfmyc
+kaWC1VY9y3FGWSA1VMtkbRgwm/jc6VOjk8ATI2RGrSuNBf1AkW5vpgXVX9XBsGGUGarpeQPLwYt
QSbjgQ85viUCd8pYZZ5dHRGK1WrEyUtEBG3E54eUJ00q3/nERMyfFtK4PDPQTOFxA1HtoBZX7FTQ
3MjyhgZQ80y7S1er9DyLfH500fo1Vz9zheq88dE+LSAq1+cN7cUU7g0U7XkUU7S9kgP7h7AAK802
DwWdgA4QLumiqcsqvT9KSQyUUcedJFCoZHMidE6AcSFiYdyPejN/3a14pZPPBKAjn6dWG+tXFC6S
YY9sHot6jAzIDd8/wqciea11h6YS1xzu8Tf3fR7Fs3OMM41bJG6m1/APADDMDW1CBYOZHp/Qqyz+
8v9SnMJAxGFCNc4QMk1jwgBfv7GHuDVsiqjXv6AuBPpoBcQ3N6vONL4SQlRivATdF00+vMwBp7nz
nq2hxrUlaUmJf42wMxVQcjrDq2eyHSTOrUzFyAY3Z/FC6aJTnPm/oFl1LFUfEZj/Qb22Yq6JidlW
ECf9zNLv5jVwrounEqLn2HreLdUGGLFU876beJrN1pDwoc2ehfHkoTaHL5y654SuJZjuTBPW5Um8
Z+xAb+aCy3xrcqwZFM/O7ZFpI+kwebSE6rPRUqZbKmWAliBCD/EYyBRy9vVANARfb8aNG3vqTDz9
JSyvSpKvTuOOSUdhg1stVs8n9NEf8A5rNbKHxJfNztrjcX8kU3hm57GDTpoSHr1OSg8bd/tvMAJ5
GXGnr+LWYteRZfNfxSQ4VGTnRp9freRrJ4WddLHQ+vh6fhexnfnBTBGfQAa1+R8dLueyxVn3k6K9
wdaiW+eFK/DotQiOR82Kw6zvmBjjbGuyGiwQHxBM+x8neI2Hr4Q7rRgVRH7VEi4sJ9mdybhw2wUm
svzQtC2nP3VR+dWJRO20IqxyQt3IoHQWiddWNmNImz1A2GbRScdCY3jqwL0J0sPnj04vk5Jle+8n
zCQn4h9yzZMO/axgjcjk0PKcNSEo7DPzzN+UxFK4wA5tQt3dDhQ7oTwJ1c5oYOlrANwpmEfU41l7
FpWIsOQsdhCNE2QETy8KpzO9JElxk6U+QvqUJ5XwLivsu2z73jT/i67FjvpcpW7k/fc+m/0l9Rci
CCnzxs3LX29wLn+g6nb9xIjFJaFwyVe9gfMT+1kajxyqDp5sOSSd2QRqh1VoIVVYza54OfVvjhG6
KbuDH8lJn9Nc6AK0yGAJHm3r299C2Q1bmPTCLw+5/5qqUISmnocV75s45Jg0Y2zt888+4Hm/L6qg
3rwu6ZmhKqo/PDR+n19dGkUmINk7+M/MhOStmsk0ERebETwSR2FsO+2m+GNPUuEdcKP+LTgjuH/9
r7hFHhSdXfG+Lu9sXAy7UsDDgo2kNPoDSGlYuwrZxhb2DtHnp3m+Tcla4QmMIukYmwBoTn9sOwH/
RqYQZfF6cIFWhH2EUAXghtX4TrCbTDR0b8PI8zxiPnW4ieYZJv/E94BfbaE/RH8zW3R3rK+ahsJs
plY+LzmVS79WYFo2jwyR9Mge3K8kVgc5GG3HAdlZjjXJRrNBhQ/RWGUvwFry2UuBkVfRU+e1KzyB
rZA5wKrttsRkcf6NknNhVoLQTPLdHJRVyLrmoOlDnRuoD7hmveSC1qh8xvESsv9CPWpZP+dRN7Ma
5gyp3XZa2EGKAryVprpmdOZGyu1DFmRw73H0gZ+dyifoaE46ASTkIIXuTtjnHvuCWYvX/GhwsIln
HxsQP53sUVY1+FqFAAINbF63VtvrtBaPs8tZN2vEjGJ+qxhnXcTY3nlhwWWEF4LEudwGllFgFx7Q
BlYh3ls++cUw+fZSeGcLIUNTLMv3w1XFm4KGffm+pspmHQ49bnFLVq5B/KVVkn99debfCChNFpnf
SumSsW36bhKyWLAduVTKElNsDMktMrXtLeM7ccYhg5mbR8ggcKWTaj1kuBXw9xFOYfeangoy0xgl
IEu/vOZeIZMA8QEiXMv2/hrFyEIkp+BTNhdAXULx6xmC74ck5MgjL3s3AjxaNlUQJAMieEXfEhRI
1qf8QdLO6GWNwrbIQFNJDfzj9lQH2yYPxMepUmkwcCWJhzsQ/zqRxsgiOuXoVn1ExwoC5U55JjZ6
bB3m9AqbN+yNKYeZV98lDe2urT2z41Oab7NCoiJNUNGcVNAAvjFiLtKvLN6O+qb7n/jULMK1rHi2
Lyuh8wkr/UjntXgLtczmqYNX091DfMykU2FOdHv9iIb4FRhzjyjPH6+/iHVLyzsPhHDB1ngVGBiT
6r3GEEFf3C/8iQweQficx+wgOX72PuU+t6GTOIRJhyyaMCj11UjLjClCp0ZySpAhAXV5T7FRqgGT
ptQTLcRlHHJt847io4et83s0HWrYwvZPkJeme77tBJnjWhsj9Hm+L7b184s6Q+ihWDOdoGt5qmtm
RoEucOMaxQyw+RROHqbDN9iWIzNNN3hmo6VOr9kM+oLEpN1KprS5lZqvpsQqR1aE5CDTAhTyDMrQ
6y1gJx4No5aDehun0YFYKa2KX+sC9ks7qVB2H2Rd7CDQohNRi5iUi7yNOu6kIXwtDh0EmCexDNT3
6J7IuKuOgPUzyHF2scvZrtN1121ckQ7bUsU1qvItiwxQiPMlX0Ku4pnK6rq5IP20KNQ9oDyFFNdH
Axv/y9+91vWNPKsmZ1Zq1R8P/ko+Xyp6qh/llhvrQ/zHGo607/blgZbScPfiQCrCfL0iPKMcvaeE
jco0nq80kvEHarSFdUYkmmBskBx8IW15Sv0JtvoimwIk1HpkR2nAcCJRz5WRu1IGws2artYmmT2c
9XeNWu/PnU9gM+6f1HlHpYhN9cXh1voE9gvAx7gsaW21nYctepq3I8n3V1w0JLHc689m3mbVBqXp
5CV2ER6drQYWFEcJ83MSar478W+DIjFN8bszF7n7EZDU2iEUA/aiPQwmib4QPMCg4QsTXU5lzunj
I+t2h79IRcQQQdeIRxHyI/DYty87LQU4/vAv7s/msrUhIWIjCl1HIZe7E1qmvlcPzTA3VjviedD2
AKw5y7riT7LBPDAaeyI8BuAf5+Jr0ID5rt6y0cpgGKAIjcaTsD/6hABITq2/pUKTyZY8x8/5EN5I
QdYVe8SYmEUZSzA4Xm5PpVG18KWhl8MHvlzgoWL3YwQaCL+QiGf0xY+dyIBOZ7Un03VisBqZ602Q
HwJT5uuf8p6+86f1mucMrFvsvfL17kBKh4WHJnI+bGXAWLXNem8qAMMGmYafbgv9AdRqgeJN2RPS
s8KFo1AXWDQgUlM49c2PQ+Ae2FN6hWiS64216UeRZPBT91ULqiAugSzNBy90KeIIePPiH0OIMx2d
Ghc1xfe6/w5fBe2fycCMofoaExqrIIANfXW5bhCHNcg/B0rH0NO2BQxTFDc+jseCVyP7u01cMcsM
hlst7G+T4GlcGPqCuymFu84gMxiqdFaLVDg/IgGRl03SK8wD06usP8LG2mjHvceOOJgmq3kSk9b3
c1tOfFAIZVKpwgPKPMpBugnNFvSH2nsMfy8Bmg49g+yuma3SprSjMRK8Kdv0cNElEWMb6cAezR7e
mS9tW7g56aPI/QWRRyAdlZBhL4P1N5nFJwjKTZ5OJGPxyvD6AvKqg+ttroiwYFEWrKdQbiqe6sAP
519pQ3TxJvdJgPwCZB3x1lb2GKQ+7dihekqnezUXq0Lutbw1Iwpzqk6t0Tm0M/kSTyLz3qsoZgNY
QQGF+N67qArzI8znXsaraRK0aVEESXqiD5I2wTFErq/ZVr3RVZt2LdFTboSJtj89BbOpF6SKqsge
yx520/PyExgNiS+vCLlqrPoxvDiXks97cY5Ykm36nMPW6HPZTYKzm41q2PMM2tQ1jJUJtgZLMzyV
Su1dHZsSlhnUvgKl4XnFgywhqDR7poG9RjscVUMDywxpydv3yE3xnW6PCv28znZHoRmB+Yk8DZIT
Ek0nZySnUzn6JGav6wFTTCzPlwvv+/aQN08HGaStdyRIQYdcyYGVIQHbb57kEXsQIcbcaFjMyspJ
YBcYVzvKlR1A65g/YSwdBpdj8tDy34pHlQ+YdfGIQNISAe7/+dhCjTVqFzIEXzDeMmzEoNjr0gpy
TR9vWseVfe0cLP3r8jEhRcKao21mXLaUSLfdmJDU5syIG5LWvzcDZQkGNVc5Mw8WjSEq2PMoH4Ov
OYy1rOln5MqTtUKh7PuZxTzAih7WrOzzqxYIvztW6w0fIbRiBsbcBfzu90AlaOKEO4lPeF+iRCaW
4KmFNy3gecI01KV9dF7Ty2kGluF9A/KJkmQefItRGRbvpxuYm+d9xZWnoAvROPZNfbsIN7NiWDbY
8htWG9kBSd01qfIDSdANR6Y9DLDOa0E53tVML0RIa7lVlVFLzPOzfDKT389vliryEpEjlTkIO690
IddY7UaD8SFn19tWgnyTerFgFRTYHFzVPrWXOOTInFoBzYe/TnrHm11MkZta1hjQ9aEN1C4CsX4l
I9tnnenrNxoodtheLEyJFsJtXvrGLYpZlXBdwqmj+K0tpujlGSEdgFsefJB1lhtmIWoqppjvqrFe
y5pcynhhSaVmvOPLuzqgX5kgKA7evRrnDyh1n5eMcZoWwyrPzUKGsG8e03bnwJsW//MEerD6Czie
t7xhYyMbfBntCNPO9oIkC1Cx6zr19KzvTPdSAoYI3fVV/KVuAg07py4Sb9ybikeWMN3ztfUeeZDM
6Rfd7ecv/ghPAvvUiPEZEycLYgwmm8K//m4Mgp7IxueGS2r+mkR1Nj2eFwqQkxZ/D7XmKy1NI0c0
S1q/S2IxRvtPJNGD47E/w81jXY4WBVxZ54Bd/t9mUvI1gGH9Unm0orh9Is9nBW+58eZRoXmSm9mY
Ukia5IwcmGddDrj40Cmh29mfOz78NCl0qm7hg46G8g5HsBSuEAxjA3egb/VpdASmxt33B4B8EnnG
dVjji6jYQvxA0wrrJsHUw7uzhMANTovkKEt70Gz/KvWHeLY1cRmhzsPI/UunfLqhH+AjpHk30tMo
ahH4ybAUqNhc8nnaw1t4xkWaOvFRFISMWLCGiTSALDGgKuX2fml4FZTDzzbNMr/NXycPcp83eI+F
RJJswbCauUY+iP2tHfBsDmCkWP6synA5gcZGTqEXDSOFQoELRx44JmzLZYdfCKz/TUgHr4jVmOg6
kQB1IAcCzFgfC83Zzz4rBf4TQ3OalCjx3b4VVphzsFDalKoVIBBtE1hgDZUb6ZVQtkA/sByZgRJW
/qwvLoKVxGkMTPhjDMqYxWB7I/IqOXzRGi16taGvR/NcVNE2vPBHjYF7so3HzAsn468x0BHPmt2w
wALLwR4HuI/gS8jGZjgRjAMOVefQPBcg8kAB+0k0m8VZsXhMcahOXjeDOLyOEcPiyuEGb1VklP8y
4Pr7kjiilyNeBgJPxBSAVC17S6UErctHqbos0xq+EMOKpD0qR9/bTvl9IoVrjMBgkuVoAIkKNoMr
1DqpdTwgw5L/W/uticHk74aR2L7DmmvCIn3bqlCFnkmGs58baaQPBJ1wkQ0GCxxbgwWRvT955++T
9ajoqhP7DDRc5FzEryjKJH25LyOl1zgktXc6ImFuw0wTDRrBb+tqV4MUArmWH7sQ84yIY1+C1ib0
BubTBOiT3iUyWQo7016bMOazVBW+Dt0O6aQbQ5TeW/wVS/+acJXIx04T41rXbOBimy6J9WqB0mUE
TcyfspGyqg+uyKa5fOWRPKnlMAk6wsR9Xt1sG/3qAq+lIizNZqdJWAe4t3jTij4smgmUXbQx0kvm
1LPPQ1oQfOb+u8KykHVtnF6V9r5Tgmr4wKSTRsnH1y4f1xlHST/LMF5LBWx/6xjEiec+TjvASLYl
3sNsjrBskxQTF7KQOnKa7+TwN4bcjDyOkP/g4DAEvwsOXXlq7BkRqz+GNhIy5HhtvS1gkBBBy6JU
qaxL+q0YV0YFg953rw9Wah7bsTC8OH11ykvyBfrof2LCU6jLoSnd8U61LUcxzf6EsPFxbXHcMsyt
dDeoYriibACTzFn3x0Dis0knI2HCQHD5s99Sg0FKjjRc7vverWdA/KdFjGFXQRDLGybhIvA0GtM4
Qg2G/ATYXJE7CWt+priN9aFOI1tiN611e9ekloLHOpRAO+wKYBdBmoZidTyyndQ7qQrTmibZwzI4
asz+ihrEiqRNNJryJxTG+tqi1GYC3xTHQ4omEz91eqLOIGiW9mwSb8PIAxYZRBLcUKrQz+o2Peg2
5UATeOu6GzYDndInWdL6saKPqcWKwNQYe0HVRMs1cRstriu4NJpBXMuKE8z2/7+6eYZ1jqAeGt5b
sD/mw6+tenyyhf6CI7bgHzGPPxIx6pJseBcWP4LserK0rbwglJ5tA83+73KEHAeHvq7P2x74iAns
QgVAcrvNVnBexob8HeHbzLve9T7FwpNAel9z+o6lyWM/bn6azngKjsEON2AItv0CkpJAvumq1rgk
88jz8P6QbwF+kdzEyu9HqaVjDTGfcDDn4x256aqApRLCPIDcDY2JvA0EI8C7MQ7IcdsGrmehfGph
Db/ZMDSVMjSHs5pPLrvwhXg0ArobUQLkhZ+fBDZuAfQnNCQleR9y5Hzpx6xBUMQDw/y0AVAxrjb1
A1OeC8mRqki4RNQUHeXQbf1m/PBhzM+Phf/G8uhajdY9E7tBKKvy+hjYmDgj5KhVG6UaEEotkXTo
IQAXfbtIEu4hnQKL2e61pBwbVV39ImB8Gu3IqXLCIbxb57tDnZkEabejGNXNjpbU0sezyGKcqkTF
L12XjSrptsblhzLHnIMpe0jSJl9k0scM8nWELLTMBnq5aa7cgOBSPPU7VojLwqsirlxWxgN4nSPj
tUfZfqQINjiwTHaWobd8bjE9EtrD+HAxosEPxfeZFlM+Al0r3cbiYkIEBJvPGeKmUUR4AB1JXSEL
vOKE2s6CrooLIczZ99s8ZHGlw1dVz2T0qKMnzhTd0AkDgZPO8pDjDlV+gl2lgb4VffiC+GbIAoz0
lv6wB5MOqlIs8YyU/KDKe1yVMHG9D1FMVvhcfoIu8ieQcrbIrkL5ocrDQ1cWGGWW879dMSRHM5oW
+AKefQtJVUEe4sjk5+K+7hI9I5KxXafF5+ApydgvQvw5l9D9LRJMirI3vcKtAYOzRAEv22IEsHWZ
gEm8UvYr3V7PGcs2KqmskJOuIvSaJgiQPXcF+tEstjaU+iZwL6pnorMjMCvrm7+1S4itzxK1izj/
3Nyf1wp9xkMGS2FOYQkjyPS7cWAlhs1QWvtbgL4bcFZJm176DS1NZIZShxs2eFETq0TO32E8AzoR
IHR6+0KLEPK/XG70GeO6MKNYd/hf4g/cWevwZ3F+FIzyAGk2k3ha6j952lxSeLhcNfB3Uc5u3+QK
yZ13LxZKXjyqWgCiJjVd15mbj2xWvykNWIkEYozlrPbDNh6TAADMGK55l6I+N0x45dwhhweE6qu1
55ADTcjh8FzXraSN6T4T/01r54Pbzlbcqli1Oog3cZ3XO05vJX/Ahk0Qc7mblJjPWild4aFMoQUC
Iw9oXI2dsIekjIjWLQBH1q7SMWpW//3S+OQc3vhh6SaGprpcujGBER3K99D0LUIbrjGk3JWP2PQY
cTSmXhBspMNTbxlgsJpa1rxPUcwBG7xiaQSLiLmZe/pfS6cO4uAFVWeOVr0GlNyZJPCnEzzPPCgo
6OnHvMMffwa93H0yGaZaV+YFFwLEzfy1xZ6kpgVpU9qx/Trh+ssKQq8tmim7Dy2N5iondkOKmPLd
KeIdUW9oK0ADWXEg0ejikq9jtq7Im+NpgZ1EJiRklFI0I+e6/BQdW7tlWVaX7MtLpbkgkXV9X/Bt
u4MhkmLoh+77n5eZdEhMrI8s5QfCKsqDw5Ie7tvAsPaDOuAh7bzvZrHlHEpIAVRnoCm80xM1lqKg
rLW4e+3pvUg2h8aBdFfgYtyq1ctXHOXq/2LOIWbE0Mn9wAmtAfWGFqgUMl+/TmMRDqEDC+w8dIl7
QlamhpUDjPODhC/ybdviStF8Y58EkDOIER1EIiUxznEtxMJ+s41XohNzGLQsDNtqNvAEZfIANvfS
QN9yl8+p48pLx82ge71Tkw15Y+uJrJNkCDnWBBe7xCBmuRJhPPCRWgovA8walz7dEqtxb/2ncvFt
JKXXFjZHUDLG5hzfbKqANW9ijiJKXVxfwc42CEiR36lHlVc03HvQtbrhsvLt4tUAT0WZKAbJ2SdI
3SFvf5js0GNQdECUzBNGEbGwboucqOKheP1CoQKZhV3eIrG49Rynu6t2JgTobZhUd6fXNnQ3C43j
YrfrUD7ZCVRJ8n4f4LnrJ3/lwFAqUiW9e2O4vZDiS8YJ9U9nDubr83E1SbrA+E/FvXoRkvKSNAC4
I2tsWyiT9o7FjPcqemvMS6Uzyghfd2NbKsy7NkN28yIflwcalQuDR+nAho7AUnSwco/2rPeOoSn1
Qk+87JDCAP6PIoJfAh9E3YOeJD7mhfyYySxRq+LLcn1k44iEJmj5NFH8Eawk3c67P7lZpX5xavaR
Y8DvB9SP6ti4b397qCh0k5B/lZI9f/jXW3VKnoqb5m6dwTaIqvh0Xu/E8wV9lFaDKlKtSu+V8x6F
PHZtxC/hPBZNYCpxQ5grNeoDnCq3h6zATVRgJDw7LiJC+RPLj+IoGdMATQIR27WPt+u4eXmUZw64
BjdKalJ5QslYmiYQl57viZCvgWnNHK5N4d0UMzOO47WR9ZvAA2zB5Wlc3G5NTBHotC+r9Zm1+uuz
tNRL3w1eLUXIuLNxSwyImn+LGH0vgja+ZxPH8NcFBUPuCUZCD2/NRVTvDppqFtlqVQF6uDEPHWTi
RJOTjHObuHXcCs1y5f07c5U7+Guy/dHX0h2tnNtEmfa5TSqrDDfc3J4FLVUUO3KsBp9/1w3J4A0e
fKWZLONVyXiTCnzVVVF2NKeFfD+ImvHz3eUgEsmlljy4Ip9S4BQZy4hgEYp0sNbB7Ku9REKr5TCY
+fv94ct0//yHJxQusWrkG4daSqDxBXMYQEDRWK40ErKC2CNpiBiUJVfFOq8JwMvX+tvyFTlOSWvv
xzWKzfzwMZOzEWK3m/y3G/i65epZAJEysWFld/fGchNYB9fiY2iJf+9Nri71BWL7yijIWlipxthc
e1KFEV0S+QjHfH8vA6TUDyn/wKn/6GHF6kepQBQccDHPo9i5nhkAof0z5kAtV0yOaE2DAR+JoOyh
mgTs6uz44WieEU90UADbHuaHxs9vAXKRBJgEorHea5JZOFMjmlU3YVrz3Vz6wv30Kn2VTQ+XZ4pD
Dj3LRGdlXsbnFGHe2KMmNzxtqlUjAWwZLXTtyxpjx47pzdn8iPQDObcpj1uDWU2TwAZSI2qRvqIF
9UJybU46JWaGVjDi+RLaEowYtHTfwmBZUu6Ia4MAmdO/ZQj8zSXm5M+nh9yrvoVtfRHvnkOq6gn/
37zTuumriEGKx5XYq+ckuVqXuLzAoxEv1ek/zB0mj7d6jU3/1pfRwk9XImgqrQocGWOMzyRe++N4
R9W+V85MOP37AG//5DFb8KTD4bI8UQsOhYpgxyILHHCsxh7Abc5yd/vZb86cpYx8xELAyJ3T4tzy
w6LEvAIKlXIKqZwZyc6ayjI5pmf6fb/Dxlpdg9Y9EJEU82L3pqNiQybHi1w0DD4Nrwoffttl3kRy
ZoCxRB30iV+nFyFBJptxEYMwiwWqGSwkG9Q/3kUZIJLaaULMbvz+0BXmq9ZASw+SwhPjNGpdhOSc
dVceUPGhtsHSi6V3HMHh0UAt2syrvnWlymkJ8PVkBH7ZijIUH5suBm6+La1Mq7SlKlC4FI2/25SR
mB90wfSY4Tvw7SqCJFiWr90IZBlX94fsgSoE9jrajFPzuH5AQ5zDdLgQTYL19CM5Fp1rBo7rRdMS
sQ5973BRir6O9HuopcPy2jiZtL932vZOfGGROM5Rav++l056WjpC96rfMLA8a57DRaSz9z14LCPd
O7CHqNkEl1dNVLrzvK7oLZ6U1o1AkIG1av+gW4Dx18yuIgEHxvUc1t5BIopQ9goiS6x4wKjD8oS/
9/RiBE0V2VSijV6pv0yOe5k762/k3vGout7RIlAUq4CmgivAdj748FkhUB1W5Zw+HHU/ZjChYLrk
biQnfWLSXOxHMpH59Hfp9243M7dMKvMzn5JZ1VVjAzDVJpdLgxyjR7L9+yPQXAksmn7r1mn78qVl
0mlpcBa2U9fs8mMrXg/Osr9EGWyoc12e4rrbTGxk8fsNjc3Sep9JKD4IdAp4yIEvU4AgkbRqHEyJ
+sI2kZmNL0RTJofiq+XCGb3M0OYfjv3BNMHLi0COGIGasdfMAbmUX9wDh7dYiDJwOMQ8hyzYGsBW
SDQeQ8LlzprumLUhmfaDqVtgROVL3jTPlB9GN58xR8GuAiMqBoiS53yXgJ6qIVhfJ4Zjvj6T/GhC
ecfj0olg5yeG8qKdptEEHJkDt3+yOQ1FU7b7KPDFuHezplQ2WF0a940FVwPdcEFo1q2mg4Me0ixH
rbh2gAybGv2YW8Bckw1Yst7iCoLzfOsBcblja51chNnK/Wdrb2gwXyqeH337IIzymGJ4977kAI4w
OVYz4bG3utcMuini+KAo1cqVVrlzwdeeFORyVj4lPLLWztrDPlrjJueS8rjHSScNYJQ+h9DtBGDU
bsHcdFhxq2NGg8C2KitNKboRwrW1NnpSA7jKyjurnDah/OaxhNvF/306EZMgEHCKucP4vFxBGDvh
8hreOFvGs0i8zZ1g611ZUbIoSisfw6UEYmO1f3E4xBtCzZlH0PvCsVertBOOG57cXXYhKlhRmJEf
11iHLQoqTZCJO2+kCiQpsaPAVNmvgMk6x99YAN+vPNul12pua/JajGSrGPe6nenPx9E3rluxzVU3
g8as0VBDj0K2dr8SS1P92E1+a9+EKMaXVplaKaHmfgKe4/8mgiqTHT+j9IVJ5q8g1GgsVMVeJmx8
L7LvEHNhlEIg/5JyCoiXhLxzk4k11V7FGdu8xN68s/2Bf2ssNer4mQ07vLNiHMlpLIOrzfRV+8SJ
+IfmW9IzWbxXVclLPfTcGf1aTQCVvoMRUctPRMgu2bo8VHPc4+o9mSw28UOkuUYfgPXux2f7TLvn
WVR87QFdcgoSGcOtBaDFOE56PJYXPJStU4/shxf82sGsJf5WkVS0QNeXBPyOkTqx3vfPZx/mfLiQ
u/RbwED5yvtrmVLUfjxGyfjthJ9sKAGMYBVNuphDtgdSxFu2nZIu/uedVHos9B7SiCzbbuvkU42S
vV43spv2lF/Nw78MlJ8IYsAVKYvdh/Gwjkt621c1ZjAsnL68uyoFvmMlx9BaHqQM3Wlu+bXWVsJ2
/EMfNbz6BEzB8D7jpV4p3BJNa47bWrljcGDw57Mu9+iI4MW0g8kBsgCdbYsujOItetJelo+oomPI
htmD8/mpXFbJxJPvZlL0UOS+bxm0cHZb2X8ntZZxL/nv9m7mkTINz1qHc8hAkAUpXh+5oW82wLjw
sMnDWHfiLhwA+FaE8fqxXlIqJe2oYlYIKS+Zf7QycY0AVNMvEEbspJ7ERGq+bF9T6yDBbO8Vh4gy
YVGRPvVBxJBcqgcWJ0mns0rwvXc9O6CzBuiehScj88qEpiKz3PdSlxXwjKf++dfn/MEHl8IoeFwM
uPISZMG3hrgdLfwFBQsM3CQ6TC+gU8N25QHNFMenXPk9erJTrdK3uFpBhqEBXJ8XGNH6xIrUF51H
DxM8cQoGWPVQj2G9Lwjg72Cr90ESmRM/K6PjC6HJB9g+sK6CaSC/8VgWZbKHpyPQvWlRbnFFinYZ
6lwRetGv9w606T4Rgb40vovkJbyK5zU5pq2pbM3hFWKocBTv8Ny6JLVTeECS51ZybkH9DezW0cOC
dQp9GZw1Odwd80IW2covNyri0Imw7wPof2QZG4r3Giuxnlgp4FmtxtaGzcK6H15NhPJn5/jb80zD
faxztTlF/bp46mhOupsrApeS4jiQATRVMsl6JLU5thyzTJ4gT0eGlBF9TJO7jBgqCDmUeLD6FWXH
eqj4Q7KVfI6V67eS4csr1UZWJ1pzTMAueGONqpkvzp0QJpya9nM1oipVyGiZdM7ugEprXZVq/KCG
0xnFyCvpfKoKEeOQsiWrXDfbGgWu3fRmZC+0dJJ4OuNZqyQckkyFZmog52oQTk8kouRh6KcFK9qN
WVzq9mYae8bq5zSIbR/KbWnCfapM25dgcFIQ/oCOnUwaGpcvAudKT037dOrqURtQTIX5m+6WzwgO
N5InFdYv2pWjL7GDhnwaG0hACEVwmOqgyUERUw4bmVtwgIG5a1c7TDhddnoCxy/ELlcp5P5xsVWp
ftnAhAMUYosIFL9XYcYczXS9yZ13t4lhu9+hgY19qx0mIEHbwvo0UKJURsje9OMTSHcMMoSfzWKF
96LVVg7h85o1sG67S79liCopJQvtRg5N9z9f9VA7uysV9BjWCxVwpojecaddndwLkIOxJ4XIXAgt
Wo4GtL8FiGWiWcj5RcX9gqRtuyt2zdue43rrHxiDaKhzp8GtyIwTmB0K2ZQp0Q7XpJDN/tPyZQVX
qFo0qEzcauFJ5Wc71vR3c4sCQr6u6OQF4R0VU8gOoT4AJhjsI95AtgGFaTltOxKzle43kIRoAYHx
xZvqrh+CTTRp53mvZUYAre1x6Ul92OGMT0PLahKkwAh6fR1+kSFRkGWmW0ss+LN0jdFf9qlfZ+rv
LpG0QesPjWQfpG2QlIK9Jt9XKQq0vz9VWBwSbt/ge4SlQKGtc9RmSZ32hTwT6LlycFs4o35N1CuF
LGpg+PmJ13usJGyHVZXjdrKIEdZsqTcZPpahkARcXN+WJD3oD1w+IcBFaIdMb12I8dT68bTCSzqD
kDYo+/n6u0b44goKUn18KwKJpjPfgTMRyL93o3L/R5LYZZ+DKNAW63wkQJwMRzriETRrtEcze0ve
OchX2ymE0Mr8f+JrYio6anOL7fhRhMIjzx1n/WQDyUEZygueZSHuJqtInQlK517jj4KPHaVZ4CRD
o3vRYskiXNoazPmhCHmKhkpYRReSRRIpqFQWO8HzmzaNugzA4QJ4VBCwkc/LsRMwyQtAYr3cq5eB
Yh677kA5MLwZNon3ur2Wc/opibb8UUB92ZoP/Y3F5K7NTj+Pxmf9xhomKbuAkE0v1+HMZVcDB1eX
3I1F1ep+3qNjXpzX0uS8T6zSrYaglc60ykBhd/f2ZknbYZNYRMmIPSfKCMmHIE6jv6tSZIYk682e
XWxa5hcR3qPM4HjNG1DpF+1QKENVA9vAr35EXVNgSiV3tNHuUIQWdZ5lpAADzV2gTi8W4Q+4Crpq
AUMZYHjQaI7Wl6wHs1Qj7X4MhAts4NXrrezsBMlSzylvxPbfeyZ9tfBqomkD3csvaVOsFDem7+Fu
qT4SCGRjF05W/hgej9M2KjL5aUWNi97c1tkQ5bdcltXJgfcdcEukM1SzQ7XcBj4+IKBtZ01NC6aP
xUoC1i1Pv6WCD0Kb9gdAwVUvVbZMM3+iP7Kh2w8Smyz5966rFmw6+gb40nP60t/2Pu1fAFiEvaS6
vEoHxMsW+IxazjBdZqOvrPcIgKFedADeaSEfHBRg92GNOFeSn5dDWS8z3y9oIDDT7VyB1Hed0Q6P
+G4AcXP92Sed0mRG1lKusr2/DjNsJ0w9KMtniX+bQsXBzbeifCAuKTOuUgqc0MzCzwMJwQmA1SGT
/ozEZNLEXB13pD1EmZhZmlcTRo1PdN5m2vKfT+2ORMkj/HupOq+oEg7FNOqfzgcd1zmxs221+7I9
QmVC9cSCA0tMMJfaw5Th3DgyiU6BOS7/+vXOXZsg99oEIBtNgAEGGh37xev71kk1Y2kL/CFxMS4Z
rb5lgThnxzNsmiKFutZSxqoq99oNyUm6Cjhkq3OOsW00WNGClZxVi2nDMYMCFpqWi0A2GuCCiPUp
YfgLmp57PdlcRN69dWx4rirbzjsPG7HyUAURwjp7XAVqu9mreNba4aV7bE1AoePesLa+pbdWBA7C
H2slQ4eN4rJw6zIwAU7An6JYJP9ROyzwcwlpmDQF8596Sbek4fMpPZCRVXlNFXtpIUq0DsJJkDaH
aLPM5PS2SjDDxTWH5/6wGdwX9ELRG3op67nrORvthtIE20LIBC+kkb/SMz13SF1PYn26IutpBkZc
//1hIJIRnyRKZaK2p/hojOEC5MvjG0ZMi3O/koXrK9zf6eaCLHwbHrXqKnLwSDlHo2Eh2PRQVnGC
2BnEU45nr3F1TpZd10KpJLCyVSVN2cm3S9YCJ0s82tYfpqwHUjYnzpQ20H1/9IZ5rbCUwq/BFRNQ
2G5hNK/elCmzMGxYE1mtefNX9xg+eLOmHUqJIFFTXWvMHbaavgVtUhafGgNbRZtPDQd6VggN32xX
xf5GhnTenafrZw+2r7VQ3Shou9RqY62V8rhlvslpEGQx4xbQ0M/VKOHY3VVgQzTMVasaPiBuF5NV
vDKe6UiwKziE4+aRvIQx21JOFFHN4z5Pu5lQP+hL4zIthG5Ibz54lWls4uo6IV+doPj6AODbF8Rw
zWks0o71LF5SA+SNh+D/oDkBGoVMuNagUZ2jDoYAKVWsLEv153BVZKqO/0E2qGaBBo6LC1U5H7vG
cgVDqgNxLHnnl8wyiJZJDKYGmyt+cyzgZitycViY1eZhlT573WOu/s0UcM75YyI8O67UaAR3ZX6a
I1ADvOf4bvRDuXMiSMa/2vXSh+x/IBPj8tiNFo6q5b14H40BV0n/kRfeq0asBAupVcoJk2FKekfM
S9eDtv8+XRWSDt7HEgX4in+n+UVzLQ6k1NDpeRSuC3kJPD1pflwXaQPd4ttOFnetdRtBmcyRi7+2
totu8EMQ68Ge24qnFGy5QcYJxO6nwlOqcjjCdnhf8nzS8shlqXMilDsbTGLHm4UK3picgCn4QG3g
jKDGHgK7oIqIEchriL7xAewnT4IdaCD9rdmhtyMejMZEg8wj9YgukTOxLhwnD3OaPKHcYNLdzFpW
qBKgQhAJD6VaEarMs6cSzUMn6/hjKCWdCK45q2oj8ZYHF8Uc5CRgYFz4fiMncazK7Xn6oSLvwAwo
EGvevLC4tegUF9scf0j5KFsQOBygQ5ZH04eFzESCN4nkr7d0AjCrbenjC3TTAdK2dNZHaaQMOpxv
wl1xAdc7tCowGDFau8kIPfaWClmz7AT/YlofoZUY0YiOUQOjhj1LQWElMe4qPsXu6nsTdBkxsWFh
2aqlBDxMiRugidUgVwoz+Lv+ULEBM9PiPHOkmJeW/KKu/ZRj3ZKaQ0MYaeH02NXoEE/5DeEFLxH/
/leDENkVZn33oAEx9xB5Des93/ZSBP9P+/nZW97qvug40XNWbIyB9Rb7RycWKvND5KGlju9MWvpJ
3PjpzOEClbE736B0yYQZvyNgEqPjkjwv9eujHJjwPFaMHnFc2Dllvp65/DMtfZNtjaVf/+I8ouYT
cA9Fi95pCQfU5aZcTKY/JsO5stAQgZV+bymu3k4QP3KUPj1sU0yKE337PINPUY7RsPfudIb8/xWk
RIioRYShPAJ3GpuzdHi4g5HZIM/MZN7BOuit2ZBqAfBYqUTWXVCoG7A/qcsOzlyivfjQTHidTzS+
z4EPEAYxIFMlO/TxJnBeSNtnrNFQ9H1+NLTNxMb/v7/GHgbWq+rmlW5CKv9vcRcrN84n+3+vElC6
w31Ti1AoXh6GF0EcEDCU6JaD0CXuH935kxU/wZndzcQYeYOkDaahb6mqlqIYyvdK3OcKhiGXgwvg
/exc1ixoxB6U1iqzqq3X9O6Rnx3yK2M1RbZg04T4/IEJUhBhI0NrLcZJppLzQSPAiqt5S6i96K6J
4k22cmB8JStiCq+xkVk+2bJWfw1vHm6DJWFhzpdxs6bksnIK2QDNL//Ch+8DpAK2so2qptEnR+y4
t9wHr7FD6dQIMN/aXo0m7hO5JrS9rfJ7bdgTuiZbNHjk1LLOMCrfZJW20VmXuq36+ZuDBdd+xU05
zilI9OAz7RmGSk/PccmAJtAGY+gbaBIZrT+V4yMwd9rAtqLD3sb7RoZdMyaA+s8fcC04dD5UoZy3
aXmSzi3R8NaXLzmtttHmuyMaJH6yb58tzfhQi5B3Es4KQpGIAQgnmgMplBBvoidHgo0jbm5ILsBc
swE0+RYVGZtv9hEpNjZy2//Ey+/wiPv6o4uk473o5Rb+ZTIsn0C64PzIXYCjokCx2SM+N+FAdLVU
2V2S3cYV7pE1NOkFQhppJPcnZxLj4EKj0azVunwD1Y7XMiXWcNgA8FX+3YBIBLBD+rJ7UC6Ve6Bf
sTGjTBVCrecIxEI+ctCr3MitiaLfYsk2mfxpQ2LbMjKwMCh67L9+HPQYeOVMG45MqPCgsg4JmzdD
aMXP9E/94HBUw68PzGV0v+HduPO+UW48enroeLg7j5q6i/gVeV0ozApUW4og2wLH2lVhse4eO0hZ
nCi/i0k4xcobK8qddqmPRwq2YyfW33OqsR2vrTHNQyE5HvGgj2eeMD2z/EqE0sFEb8JZ2Q0zHNQs
Y48KLe9IAURd7oMOggmVqq17uLUNo1PjHgYxymV1d0bwKfPaUMg3ofDoqlPHpG2REgfbhuuRuqQq
QLYVFO1Ec3cg1bGlRgcdlB/djdTAqv4dw3R6BCGdILT1VPVL5hPsbWlL3/R6PlpHVnBjoBXx+8cy
XvdldwooknQY1itdoLyZGMZxj/dsYmF2QPVqdSKjm5jKx4oR3k4HSmIU8WSRsyUqBWHMt+b3ZrO6
DQYuIFxtQ0XxQO9Lfg8sCnA0oNrP35IuWWYkqelSvWQV6RQBtDOrqdvv2wJwIvFaz/lpc28l0KP8
csXBKe5dJdq1dFEBV8V43zHhGxN835LpTHtzB7WiW1xi9KiePOSMyhakmPSRINqBMy2IzguGyI9Y
hS9eL6U0qNVSHN48Q/+5BPEBixhGx9OdAwL+f5SHGcdilFq+QsSYD5UCM67ROYhIs+3d++CoQF6K
x15jVZlF9x4nC/rf04Z4pmOSOUr/kHYy+dEAk0DTKeYZsLTZLOiKTWImatszlYBdsSv47lfCijdS
zJf3KbU7j6OyNwamCN2daDYDW+hMafR5UhZskNIZFKD/2KEeHWh4IGZ9h6ZrRWoFVwNiZwsdRGxH
TDJlFdRuoa3sXClNlSbaYflawtsL5xohXKjJ7O7KQctJYyzLGXJP1ezx+v5ZQuoIHNjWwBM0T7NR
DVi0fhPfJ2gCH2fX1eGfaJoQjzUQ199YgOw9/7IZnRGrJCCnW6p/0vk5DY+w6q067SCXJS5KE8/n
NcOfjzBl/y2vqbcYPWBSgCW0ftw0ui1kxBJBgWzF3JHjg8AFjR4M+3WK1gqA/hwakLrmGOB7ocGg
v9Bwbeuy/C2JG4lKkBuN9sDFcn2lWhtOykyuKqi3E1GBYZtLsGSCMZAEx/coKItbPz2i90X6I5L2
Sl7w4Byi9Uj8USSIXWXJNYcEAoyJ1Vbx06eY8OIK/yUyI/lRUBpvNlLQ0h7IPLt88GI/QoVLfxgi
VlcPMgwBvMbZrCLy5QOwLlhQmh46PKN6brdIaRuK1c7f/ih5bMgPfmjXhmihCqgrlGV74ZMrgaui
AJOKq/QZI+PAeHE5+LI+ye+XNOa3kC7vqO5ZnEm+Hm5cAVGvgLQYXxcjYLTm0soj5+YRokI9yVo/
Uv9l+5IzYXMwZCbtjlFmOav7+42pl9eDLiZMY7tbMR4r8nZyAOA+Us0zo/G57J4BVl820KtgFODX
X2U2w3jwLfHcfAlrMtYh6HmI42WPNoTbbpCjPuGq7jdYcdcouXvzFoeNGVBGp0Bw+XpPjaWL9fEO
YBXKXg6m9CYBoVgl7sExb/HdwStmM9UhQtYiaS9XzR3uGneNPT51gy977xvB3V0lYZVauVVuElH/
dO6azZ2mkRev68WVA+hrXb1M8xLor/LTLnnkbzlk9609HSdcgQZBUfObNhPmar/uu+a1KoFJCVhT
3hiMwtQxruHT0mLgkdlA/rF4O5XTSCBs494ONjnTppvoVVSz72pH3fpaqhkpd7QThHgDEAqjALYo
81CmH94ZQAjiN5vFI9bF3DNYwGUIHlkGRvRMZdfNYMA141SqIF+hm8OHhqlhkMIqEr5Dn6MWRUoO
Ct7LbA9dZpJwNJiT75uQuMdMMvZAWpBkM49ljSOa51nTFQJaWOCjfcFltbNGc4gEloq7Dvl1AVX2
d9+q4LzzjQBTkEuDF47jJ9clqCxrsE/J4sNwZ1jsa9Lo0nemm3w5Ev1nPolHfsHURt+HcJqhFbUH
NA2r9COeyXIFXy7C2qNBJX9ae9pfyz+UyZAPl/lS0BLi0qyQ0EFV0EdMIeZOFxLSDaTGdSJKt3k7
yOhlvHIJwtN2qv9xgXnYy0nM5MW2txH5RWu2EDZlpX4xYDbaldhjSCbNtPplZI9HEW1ORcHvrwx7
CSktOIsXodmxxyFcCVsynva6NxxYTmHE+Anwq+591ocPdBW7Rq26culLMjrOAN66bAzI1IuF/b9p
SnmgoHP8WKRnwng+XSu2u0VIY9aW5XTXDYyQB31bBtWDjCWtT91asngQgUP/n3jpF/PHiDg66Uep
Ud+HreyftwlgeLsZWtDs2efzbumWT4CqUcpjHedx3HADtBc28hYf6usDw3TSMgTxllvI1XU/AlrC
AGO7CRcNxQKFnvC9VjCjIMCqMtR5XxfKJqYBXsujawkF4blT7YsHoUjggJkKwGIffRi/3eOqseS/
a/gq0UUqTlBLwcmgA96gUK502w+rv0JQlpvcAh6JXaGAwLcbIzABvjrvbzdYXgWzTgTndKEDSK2f
29wjqiWTFHAyejjoIA5COLexNRVHWkNR9ADqbWH6dHaF64ZRcEFAwYveMu2OI9OIB0xE2r4TmCU2
RTD3fS7ybJyoMRZ8WYFwhamsS6SNT8TrEuVlozgECtHLJ7SFHcpChoTiYyDECKH74jwrS1dMC3kn
FQGnrwb4ocEAKtvGnYLCGmrBcEph2LlyNKfVUVMswV38KJrxftMDk2Z0wIW/0qxwDtrxdAfoYxgE
kITSkoVcDsT0tVmBlQ+q75A86krutvJ1/XjqO59h9874nOy4bMrFBC9zGe46zckwZQi/0M25IQ3t
qmzwaF2+1Frak7XOisSbXi0rorzNgLKAKXZa5IGmODNAv2yUTwq8RhpuaeriLQkRFJCxiMT0oyTY
2j5gSPlBPcLa199leNsZaQIlZsOBO5R5GeLOEZl6xXFRC758K+y57PlghSMZWMdLkYJrPl6m76bX
q3xSiioCD2m/Mc2ZizVlEp7nXCIClXFbZJRxQqSJLk4z85bJAXclS+17xVSYW5QFLk5tJ3kzGuu0
5Fe7WiYoVtPi0wPFtqgrrXRcZGldR2ohZoo1WqHKMGplh4UI52/V8KbYQ+DXaXcNpXXiwQNvbzVw
1fte/pfKij7BPmUjs1wOumNCKtpeGrAzmMVCkmCw9uLIPf5doulWWwjgBKP74Xr9S0z/R/v04O8a
27X66LiNgXcNqS1QjCoL0UCHjPxyeQxVJP10njdKv5iiL4u3qIQS7N16CKqNWZGzyGjoNyZhntwm
xChM/Ap4TrbDweOZdMfvvwVwYR1rE8PEfdsV2YSP2qDsbji8VyBwuAMHMsuHw/5iJapRizztGRKf
9Nc7t3iRoMWxDKzUudb5DQfEPrH0EiOuByCdPP63lSKOtcwRJadF/kfAoQYQvTkVcy6yeJNiN4/l
QX9xoe5cWuJNTttLQBoIF4Pt+b/sbKytcz59DJd7TUw69FAAv6AHmrFBNzNcyXWSwOcVEO0BXz5A
2GNG1QB9DXvUscJoz5H1irD2BXSyzOwSNQCc/X7TPU7Hvef6feHDq1v8ljcU2mYybij1S+AtiQj3
TMnze5sPQUv5o+ni2NOyx6g0cS2Nt0QY28Qc/dtFtvjEBQtWjIn6tq1aryCclbjxVRXFkQSNP6h0
zOwNgdu8FF0VUR2VAEBi5Fe5V+n9L/YAQrDIEbJIRbSa0pOYmPUvUklMU+SYcZF/ia/OO8LajJfX
0vv+nUpKohueZEOJ6eRDwr1Er6v8Rp0VNLdl9tqH0M//PhkVtR+EIllJ0R/o3xgw96EfXC6zptbj
I4KqVeT0FayuRlMDNnhOyBJHpwsjRdkTH+J0wkjqCAWT3ZWiATxS7KuvCsl52E/QtTnteVwalVgm
mDJU7p0Kg13AtgjjcAYQfrYFA56fxkU0X2bE9A/tva5xOXe5wN207Zr8o8jB55glmFdND4otOff5
JSTO5w24JVj6HhOShDqb95/u0vCosEaonbr8wlZDSGQMmvSZPb0MhAbOpH7DyjffMqVBX+VE4PFh
Cs2GQBHd62E3GGO+q+JyU2tgXKAdnID6dcU2h91o7SVyLCLxGVz8N+oj6Om9gLe5g8Vr32N75Zo1
o+ZwpzNtin+w31dE0EstKbR7M4e13TA2ejr7gieTNRp5unhzWicnvYTVCWNfHXdGGkyYIlIkENCS
aYIxLkDFSmEdYN5EeBt/swsEtxCAkHt4/Ymo8AWUmmVrMN0ZvAwDepDfcEcYnGwnkpuqRims/ewA
Mnr3BqTn0rOJC3s08fmH/msgxIWDrrjm6FoQfhUh+AAzcpDAb2fnVW4SGRTFfXl1cfQlZXDfV88+
TCQfFvps2AitAV9b0Yre9awPtCZdFk18lf9xQs23p4YUtiV8B3QuML0b5dky1CDfT6SfvrVjM8RE
du4rzgXF/XxTYPXGrCSDsdc0YPEmO58vaE8/gPEnAOIFByJaa5caj1h4NGw2aa60TFQ57m4seD6g
vIZIACVvadZQPl3vHPPEiRXOWUxfgjUA+KufJzOes9g6a40PjD40lZqbmthnQjsvTm8n0bPq88/J
GFR/WLaL6sAeQ9yiVtD8w5No439QZFeGu1zCEy3oJ+aCqFk933BMJYspHwssE/Qw0e8PGvix9OZB
h9BLURqLwOE1ooa5PuaHWoNEdxh23fGziLmemG/Mxkif1MjpvkRv6Qs0hcnIP4TWyHHLAyQvWDho
RT1GjDzDL/rTNaR0t2h+gKJMdORIx5L71uDZ8loavCPi/Ug51hjbF3+PAIcs9dyXtTFL/HAzfFX3
ifDH+FAh4AecylGddbj8O36bnX7hMX9lZJ+bGUUrSO0IWlFBroKhMrlPKu+pheu1inUFEofuamiu
bxW7SINbVjhWsUhxx2RHZi1yYgNmm+pbqVRuyDLIerowITv8J6noSxb9dLaLIzODFYt1c/dFFJg6
SRy9njuxNARdIxmJnc6fyjWaLM/kGbkQ6t3PgNwHmxSuuICvxh00yWg4E9YaWH1NJflYbss/sYBW
JxaU2hTar0zEl6/gsVgbnt5gPo9RoooM+nIJlZ95VFBR3YEAlJ6AqTOh/lYpR4bkLKtLQDXmcWIP
9wDucLMweWoofoTAzoWqv2cjRzTsyoiQUkCiwsJ1EgzCK2IyNkKhsLyt7zemFOaRY/iPg5qpOFQB
iBoCNa6xwzAWLB8BZrVrUVHHQHEOi7o2ougxt9HyMTfL8o0fYzOLgWYMu7n7U0zIiBuqLmrLcJCV
jHIQgKLzS0YW8WH4m+vG+ClaJWJ4zVAebUwwIBBbR5VhUv2l7cqKz6KCkD/g1yOnEWQGiTSNWKiN
2Qc+llsifVl2oVBdnCjZb54kX+RwaWXX9Wq5s4IQzMkYvDWK7m+42W2M+fmWg1WADouh6OmmuYpW
w/2KM8ghOyKyDzTcU2oQBrm91RV8UtLNCx24dSWNbJ7JvHRaora/HYElzKmP4JfTEtnPBBHJ/pRx
hOhIrIW6XZ5e247XZS+kTOR2nDF/+ZelZ7HTPzFeWpvAuF3opLWpGqxGLz7Zg2SuFfznaiyclUA0
iOqUFe5TZ9Ws/7z40cuO/DG3Ll8rUfdPZ+kgcTvCWBQMgTVqKFYvEH5agltJ1SS8oh1c3dlCpnHn
cIBC6NscYDYCsz65fEy8O9R3r+hrxiD6hVZl+w20KDZwUAsB27Qs2z8ViORzc1RTK9s+WJAVurv2
0ELpTvSok2+81L0oPip1KhdnHEwZiM78G+Q6/TcvBE98liKPSjlsJBkkr9GKYr54+cMzKwcdS1Zj
CEz0w0GtZ5xWcws4XyPz47K0ci6OMEQV5R5UqqsHzI6JtC7uSGp88bMkiLlZv/v8PTwPlX45MfsR
2cSDo/boPk+wXj/RyXqO8EWkgOfTpIzzoQOV6+Fr5F3gQYfvJ7GCtpDh7prX5V1T5Api8K5G5iiA
Xgk70tuhTOm9q6io46vxcld8YlogTnr33PpFdhTf18tUlk+GM0MBr8ydkyDpU39zznNgRokmSO+q
EtinGuzFuKSxqYMaH9oyqDNFeVesTh9m5oJjreg2oI4Dff0oCBaKOjxj8ny0H3dGXPjkHiG9JUlE
CSbnp+rxdpK9G+nl2tf42BZF/i6f9Sax74dwUm0x6scGJv2DyAX6bxq/7rqUFX97BPFkt9L5TO6b
53U+4b7oO4XYSD/Am4aEwA5BUjJDOwe3noydRxbfCqzZX2R3/eBm+jr3pA6ZIkW9kRnBTff9964G
gy6twrY6YToozT22BIhakO5Xny52qgIySTN/lfE52qE0T/dCGtUS6tsLpX/C1FmbcjDkn6XHqCTg
tx3xcy+CmX4tbC7bXEc0LZg5KXIv7vyb9qM9UjaYhHNuTfdUlCIMzmiow5lbsbuaNkM/mdsePsC4
vvMNgMLzwKKL37FPbPj586atJDb2qVwK6Ir3h7H7fqdVJKiNA3G2aJnKr8QLSKlx3YbOlmcwEE9l
3GweNZ/Un1gtI/9Z2wPPvzUyWIL8RISZPt8mues27gxMzq2wWZb5WXaraFJDpvgr5uOVEBxPDGV2
fsTOwf1D1ru4DTqPCFWd5Ja7K1U0mWWWt2aacgWWmGrFfBWp69eZaJLtD3U1uYMe549fw5wJIcRU
WRdRZsdAY2Iaz3DX3QFXvONVord+FfhsDhX/a/zpJcT9pUhF4M9nL9kDXz91XM/Z1wHCHAcgedxX
sqNsMzW8EEFGRN1m6OtE4e4RY0eCoksDdeU9y3ARBhZPHm8Xuv3On2tMMqS7wEF5IEuSQG2n7cIA
421TKoGpku2tBp7xlo0nKBiitQHsebzx2U3TqDQBsTZxQR7YfGdGQgkpjs/d3RZFcG4AHHDxZCCr
AhQO8fkDO3o08vPSNnuq8fCuEFwT9XBXX5GaO5ZzrF39+M+PMRWX+P3eJN6nQXrJIhyucT42SNYD
ClOFVNKeTRDw59n+SFN3se4a19pFKbqVxwomVSzE8hZQys5tAEsQ/BkR8EqBAvS7S67C24ONsuNX
CLl4beCoZVMzPIi4d3HcZ9Kyv6BPSYU/31hzhgf4rA6wqdu5KkJQCzGEqQo6oAkkr6lW6Gj4F6xT
kvQz+F2i2SZSZTHSQAj5O2zeW4+Dl2AMWyTJf8kxZrLdu0bP3qC931SR1aFVe8B8YoW4wgDSHzml
n7JlnGs54i1l75vJoZ1oyl2fqdG4nn1E1K9E0ChuQZ4ziRHB36J/DWGA1WUmWB4arBQs0Eh93RHF
Cu0qE1d2eKSlBtRUuNzRnNhPYN3AQ9PRPAh+/S6MTJsStYRk21ChTiCsK2JzHpVDEKpIfmj9zDhE
SzI//mnpnBER7V4NoQLVIeJgWxXyhFsxE8fGlwzjOXEt9HYP2R8nhmWQ2A7oZ4icVknSjKjyRnx6
t1ZPiUw5mOgVpcLLDi0RtNIGVZjSK6jP1br9GOXxORtmPyuQoEsaN5Kb+2Vj2a9lIIcgydERLgCL
jC7ty3jlSfeUaY1zrnV4uiRcwLWXItIi631JKTNFiDSZ2mqA1FsV1SSVR3+MyMi9O+YBiDZPlZPM
gUkLAaqr+d5yWHJl1j4Cd/Bc1Sy2Iwn/HdISgOfTvIBoaWgVah/BGg3mlUiMqPrwEE1SM3cksoO7
MI1y697GqaTK1pvjkQtc7d2zuKbt/WFv1SYZENPLHgtsYkx3ly1Wu4OoPiIMyjPcVOKjD368tVKL
CG996VKh0N0D2Br5uXmartLkcJchFN8rHQRvHs3EXqtQP61kSBDymf/E1Hb1bx6f2KrUXsJlUy4x
k5AwRUyT47qHqo0qnZSqO8JRo9FnrUrUMrpSHAVqigX20Hn75B9QG2al5p9XV/nXC3slA5ZCxYVQ
UutuA8PCyTT0Qp2kK0rGP7dOhRAAvF+RbAwbq+/LfRm0IfnDUlv9GBCNgRV6t4k6iC0Vz3mPeWIr
0k2NIxvbHIDVimWiA44XC/ocbpJtp+0+IVAzzktQSEJO/aGMGS8T/Upvdmgi83p5NhPz3cDESauP
GrUNQ16sIxXm3bMEJYVnR3OCg1Biw5HXSe3SB/T2bTwmxxH8JIrEb2FIW5mIC/FHeXxAtwMFAn92
9M6HogLuylJoWyGBv/pO3CX50UFYK1tzCFAwf8fA42AjwDHb35yTR6EuED28WlaxCbb3RwdWY19H
0ewIV1tJBZhPueZr6bixWpbOSh/+zEfwvR3ey+8UQf9+pg2l2s7AruNCJxekniU8oOfQYGe3GrdJ
g25gdMr4O+Eawj72ouwBW+pnWBR/Cl20JRmQvGnzbkE1x2oXjtPW43Vjlmxpjd64LIFcfjCzKJ0C
K/IGBfYixwNTQxo1AzViepckMPx02SQenHJFfkxsQNcc8CzxcPUHzx6jcciImBDbjDbPqOC6Yckw
NPmniCUTJEvaGr72GZu0/TgBlYRaQ3Jz2Dr5jMgtlh+BRE+SbLId4L75dQfcS63Inv4UWtdFl4DP
UUgVbZQoHeYdK4NfDDDdK6r0WKOoyTkgJmMNUpLlmZHsbucsTTxuTUkVZTuTDUwde2WudTTdA6kw
DiNOe7pR6n6FvmfZNdCsXeaYZjAXjOa9eiBhaLlk1OwZTdzEG1Ar45u5zReZAElmxuNXgt2OLND1
m0Yy+ouQLskhvEN5Im/AomFChk1V+ga7Rc0ZlsE1gM6adLoRnpKy/cl/WpaEB8I2zGUXjndEmJ6J
dwx1WCGd4na1wyIb+FyXmB1VSmwSQeItBwuYaSgxRZUJca2AQc7jhsYUWLSfQTIrxwKW/34Dm/st
cRZdmxQKAZDcBBcNinMazFp1CAxPbHQMkmoJTrWVaDvPeOrTbU8uxflKKRvBgqPwWHfBeGm/XtrE
cUS4YxgmImrVXrICI006TONwpfh3Lacwqvatvo1dfz9ioG5EKqrINAgFf9GpmGZzdwWYqUbdDfaL
YJk7oXkg1CGhHJbcmjM9qyh6GDrPttg+JGCnQybjxpRCoPdiCDibwkex8AEENyPbhjQwgtarYTHw
E6fWgaAp+48bZQG/Xa6XPAqb27Fy5v71ozq2B5mhvXsP2tL9yFQnvueJ2VU+oqwEPq9SWK8Hfg9h
LHBL7G3bqed3d5FWcM7jphuhuXtqAUoTAmaSnrZrrrISqGT6MqAZf6Axog9wrX0Ww+PsC95nmLyg
sJy+vj0BOZlwmI+qAXGnMVHLdz7+/8DUrLLoiRQ2ZHQz/4sKLIVocZ5zbNir840d08PhTO2fKI5R
PhMOLf46mzXZ5ApDlopEgzuhOWeU/Iy2IObx8+E+Ogb2XDBhrnTd/Mr0mVWviTRU00TEU3iu+0uO
oM7oRdiCS8Kohi2bmEpJAVnXoUTxzJAeS+oRCFh+mMrtvxdK/rZCOeTD//IdhkTzlRxCKwpXbrqk
3lfkOEhyuPJGojDrdufUCxLnjt2Kggi9rC745lHTikFVloI08w+iIMkR0lvnGJVJsAdUYfCGwFfB
lZnm9+h1CGs2l53vh7cEoDOD3R+xgudZdm3mXhJGQazMHXBjr5UQH55UMYdr/fcpdFo5SUMkjMcA
9a3X9Tufyx9U1aNIb85baxHH//QHICMZuhcTpYDEo2WyJZrYUxFq8nS1oRdprS+abcxv3QliK4X2
B/LdbEe2ysMimXQcg4MtcarDxAYfLx/iWzbdw0sd7dlw+y1ZlU+JN/BIy4A/1eGQEXzJl2Kc2sl3
bq4UnkvMpI5iYFqWeqeAxmn1BO+iwtfzsvhxQ1p4U/7w3RFl/xd21Dffv74Yy+BahRiHYLKfStih
cjcfL2kA+P9fLN/7ciEEA6J0vQca6m6u40pyk3HXer9yMqN8ijGOqObdva4gP0ZONt1KIjZ2X1JK
Wt27NsEF52IA2AXKbUf8V0pTyYcLbvtjHp2VtMyjS76EENG337eQMYif9+qN+KHtLxiVEyaiJVdH
6GElmBOdhebznKLd/dsi6dAfQFRtUALQPHeWHIeFsX4xS588euOgY0sMhwWKhyuycG4ERXjif1Vl
cKAjK5Kd+HZ8SQHHnqb6LJ62N9l/XruL8yfYLLRZCI13PbWSJ81S1ehJgnnI1Tc5gIGu24hQuyy3
T85vZ9YI4ZsD5txqA5rF3RkoyusH/OfRxcqtbZIznb7LoS+5mflAzmf0453VIQwEz/3LBL2xKO3Y
HC+DbfN8tM0aX7o0HFssppv7ZB+CICi4P2wJMKngSJ6YXEdvUK5lIpnYt8fLCgxxJLx3gymdVphy
meyGwULP2fR+GhR93Tt8+fx37CDgoOdNwK9ExKvSmMWO8NOIK2zMnIKqqR/+YnL5gYrjQ5g+ATTA
DzHpsPAGDDMLsA8EPqfgLumfyd5vyCAIkEQMKXvHqfEEEL+r7j62AnmmimxZ4as7liLVXN53yM/g
CcQRdYTd6suUqyNF0aF6eBsE6vBRUu1JDPK/5E0Bpks/5ABPKdzHOmhLk4htYL1SLTFyzygrzJhB
tEZMeWxQvkF1wTRs+XVXFrXGhU6gR66NBK3tx6TD+FGYn8ERxqpmS7QmygBFJBFerrO8IkOs4svQ
TmG0HB4okE52LO2cMeuayPU4y5FwolLUMUoTeCvlepPA1WVAYClGrV+WmqOoAQsHN50Ph1BPpGp2
H0ptdY6GpJkXuV7JDci7nqwq1XnG3b41ycbCo+vwhc8NuQbZWKIQpBtWbbETRIh1Bn24JgZQ+Y55
azPrwfhE3hKSCw/uArAhUuiwrLdsNSNul01NtGqLVkzSwyVlc10mqaywv+4vWxNhbloF+x5VGUyt
k//N7rPGB/enJB9y74cDWtKapCNPTelRrPON3uZDaTe/P9qb7fLfCrVzCqZ9peJ4C9sq9U2iabs6
uNMOxN3nqKcDgu/l0e6Le6zpAs3evpcJ+qiwcQjqg6prulEtGC45A/Uj/WH+xpK4jCqbeRb6c2r8
FPfHirQvg2q+7dqeEbpNXB8xDa0vd1ghlz6/uMMAIU/OEzn2yeDm3bqlvnepx0V6vbLCtJOsrIJ7
+SJGvGWL4XYtnH2Rd//tRwkkoONetiPrAdwcGAxxoc1L9cqRJ1Hz0DUbw0Tc2mF6LFOBmE3K1iUu
lGl4Ic3v5A9cGOIBBYgty+qq7BuwXlunGJ5tXSr4rrrhYVi09UH/uaeV9NjAbFPjKmlgbFWCGB0a
TMtniHOZVPJwg/kjsMBtHfaQOvkIDj+0EauTxehTKSyy8QT1cNr2Tqfcz6G7eq1+90KqKmf1C6sg
nVQKVbxv5yE4+KgAc9A9jBcBFkZr7kojPnX0sR+8geDWtnrb4huEPe4/n9cflYFxyLIqxMp4mshu
h+oISCbzzBAwGFT5k3j4qeMU6bOqkZvRWt/JXnk1jJnKPAtLvyYpKF6p+vf4vfPeP/squuxlrLyQ
0NryASP74gQTX6GgAfV0gxxkA3GO9aVU+WulOfF01aVhaTWa7yecdvmtbloDz/RbI0h97SYrWwpY
bWfQryTaxgDJenev5VYbeR2G468e25+2cW0MqiPod72e1URhXBZBM5p39bWXpvCwHi3xJQNZKtRx
RQxh+jsUEKnwcCBGp6mkKYigQPQzDRGsTldZZBICPpWpqXURn8DHrqp/yCpeO+JSEJQK1vD9ozxM
U2edNnugV7nHIHN/XJTzcKM/XjSfAwlt5j2Ep86lVQ5fdCBU1xd43p9g3Hl7G85sR7ANMhtMJ8M4
1i6CCJzePOPDNR2tOz3uUnJP2Xx6lHo6HNLwJGIpYPxjz45Xj5+4u766kDoC0JfmRkazwPN8X/sK
yWPEnjjt2KWqNEMwhuXOLriNpJWGN594225HHG2r73HBC5Rj639xqmjOCRSEqJVbiM2HcKy95RFl
FrVQR8nqTYQD+CnhnSlQjnT95kbuHEpaLSChL7gVzkt7XTFhXy3zFZzxu7qrtc8cki1tq23xweMe
djJZeQvyarIizn6Xwt7F6qsufWUlCFKBORzroXbIWiTzeIESJOBAlrUxtMhYTGxy5yi0zlPvcJEe
w4YMlmbd2g5m/W+fO7Y8AbSyg9toD0Zrx1UdPqrCTI2KwTD4fuDDQxKFC/RALU0DGS1Wh8FGI7jv
c0xRTxaelWQZKTYfzf7E4Nmzx+pxSyegAPTefuOQhEzD0ZP3EPDk28jQKQ5uZVeG8dU8s52Ma3dW
fmns71yNnl7GxBzFS7XjebrYAUYapMjUUERPkFqXCGYQSUqMkDDQVihIM2rn8MvyHv/+pGZuXJf9
cfFmBGnLPnxtEPZ4lxK2runvHRVq4Z9upiddphIRXAihU/yutmJwBbLViU1QMuV9oWGe80JxakFL
yLuaKWC+vuf5Vl+fO/vYs5DH4jV3P9Womq5+WgKCxsh+9OfWFKln9lzkn60rqbvVHYE+yR5YiyUA
0ncfYfnNZwRzjP+HC2BJmJjdtYIw04F4Nq9F7xeGzR9vBrhXegYzH3aaP8Bl7H9fCq6n0OUUgbEg
QSEmivbk8zkAEjnPaVSpF9d5L+0ix+IymeSAeW+UxHLpHaxIFruJvpgTxVPCksIjDrTvfkI8pgKJ
aJvJGuNa0JyA/VSNYfGOTWS/fygjWzYJLodT1JjjE7QWnIvgNBmOaWPwd3zHuSrh16EkEY63JeAh
iGiupE29Y1ZLl9i1BzX+8XbAreUwJWSGARMazKlOTGxRJzip/GQLRZhyfJywO0Mbkmnsmbx2GL32
oPah+ayYtBPfU/nM+gpgcWpCLxYCOcPoxNGS4wz9TjCVAwKa9dbuuK/5E1RS/Sjif0kmohPlf5NN
7C3esSEmOPbNGuZh9jiaSi0D+PEdbg8slVO9OQAoMIQYc7qAIHa4RuVBS6BD5d4Yd6aKTx51m+S/
r7ocYdOTJ97c8UtmdrfYgUu9ialBjhTHQZgdYXZICp2Ei/a5CiaH9lKxJ1+xW5hoGnrjRlwe75jM
IM0/1hZPVglzfc5/N5iMGTIrOTLFNDYoE5rW1nIwaOoCExQDMkOdgwK4y+s0AVl6rU9WXegtHUot
5w6eAbuSfaMzpkUFNdTSoiz4swWxDDz/0QtxuM0oQQawHWTv0KIndbI3BdXGZu2YT4sTWxsL509u
lQm9w1ivU5xPFPJ6ol/dmD/VIsffUcsH7KU5cd9K43/u5BtL99cRoFWrrWzAhUnlZGwEeGgwlHgw
CCD5NHD722mTK/LgGnlJDqoR3vydS+mygdSTU+iw2nogheChBjjhtHKfqYzp75XFwIr0rxiyM6vi
LmGLQ2UXZw0UUxD73nWTW+/JlhV1BF0UphJSOP0Myt/Uv5v/m9u5iHkv7Yo/weCiLMPWVOYLK+9q
BUg8rVH0zqNyQWKus1LB8C34bm50LHT58RPiJeAysUsAcWhmpN+LWj54n9P1t7rEknNcOAYaHF5b
L7701eEt0LGzE++HTMh2n4s7rVAxH+5FQJYfL3T0JJ8d54p0agjuFBi0uErlm/ypc1af5l0GklBZ
Ce0R72ER7QaWuiY6iYmi9+xyqtxHcJWqj5vs8X18d0AwIneqmZQeIv+V3HVuZMBCbeemNoQ+1VJk
4PewqUxLwo1wYfxiz412/19gwNL/9wVTuXCw7QmJe2Wxdaog3OcyKSUENvvODxuR4LfgQxhrpJKJ
taVMmxRJfBtB6cdCa/1BNhm0qrI3qIx9J7oLLQ1qIHbwNNIXieFZidlvoc1XqM+nNp5RGs4ms610
g3+46n31ZTW209mrk6R8YjseTpQdJ5Sgb9MKHZ7Ftfps90vDb/jjzfjLqbSiU1TVE/FhGkTRc70C
SyAjhcINREW0Fj+ljyeiotoZ59VLv2VWsurUleq5ekzyRCha57gGzzQwPraLdxi0wL4Jq7rFNmss
Lqr8BCHkFwmrqw16c7UoRAQ2yJje9uVmQkktiBUjAV/PcJK7M0Q6WJr0EC50zckc9cb1WR72aD5y
EojQhVbmauFaZdsKySI+QeAj8tFgxyz/DOci5KcEfIGHya1FhExDrob1tyIvWnFQTM891dKStjt9
tc6hpOre5sewfOJu+hL8xuzz2sWa1qvYZaLTM1g4KdSG74waXZ0XL3WndRXlqvfH50s2sy/PGb1O
4MbXPh1ZtV7ZQPOuQoy7stJ1Y5FvQk1c4jx1eixxKoOj+XjW2VuyLkhXmOmK4Olej755mxPMARlj
grq4IyZLebr6dg1ld5q3ixf0ltYw+JPjKCJdIMvAlLFyWAMYqMxJeeSSFa9w/XDu8T+Gi4c7tEUd
kZsatR377APQYjsTwYunqrZgzm3geV48XjzYOGGtKQEjUPLjNCboJQTTkedlq1efRo44OlGRy8bv
kCAKABVsWUIVrFUTsKVchhnn1vmMYbFBfjGfIzaFmPEImv1gmBifby2VYkLhRWl75rpOnuK/Vovs
5obIy3csusJygSsKsw9y3sVSw3Tih0R849K6iPUny5jsSv8Kkp9WH18CryFpa2XLzKM3VVp4bVBd
33bRL6rBeRuDipjwim7lD/4bDHS+h0e4t673agYf26SqGZwcXRjlekqS71mDXzCDqFFHFBe4ybn4
4LVuAWtTKNi8AznjJyldEd+OVuSDVpEdLTkQcROB0D/4XeqloJPuMGbbZ0BF0Sgrum1CLkWp65Wv
hhaQFoWLyLLWLk154sd1P0GkK9Y1p0cZhbcvDVJ6g6q3l4D+RtQEnDR/RRONvPil0S8M7SeoaF6K
csDA38Y5aoqSItCd+If5emnk62TgujguL23RtpSaJHrA6shKSs3QNbS4u7iG9App7z1ZnZDx50IJ
JsO2Vw6Xj/EK+HeakLd7SiH6j+8YNJIdRWRpYS+2o7pjolS3kGNoEaNhVZOMu6bNLGuEzWTfSYHV
Sv/b3ivoILQKtA+DODjPCAD8r7zlZmTn4usnFCLwlr/6Q19nnc7GwTjWNlccTiqCUGecN2lcR/k0
Y6lA5YBBK4l4hNjrSSaXX5ZhUZgUNxo3b4jnpUyeTUeYFPmQOmXz2hChZlbtg849mMr9SueuobvN
/pBuV9UdWAjz9JUnWrhJa2d0igSpk7aYB0NTW7KY+nIniCZeIkjrdM65CCRYRH+q6WuCbqe02L8N
nkRzTsoU1dnRR9dm6u35mFaPce1wH+51lo8qQgPbthkEAm/sk5sorXi5zDDecpH1LyBMaDRHIJ/4
m69iYUEgJylH3djHuiJtrX1yPZCmrzDX4UGOYsgeldXapw07kejA8F8UxsffweorK5qQxmS5mQK9
ycXd1E991cAbOOedsW+QCVCkmkXJwgY8bXlWnF5yIdtENwG6o5x65hq68YQQ18Kb13K20+O1cdLt
h01MmLfyfg9pwrjDKlcot3hjDT9t10S5obKKFzpTtCda0tjjkzRnk3bmf0lo7Cur+PjdnIVbEs/8
eu99G1GoD1kdkd40AFxjkk0iOkBqXnzP/N0SKPHQju17ijyBmJ4dtLXpIi7C6iZ55mL2jhPs5p+r
srp9rAEZH56rmpw4gtNEnmrZdS9q26N/E6X2IPhPAYwdSNYEIE2UaFhi3Fh4fC3peletFM3bBkLl
TMerAcK5X1QVbEpTDBsPA5WQb+cWdzoTcuR+xNAm7xClKMhOukz3fhX8Le+9uy6mVzu66fJpLbdL
xruUo3dcY/dZGcGx9RvTY+3OymyHwNoweY0zCvOMnA/R8LNNR4EXxV3H6NXYk5H7I40OiiIQIBbA
h7yMcG+XQy7sunpjX9O0O76YjUpFJP4tSOm1xOnfF8RoqY3SODdKlwxnzCMJ/hR559UcIKKBD2W/
McADkOH3X+adtPGEChjIlVj+Ir31USSJifxgJhMHVk6u1nOx0OuIpaERKFAFpP1OWTc3YJQ7wxwh
22TCVHx5MC0TICM5y2KpFXYUp5v1feaRLuCD+8dC0x/wrd8h9p2+Pt4A/uRcGUQgNa/6Gb3rKpEJ
KWu8LyRUBNSJZqVbCnPH3ClrfNMF7KXl5vTdD7X3MsPyXQzCDllutE3FM0gl7ff93fRS91GEN52z
EblpnFI2xUAdFXpiQ9mO+fPRJv/YcNiGXrJ081sK8Px9DcAFAaj2xxdNGdqpRRfIYJoTlCBY/Oo7
Gio+3tegM+JAlPmc5juADaIjSkExFMnbeCG4n0b3aauaLDWxY2bJfxeiKIKQV4lD46OtFAJd7oQ5
B/+l6ClCwSXjyWGlxN+gNsSZvLs7QV7Bc2R8FpN/XdPr1hw4vH9fe13+aP++lXdFmu2OvBVmE31x
zTnLE77JKMVNfkoEVFSViYFmw8D1hjD+KQUx1/jOv8AxZCcvR1bUGn5DpGC9GsTBDMGVo2XsmBVP
QzzVeE71lpd6aV4i9zTfSWMxvI96TWSLyvzDY75lvzQUw89GkFFhhHfY69bxVDHe7c6SA1xuRTR3
yuLsTKRdm8NP+pSrrA+hMUwm3H6M4RSJ3707N53ZCdGrsuytzgKEOkioFiUEOAYwuCnvZEwFg6Li
0Knxt5/KcPquq/HM4uCqqLGnCmEyFJXkrX8CtR6jlnqjlYnly8XBlzW1pFcrRk7o+43yf0hz2lps
PcrthnT7r9OReTB0+4lX8mG7/1sIHnM7H8iDcchFZQTKpIgrfiozQfl72diIpvlp92Bnrt6MpjV+
/h0ZzGBGwIcpxqvGFCkf3VxgFBhNVgQIyPg/C7HIkHw/AVyS7vK+IKNSFp7mG6Cq//5bQ4QC/EU4
Dym77dj5b9gyme8hiecNbDsNwE+HWzaISmuTtxLqtogC7XlH66y6EQlDtuxS4ScDekjWms/cXo+r
YsJ8CZ1vRsU9ch3r5eQ+RIbR1QtuVV80Q+coPxW4IqaoZKyXABQMgkmKVuDUuifpyHjaZh3mLHBm
S+g2cxUltqkto4Fo6lPPIR98A5kGPCjNZwbhTOzwChQIs6wXyxHW4ynmIv1G6DXhT+OdD+Jojiag
T4BbRR7hrv3vq9JHmhKJbW4byECm4fgZ4EGMIiUZZU5XqeOBiyBMihwK3pSxGvOMkAq2lLweUBd5
ZXpm7aM0OTQpeZ+35mqrT03yKD9QVs/6w1FSlvit4W1yghAknDYrch8KcjoTWX2i287zFRuWtFyT
NCGXdR6tEGm8HniFdf0wiP5Fiq85AyfjK2n/loUlK46A4iata+CfFEF01UF2B5tDBObRCW1djx85
l9qCOIM6AojMaqXCIZOvN7kssKz0YwKhIy4R9bJ82wblpYD3sQUCwQChxHXyrWsfgPAAKqr6Fhhq
dFoFT/T9y0sJ1czmmv/eNEYrjsczcWieMArmwQ6XGgrFSJmsQPQGc2/Yc0hGaXuyNcZL0kenyieP
jOilcQGsMkLsro6Kw7ABs0zDhX8Uc7ZitTFcmtfBiX+soEPnjAETsREnQhAJKHb9HYKMY0v7gfZn
o1iF2O6V3YluyjvmKymUfi9f/BN1y3G94MXO8zIcHRRiBJPwKrDyPWT9rnq6HBtdMVYnnr0+k0jR
Tnz3rbszwXHru9RirCWjYvkgFUACBm9GMbXKI2h+nY//Nv0V+XzdCb/V4yKQrM51xgpzs/HS/jID
ok8EA7WX1dETQcxtJVBuOj/Pyrodg7hjY8FsHb+EkAUXkkDaX/PFedBggKiM+I/L5yMbx4XwJppB
Og10hZtK91VLp3nSjV0ReeiAMRa6p46CmZw8d900WHtysaof3rxVkAejkzBQBI6zFa9SLAZtSDa5
CLKYO9pDQ9ydpJgo6HND7sUYBdCrAmvus3oroEgy2gbu+UzTjTYixqtIH1exrXPGObIciUujfEaa
NExTkZ9tJeolFrdsG9vGgomhqEbCxgdOZ+JUbAcNaWPNGsM2G+N64U0x7IFGrPtZo8bgFLcyoXhX
DUyQ8StvhnJGwqTI7NKLrKzuTcgC7MDBCuIrYo0jyCLdX02EnCCxR3oRweaNs0khDeijF5aNVGRb
zdL+iJBAvj6hKFDEhQAog/oBkHIt4NJ006GRFqaVQvSH7+bi5c3gbn/R/uv2FzlSVoOTb8muASjs
oK5cx5BD7kQcY2VOPAoLQnQHxFJhOFs0Q62XYiLMYf1GKtJqvumLBAAj8Y+lxt5y1JNLAKXVpjWY
hyqNnVPnMm3F9nMyPieCSlUbLvA85KNRLmD0Vhk8DV/pQuD/z+X6bMzG4leywZwNWWm2BMvMFVJ7
t/Q8/458sYFk0ePjO2tnH6T53pQc9/zyrbj6qpLP8Iekfiz4/Edr9suRNqhof/E/py44WZoRx86s
sKP1io/9GodCfL1CBAMMHr8bvRcSsMxe6Iac9l2ttBBSPyFWlddYTrlPLoIsOcx+A7wzeqZmo/2B
r7q+BGShE8x5SV6jQ5aPjVNrJTF+iqp2dE07T8y4+/niAe59DwLliiNkAHOPr/HBMw9dkyM5B6AF
3bnAC7aalLASsnzWPch8gAy/l9H80QAWTXZtGdxynBqzcLK8V1GwsA1+xHlIBCwwwbMbq1b6H3/j
FjZjsIGUiSYW/1tvw4w+I6Hr6voZzrxBmraylEbtqzxwR7Ww3NTIsFGgmWi2fMiyslUKvkdGp6bo
mnQzJfZXoISbv0c7zUuAj6J98+MbhvSYikqNmd/mmYIJysZh96279gU2xpflX+XJ7jEdRV4pwBqt
F57OSGrwyttoQ9zVCale8pHtQ4BZosCObPPkZQlIKxiYetSldRvvZmx8XyKNVG08CVATBIFnGxVA
VXHvRYyf4+6wwgxFD9nHAnf/BApxs75LoisfDTYPk3qetoxzGp8ihWMQcw2w74xoBMqVZEE+XUe8
a79iitjEPlGsf3ALbCnmKZZ/u1PEXiH3Bg6oaureuxAu494LDu8pqzVT/91IvmThR8d3c25qtwb5
uTelU+HexGPhBqYhZbr1rtvIBU4yBbVre6II7OYMCk1sMRHQ66OhfyoUFHtzyP8ZwEVKmvrErVMO
dVGQJ4gMmn8OZQEIwqHekOo++mcTXWP3w38bLrgI3AWpJkpkieDIX5zU4bvKbulQttuldHqijAzD
+ZmxWAxf7WE8VjUFYg8uRJW7A+iV2tHIhT5yhvIvUyrvjL8171Y/Z8cIQ6NghCuUppTTX5HpEp4y
ORPk+k08t9Gh67H+TngRryqucWrBypKzZgnmYsU1jtB7//MwUg8UMgPf9jSJYS1/qI4AaraiJDMA
+basrYRumFEvgcojTugwO1MZKUWHvaudNlv2QoiTqEBFgMURQtP9Rw10ALnmXC7UrF9p/ljbbd29
puu8rNEkgFrUCIqOO7iSldJ+r+IhVgZ+Oq9GJOkDW+oJKTmz/ouxAO19INPW+lh67iKfLfFJ21rF
srzgsyKbqd38SUfUIarHzYZNX+ge7qdl//rIpEh3KpCaXrek23niOfpmEx9wccvznesKGYoFCzaa
TV59uu/MDQJTlSgeSSvT2SdYIMqELkELLdzNI4flWpNQFIcbBl4RcsyAqTQ2PPUhMKGgV8UtnKBM
x8zb7x2labPGdtJu0bDsm25zYElx5Wr8XDlYLAiHtxAhQrMtBM1eMo0W/X15qt9lxar0aIjeQ/eW
LWrStpEIjnYGiahe7VOar+5iLIhXT+fz90YoQhOdU2AzUFC+7GUY41FXsEO2aPfJqECep+vbq6G9
z7qqGxjU96vGJFshXmQQ+gL4QT3FpOCmxUuvJggecaezTCAjcmLfyxbkCmgoHdVuqMZZ8svLdRhU
PY6e8uIstOJ56AT/Ld4N0A084S0pldv4wIFXo8y9wEfcaCVE6yA9YL5gVRFApMvVS3mrYBm91ycG
XruLKoZtQTkDOfRlatwE+Iivk1C8CFqyp2pGx9uNlCKbB0FKSnGp0lpzK3y6Y+WruftZaEgSG7mD
FJoEPlEOTSHTkUXcRot7m0BXuFeOzx0MHqLPyKKHvKOJoIoFkkpfYdOK2lk81aX6ldJL2SqYKfDP
wsnrYsR77yN2auXLIuYauDy9CG3uCEZ8psXURucd53n8sQ8kpSiwXFiRZzlB1/Scki75A8wtQ8Xf
ZAb0/SUvEmmMWdeSFZCpr7kWEAX9+bORaxFK3pBFQFqR4V9Ht5OnLGwy52Am7KOr01A0padB/s86
RFmdXTEqByeJLieY1X/MqGAjkB5UZymicvzb9nuu4oHKWxcx0OiQxufB3z0jY7v6TiRbtT4OfBDc
tlTk4L24VvpxR3VuhVRoLwyUwQffN4lsta5dgKMXrYOP9NDjldHuPjQX1Er1IVQ0ZacfR9bcpFxJ
S75e6QWDidchSkfB8EY/CFc7DQbyQDldVI5j35QwJWCPp/VyalEZ/HwbAAXMivCLt2zdTDH/i91a
SiByDlwUsw6w/jr7VquyKJwPqJ67NDLOqc/DCDa6j/xdbtg7Fa73CkN1FrWoU3ld7W40qaadQmoE
EHgSPmrS6BTYukjtpa+Ih52mS9lqvGhSw/z/SM+ytTk6M01ALIL/MEgPCuq53K+d2e+ygeAbU+uv
oYSIAsaUKCuOdAnLLC6oSNK68RcRf2q5LE2IfuYJQMsO4epYBq/06JxxRYYdSviboWkP1flHecO+
dkaVCKsb9Mfw523lQp/rSsDzxIOf6eeM4qXT0n+qmf5nE9CBW366YvIfkMTJqx7EvXbBRj6w3jgX
+73HSpPX52A1ImOiM3VMl5g4u1rKSwuIJFIqEquwBKeqZA2qSKqRBPMKD5sd9mX7hk2wQzeSNp3Z
2+8uMng7PEw6YuTAjm2iFJmwvhQtk54gZ+D493CaYVoL5ow4boxttziQ2wnpwd/dOXcPszo95Lis
k4Oi5Mc8HJxg0WLyITEyp+JezO4abdZFHoFqsldTjTc5VXEvAOGZixqfRUZRz7GZsEe7RLZG1tKm
Jro+6AhkpoHTOSB8aY6HqArGJ2fUO8/aKuWhzBIuR8P0gLqiagdxXLJvRo+YJPkVmk+/ae5cPZdq
KtHjI0vQune+wd+jjLgg/K5ud/loyuGqtF60aTV9/8r4H+UYOetpRGkZLnq3ewtK29vWTSiw55SO
lcizrva+d7UQdhXiYIk1Sg0iPGETCOY+Tp5wapftlRmIyZiiYENocTV3m0Vq5Nq+DYJC15e6Liy/
wBgqhAbMSTFdpxyVfFqN6aHvleTm9LYFGeb77jf9AG9ROZGFm09PDMRDCy5NZs6cZtfZo+5UClIW
TyLJiHzGsjFL0oDdGBCLTVLlaMIBfCgVtKF4JfbupIwY+vVuy3v/qGFOZKfyugbuxqXyT0VH7eHI
FHqqWa6m0J6hKIpI1aKayDfwRshOxY7/6cZ0NwUZdtKzat5otkqJOnsIJ27IV1amQMvjEbznxV0B
1W0TFs0QkFQkkByNMXpAJMm6/NqO8eI3ZvMGWSsJb5lvA7n2IOt9lhnV8dspZO0cG9W4YeiOXegt
w0nk+/2vnf4Uvd7TTTtKswiRSbdkfTXvbPneZZHQoPBRkLvL9oLBWR4x9OWKFnoLVyI9tokAu3mF
FCfQJCk1XVZstxAQBPcfBbckSMV1K2PUBIJwprhwFuFcLPqDU4EdaPif0kxsd3jHSzHIbQRfeG/1
kL12LGun4NGFvZ98xGj902jVZh4+hk0Ph5aL2rb6Hg8pXZqbbGHrNH0VqJYwUG0rkTzXg36s46c0
VFWRAnyD8OioOQokkQC3AROJ+kiDRQ8ff8xhB2jkaQAsdQv65vSdIW4eozlc2IyuUy5r4/H4vksM
rdJ8Nd2Z8VvhCrT93EABmh57D+ABHVMNoKtvsWCtTwMJq+gyZYa7ead2w4CVOv7fh+nHBqmjCZjU
hXiUq2x9pzmnjuSAreO9LddwKx1XBlALPunguAsbkYIL3geeY0sn5SHOYx37p2GRnKE4XLEFdTaa
I7H5jMneCq/r5X6oJsaykvgJtO8Ry/EdbFSM5kfFQgB9qZ60cq3iBDDI+vgPQquwsBCdx7W8oSYB
Dv3R0OpBVe/bANrekCyYXduslQhVGcpuPyTdmM6mU9EIvIqFgeDEN+mSUrbrlyyMafhfQvwYzUQ0
3OGQv5jZOWMayNBPwGpEgcYm3lA/K3lX0V+2XKVsP7gowZjoLbt59dVopovFNzcUYa0lP/UKoXUc
10pzljGPSQLuILIvc143jbC7pGNLUW2sGHikGa2sbcD8zTTGqxDrN35CvvD7iBwdvIhTYDYVnp17
NEJjzi1GzKPWlG7Sngk0bmL4zB6t7NCJ7S6Ch9tlhq67xC/LeqY+1/dNkkQ8tbrYI76ywaH07GiX
MWRCV5b1Eb+X5enuLf80gY/y9paL34VBRCe/02RG2t4abJin9RIDT9eJRD6EmJYGAWTjIyYtbv+4
5EERdAzKs+SQPkNgzobQ63g6FFCKyLoyAwc3JTnSxUyqwzjuIw0Scrwjoltd6tu8togsUBo6gJyl
lzXTI5f4cuUtklJY5k0JoOe5H1C/VC48MHVHpXzeKDLJn2EK0dYqCCTlrfs/9gRb3hXIJjuPp4Tt
jwrR68i4psrvBYm7oGDOAGhqzcVqNp9fxMoWIbgi2ehDsC8HGG9X2JRewMPEIjgahhMUKOaktZ6g
JBktzsy0Gn0N/GKmTryanK99xqwo9V6c6tnFwC+NmFP5XUp3zykxxqMUyZN0vAnT3Pe1/ir7NUfU
6QkAiIY3YEHJPYiHj4RRH/Fg1pkMqrfdGJjGSAhHfCLQKACxUNmL1NxUbkEu2znHEjtqInCItWp5
40uZ463mHax5DtV4zfv+QAWxVmLJRD6Hc4Wo8Da6TSYtmEp3eakokAQNjF1DyJGrqo9yBpf8Y4La
sV4XBzAwxDA8DTT5ek3IMx0zq8DXF8culuW7M5nu6S6v4Rfp4Uck+q4gX2y1ndSL/Ehq8w3kFqwp
Z19/UFOcHxIvLiGWGc2siQ7rvu+C3ehDOKDrG5YJ0vPtQVvQXbbQ8fyylst83F1s3B0lpqcf0/jI
fuxBoXMGow9zMFjZLakO33E1aUquJAusVB8yXMhVY8Hf3GIWT1eFOOdO0GvfK3GLk6fxptKT+ylB
TIy9s27ybRjFpi1KZ3ehETHStmfSHsvcNCaNJcqKilOUleHl0nFvkyZiLkf0MohkVltSVBAezTH+
lF2IsMmcTZOMMCIns6ebvVqcqG1yRJ2hQdprSFKg7hoX2dY4JXW1LA4HBBIHLV6JfquvaRVAkKRB
zFxeqtkOuJk+3yp/dKAoH+SB/5nqRMuyttqC6XMxLiJmBB8Jly9Do505D9BSwhFK2hmby486V56C
CXL8mEVmhMYNVEZmbWcZ62+AoEvsR3PwaSi8m8OIKkGWmOkY3arkBG9aMMHLEl60XUxZqkjD1+SM
y0tiSdrcm7pVjmq00pKehdxpkUUcSWU9sscPqZgWF6wMlFM2y9PXhY+6A+wzsmqwc0w6yDURpa1T
bhQClkBzHgfNv7ZUfb3zhPRxuuJvS2pS+Yu8kwAspYJUfV6dSLW49Jt5y6FZ+LFRh3/TWD+nAnSe
tjXhGapSjfkU7qKIzd1FpfBimlqXLTBei5qLi+Ep3Nep2+wCWbBu+IwanaevWvgwioE7G+KHp+xe
j5Ry8M+574GL54OCbnExz9h4thLNS66IdoH149YYbjBg7frTYopuOCTzPG4hYALT8uThe6uezstf
6VKq0pPiS2as+j5/UMhtebvkRakwsoRMqqMfHGlTlNRWS1puh+AUuni7A4ZkzA1IADjtN6K7/Iau
A15Enf7h4349YHKV8VmJxgbIW6E5Vb5SCSfznlCR+NIr0ox8qknKabZMuQVztpaI+nuQeytEnB7v
6VS/HjiKoJhYUrLTsXUzJGaPiaowEjcIkoQaVtUsjV2K3hya5fo0fcTPKrITrDH2uJxqVdx78JXS
U6ouGYl9gvGyFOcrGwEMpxTC7Iwt8ux43GYLpNZwNssu1O6avMIVxhIc64B9ZiMLUDDSYtZnouTD
RzylN9kl/BvLid6syh5CNPRum/iq2/Heju1+GUh68ry27TUqUCXMMJ+GOBSEKdRP3rmEwwLCcpZm
y90GmbkN0Yzr/4g5ra4lO3MuC5tzuI+gR1L9M9prYD/1JaqrS1sq9OsJZJ6cOoXyRAvlHrhaDwC+
Q2mrzvnWM2VkzU/Poj2/rZGp3ztIbqsMD0/dQny/qeXZMECef6G6W8VNJvg65S/m/DTB88xejJ3v
hFOVG5A5xHq7bBeEftNePQUJx02ehvuc3eJKVURXB/EPUVcW0i3/cop3xWmJr+qkVEl86fr16dvO
eNiAlOzfed1j/YJvcvU4M1x0chHZP4wwcVM2wCTLcQJBTjD3P2iIolpTUzyDED1V7lzeZQcG7KRe
ErhKWsbr156jGtY/DoT7OUoIQdUqPZm+KGLKt+8/3RpZgiLoHnmEAL+iK+OpynCgEtUJbca7AwuI
m05KFx/3bTi9+PhEp3Sy4JBnKoL1Jqc0h/A3ICH53N7RHSbdo4ksadh/RPk72k+J8dFeFL+Cts8Q
I847PfxFLjfPQ0DLQ/SBhDv2SFgt/woMxyHM7tZ1OxT4uPsK5X5eA/xTN39Bhg5l86Hk9fx0Sqe3
n4jcNaLhviC0LKKt0665WF7b5utcPPIV7GVwAYM2HQobuaFzIzfzOnwH6cJQe+crRnERP6adQyLf
jQEoJKbk9kGXd7DeeAdO4l1ge7gQcDiqm7V+q1ngxTfgtDVP8FCOlvzvHwbMG01zG5OVl2XRl4Qn
5SKsfjuJCGIqx/ilyb3eRrknjzDIldjTskMtFVE/ha9sLuR3MFyN3me+JpyQWy+tDxQmcuyjhF61
yVXHJoAGzG/zj0a57uqyy7jaF3XA4qmR8OwiD83OinSw+s6BGUw3mzgW0HPrSHhHv+Af+u0OO6zZ
UHiA2k0ijp7NuJ1iaWgL07mW7o/HtvZLjGPhkmt1n1WHd5ouf3au5UX8Xqc6RC5b26aFJflj6zeC
h2Mya6uIz7Mvty7AZs1AM3GLCi8sI0gpfRfulw5CpUaEsG2bEUF/TFMoPEwqpoUAxc9/lxbml0lB
MnfLudnmz+NOqWQ9HSh5clJAzJyyV0ukBGS3FY6smuNkb1MySVXTOhWuTP0cKLlFVK2vFn6858cc
S+pvC5/UABqAldfxMHDe5Hb+F6WsrEQBmCG4jhTIHvUvZuKSV02Nv9K2wgym8KGJ6uP+B0xSD2FE
cF3xNcXwDCiYw9biajuVjxcza16DK3iy1BuIfF1aaAUeVXjN6e5PAypoOOu9qkhKleGOHv+NSE16
gUiYQhCcgT4l4E5nF/JidtevmowjKLQAnN5KZwM2cetUR/op/+E0Zg16CdoWMVQtBhXlHkHcr4Tk
1nrxbIrSk/i07c7/13NuCopBsRkJNiDnPkwyQx4tTqjRYzrasjf0iCLdSnUC0LWFUMARFz1W3iYD
apE6czJhyJDwAYREokIsd9nGHWzVD49izCZ76jkSbwpySoE9IiKjonTv6xgLmO2vFaHIhxveIWAc
6b+Fmc/jX2qYwAKZOoyusD1aYjETg4P9wTmTg6PCvJ8SdnB/p+2hCyDvNBICgCm51gLvyX+5YIJh
ae7I6frukejKeih5y17KnpEsPBTdHyZZTykvByG/aKUReMTlliOXJI9DVQDfePbqYrfCPNyCErYI
zd6ha9rAex5I1J3G2GCKoQfEmLGXXGybvt+KrU/1EfFF0Kv/dc4PpOlbkzrdjU9g/ZZnJy181yjN
jNaHfs1BiQueriKNINHDFtVRnOT7N5YYJrdiZOOfHJb2Rio3YSNMcjwxAgY72B6rbQWmMsg8kCDv
z1PX3O6lC8sI4X+lD3Ce9a9IJG4tBybdA+mY5XS4YszyXD5G14opYTX5S09Pa4N8K6FiOoCAIj00
9A0mHAdjDY6vzz6sQlpuw6hLjisCLeyuolFSi1FqCzR3G5xH1I9hyIJfChgLgYYWYo011xJdFqKx
i8MxNDsEpkRF2cvc2hPvr4i07S4lK9y159q5QpACUX8pVra+k/Gg3CVaBpdsSyjOQZCJbCKWoGAX
b+ISMAbYAMXM4t9i+E/95vlmvnnMCsGB1g88KfhmvDVpXfgzdrYQBGIvY7OQNRN1vXzhRC6o2pbJ
Q9Ds2vBPalrYcIpFmUmPgSywn0koDf6YwDblo1rkv0JZnvSYlL9QUtPoQRGvEYDsnO6EIiWTthlg
u+BNYeySNRoy6LEHIz5V2N3+6T4NlwJ3/Vz1g3EHLsK6xOJxbXEyTeFSyg/MwMuyyIVMBJM4w1ZK
GEea+HOiMcxvwre77KgUFro5XpC0ajLkUc0/ku+ZFNGBj9PPi1En2WQsX1Zsw+p5KRBadX3HT2CE
L1fXV8X76vxBoMWVQPI39cvtG0OpK8wLrxJ+IPJFIdVXIP2wRIrZoMTzmRS2gYQsWGvrQaYDp6Tn
m+XusiSxJg1Wdf4cDiq4K8MOJ26bT8i7XrTm6bEX89QwPvPeEuxXNkKvBWYtZs2iCnG0O1cf3+Nv
KSKgneiimZ4EsAn7x87MiQs/QMKs0Hp1EN1LVvRPrcRgjG4czGOv1qRz0tM3pjd+E/y0AsbETj6g
MmMtT+/5zvO4X+hQxXrbAGyURKTyk1LE8qoLIuQfKh6SKXU1srnWkXX6N1cBhYvfM3MBRuJ3hCs3
B+k2v/75K9LPVuMH0K4znUkqC51LpiUICxqLdnRt8+F2SzoR2J5rl8mBU0x039W5M+/Ernu0LwZ8
T13nW+yqqKyOzXJGmTb4iD5Q0ZLOdh8p9Rlo9TSmQY79g42SFRaBcUaFZfENo6wcQBShaEv3QCCR
M1BQShtFJJVIbo8/BjEJElTOKxOLXFE5Q/fQMPXhMXXZxWI0fdcCC12LqjN8vuesNpbsmpyk5gDk
rNV/VPcbwc5nyM0itAjHINAbthcvm/wc6MXmVz4Ga+t8ixD1YmeI4DIXo7nRmgvMpY/X2HME0xUM
peJI2t8494ZCZu/pC0kS6vV2Zu26kMZsZLMoHWqahj0om9YrpZMqX38Pd6Yt3UhT0cbuOuvxWbNt
SGAgDID51Ur0wzwg/lOJPb7EnzCRtJH2xx2iR/cCPWb8VJL/0MU/mOepeo/8pTTPHlcC/LvIot1I
E8ju84GzdAbz6Fq8Eiv5LUeclCE3t7DIiiihioVdyHCWOJJWXPLoxRkB8RfIazUY1iVi0EuCTFB/
XF0FrDmiywP6DdK344lmiRBV69u6g/772rPV/y3OhyyZ+/ojxAkUuEd5OyYYcsnf3v73TCQVqyOL
dRHpopK+E+iiWUESzR55IGKoqQzW92MT+FfNApGve2pME+RW6vg+GVoZGCSgTwXkDS+cb/cqG/S3
wBtS9COXTjyuHO4ABDA28xlNaNXzQ0lqwT69fANyDSPqVpXqO5WI6iPZ86T4EeNBcCVFc4DSIxfq
CVFEOlqdxpeFJ2aTeZL1WrCzOoydUjM5mQPZwXfhNsBAu/f1Qd/J4JN6E7NqTwAtctcwuTVDnBdv
RrA8RfU2UWfTE+N7DhuohLZJTNqIlaVs0QnGTvx//i6VpkLQ3W3D4Dlokwh945OK/mqMg5VXbjj4
p/dlabJYHKnmpjO33HqHAsYG7M/LvI6QcVfJIWZvOVJEyrIXuPecggGyCrKFBx/MITic/FTQcxrO
QT74fY9iDszyEJ96uiYmGzHmnJ2UE/pTrMn5aDM9zoOW/SpFYWUgpJeIwdxtyYi+eeCWtalVT+5Q
K9iGwWXEU0OxUVJJmwif0/p1P3jZKGaNKtd+H3nvZq9MV/Tuw6b18qk27dKpcRx9OfxxDlvx1m4Z
F054ia093Dj1iybcbCXP6isLEeoCSFFxr/jfhAxErPu3wNl0iclLGYt0SkCYg+nqQb3+np7z1Jmn
c8h0ml4mPMSdcznoUvgJN5l8cK4HgW87fgBqqVALJHanj9/qZBt7pa626T2AwZrQy3UBNASoATVo
0oYMMUDS3sU18GI7caP2FiqZaFgTkf21uE5wfi3r7fZwESzEImYXzmtRmb8KTAyfIBz7IEWQ8Bnt
96h9skuwov9gvium9TniAI061S6Akbn3Beh1Cm6nS7PB302jtg7SgbGn9dbEisNDypX0y56LlQ8B
hS9XF9v9SmVpgYa12xPJFFlBkLGzXEPyHEvvuBzEdQS4W8fBeOC2DcEkCWA08gPEjqxNlvsr+T73
7elEjmKMwrA5ONVfI7aqA7mNo0m4YWkdbktnyrsD2KKu5qkSlXQkCY7oL1kl8BbNsn8Vv9ODqybm
vD2MakoHb5W9LIWxHQ9UOMtYmPfElD9L9+7EBj/SLZVL/YlE9mVRRQZSreU+Fi7/rKWqE6iCX0Yj
MgwsljquOWSlFkGRTlZlvk4Qf+4OKmockizeI3L+dy3yscpfQUlQQhM+FtKlW9NeRQAqQWCNzMMs
oius8CqdsHRTltvnqcGmwq918jV2W7ChjeY2pGApDJJXbT+zsRHlsB9JO5dRmU0YqSf2wLuOVEtD
hq7SYgMDeOzWUsoS7gq8UMVZ7so+OsY2QDylrk1bfnUOlw3egsgtfNw/86kftDjVeJM0AMyfOBa+
hmWxSg51LiohYJUBPoJgF6tAiVzWuy80lsxOy3UvIU+Drfb5Lpk6mENeH8j8Zl3uR5yj8Xdztt/X
dQPBYqbQVjAQfnBI6I6WLLs05BsFSjRsgiJfAfHBAzZHv+cCja8F8c5WsZAx6HLEnYkkkzBRbVyh
4KBa6Q33zkdHtEqNYGM7XushGOoWdDuuwDCCwjzn4uGRf2zeAfjTVfnaGyf1KmFj0hZA1o5iuUhZ
c6cClw7aIkjrXWNYWIDjk8lfi9ZFY2t2AleRZoGadEZSowxCr0Kioq1fluTnmLyNl6G3ABFHOowX
0qAnclFZPqdcCzaiXdKwouoldRW2t9W0MY16vUZwwEJzMPrhITnkWpD3hCtwSRN4H7kFsNnIBUF7
G+kTtQRWNMRRlMEwmXVftipUZVALqKTlTEiau24XWTDAsuVTeP7LmpsDO6l8V7lmTwTs+1suFODZ
gtRWLitcMK1E+6fAQ6Oa1ne/TdrJZQvPTn8K83KRrvzeVO3X39smC5ieGGP6Sa3jq3zmDP6Gjt4F
kNdDXdFLZx81wjMATjsUSqgFPvCJSoetA7bAueBGzqvqc3yJbNpvPhtHKa+EAEAwrCWAoLAGru8n
OT13Y3Va11c6k+xfEDxzdZWqshEvAzDJdBuQMffgfu++Da+QtsTUeXznpUZ9BXw08/y+KfNimsRI
tWW6WF4rKpFcRw79P//Na0lC0ikJiA3DTTtplaMvD2f55jsl63oVwZDpI/YcAmnVazXmTlNJOm9m
5IiAU3/3Jpv08h0UXstGPxQQJmYDzgMb2lRXQQ8I+Mu6NLrTMcCXc63KlKSlUtHJy9N2p/38u4KX
17dKu4pm9u4xgbAbJUiEfDUa431dEa+JfNzlAgPElq3rfUdwDs9kIF8wPBC6VGUIOFggd2CV8a6a
YUuAEeWuf+9LoVK1+mFHedbX4UPcWZlRlCIwWSGw5xlRtn10Oy+uz7tP47RG4mQMpgyJB3VE5E5u
jTvLaTGhUEQasjhY/omi9z/082WPSxLSzMEzp/FmYkMQEILaf8vXVQ2+FqeMz+Bvyd3a8/6Ti33G
/gtfTHEKkXP9fZV2FZlSUEonm1tHwDn7qZJnMn0ZuowslS44RseqVtbW2kroBx1tOTtknet0fKu0
yrx+Y0P/D04jkOJHJ32WYaSag6ZNvK6DyaQiYDElgR4SbOfoYMd/QGG8oNHg2HRBS3wTqqXGtEAP
iFonxXsrAHzhP4kiYd088vodBCgR8tsllg+aLPItHgLKtldE9ne0nDcD1Xs1FgjJghkhYMINgoW0
Pg8Yztq6b8u+EW3KOKe/I8+Zp4QZDLtDs70hf2LRmkhZ3dzOak3R5xv91iBUgsK4YetHDqZfCS93
giIwC+pDBwHAOV4yH48GPtCyC+IyUqbYxBu012rYw4rFuAirCkiDsHQva7jJ7ZnI+m9/zCzNIDoW
NqchUHAkeyDsDKQUFBPehXv53Gfkg+UryRXzFSi4jkY2wa0Ux79qXBUk28V1+qDdsdHN09cR2Yno
l+ps4AchkjPGfZX6JqwOJgeYYchFz7cVbGhv/MpsVThQqcdIY8/Oz3NC0CwknTBiGlECJ9JrZHYF
dSKS1QHSdr7LydCDPDPDg6lvoVcowtQzLZyLl5o/Ab+MgaP8OSQJejveNbya5AP0jBGEWpbUYnix
hpx7U4rfjZG77RbUr7WP9tVTN7js45sO6JfBhspUlUf7uiJ94WBx9BpzYuGvnv2hNLRseGfi85WV
zK4jeDbWpOOjOfhC9VGWLN6dracnLrMGXBEJfbO2lu7Z4hK8eKRUd1jJIUeL9y+gp/ialJ4hj6mx
RvtDC7hhIZyOB8pLZSLiq6g5dF5p2FWHFAUTpL6akKJncoPNOisJbueh4wsR3C3fC/mzviIAcGKN
NwUocuQioacyb4139cKWL9+VybQXWFS3FvDzUF6gI15IKAz5Ed0S8jvZR936RPU4aYSj9ra6CG2j
hR0PzDswu+QuRiZekRmWwrOL7zIAqmUmjQvc8TOD+X6Go9N1EUr99npydk9VULsLy93/4Ls5fTwQ
nCr9fNRkc5vJsQE9vjBI70aLUhIow72DToN4FlPX13Np2pY3J35r/S94zXKhEQZNSaUTKODRYKnm
tBj7HaxDG+O4dUY6Sxqp+nMWdtdQM2BysFMS1DXdaP5NWK5qV4B217a3Hv/8jRBXadfnHJMc6VXY
T1mf4Gj1Hi2R6NNCP8ZNaPHbY3IfSTUUqocybI9npCyR0OdKqeMnAQBRqju/rDjzLnuJ1rqApyI9
R5H9HS3nfGslZ+DGaqaKZZlQojyDyrACQVIspycgErxaXv3gAYdAw1+Nr+F8iISCFtMOXM6mL8Q5
mCAr3QJ0WFd37rToc95Ws8aFIyfbZJOuGMLz6K9WuGUHwlY57aKNAUfLGOwq7jtBoR5Vk3lESojH
L3/PxW/4OvqeAk6mnABsWLLQvFwEC/zSyu4N5vFQ4KbwP0J5lTG7rylShYzoQNSRXN9rmw6xRcKP
yPjJpYuxnWz4ap+7wzC7VSnLeSLioyfYPdiM/D+JW9FigeZcHuNG69sdESnJYtV3yhN0R4Nqw9ov
4FFH+FtKd9zcFePx0tEw0A4vmMuXW9bcNas+DsO+sA/NXjPLa0SSOiPRn73xRHmR+YzvnoGKNKCg
ZK86xiAkHzhbpviUi/ssmgJbOeJMmK7h3mnNvKiHwk+StDVlzVlHHUi2t24IDxS6qdTJoBh+2LBW
1Futq0PFTKJmQnFrszzUT1wLIP78d6NtztPGZ/VtguOu7+OY0HJYeDlBFxRNUHMEsT0588sLCPve
+zJ8TNoD2leky9M0QXzfVkjZqqIiY8dtmWX88i4ghJO4/JaqRVumm5KcsFJ2ll71Jfcof9e/r0YP
3eLoWBkv+iS7DHtyEn5+EQLFOm4MVFp6oIJ4E7/hwuD4yeHdDfb+Y0XAWu6/oz6b2GX02pwGssJz
GopsRMXECl1fEyoVsGCTMvrrxGbdzwTCcJilFzt/Psm+cqhOeiikEm8kSvpCyVOXiLo5WsZeaHkg
fkkFMGIjy/tiW1Fe4kNLjIatX7m4d0x4gyhGj0mjkdhemvV/6TYdYLtve8iUBt1xEcdfmntDhyOm
aVD0XolIie4fupi9ZVzezkKHfD8ZqwkSJFT+7Ux0jQl2r+ILf1CV+mFNzxv6U4SihgWb+A+K8/0Y
2F5/ICvFPBjk8LoXIc3w5jY7JW1DySm5kdnAOpZBQ3I+sWYROx2Pdxu1DVhSsHBTwLlDr9eLl8iS
OgP+yPFTYcTPU+qZboaef23Sv/xFVw+edJkl7ExSfnVrbq66BvSe0OyZD+h5q27r5I78chDccbw4
O0BAE3TYYBL4Rx3xyyeqFxnh+N2EWvRj9huAPT27uslB+l8jHrh48AFJPqtlmfMfNiZzW3Wjg+gX
Z9E9AyCYrQ3fH44bNPpe/RCp7MRz4kDJ6DsNDlfOaA803VDVq+N3NFyKxOhXCI0Di6l8k8QOcAZV
PwrbabIobcr3CoJIPD2Ldk7yPG3FJwMA3nyyUhBRSNSR1WWokDMCguFTyhQ5QrlElZ5Sl5Ij3hwj
Uqu1exZ3GVf7JCAz3yG86vysErUzLF+BVLo1QJap30SaExyrGYpDeOlJNcTHqDANU215KGMkihoD
N/4y/SeHaHPiacpgUyyWNUk+5nPXKHfTBSd0NFTWJoIN6+Z5PxXRbTxsTBFz8eVep6AO57IicZLG
Ae7ZuxrgdhSQJUsfEnyvTnxZjatZd2tPCE89IksP8nGJ3ZIdx14X/VdO1lkkTbI0YnpZjjIb330P
L1GO5AqTkRIuDwmqLhN84i7uO853GaB16H6v72ISIbkcWJlcP3kw56KEovCCzLsjtA9RRuvAOkL9
7rfmzdjTqr2MBK3XvXNQjMIQscvUlE6FFNQ8fvcSYaOdZE1T7HKiOSmOHYHR7m+Fc405AfAu7hOu
36cumPqO56cdYnI7dUMaRK/WLbHjnfnpL9XeIwNNQMQrZRPH8hupvWTNtkafQ9MRpXn7QUTl9tbp
38qi1WJu7N4XLtGDxpq0f2oAW07tGM0g6TlLt9Yd04OBMfIqzmdLaDTZLiF/2MBr5Qxs2X1bK5tx
Pb+JdwVjwnDdhN0C07wqhWtMjaRnfW3WL1cFkix8uu8pi5K2HqMD3mN26nDId8qkms7TuMqqhmDL
kRlG//PLIqKUa1bkiKo81CjvJc+QVXZ9WPBFByf15gPZ9P72XGty3DU8Q1by9Y5+GtxThC8K1CAk
v1ik1/jU4dR83nJqAwZVEpB4NFEs5ybyNr0S7lfEg4wSix1IehntkQMUemiSBsL75oBEX7hLsVOG
Vvog3zPr7P7WTg0RfOq0Coy56ZYyFxdvM1mFHHpZl3O7F6Ak2O9Z0oghqOjydy/uI1bfiONV7ex6
Qnu5AUU3XUkQQnbVDkeuplGa7jb5qtqL7zTTtj3JwnG5ba5iyADYh4oRehmqvWXEF2kH2k7iHZnY
yT9uAEYSJj8XJ+nXFDQb/2opu5R22asVJSmI0zJu9uWvyyANLjsCFPHfU4AXvJxq89wDxhhpAZMj
NH58LI1RMXpi0yeY5zB5eb2wlK1i7FeOSI9m13JZr+8+iAFxhgtb30sjiWrTgWwJftSCIzrSj8dK
owT2L6y21eMkWgTlCEf7kU3BbYlsaCQj+Vx5SQ8pcelqCsbzjjOWTqu+856gw38GT3r9zsQQp8Jb
FV1ox3EDg2ZSo6AeLu3cGqznyojB+lR2oM4Vfka/g6YUmDShYnkali3yomuv89PIuQgnkybaoKlx
J3fpwoTCQjdPDe6Cd63kWL/lnyKVF1TQcDq28nTo/153v2mpsaha4XcygDYI90tEoQrZRgVjqM7L
KlKdlecBlsA+TdBUE6KM5aHcKlvauE91Qsyk51ls/abueB2vfZECU7K+eNEdDxhwveq5M5jB1l/F
RaaS3BUStCajP842QjYEfR17ghJdWTCyysCiMctXR5qj05Tos+8uCTAqnEQRjgMS6DA0KYkVbABS
KVM9ez6v5HWPQzOYrEGGvANtzF/igDs4KPJmrSX+ZgRDEhm+cheeWyMPyuBYJYIuRBSVDu/8U0ge
z+9t1VKtUSr+E174tI/JZT16iS/5+LYmowEGE/ODvQHMOKAhxaK1Rd9J0V5eEkRLBrkBY4Ut7xod
8KhKzCkHVZa0/0qUpGeSq3DnmNB/0yNi5KvYbae8mnMhok/x3qOJjE8MLearkQGqGxIN6UTov/st
lJg49hreHFJybtqqdwpaW6dalqOGUkHVnfzWiNcNLEu4RQoKFdfwwjZi58ByzC0J4IoEoFnSaG4+
Jv8GeyEFfgIfT9Dv6Z1BcuWEeP84+ARS4JYo4apffuwd8lbAs3EhqqUDP/R0D2Fl3AjQp5dChAQQ
+qzpj6qc4lAS9vkUSmRNdBu1X2F+FMDRNzbIfcEX3g5dsFi4W772BipTtPIQN/HLxPI5De89cWx2
Htw7z1HLtBQE7mZFTXqI0q/OoqKobLxkQFKe5F2FQWoRjkSTSF5brJjLE9cOpLyS/ADfy+grD4gi
2V4t0QtHG+sH7C4tOUFWuoJ9pEV7OylFPH/WM66n22NZdMNPr5hcXdnOS8fIjh7Mv4KB57fSnAbU
CkktdOIVlw03HL2Cz70WwUgBBGpXYVesYwEJDFHIlAPmvSH4rXxQNUbOgMtBqQHhijdWVAG4xSA4
QUHc92DiI4Vuc0Cs2lrg2YFRZHCZ0B1C+AhPF5YgYCKoHmwNoH+RV5PpwRd4rx1Bne3Z4B0AvsrS
ttJo80rWf3xEkEQlcIJXnt19nkKdawIFJMXqUeokDRNWWyVf2wy7eYUkXTYHFCNPq0Q0Euhp9Kzg
imMYwHQmWiNITdtd+B3uSO0apc8dybRR+02PV6h8UTc+e8eEcQo18Q3ejh+04uJu4Up/wXK3dXQ3
tUE3eFmBLVn3OmjmfKoqaWj9WbWn3Rlygl0ch338BwcSUvmXUZeRplipAtUh/c/UcyaHRO7kt6m7
kZFHc7uce4bhF9C+2OCX81Sysx4UwWDalAX21mYBhGNkeXw6VDydKnb6jkvTPBej90L4J+op8hrX
gjVpyZsEuzMxUBL2i/akLwtjErf0IOXKHCabjQQEFzwLX0cuZ070oyZz6DuPnOkL69uMEjtrRUea
MsrkMUICQjrPgZDozVdDO5dVVRB/Tcj7kuiwkuPkn4mmTiGcetYYBnNDXUcYbIxy4HS4a7CW75CY
as/fl9BnPLWiRgajXDUzUl+2PqNHHRkAjfX3icOaK9RIWab6tRy4Y/Ka6hdk38uPU/OXuut+d1Xf
zvNW5LEoqhN2s91SHMWeh3rDs4zwI9hRDj6pxS837KOxvvLwJWOhK5C0O+7Qc0+7LmxlhsIa+yzi
cIXGeyalklPXx6Eicimu6NN3kdZOhj6NoAm+X8+wPOnaNQK5E3KYxFuTb1t85wSqiOg68sbnsg8n
bp7bKsIfhwucDqXzxn6RqAJqD/vjQhwQWXXzKzkI2RJmdKP2MtJgCRa8j3mVkhLrGbCNWEVmGuaf
0bnDzKkU5s/oH9cRXhqCDZNdNYM4/HjIbTchPHqYrw7wY7kKkZs5Q6dcrQxoUKUCbQIjs6napwHU
ksolGwTk7znVhIWmYp31LwPcZjnnakrRY+66YZwqDpCRlxejf632wnArUDL1HTh/aKQJBtqfVvf6
y95XVHx3tec1wiAqIBvu1gCKPXfT0okSRSXMHNwtVBlOdYRF0rrcbX4pzw5YJWdWtpevT8a1UsDt
KR9ClJw+DcMic9liqnJdDHGdUaFqKtoDQMX66f9xK/jfCUzvrwrXaJLKGpUEdk9R4S/IA8IgGMCQ
R9Fjx8CHajGOCf8vr3P/yUljtnhg9YhLM+2agE5T8x44Bo4Ayiu3Q5B1/O4541r2T5eutIrrmhao
z2uRhitMFJGsgy9xLFC1CS1fThVqVSPctaqeV/8KSMmmRZxsVUvmGPii6eNCixW6beBOvO34XTOC
96k2DyGZA9PPUwbo+Z0d4AAtycNl8TIWs0kwBbiMKBpIhafucXIkJXka6aUG99rlzmw2YJwn7x4V
iYT11/9vt3TP4dwsMFQVyQD+7jUd2RV5CH19iR4KvZv8vUl9lDTtaHbYiWVMkwO4qQi9oJRU6jOJ
YMcoQoDBs+0ypGxnfwmU8MV5CUNe089QhaN8+sv8k6uCdh+4SXi1o7mnrc7f6VvIaVVs9uJFXHxK
OPtnIkkHSozugI17Sit+jIedPPTL4SIsZWQ22PW/tRzhZW3ScjvZkv7s+a+YXSAjR+yXD03VNMN3
Wyooan1VuB0NB2krbBzwd4tCQFp8kmw6Kh7AEpzHNjR2zkXRyZUaQUn+MbZVs3gK7W6lealcnMkV
Trhw7kO1Y1HYSbyXIWDTGMFhhIDCNVwB79CuCJZzl5cHgvNboJzvVNOOwLVDdKNvdkSLE1wMdLl4
qbTNo6cTcyCoI8GIDn88d4akrb+wpHFuzL9kfWNvfCf03Jf24TbCFI7ZlYQO/6PIBVzaud829BdP
k4H+czEUGse3iIp05aESmN3crEkrxY7Eu6hmQGGtl/g8z88pmwPLWDdtrDh6z8ilXtY64UnKxmQj
/QmOPxIH470rqyXtdetg1UIHPPYWvVGrptFPUrrJk6fg6Frrf+wSD0caGxXVTIkYZTNhjJkPUoAQ
6VFMsu3LqMNAiGiBZBICjGDafBiD9uQd1lxYshMjKZZSsg16vyZlImLGrnFKOxCQc3/LFotT7rKl
YBOmeeN6od2OS7otDGrt5y13ul2L93WmxNrPZ5ZJbrUF6jwYjEUarPy58iUQ6TILIxXeVG12jkko
tOu+qJhNqLJ/au2aljj4klv+HTmS6LJUi6/RTgw6QOsUM716xktSOClW38ZKcaFnAm/gczjmJS9d
b9UlorOwCQBSFPbkzNNKh/iuMxG4vmyUEs87qb7nXPDxCe8Ik9dx2MadfNhsUqti+pv+FEN3h/FM
CUyg2if4YbpZFZT6RfmYCHBlpgbeJrqdiJ1fgUeQqFK5yqadf03HXka91fWLG9ZaQjRmdRzZOQ0r
UyyEkFG0jbXoRTG+jGVfA3VKPh6KTXI0ivV4RZnsbGYPvRHGd3Qx1EnRotZT87f/b9ucA+37sC6K
DminJyUY3qjeGWkxWB+OG3tI0uy73+2mXWwHa1jH0cSeBzY25djIE3ijwKJNTSiolLKlDdwAE50s
N4pYrHCSYsGlcud91LxG+9XopNM6p/9GLZ+AZsScTc9pTR3G03qTFSoGuMypqQ2juPxotL1ZN0Y+
gMdRh8lf/m/ySAZGpOntKgFwm+C0g3l++l699oSz8pAbaeLateca0hbKS74Y2zf+d+tz+dCjpanF
WjlXmsOa0YKLFVEkgOQY64KcAlNbg/5R/3ZWjGlZqAF6MteUDLYfNoUXX8+n+WOiWpXptmTyA/p2
6TInpSb2Q9QiEWea7duSoeyjB9J9qOJy9BA47iREs1jXbfwjEq2yyy8YIiybOVReFg/gKwgwBZHx
dGeiPUms8RlaV+sRVCQdJXUHBGV9gl/O85vXRahjBKgKwPCpOvqiRB7tgb44ikUl3n07wmr0Y0eD
ObDvLMqShgjEPhUDFWwKSQMNbZUsGDwjezWvVvzJpZZ4Qshz//l5cz/cTKieh2n+I6rEfN8Y4xeo
fmbbIET/pGt2XI3RZV/EUWllMFz+tbZZxt34e7mMkIOkX/9vcEMLIktwBVXe0FgvLJ/uh+tH+pIw
WDH67tqWW4gujoY/YFouGCk1kO2rHpcALmUUlw9JVu10eRSCkPIWhKXJik+Q9Y3zKVCoFXBXVATT
2BEzBPazHAvpVuBEG6f/4IIOl9jZao/vwiLFJlJTj3kmfmtmwKvAYUSPM+6SpbAfVxKhjDSoaxqe
p6eRyVaveleB5lxtxgDtl1lCdOUEgcTBX1Xye5NQyFqKdRcJhZljwBzjVUIOoAn4NsaLGXWMv2lA
Pio1Stay3OlHhzRST1xSRFM9EGutfDCYH5WJBx/A1ffBpbqS7gIDX+55rLRclyS3J1+xUFHfPttO
+XOdob5m+sbbmPUMO6JHPJhk6mRiybcqoOQv9jXPXO2KIi2sW2gfDOex8tyTMV1T34bHEVnxcFfi
D+8++I+r3BPoxbJn09NMkJ/6eULiZ9WbTnFaQLul5IcraPqcNMcwwWHtfts+C004Uf7BKqet6j6A
2oJLrdJJ88sZ3NW00ctsPRVOoXNDI4NJGPJejAl7GdVOdkXUQLUA3Y5FGArEv+IVnp59AQoAwRVF
0I0O86R9EadON68qcYBM/3CarpmC/QmfptvLfE/WK2FmqEBRmms6Nz3oYfb+F1eyRacs8Jbjc4RB
EzzVanyglsLC/1Y0zK5ji33HY4UKZptj/ObAt5O1VA+y7L20JvRqRYqwa9g4E7r/aaOKzW1yr6Zy
SdW1C6RT1JLxKnpY6tt3qzfmK2Iw5m4swCIXUomQMZVzBiiilfc/CgjNlAt3bNTgtQmby+eYI+pe
QDrYKDVM0lh/5LxXaa8B4K4bgE5lWHFOZSBL6jvmCaB0umHBZhlwHP8el44HO1zdL8lue7Q7Pq2b
bJrk+QuLgf5EQ8zDC3tgWRAHYoXsmAlOsm42s65CGA395kwo6lzNdaNu/VPHC433ZfktuqqeCgk9
TYypY6d2ngbBP7zNQfey751H6wY3VXckzTLbIQdGuHu98DABtcApDe8guTcebLjfAeiZK4PrnWqT
4ZvvJo+sksjgQBgl/z8JgAKWyHPX9FlTgCKXT4iqFTs+zKuobFlNhmyjdJYh2dEJExH2lT9+gjSN
nl7YU+NUnTlSJ6L/aF0eQcr6Z/OuQhfklVFMFbO/25uCvLNdmw1Zv4nLQEXOLD8a4NUauqwBurQ9
yC25NZ86b5XcKh+EO3jHyl/ffD9zJPQKWpgXbGtR7WcERVK+MWEln/6aieDTRAYA/sMIoOlNjF1i
fTxoEa3hB3QisvZRDElFjUZvkDNEAgqwELUFsP+th53oVRpaoYtwLO1yD3Bw27jHTFDheWNPg0rI
rRhmwRyTN3xLb/TFbL8WARDtdu8fO2qOGKI9cjhdjMHVDm3cARnQFsjDVywfi1WgFNP90lQ3azUW
/u0uteK6U/3niboFidtwFrGl2HfhIhrG/iegmyy2hkPOleEVX6H2Vv/apJegw1FJk+01O8wUuswx
8hkMwV0ZQ1PevjbkbyFQWN9tKeyF2yRi08Qcx3sD1GJ2EpCkjFtt12sogOS4iktopZaVblL6Sa6F
PGcelvryaUspmNWrYIay/H74rQ8b45T/QpUfW5+ceEdFL+ourW+24YI0Ln5LxnVy/7uLMOy97kq9
Mmt0cwnYi8NKHjloZLzPOU2a/P40GHLYvRr2/Pc/9SaLLW81D/gRh4fPZuEWvH4a07JsEctXwemb
OPljV58C8pQaypqjOovloSO22kHTE/qihOiQCtfb74+AnsuYJ1HJWGffiAJXDzHvwcw/F8dijBo+
9HkQCiMW0BmkuVtoUqYiG8+u0fnLTeLLGr5+Yy2QelTJmOC3MuwuQUrM7G+eZPwG5RKCpVb1aQeu
LLwyjopl9+vVYL6qbPZBWSR4UR7Wl5nVaSo7s4P3lWhqW7C2Xh30UHLA3EsN/u7EBjuAJl4vjIIn
A4U6dgnTjLz8ge115JQ0W8pLFZk4/Ir5hfds9291SX+eAPmgMBirTsdazsDR7oHanK7agEbn5Dfp
qQoVrP2b5r2ER9AmfawsAZk9oJU7enDPzN3BOi6zfdwp4Lj4AGJLvzvI0d5Akwq9QG8FPXjy3o9s
1uIAomgWRLmOj8NQT25ngvUwRx40aUp/WLnmvmBEjNHMvxe21svoWVjSd5Ir+KoavJtw0N/qhgD0
vZQndhd/VLZkWz7aElJ3DqxgIKM3bfi/7xWlFxumEtOCnau5qZTDi6vXDPqLA5cdWU0YmjbD5uQj
B6SbHuCVYrKQwT2//OAuwKbQBdZh43fwjxhnIbHwOEewFfUAC805biHz801ZV7urpFQRR/WmUeBc
ekV/BHeYu5+hXxCd4ZjZrIEaVS95C40MJ/tIvbGpCU+YFxSo2kVhBXfZoi8axrFXwaZU8/jJhksb
9uTCGCGoRbS6LHRRw9uo7Y+FaNF/FBEF0X7h2/MlVeRVQHJKArcq4phInIpt1l0IEQe3I5ynb3RQ
oCX43eOXTpu8gPlO04y86MLe2zl+2mkCtCq1Xu/+u8nlb2FIn4I8KgBqWHp8kzDg2XaglwqQWvse
kyqEGy1B+XpKZhUA2K+YFX6fHn8AdtrRkUWQHYNI/nuVTqZp1LWl0zy8s4icEVIKImbGmWhR3a09
eoFr0mWVCbzpMXVz0J3BKWaG7aBVgdIRbNt+7s/buRKKGcv5q6zeu9inDuqZPzN2CIcy91I7ttP7
GPP5zorP3Jz2bTf0HhJddPeY2FlRwaqDjonsO9TurUtojQYBnh5mpgdcvIrCVLIlPYj2nuVX8SPC
NUYriu/1489RMfq9glF8FXeKa+WrUl9ZyLJcYh4ucFPVfAxlYwm5kNASEUDRZSPiyXuwzxNOmEzV
I2bpZfRhxmwCVSVDInfi165c7bBKBQjFjUqkJV+zFh5uH2saJI3WhZOe7x6kgLNWMq7cG1CFdd3c
x+YNAM9RMAaB0d9ZPijcFUfO3xoXbtwXVmAKeTcbgUwuXLaURIJJJ0Mn+LhNj4wwLvDzIK61+1Ce
eOvirwwAyN8Ly/rrB+r16U+oJGH/1V1y2ORBKwly7s06XLcdvPRWw3H1zYRqlkiIwPZ/X7YRjf56
IsGluWncNoyIIDgJmy8aiiV3Lfp/6NpEUjjB56K53PKwsdamn/GyLniIKpPAt4LtuTwv744ZboP8
qzdwSievbIOOv1DbD5JTT3KERPW/5h6HiQMgeEzxORB8tefD9DZkZqVfvQhxD5iQRC0vD10z2uuV
cr4lizump1OzzchwsOohqer4njybctBXA1wXCjkosxlGzKhz1MLWt/s7ztyzwF6WF7OFI8KrK3K5
+kSgXMP/36oSUUgbSjdyarJiCBMOZRLWk+lMcSumryu8h1r4lTaD/biE2MM4m1aQzeniRvCu82zE
sgVfnMiOzWEOo01ibiAeAju5j89Lc0Ds2qwlRRGs5iXxBsGGPBVe8MJmeYKuAyEd9LdF9THUYOhI
K9MNeJnRBbh32sXOEYX8m/k/aq4McDyqbDR2umxb1OD4pUqKYgBchI2Ju4+8HQWjG8SIuEzxzUv0
MOA4FACrUfH5CFMeXyhyBxIyPKzthnJsIipBQP4j3iBkT8iloWZsKHtgKqIAbO5UxbKqUjTD6z0K
o1wcdJXt6GFAYfQE0DQsWOQLlvbjfAMh8uwX6ykniWXLLsTHO1RbiI6TkB4qSVIUJQ5ck0cxQ2Q7
dZVHYnomyVtiqtRnkPNzWh8mjMCRruW3jGTgTCcv4KwI/duMdKLha84mlXAiAN+80nROzuyhQMWk
mvx221V+qR6GtCUsMvTLMPHqzd19YECY/kUkO/brdYfo5ANZpFMFldGh9l40qEij6enGsZsiSyHH
AQOmhK3QgDXSHCGspwXAHJv+FCbfx7Qw7Gqiv7ls3UAUXdSGU17jugtbfTa/Te7Skbde2v/5mu7b
STuBCp+IclBClIODVDCb0bfwZdnQKCg8C56M/op0WV9r0NxFV/Blj1WSu1w4ayueaDSXuG/f4jj9
XX7NnYCMtbyrA/aLMuQZ2n3jLneajOf+ryPjEhuFJdUtjG/KyepdWbwiRV8aQ4HGZIjTaX2xg84t
D7t3t42jndEcfqS4tGN9dwz5xLxSZER/dqAqTeHzpICJFMVjS0MDPbVSA3qAOP3UV7dKPnAcJnXG
U+p53RtEPOHcpD07NNS1fbYE8Y9xibiYDjYCqafWtoEfykVKPEvEZIvwMp+plhaej7lrqaVb6yf1
0T5pHy/M1FwtCoy0H/51z3vVEJlzROTLkn682KOaZRpTEsi2j+E/dzCMXWxVorPY37d/QVXauoEA
F4p4LdMKYFQJUwehxDZ+nq44DOmNsgGWMakfw8jxLxx9u2EJUxkuf843tU1sU81Me4yfFUpLwRnb
K2m8QEtmVf5B9WkmWwF8iPK2oqKalqNmdgXFiFlSrdWJIBO7yCZrxvHcId2ahT6UqaJ5BzR++1ua
Dv7BxgsFItImKfJ4LxA77nx4wwgX9mloC8CtuA+1KyYnz5hrh2cRr57foZZnMiLH0CbRrc2tPsg2
BKKi4UYyIPEJPlszo4Szl/fBsGisLMMae6yRvJPrQ1Izh9P4lfX8yZRp3a+LcmZEteZKbAd4vaAO
lTPU8HDCKPZpRuqnzlwBlXY9cYUYnFg9pZwx3Y+UkhJxsU2LTFvuj6ZLJJt7tXBB5JqgUEENqsSP
1GKkG6Iq5VsQvi65thReJFgyHXt9Horg581cxWagXSzXw8Jjyc2Fiv49BraMFdVJzxlzx2EKGEOR
3bLk0OMkHGb33Dc18NGsnMUeaD3REmXfyWdpzn56d9jMFIn2rNeVDMy8R2B3xDULzgC/PYkoQ3K6
zw0LA59qDkU5pNPH96o2EYJpiOZSKGaqtpB94IQ8gRR69LZjqDcG6M1//t44vhQDIta51xyACyGd
VK+X3wo5xQbe5gN2QWlnEEc8NXvLyhjezPbzWX48a9norMQoIArJwqb4D91mNNmWFWSAiCs88h+s
6iVufrudnOx1ozmIOX4NWt82rlZI5dzE2QOUbEhu9oc860AjlWnWHDFKikR1kRyiKUFu/fbiVQRh
tZ5a1nrjjX/sia/H/w0QZ7EyH+WR78/pvsCyBP+tx/1apMiMqgYn6T7bjEmnQEBPqyxRGlSP1TYr
8ERhEfSII9oKr7GvUK7zHbserPeywzJxUbnLD74S55NiLkrphYObquUSHX0McZaZMshrhHtVIiFV
U4AxZEjcZYXIxDq05fQVFpk9UV8QBKGlw08EshUWB0C8qBzMRPc8HTba2q/u7feW+kopiWgHGLT8
R9fkPkFzIv7lHMI1g5yhoOkCZXqmVG12Uz4APDhRz3TMxw+L/4/8Ymk+s4ibkbjY3iVjHzOefK1R
pwSXPfohQAV7EWrpAT5VFrAMy1+6nzI1Z8qKdXOPXm8OgoAxsQAd98diBej+Ucpg32+0OzaljmgW
l3De5PFlDJsZDBIt3tC6QL+wzjgutffPP6IQt2VR/a1tIX0XsclnlGnFrviN4xZbNTkoDnttaABJ
KmA4kCW2t0EBTpRxUMLvH5YFsVOZEiCa3Qlpeaypr37oo0nN5hDGc0tN97digppdRbhsp+rM6KJm
xh45A9jMDWdpUsDH9c4GuptRUFqGAGuv+cFuH9/feZgykUfS1Z83UBBKXQcgrs7/X8Ht2XusGjzx
zW5KPm1+bogNK27L2DlPuX/y34cy3tfvGRJfWv/io4ZtDx7dCQq8xTQuDptkC7iaFMYCS/gy/ww6
xPZWnrsl+HG+CvCYxHbHrEL9C1PNxFy3Ylu9IIIR/2fcruaeJcN1T4tUWRP/RNggAMCEtEup4aAK
VEvoC0qd1rXXk6sL3hQDCfmvW3dMXZJzMkqtvMXxMCh/8MYG1msCEwlqtAK/LJ0iAHTXZmUZTrc0
WPOjwIDvIpFhtdaB9ZZ/zfMLMAg9zmWVXGhUrKxZmWLtE1+t0NfSn4jcRFmqTAm2ELMvZbTehCsM
rBWAtWMX2Oz0kT3iUCldyGYzwKuMvajxPQt7TXS9+sc0CorT3/fXJWYCmwCaR8m4zW6ZCmmvKawZ
vL9DhfRIerY60SxHz9t0olFVOHfOxvLdoD2uarsrWsWziQIcB5EyKG6VLWmE5Pa/mEVVMJbjNqd6
sFQwF4xrmyWowtgVaUraCWYDqSXZO0bnQmFsehgM6aiMg0VXwFx6raU5+iSEN19yByFNpTwQmIL7
vTKslQ5z4+rJIwT9z7+9PrSa5KximTxZ1jsek9oQGBVjFyEs6LwhOR7kIBUH3KmN+Bloaw9MC2ON
eAMKp+ovpXK46Tl20xSL1XZgwPnxQhgcvugvwsObgMd9mPWzZPQPeaQfLbaAZS76zH6KRYp8M2Rz
nF3hLabzkNAa95fVnVS4ie4FLfqDL8G/zlKVYmTNnvJqCCqc1Q8T5Nba64Z0iIkPzOfPLxQnQ+VP
YzZdUFjxCDxF/vi7gkC4uANBoJDD/eNUFR6ikU0+wcNLlkv9Adu5ovlPpx+CpotzNReTi83OUx03
VgZ56MYVl1C+vEidLTSfwihSn8lVnXQGLmBONI+uz7H5LJDyDqTh6h/ELmp/SVwEHe5L5cUiqfud
IUBMvlxJLO8p01NiovwYO7nn2rmsHgObb23yJSguIt4OrMwLPssI7zOnh+MK/lXrdwRVVqICnGEC
4xchfvGcyF5Cx66QZySRm6tBXoCJ4i5a+G+/53MezzFmQOXsPlMnSc+LrRcuRh++tsW/nyywDgMl
NRgDvCEH/29CszkMt3ydO3Au3jYpOJhQDY9sq6ioMZmPqbVpe41ELFn6Y46I7PRbZqB7AfOyqi7G
qtgfbIPBFngSi5AQlmtwmZzRnouMUM1KXQA3hX95N0t2jyyaGBY9Oqh8Fzkdk2qO1DNQIilG070U
rpiRE2e76orLHbPHfANlsgTWc0qSG1JIaQf2f4NCbAKoCgHLtQcRWP7HgSa0zWeiALXR7ijawEwx
IGjHZf0RH/a40JgepANnRzxEx4yTeDFROVfQa+HcT2POUa3lUrXDT7ZCvy1pSLewh3FIBV+v4tz8
btlBEKAxBt5gVk0W6WYZKMrK5uecFu25izjpjIjxqN/39Hi2JI5xp6n4oAwR6AHoyVt8SGHmfQkN
0mSiHAhTrFwLgWS52rXHIL2mncxDb4OJmJcRR6+Q/RKYV14zbFfkco+XdfJfQX05sYkXnhA4wa9D
O8JDniULRzm43tuUG1k0SIQIqQynOr3XyJs8XEMBODd+k9/RxzSiCPCsUZLMsjvIODmmmJm7vbZg
3ZfbThKBWSZbs4Gh2som+hzyRoeSulPzpP/KUP4Vxvf9Eoydr3WaAVaWEcHyaDaddRva98jpcsLN
6jce65lD81HTW9QYPB0FWgpvy2nsfCNUJ0RfNFQH9C0hRCCh2/QtXLxGWcxtgw4OheKE7jDgX6Kq
NjWg1Vk22DY6AoMHV2cvwibm8YuSFBtbmyI6ClRcnbZ1LE4CJAUKtkAeB1I0QZsuJJFs9zqiY10C
HX+eBXgV2Bw9GOs1imBjXKzrVJ8+pbCuh0LO8+t2D3MQvDFZA6zTOg97YeVgElHEQ6SDEN47JuOv
Bfz1KkI2udHBwxLkV43+U+2r+ZrA2hDkkrpgb3lPFkZs94yuKs+ksB47qCjDrkDK0rS7lREqKD3/
7l9jGARRhyLTCDpuclC4/Jejn7qdLxvkv2tdMLC+G5jxatCCavLF01v4l9/XC2KlPcxOZ127U0+r
KZtHZ6d09BQh984pcWu3ecgcZKjVoJoWvx4q54NQPmBR+uBhBvEHudG2wvMVJg08WafWJOGmqc/P
xsORT3luIzcOckkZvksMcKyEXHl+E+8S55Lc+mkAFRwspBbLJFQF/vxebijdszW6qMozYtt3K8SW
NgPS1DQ2lWEqf+scvd+bRhWaKBYcWAaryF5iZOh65FgpqP7a/0xZnOTPw52JrqYABXVIecSTtYTv
E6scxCNvfv+TPwYjQdz5VxqGYmLSu5A2d7KiRz5XIq4Tdg5/s1HGxIjCAt+ZLblOaTUx8WDOauUG
QdQV8kTnfHoO7EFAtiBdZbxp0J6DQSkka5A9XvICp4iZjjU6aav/ChGwKjFhiwR7qwJAxHUVMjsd
Ftsa3/8jTYo/Jxkjmf+srJEpcTVJOaaE3nR4uiEt0UMVtcvF17mxBTUM1dDd+IUV5ZgtJOq0mpo0
ORp56OujwNa02xXf5Bz1E8OUrHwjE+Sl84dwSEnEFg1RcpZObyJWJMIhW1Q7MGDXjk9C7eYmoZ7O
n7LmXZtE3qWIlXm1L5lWgfp7/yBYr+bmhOq4hzJOog/BvEn1cWMyuGja2osz6zeMOUi2TfGaGf6S
GwuV/3zWF2zJsnqNDfz/znBNZgLm+Sb6BJRtJhpYJvVbxF0Z/N5n8CKnwtunTbaGW+bvhwJv0v4Y
9NjSe6JRLL9q90N+DJtGarQZxuWeEU7d7Q8v6TPrsPC2VJRfFfTWzG/5mmr9ZmLGayeBo20xY6rj
bafmG6Pepi+4+pmb2xRIz6X4iu9ZC79TS/vavnBbXEzmuPLQLxl/QygL4LX6iHghqdlf14ASTr76
xJfYwCo9V9eajU7NK+7+/eRhBTnaYZWpN3l7Gi7F8jBavdb8Nmn0mHRqt2jw+s2HPKIw5buF/VQD
qegHNMd3Vmacw+HdiZ2MNpLDGINyQk+cTraz9he3eoie3GX3wPAqBVZ55AUJr/GglSBXr1I3j1Th
VYzr0UwsnlGTgnya4zKJckqA0on+FQavGSrH+l2fA353URW87FJPx8bn+KTjG2Ydvzan2eA0ZTHq
Bjk0jv2/3fWJLZckd4t/0u1C8W5MyERKfwhMf9mCEmEhmypWXIAJoa8PFQgzHnuwgPv90NJfLwBG
dpg0wo27JA7bl3pUHvvonR/rJ0Y7olSlKckgTTtQW13Uu3lT5tntm4S/od1YYeTG7fRCsA7XXOGK
alaI19yFuiiDTgfMQxINkhkPzkz57TYE0+WlwAciKG987B2x0Bv8z1O2rzK+KcYTALfkk2V4owaR
aWqT/77Yj1We2SEs4Wzv/KPYcpvysqRctYxLBDH4wjBIWQN/GMF6gSJsUoGQfd5gwztmrwxoxHW8
S4sF1nClHk4wn8UXSwKcSAudUryfJx9jBqV9pLZUwo4igFYTETQ+rGhNxrf7M9D9IE/90ck2LyYl
rKCC64RCe8sIfA3gHlPGK9B3t/bjXBCHe4ODJZ2tdmbo14jw+nThoA9x556pT1I/7wGI5EY085Ys
Sj3OsF5u1qtvXQoZDkFVd16MhGRMkXVRoliICrJNwVwVwa77mMwF2KPIFqJCmpqu1TSwj+BioInF
WIvMBIPZ2qNgp3s6CYk3E5kfVRo4mjW30xzXkHpVeYAScHfsoR69KYw9IGuRxG90ZBThbC7vmEFw
C8XN6zOIAJAxu83egecBk0MnFItpxzDKVpCfyB+H9KsAB7Es5nfiaqpFpJp6Q8QvMDPdD4kuP9Jo
uPHcAVG2Wk25/XHKfR2OdWN+f2lWHoORY6Hnfp95chXgdU8+EVuPntudCcdiEoGjNhvRgNwJdksA
G/DG4utu1fXqhO4IFGbxN3ErWzEKAxKnOkdxSizvayFuv4WrzD1xQkEXIWrFbiYpAPGQlQIddUZR
K0REN5p04itQbv78sp1MPwYkF3roJnI+qqmbxwpXx99DNrlp/USrETrjkbvfCYd0kVJulIRlVMQu
nL647mSLxtA1JEtZqJOmpSqtafiD2u7WzV582ICphI5gDX6ciif5IUN3AZTNW+GUb+HYSzCHT4oZ
nKj8SjypeYnPdQZ6vfsGnKCXLHMBYo+w1MEjhcY2rFNt+zZLINFbBcpTwwpp8y27s/9oxJQ988XT
J9tXkFdaPsU99zbDDilwR57JRaj+cpPRD2U8lhU3NDzrFMnIeKZJcxlobTp38lWbyyAtqsNrSpIM
CDcx00R27ZG8nINDQdF3PYJ3aX6ZCg/CGIQ6GgUR1kKK0YG80D6K+3FBqd/+zQF3agFurgqa1qiI
rRmiVLRCBO9haMbgvRTUFV+tKxCp61v0Z2l6Rt4H8rTI/XVNFRgwWAqtTLk3Oq5MZ6G4oILQehH8
+ho3r6azuMMS5XDFInbJv3gtLsvDMjyU70ZBxJMFiX7sjS9Tc+pb5oG+Uet4DDly6EwxHGYnBUCH
6nG7/4nzOnZ4/pW8+6Gxonzl6ofENqbBcZURNLJsxjBoJwpJfyTJKjGIbabinlQwBtgB2n1faJJZ
DDvoXRzD8WMVVlVhJn19+bnS6k6Sz1nRZfQSNZtB2c7UCMB/venLsj93XftHZxBnSuk6CDaXr7+5
cdVCzBwXfaEpfLIdaU5yv7WETI/Sob+HTUWu0zyoJzv6zGiFV6U3AQVF+IR24R4Lt0IyRLTbE0zS
Gq0QLwtz4XVOE/AM6q+01+YLIMjAUNLAbU6IctOSUk9692oVazPGcYwNYzEnuPvQokyOYrloUwFP
XXlTDSxSjTPy8BCB6agY2AsYB4WbkDdFnWAUXdwCYjCHOplJtzafs/v3sbh1UPNIGYxquvDhY8gB
/HDTXQAob5nNevF+QWC7+YeayantzhA5qII1MtdgzhwTWuLva/ZAR6n/TTlAXOQ4w7J64moqh+j4
7pu3e6l4xoMRJ3aJpcmuljwVd0RDBQu5gbPOuyMix9xNF2QvJg/TzABClnLhrpN4essKMJSIxK9V
TqnUEZAp3JqMEnmsjvrieLS8038n+cMjzPZG/kUH9egvIXpSkaaVQ7O/u8W1RyDAa7oUYAy99DLY
1r91gYnFeJIwk06HkiKoUQI+jSuBnP5gXCRXMxsuczttFHMYeg95XqMIt0mJ4+KKMlFkDrGcRw7l
eILevav+2Zq2P2pI62nLaNWMnQaE6IzgFkNc68Cm++BeCT5DPcKkyzwa1k1f9K2BobdeYZ5AX1fp
Cj5F8xaJe6gyr/vRtMPWx7E6J8aP7mtASZwwJcpBg3UaqYu+C1mRejxF/ien4AqMV0hn3dDXN+6l
kZCWl1NLSryjIMKIQf6wC/lL6a4RuOqEzPi2n5g9O5cCJe4vE/fk2uZz0+DqIFdRg3VVch/lb8Bx
mzM+jLQt+M3AoUzNVbAzLpxBDufpcucn6ZXnT8p+fj+elfIfoC80Zt5VSXJeyyulBToBG6Vl3CUl
xZBoouDMEBtLzsRb45K/cLPa0wcstHRzTU8g4jaG3OtMFVPO8+jKPncrK6ZwZ2nrYgOOC3UdJqC/
hgnTQj9dfJiXj/rv2WUuT8JwfXT4QuB/mzBNzLRqswhphSamqAbYaEgNArQOuXGRwYk434S5IfHg
AnBSK5NlzCVGdlFD3pxwYJQ1Uasl70WjFwKL/eH7Pk4rhm8uqcwKJuX3H04sKa/NjXCtVNRsGBNK
9ZZR3K7I1JRJFNOqny2fEnSmyepyYG0yYNC6fSqz1P/9PILQLskqlXypyrrRH5rp8UKF32GDE1Lq
bmUa9e1EbkiWgccShT6Db1H6IXzhu5DSndlVK6oh3NqWSSAG+GIT6t4E7FB9rRK25E7m4PULrSzg
7+IdXqFBZRwKLFtEM/c33m6Ik7aPH80CVt9uzay7j2w4AvnKaIqAjDne1OzTSqoFSmYYrWrqyqQK
uku589VWjS9Yb3an1ImgR2IKVNRRLE2omuOFYLVV3NgQw2oSOhRhLkWKGa/MGkIaMBqIb9SHTxg8
UdC1CvfOwsqpRJOTukq/ufrFkE32EjuntSrtTLTHKfOhzj44bumfiK6M/hHei28w9wvUkiZMXsnt
12EhW58feA3XyrvR4nshFvi+OreCBOAGmbq5ausW8f/lSvNPr/wVa2QF/Si7Y82ccPZz159gNIhx
Qciss+7Z6ttGdCboTY2OlzFzQPi7XjScibRNN6uuEBGpGjbP33Vkv2S/BXtNYjk9xhyGWKkPd+eQ
j5j3f4BJRgABpJKqP88ulVwA+Ssl6XhzLtsJwvE7GGEc1Rr7cZ6ty5lWB11Zd1Df9Vgz45Lk6eyp
ZLYOtscR/+WGaRrPdHQj82O0WA2gfjyLwK11t/Q9tvfhFI+ittA1pGusSruM3E7buv/ivt4R/Wtf
I+ziLKTGq+tqGxCDdkDxOeR9AleAeSP11cRseqP/eoeiWrrT+nk4dgvN4ceaF1KEZovHYr3+d+tG
byCRE2USRMvSDVsIVuOUMEmPyVO8PybqOygr3k+PfcMDltyiLg9XtMspTn3nxuI0uB0vAt6vKeh8
Cwj7WwXXU2+qxHKxXc/Ia1XWle6TJPBmwelSubQZQoN4uDGDIMX+bhLsOsIBYur8XsDfoIYyFvT9
uUvYyr5fdvf+sO4d1wu8OCjAgtW3cQm1Za7LtwyEXWriPsDrNIVHu6AZg28ry1+MN3j3TZhHKsWm
6JDK/fEnuVypRDjYXL0paPc8nWocFJ26If9+XrKpll2t5nOfX4Fg3sDNqSyUrMgSktAfyaWYk16z
WQL3XRI7m2Wd7lbLgHSDkfYqp3VL+ILn7Qk9x058Tj1XMaJe+Zfv0fBbGDtP/rDGUr8qNPQ2YAFm
WAejMbNQF44bZacgf5aSn/TQDf5pDQplRcbQgD2REyChTStKOQRGs8WcDFgjEnKTnvn4P1v7qyzs
y4R7VjE5bJoEBiMyBDe74zXK+Shi+SmGMa4ueHvVIIJqS4eHXLjW4c6aXWZUxx5o9HNbK9rNwbUA
PsiwbTud+MLJkukuA80OkEKWBBoZKl0demnnZixFv7I+wlTQWDM6DXKQkgBRdAJ6MLZ7LLtx3QFQ
yDkzw26fuVfDVQKXpP26AGdIv8xDpwMHvmAGRfqnmYK6e0+eC1d1rANErktAVBVRokhXBBF/NFRW
oDTULafn9Wm/++zel7QWVvXwBLWDVMnCgcyWBBXqDE8yzWTQZtaGQznMD2QWtomhzAjDhxNLPGgs
KD5lXLauyCKSKzHlL8TK7Cr1kPgDqRpCiFexjiWTroUS3+HME0TYWNRFVU5/my6eXtCcyJ3b7N8G
TMjuscNPlUjE/XXAx20FIp7XuL216pRvH0dH6XuPGVirftldctQOJtMQ2CuIrP7waSiv093WdeaL
fUiPVi6ZX8njaGZeo1pwteuGPsLETCVAlRybbo0JLejJ6pgSr93J5AIT0wIb3M1uC/JoKKTyT2Zs
kRGbDYziJZPI0IFQaUEXxGcY+3u4wVNw3RUOVm1oORQ2xnSJ62gsQ4osfdpZm+deX0C9+GRjuc24
uZPf5nluHp3jv76+tG9E+nr6QU/PX0D5ayRXZxJBflfoOY6tEYptOczBcKswHRBd5FbDPE/kpgpx
3zZKThtyvl1JdvBKTSj/b/tJEW4Eu2ZyAxZPjCz+RGPEqvHnQ7ZTuyg8jR6Hh1eVZqQDGhUN+Rek
HelIqx/xl5xT1KPHAmGoDj8lShvGWvynbH7fAGk9jFpJZkdBg5B2cirYheohbyR6sl+jwk31IxxM
zpv16twIYsh4AT97aBODjz8sJ9YVb4u2lZXg5rm/cnjURN0OHKqT7ctLQUQVf0dCML4sP0cvOm/b
ud5h/vWDAdeQoFS/LAJ5S8qrkRA7+Hfe5YxE0gpC1l7ES6QskW32NJ76Pa/LS5RPROMZ6Rg0VtUO
rZzOFDv96NjLlvLSjckKGOccMiNJ//FT9xH7IPWUqsNc9RLUqYm777fFzrAUtiDJXsJukN1hILqK
agVVxC2Qc0TlyGp8B+jUYM/7QUu+05RYkXMPstrOm88p6fKPHknSK3OaW72Fp8NuioDO8/4p9w0T
DDsLfIY9dkwTzqbiX3X1esDBe7tC1zDCakX8ekc/xH3XVLvwgqeWvioHnsAQneiStYnn7Krw/8HA
UxjmqIQ8Zf4culw8UTpBmhT5TmoZ2QZFLv145MyQGXApTD7WN61yovu1SyrGWs91dAoJHP2VWAn0
k70n6WPmHr/u1t6eeXLCGC5cX2OjHHjGcQiGUlTwX1JOySfH7r7GdNxiVo/xmzRxX3i3lcxpvqiV
jfTE3PkSychkp6r+1OwZ6ehRo0u1UT5G+96mGbGCYgNHktVHhoTJb6qetXYRZ0bscKLDlGFV6naV
cxmYGzbxmYMCjOgfYi2u9SYrhmZUt+eWHy9JJEwsEcJXVFA2IUpxq5ZIiv0OtxdTN8MixaCRQ1Gn
Pe+p/gafYitvAc8LguHk/Kb++PNiiOD5bNJY18Mdspn8+zgKRxFSCsEZm1ZUHBAsCeGgDMmoRpMf
sYLTm0MR/amZqKbtrbG7ppDglec2fS1nqzoOgdWMqQ/GaxtmP+QRsdDeaPojk7o6KEGOYXKU3VnR
Pp5gN9klSG0JSMQc9MjRC+CZmGtceEle9G0zTe2dPN3Dp+eX47o7/0Ka0FWhhclx/ZUR+CM3cRqm
yp4mzwai3Q1RazzVwjQCTQrIlLO4qelFlhI0KjF76iCuuRCXacVpNPRNJJeykB0Lf7nrQhb9MUG9
1+oW5eAUTGvwU73awmwFTkLA0k2hSJUuyU8gwhjqv3l0AFntO95XBcE1mwsp8ElIzwelylQXzCp7
k/15GvSWArrp7trga367zoy7bU/BEfE97T2pk3t8O2LSdn2KtzR5+n+lypXKyqC3BroQdqU44CFw
SyL6RJGEKeprO1iViFT333PXZ8j4UXIcLIqzG4YdRpQHb5kSTa0WYbVtpwO7vwer9NhRg28GeIBx
VGDVYO+dKZNOyjR2jDRH3idh/OwteHKFwyUMVN2wZj0pmnuRWvu+4XVSffue9944bfRjlzjBjd+n
Owo1+WLXzrlkOFdAda3dpgoBsqxaEcnpeuY6baaDmxA9SMwZC8BmyqhuTY1L6mx4eWf8c+1Pnt0g
5X8smLg5qWu5ZigUnmK7jMTPwx3zSJxVvHG+Z7ca3Zimlocg79C8SvkX+3aXxCf6/ZQn6KJINnHp
d3VtfKVDOYSxvrqidKOzXn//QSjxruBxPkFfvfF1im7rd+CFXyNz38rFU9872AMaCXUJBtZS/Yxg
iEtjTRwU/2epDT+qkRBDbTw69t7oU+cxW2wvf0pPSnKvYPmqqF6Uk4ImKcBw3xP6h+XHEo9qEAYw
9JJYFSv2YHZivvX4tkJPu4TIs1ys9OUFHBBOLbpvuKgIhvuiMbPjx+GsqSRTktkpIRI+7i8lTA/b
J7hFCVwXi+IqLCFTD2VParlaK9r+eI98VB8+tb2WFLS77KHTSypeugm3I0xa0hfH9hNCEiqKq9US
grRQTazR8hN7A4LZN9Dm/dHpdtnJZzy1Khs5r3iATovwRKKdCRA1yWAVKD3qsho7X4ULJpEXik7L
IWuTEg99hipUztYMmaG9HIs1i4PpEpzLlGcfqdP6LPLp0TSsNlMB5ot3VmIPpYyGB+6VyjwlOs7n
dujqLeRfTGwrDSfSweP4EGja3vYOe1TADIvd59u3wWza6y71P6EkSqp1khOELwf7oY3qQgn3KzeI
5+92iEAKk9B/F8ppd0SqXCUyh4irKTCmCnitlMOANYzKypsZQYcHcXvUDjU3zlmMwl9jEXbnkeXQ
o8GVkvoJmuFBUwxa1oYKnoOOcEDm6XxL5SDXEylEd/5Rku88TiUfDHuFhxCpPJoXzrzmf9/ssKe+
jNlJE/NKoYQyc+N7ZFQDWbVAXPYOg+DjhxUKWdzopQR5kda8oySuEzn9uXvngE7MDrjoH8/G/CtL
ysPVRuyjQttsdETh7YOOjafjhKzVNrqKBHNr9hgoWNR6aOH1eS9I8cv07wofpC8utKHA25qn7sBx
KMrpPRuccR86nV6kuv3mxBPO9BvFsw56AqTzAmkK79ITHJAC1tHhFkJ3fVvzR7rT1q90kPGNC3gm
uia6NsQI43B3IvKz0EEMOaQ9kwCDOY8J/s8aBvkjYQ23TqZ6uC/fpKDktliWs7FLf7nCDFRM3Qb2
2XLgGrBLpurRFzvlXah17OWCHqED8rWYJKQNc0JmtH/eA239BTWNhPygc69mLLmLZcl1KC8XhKDT
N48ccQYRvTiVPoDpIQxdTXC9ZloBPPmCNGJvHtQfXxxfbkVVmXByNFFLVbrOxlFjxhYXum8/k6ZD
rHY1zoACDabH8wrsVZAopUylcgmslQK8sQDoQpAX9VXhXT4KrRI5Mym4yQRSyc5TXemLujtX36X5
YZRldCltERCuKpU08fQDeWa44LW1DGXuG2E/YkHWkUwLY1wTOokRL9i8jKrfwPWmZ6m53xQoX00K
9dui4OWXPBYtYQhxLNgbJrPWMFwcLU/onGhLY5iGdghtXpt1xq3oEeCMXzGZ9GFon2easrZlO3FL
7iAxBnc7g2SOEke8tyEA6QEhGEXSQmGegQuoRdJUmGTOfgibk11Qg7ILoPBdY6ePZzQNMbtWef/J
Qtkhs0J8cPNVA5EQibjv27wSLxEdXYPS4lj394wTm9Alf7++PQt0QWro13RXPoDLwOKO8Oj2dk0S
Ul/JpFxR0Kr+CwMwD2USmJlV/kzU9iVym+nfHN7AiOWZKcHfKDAUhpORUO4nM12v80xkIJnLbCfD
ZqkF9LG9qvSA7hzKaNcZ08YszwBd/cYL+LF0R2r6TXbZPSrSppdPVotGOz72VUb6zrjVEBTm1/sN
9ULYfaVeW/nsCXAWkwsPra0hyUmhGMmCb89rvtyqgxzZJNYoRBmFkEnUoSg8J4D8pVPRe4ESYqBc
92BUtQatsEO2L4OB53bw1XzDQhWdgwcZg+6MJWWNqAcnim/sMXGC2Te1maqVwgt+2gA962272hOQ
gl19/xU4Q2ria5hBeMJbhG7Rf9drZrlkizxK7pimr/FxrUDnQ2DU0Ss8cfhdp1BA+ogZpfAxsvjO
mjTiEGzx8PqtCOlCq9vXDYpvHy3vWuXdMc6V+RDjiRj4y3Vc3E+3fiHzOGiC1C/oVbPDeED3xIE4
GcTbtKgcVCiCH+GRBeF+jR8yd6RkO4uxVOnubYTYrYUYSO4XuFOHU+eSwIiVhZd5BFQbb2ghz5Ql
+WnrpsnnmkngvZKda0y8n4rCJxqoUrAuxms5aW/aFZbcVU5BsB4WMPByuHfZzruDqimZgoYpAYvS
SLGAGDcHlEqFcfKKQ+iuuho9zyAl/SE73LnH0GCLKEJmha/JQp88Vd3BJlkgLTht3UKqzKxC6zlc
AKZEVtYy4QrsNTHB050aKNwfuO+Aam8PUI1myXp2fuT6dOEoSLqoRUni6n6+LO3Mx8ZiFdkOck+I
Nz7HatFZkJMH8DqcttdgJAZp4CgpyyppP9FreortivXKkBhxSmDi12b1fyA3cF8UWZNfpWrRaBZt
ZwkbTD9qbCl2v873YyRRKkwCin3bkp2McjfTPD1RJnAAAZAgCkJoM/9NeoZQLRrf8BXW/6VND0q/
ZMyuX2ZJahueQytTLLi2TiF9YrQ6dxLajW4+eVgUdsxyrhTBNdqdeZzGxc9rUH5IZGiMdyDw7SoD
ftAX4FN+fq+HGAfg3KS/p9Pml1MLKihrS7z1Lk7f+FmkZ2ItkOo58fd6Un4KyGco9RXpwayQ3kb4
L2SEIt9kZUV7lMjYPirkw7ZTMujTu1Ngnq37Nc8FO+r/N2rboWKQIOBsxTKjAqh+tRjF3BgiNjbo
p95CKcn0QYGQnizRerkqcZdj3qKHUYQU07D9gl1gKJjQfSkzc1Fykp+L/9NSYeQ2lKx5sN2DTQ4X
zpyj6k73c3S2vfAfWxFH1Uh5HHtARd3Jgia9zj4+qJiZ3yPSxSLYmJBQniLZeXDeKfT0pAo2uAqd
hy4Su/J8O6NY0jdrP6RfbmQ+vijBEDddqdYVlnO55erMvtVkkdIXcW+T+++HyK0dTtn65hx7QpOC
F25i9nrDkCcPQSqJYXOSWMW7xOxbl/3sVbMmeG62wchvEZ1X3O71T42rGqffUC1iaxK5p/uMZg9T
e246JoGjbCcQOP5cuvR94c5Jse+TofRts+cLCcRPUygmYGHlq4zlJTKA7xw7rz88By7sIpm+Opwe
IYJ+BjWLaCafLIkKXX5fTRmDQKukWDtsLXVzBJl1cb6Wa7Qb6eKC45nZzbkKvoBy1YGwtlq09EX3
EcZw4kVPK6A/LQcV5Fb62GboO09ekqNGgkCIaJzcXs6ZCg/3rjeivCA2IyR2cBY4VpyjIAyeIZoY
F6nQz+uFLF/sNdSiIIkTa0yDsZl+vklbVfRKwV36O8sytXBstKyONnM296RZhXhJWwlPhYb8P6hL
+qaK5cWZKNYAsT53BBf8ciWLQygSQXknAwThsQwgJM2Llj5cURblwri0yODEhVeaD9L5KHLgFAnd
jA8Xsf7IXLyLx4eIJ6h/PxDPKQgbYWnF1by0XU25pDawF3xVqR4OlJM+bymuYk9oS+RhsKaOO3tp
mEsFd6+nlP72tuBkulMLom2uK1x4HOPh6jpyxXg/SHIhfOy5KWJnCMa+BMcGMtAwQvxN+KDxeUSf
x0ZAnZVvZk7FTJkS1moFcWJ2DnClegcmFQ6Hdi5r3+gb57s7JFhkMGCMBsIlN7MNBgUb5ZxTOw/+
ZK732uW66Qdlsl4dhzmo6qcaH4JLU97N4pMKNWzXeajhtbQoTAQfv2WVFbyIcnn7WCxfkCp02yAR
P1Wmj2x1LdrgjQaBgA7RhfhXZ08PGEvBqas3POLn6VaC9/svSNlrvM0MNG1b84U2om6uJq3964rf
sYWQmkfPUbYSe9txagkCjG+USzMFG78oXPJxucoqlVAQa69W4IUNWcdYZVFiBSM4ReWlUMfH0fmQ
RAbrFnPQmx3YM9CXYKNb5VY/nsXRH7de0x7qCd90Hh35AUYvn4Eb6ceDvdr5Yhlxo9jLB6eo5GFe
MAvK7js4u2GjoCIAh4yY9MijQsE8aq8RGazBSU/3Xu8CmpENCDfp/dLHUFVCIDAm1L5VlWc60Qg1
XR1u+yJoKs1Y2fNRRk4MKgglXpdHKJJFu45oy1wk2mUCSNsgn/TgzA9nWNsQkvyH/w4NjIwHJEth
2TOeI+WljXjBWzoIbAKmn97GX7iV3OWBJwqgUvbIj4C3zWTW5Nk6HrrUMFBnuyYfrIYHRN59FMDq
yiu4aRCwvvXMYhfzr1oMpEu440Csd8eCjKGnQdjWf7Z5l42nVJWZc/nZDwO/LA2E1G5W7b7fq7RM
eHRkFBuTJTtIJ2hEFnGjmrd157ubDqgsoxITd0Sm5YhTI/Luq4kUTemREV9A9xbCTAo1waJXMouW
IQUgXlWh0cqR52o/ZqxdEyty44rUH7rN7DCVt1RE7JnzRVNH8DLsTxOY1JHWdAoAGYRqlerKenT2
owIqGsB5/kRcsCsfptU9BoU+NxZbYt2xeTnn1oLCypTFysTh63Ci+A0TtDPaiOH2d1JT2TrGiTI4
0gPySvMfd587RG3ARUtUiCu+As4yxQ2VL8uw53kbjd0euketvSi7MLH2SOEtABHtLRwhZUiburtN
4K5brFN8+GItHKMlqSIIsGIN6TxVXVKhFx9JgKhbTN/THKsDPgAufztAQG0zPDl9UMl6BvNLfbNg
zIoVtm6wSsvei/HemLHUYYB/BFe2kYXKRTiDNOGIjdWDfuui6Lrf+X2i6iyrF7sIy3Rvxj2q1sUA
NMvKLp2yQBH+xHF1n4ijRQU8CujX15OhNWfaHpebHx7FjAc+LgT3P9vFaxb4D4GaXpTB9UAB7Gec
2ixiBpLIGM4mJjLyPQYA3aEFq85LUZ2+eS/ZC/qu+JW4YTrMN8AuGsRF7vKHb1Kjrf682dgxePX1
XnfkwM3VA96fkBTBNOqTHhCj2ElT5cWyzZmana6X6L7RQB7Dew0DOqSHEb2mcX69D596FnSRlFjp
8YuaxxopeVnNZko30qPE8kNuUgKBDzxdxpZZOkSz4IcNSx80dH2Iy0JvobxnEFuNMS9guloOLwwG
BSbtqtt6jV9Syoc5mpNdkfogeu3goXr9nMIDlAVLD3vDfJkBe6Se+y9Il9H4whPXvEBE6yy7xmST
QU59g9E4ZhNRuukPZuA07oTykcbKMqyQ94RS/ox4gP8zWDk9haAZJ6W2SecrESUhsbyM7PgwTI1Z
oCj4+Mvb/GtjvSyBmluhg2m1mvrKM2b/8WeKZSsqbdREJF/k2Xzo7Tt7MA7oYrBUb1WwSC6JXjuS
w9geVhBY4L7HTjIXbwwbXeRIyeZdqF+9AuR5haZe4fD2aYyU05sBMEC1RC24WU3qQ0AaiIFaT4Dw
tZzj/gR50ukCY8qBlRkG8jOIqOZXlSlE6m4GYR+Mfs1HZ6CJCy0MMr+TY314Qbbh392cvKBL8Xif
/KZA4q5rCMxxnR+GpSgNrANUN1ycZnWOrFB/ZYYD7nxNy4nXQITLIXAtERsYto4JFJMw9RRO1+Ze
E8wOJHQNvF7XNXtTG29LV90GaRZBdWUXAN+8BgszGN0In11vy69qD18CS9hPGW6tYWmyHjj5p3Fw
cGr27TSx2OWPC4UDiVaaQjI9Ywq9xhv4wL0KQcPj+Cf0zRVdr9RWbzDgB+Oe6PKW6G4Ftja7RM5b
mey+rpmbDVTS+iMkpRmAGgHKFIx/vkJRoUghve89NeLWGL0DPbMSrMdHGRVSbW/c67lmAO6NPrNP
juH/qpe9CV44lSkmWLnw3spUqEg+f2Iod610+kIX/L4vqq6VWKS0ggc23AF+1I/S5rhORtOYEyTN
U9Tlgh7fgCbMp4p3WipJRP9FaDb0AhSRsYFPMyCSD6mP0RTDk7EkqadQ5tfcVlD0J375OunMQKfm
DAKynwcIlj5OvSBCQJQLYho2VJ32GDMZL/nZsb6SK/vjWetSTdnKQD39Wf6RZy9GbDSJcA/1JFFN
Z3glkxJT/kPtfih3On7Av9Pj4PEHmelS5SBb7+/YMJmyBY80i1oxu6jJgRZMYxnK50qG/92wOJPE
jWEc+jfNdyHvJ6X+jGsXnf5JfdcfZ/k2M5qQDdYOK67gS7YoUUo2yDeWxeOjKoIrHv4wfarvgTmb
rMDcL2dmabxyEHaTpmUj57vezWxaFJoPRjr+fongMBBhMV+Rhtij7d5qGbYEiHG0PTv6ieQN7emx
r08rspEghJ3FSMxRp88tn7+lWyysYea9b0x4YO7GtgFp7bm8nbX6DosVNGSDMAwF4yfKFRa7+Eqb
TiPj50Pt34mldGxlabmEL8qeE9IwXX8c6o17CdiXhhoqVAyn278LQR+KlV63TP/ZeLFYo+F94+px
5SdIKhxH+BIuszRWGEO351eo0kGgwKc6xjcRHjGs/if4Ec5Jt9KABI//ZQD1xJwLJ6GWQKUuuuWW
+x6EgQ3kQvk26nA8oo2rPjp5a3pGZM4uVGvrYV5PuIikXpj70c1rc16Ww/LrdLr3mdYel1gb4VAE
+0w4KsuG5Ujm6MVU7NY/qVC210CThsgcyAt7Dl9M4S4FFWSTvr1HFCBPHE12s/h5vHuNdn0SaGLg
7vFwl70myPLXYTHxQi7GxqijHJ24yYJ4zuieyzZuSXuwE6gS7W+/M8LSx+8qt18y76LiKS6n+rXP
DODUkFQqv0FkPrqNf94f9sa9csoRWmZ8Dh9Ze7EBB9VY+ArQTBUH6b4ubaj3oafmq4IMnf9j8kVx
U6Qc4LzUT9eHQ7yGlj2Ynh3FcxOIfi7DF1CgAXshvjzrnapBiPGy6TNGr/lgDdSJqC5y0XeGy2RC
nyRAnOYO+ZkLKMeCWicrnLq6xGQqYZfVjAmegZ9ej59xiquBj7WFOBKw0xemAXOgHkTYyHISlnJu
MbtT9PS5ixWXcBwsl1gIOBQtilyuWZRygwG1FSveuYBgp0kmLFyvXDeFY8nbM3j5RM+gHadY2Kxf
5Oz/TAqjx74mNaESIvuks5731SY1LuETjBQzmmaVE9uS7SRQAnSNN1ByH0254UO34Y3ytQSB8vv5
G0I7zN+SAfP18hrrVnFDDWkD22e320kaujNw8GLMieyrJgFIWQJIR3WWfQx6jGwGFlM7ptrf/nNO
/ZPesAYHsherVMjDGC5setkgktPPwRAk2PL9Dykh7iFTh6yMQWY9GQnu4XncQ21hmlrWiaTaebg7
kRwHVkcgBos+5tTozNz302BzY9zgq1GpzsllQZdmCPf1z2P3OfaVX/fRSdUURA4mlIiXrTudeizi
pNPtOKg39ByBXPgS/85z+gACzR5Mf7GeaS10ERMEYYy8q3ARUVxYW98dwZuw4zO8UvWIFdHYUFl1
Hy88Uc3Hq1rWprxYFg7t2ebrCp6PoJq2nYaIYekPBvvFqClCSvK001pUf/YxxhExMPCMn7pvBZLu
SDgkEXveZBdTS5jJu2Y1xSFhjuE6xU7PZINPOt4SVmb63a9Pa790KBEL6lUAjzFYFLOvEIocqzaL
0od8GQHXYjvpcSX3E4/1WoWsag4Ep1sD2e0jtTDhT2MoOVlIMOj2xIRfY0j+SJXOlSKpeqKodpoR
rJifDh+BBYfLwASCBvBBfYBWV8oOnh7g2z5qlkRVtd92pen+EV2clcqKh1ybj7skQ46LpJoYMqNN
B7mCaiNh/pWBlpXhFfTsOaQZoyz7sMIB/kbWCwqCPuzlvOzjrJtWFQAsOHvzK3QFZar+2Tx95jqP
ZrR9nfEE6a+H2STHMzuA82z6DfX07k8CRVQZbMURlkKuxJtTONg0Rq9m13FbJVSYitZe4QrggZl6
AdFGNriBjkFWfoiIGE3gUoKXu0QjEX8NWGwkSPAuZCNlyNhInCav/uEu9JuQKzQczPmxNbvkkou8
JKGXNQChpFxPCBiAYSrnkif4YyrF5XTZBHWybGF1wPNfRXm7RX9twClj7Y5oD87KNKQ7Q4jirwg/
UUxNphYkeqQifTu2d9dGkb9PXlZaQKsXkglVh/1Qd73NIXCBa5DjXU7yAJ0B6V8p3Ny/z/xf6w1G
QB3CloNBgga6e1YUIbznTS3Nl6X5rCC49v2MSRZgJbzh7vG00ClSJAx38BgEFQ+l7yMs6HWxbF8X
/zJ7dPIWirKi5s9lqQkvQSRqg9WZs87QKcPL15I2uOXO9TFYoWVzPlASSuwke/QdpAR3brtoBbfK
wA7X3XJ1Z5O9b96YfpGnYLmfchTnU8iTtlkBeTqXzM0vjN3vE2Z3BNW/oVlfibca/9FnbRdBSbH2
liVfaSpZta9sl6LCLqqZo67Hm7VO+u23+s46INrpbGMvBk4muSSYFSCtVfW1nLST/DO6dhwlvW+G
hD5krth+vcIHUDvjJvgi4M72Jh0qsLgwwe15Hg6RvNC62a0lBA/jcJOL8V1Tb8oInpiMNmPJ79SI
plyXAQYDW9wOzegEiKTiLf7NBWkLbWhYzUGjNa3xXIdHIUHCXhCp9pMmyOpWKZZd7cZ6V0zqgV1p
/DNNjNSuHHY5Mcmj+0ZDEcTa9TJ763k/lroZwoFzym6uWMgIV9tiGtJY0PKYZmm4CNORZSzcuNJB
XmZxSttALHsKEKj6teQ1q/aAnqccKNRhmWtuNBdJKVo2kHczv94++ks+3oTFJn20hVz/9y2UA97h
CfSiINMmF6qh+mVvBdUKDPso0OEOFS0rMwrB9UKsK0AfWyn8LtA8pINQDG8YTQeDYO9cFob5ZgAq
U1a5d16KCE3BGjxB4HeuvoGavJxc3vJhyGArjbAHiofYlerGg+HNMPQdXzgEPVK6rtlcvKM/AWpH
6pwuhAwIKFiYY80f0nUOK0tC4gFI0hpClAJiQ1uJYnVDIAd1UDZZJD3pfVBFpCPzvMuYhSrigmet
aLTYSxC4zJf/YIl/upoCNy0HsobM+CCW0YjoOpX2ruPayWROcIY+lZnkCHX9iz8NmySjfihS4l1P
p6sRfwZaJglz26E7SzvsfHqqjTO5t4MiALwTuhZdEAgLIGGAjl0rc7Rj60lYt2oOQv3196Nu8b1p
rIglPbQeWQOyWLFTfrzotLwe67ooDEs+Hu7FNnpPSsnOqpetaOZOdVIOSAMK2cDIEI4vnn2YTWFr
vZtmHkt0R6tF8hiqftgDlFF8nbsMUA4Dn1jtcf8g94JLZTEkrWr5gAbmgG0/aHUUbKfKV/E2UBL5
/TvSvH4pNL49a7Ucdq7wARVsEb/p4Fwjyne+sADilfiNXAgROV350KlbEgWJMsGCW9dc//m7BYUT
DmiqSbVBVxJ0c4kgQqzJXIHwewL7kPx1+6K4W8eippuLDtzL1wXgzFTC5e+YvZMssHYz+xR7byI0
nsFrWfwvwo3WI2BbCVbj7SOJPf59yN7kLX5+hs0nKmChq+SFqM9K1puSX+1Vd2u8DAlomhG6WOSl
qm3MPvyJEtlfkpU5UflQ52mivr7y0tPeGqUGV73fE19a6fLrYPntZ1yeGawceTYGufDK4iyKflk7
59B9EZJDvtv5tEPULZBZvzXo4aGLvi0n8qB3XbtqbKwscMuZXQ+wwM+XLFQvvBBWvq+cZpRpmcsD
lAQs418LuBuLq0Usr9KKZn0SEss34tBtdECifRlBLImoVgxlrj/VsutC7IY0NBrmE8VSMA4QTv9A
30gP5ZnBHJUXRlksALt+909WCePDIhixW764WhvKPhjhnPM5yUt+OAQnpJxwI+dSBHqJKWbjHFPd
RZ6sZorZI+sTi/b/SVHYE68QjTJdtyiTKNSLiGv6I3WechVCTt9UMCoKiRJ7F4D9z3UYMJi4MQOy
WzQqTvuQn3LsgEvhlOHcgFX4uPbFm6evbaSvNFxhrF44u0Snuuu4C3NmwU+dqw78zXq9/ryLf9l7
ra8/2DI41HPBGWlaEe6sdPMXaWlH6Fa490lrNSV6xXVCRF4t54qbFANmxMa1Iu88VjUl3Dx2Xv2A
5lb8Uj/nAAimHRepdcR7qRkLLRr4S+Mb814nFuCDWvB21rO7ZDy5fOteTpkEFQv9YoDvMaAc17Dk
AwdFe+9EHqmm5omEGTOtRWiZT590tN6UkmPQQnfn7d4FZ+gIMWPAUtiEmWMUp89AxC+1o53hQgER
UA5hoR2YsBzAe0wQF6yYeUeUb7c9FoGWzZl+kInSQwyF83g4U75yrpw1VmBiI0tENk+av0oY8YGd
hrDAfYVsEt6FXhLkCN3+LhtxlSUjLjamhzaO7E4pHhpYIEbK4O3eBM632VU9vCeuG+WMPRNjxj+W
7TW8Mrh/I4YpDONpSAUnyAg3NxhopxIc5VfMNJ5dWiK6otPCXArUiJ//IvlZifHCGxe84yVrd/42
dbLePMsSVaF+eHfbXFQEvgp5JFXvlsTCAr8V/CEAanVdMUQJ/4Nrfmq/3dYx76uvlV29YZk5jq4t
h/kTCRBXi2U+BWjudg59OjeP59cSDTwgoASUSE7LIFmqd6Xcwb9+5dcx5FTyXc52TzZBcDEkiR/s
mxSYVrkxYWxfXkPh4fjM2PTGokQlJYN3zVl+HP+M6joFtZ4yLbDK8v2hBltiJyCvs3ezzAkHKalb
hLSpiMaIG0n5PBo9JGc7TL7ajaRzxdXS+J0nFa0SjHxJLdkjV8bO67PJwvWD3qh/sk5BaUcMwyUw
QuttLzHJTnBRqIAW2vQyOhGA1DwB2ZjDbgXwlFob0/mvmdcpxM5ZZzcSqz3bfDbSwWNuoaZ3uQIC
SHYbOw2x5n0e8qcd45apyAUGemoE5SaPzkHyDp1pB8Vwt/4YTLsCI4Pvvz486eUESVdYUHKYD9By
lLec/vf6Z3cnOds2Th9LIj1ncUvf7R6u+jeIoic/s8LcZNgeZBaar1AYFJg4LDyqjIgO1CDA4IzV
dPuUDZr84UBbzGlSEGkZ+Q3OMWARM1r3GA1jBh3uysqruR39H0A/SUGl4Im1BZ78ZFuMJeoRnEr2
+gqTFys2UKdu7Nme410HkL1LqkmND75U4ffSKONBJaj0YGhGk/4/BKY+JnvLiFs+/2Q791Yec9xI
ZcA6S3GcW+D8pvC1xNTf9s7wZKzIUKPHgp6IkxvG+NUiUyOWuRikQri3pQttvGUaQTrZk/KpQQ4i
vxyJrvNxTAwMLewrJ3nh0+2Z7mYRPVCYIaDstHxDc0BtjX7oCE3ofmg0mdC7xo3uNSCqMsK8AOaQ
o6GrGL1irQAMXOpEyq8XdTwCGjMjEtgaD9Py2eVj1edKecppxG06iCxp7dbFAH5KDTOQU3l0Nrku
2+oiEfTfpCRyiN7cihoR1GSlihIOI2d6HeXgYod9Fc0f+t1vwrNS+zMv0YNhDpDI7cmHZ9jJq++d
8aFFUdyORUNPHupdiMIFn+HrTplnDSKmSKBDZD3XepQfWMZZANJldo9uzSpht5/QMbBRH0hdxkVc
KrX5hpFPQYlnPvYYhX/DeqMNuZZTMMczYrDVh0+hhAyDC4ST7Kvg3g7q+Sj6AREYGi+eoSLHnyOB
kmmvFMvC3ems45rDzIqltuQ5im67QZKXruXwfaT66fVIJEj/5GmwUOrqJk2wBh5U+eLk5rFYSdIR
Y8CHo4aDOV0vwwx9o5cj7gbt8PVeRWvo7huOQkvRQrwDMV+WuUeKgI9FnC07W5wAfVXNS+OqgDRL
hDYU6b8FNIq3ryHpgjkSHHSld4sGvYhiwJ4NFkKqolGVBpRrHikT3v79d0vMbDhm41exjIt9K8kc
J3yjjHt6PWC3wZbjx3Mg2j5rerrLEwtD+m4FDihtl5dPa0spRzf2Mqh9dTWNv5bpRHqfHZHyEVB3
8NTH+apS2cSBAvoUAzkNOFYPXMdXave62fRfM/yM3oJGYHM7uPuukstkMNKVytiQZOxLwsa2FPvb
RcrYlwxfMeWOdDu+OxzTDHFyXeRXpPcIiy0Sx6qkHvHFIlFAe+P7cmOIseFAr2krwuW6CSBDKz60
DExN8k6lCKw90iWzj3G1NzTZJpIQJ6tZpb5X//7+fb65z75ELEvb9eU9F4gupLolOZtmzFNmT3VQ
EUTp9NK+5ZzyRNsRnQuWtzylqKLtqud/HxfjRQVZARC9dnPZsfuUi2UEX+p+FkeLogvs4zd39/Kl
B/4qFqqWZxvD8DmDes400JJ/aAk7T/Y0dcsQOJV5FcZnygmw4nUQ2h47ROz4kbF8I0mzE39SK109
7qTLxtW8M4zwFOY310j5sUfWny0Zj8qEhtRKwraVxGmMilB7BhJEsY4d+A04F6yf6mT+lRvVorE4
Wkwu4JM8WTe3ehse6P8ROoDSESx9l/SqjZlaOD4h/OysSK6L91tkXL98JyWKs2AKsvJAUwEDmO7r
x69NiNylS7OR+6TwR284x8Rq2eBp8YjFfNvYUNEuBUMUqu37TuYeLkmo2ennPrMqJEW9u0wv3hKD
h3gUNVzRR/YXQHk0/6Po+aQY3s+TXHZtdZ/QZluDccleotIlDQpDXM7qyLYm/hYQVLj67nIu9vHG
QnekabqLJHj6pRN0EGihi8WJLFn6VkHIdCE3MDVWBNylxpMXTwLIDuXRr7OT8C/gHjNZYO0w/jC3
aa7zQXPKIc6swT5M6ViQ3NKClgFrLdLGUsDVabjyjg9TCgJP6YoW0+TUkS3HPMy+EZ2cOL2S251B
tquM8ikS+zi143Th1AG1RyhBJKUjYT31MPGFNQhGgVgDNoDCC2bBTkDjZbLaltZtVfxURwq4njEo
dcX0jcuBtzyz8qfTvm4/HzA8c1VjX8YB7/rmW+4FOBmX9Go0kxD3fenn71GNR5uZlRFNFsLklW0r
66/LvSU5rVlx9nMYg6QF9qPcvp5a/3tWdE5Uy/G1EbYjMuldlYscD00zhsq4mmtKinXezjSCnStw
mV628ZGtgjJQFVDMO7LVLu6+t5rGt3jOcr74UwKKsBZ87zYRIzORZK0OVscUJj7r7KQ7vJDixOtA
hMq1mEVrxt2wby2p/uVcZ1I/P0esXZiLgGDajnc8fWqQvrf0VnKphC9TjukUlgqD7hqIIoGXQFO6
onF1X/Z/LZ5pq+3401Z6OneaB352z18hbN1YqPiVyCP+++gLX7qxupjuLIwnq1u7gQmoUhqTdr0f
JfBo3PToFha/4RTxYe2g/AqQVpQpW9WlOT3ghtgP4igt9BCHgQWgtrO9ucrb+jn8phwNV5EPUnZu
cPkZLrWpUdSG1JFAyD5zuksk7p7nKqiu51dPB7zemC+4bebx2u/XHIrn62ivdv1NvvSICJBPyEVF
inIRR2HbCp0FN8kWOZwsk8WctEXXTntpp4fu85j6zeMqFUy9WTY+PflZ/xX4OdBnTZaSjIA08Ph1
fdaUY2vXeRH4Cn/z3gXhvNMvZ2Ygwk81p6s/nL+aiwd4aKCnW5ODKf7cGUFasktfGpUkxJWDUvuX
4GKE/MwM+OSwqk0fDngjw/Hc3drJfP4BZKd5e9QFDMlETzFNQcUVZR27zHQi8romDxHqeC8EjsXV
251fwuTDm6L47uoZsJBnmAElbexMednd0U1tbQrXVG1uwgxdF9gYuf9cgcfKawuBtrkf3GUmp/ev
ak8JgGrN9yR4g/WTLnUHkrM0BgWt0Yc6ly8JeQiscquFnH5V9bfYvsQvQzylbq1VcCYkcD+ymxru
leatMZd0As05LCa8xb/YRMqMXJemaMqkBlPqhNR2h6eblIcaBxX0wJud9IJXOP0HlM/VpUgdzdF7
hVvNUzUHlhiIU+Tc35EUNr1XvzGfaby3RVDijWhvRZbndQwQOl6o2jcmT2trySnv+xFxoRtG/25b
dOFxPuBEVEpHjvE9tcO8QOQFPgwQd76+k5ysRZYQ8g7BWbACrN/pCAxa6xx+CMzQowQ+y6+g7rFf
tbONJ2oqiFImv0J/HH33TYhBJ8FgqNk+SYWijc2Qq1rKERWDiq03f9f8GuoX6uIpGvpCDZuOCwXS
mpGIV/+ad6DnjPPHHuAbIsHwM/IKXRb6tFrGkm3MYPi7cSdpPJ+cpcOTgbnPZ2a7D70Ww/jYGlyh
aEkTeQpXmOrQ8PTyKiQTNo+IboDWAhox05zbBQ1EIuXnaGixERb5fedFOJfx2NZs5DVG3NTy+qak
UEJ3DwpVH3IPnKFmQr/WSZhwp2ZcQyXT7n48fITLVt3U9mFyaj68tuVllOBpPgkJwEsUCXE073sr
/s7OljB57IgddrL4x8BJomfxStFokh4SL9HxMZeeeeouuUjGx1xx9PSlP33VnZWlI2f9BD09C+QE
NFwhhzuM6lLh6BhKzB+2/5NcfZ0R6VMBNRshVUHLTRplMVrsTRQZrpLtB2LZTsy1lKuy8WZPmvlF
NfvBgdnUIod2kOhfv8DO6eiEnyF4TPdyv1E6vf5AM1NWvtlj3An+oU3jSWbxP5xZ+Q9g0K6v52WO
3Sbke3f0PVQtFiNXFxReRcezrtnPGeLpfAFY4EL4Tjt9IJz68ngaYxQBi/kOwXQS2LRXCwU7IQBT
1EzFGOE7GteQ7n02u2LcWNm6r/AacY7u1r0QgfS9fKWxcBMGeUxXVJKUvvvRgGGmcmiFTpMObcf5
tEo0xduu9SAD5yjVCw1qLfH0JJBketNB9Ef/UvqHP/2UQt1RMVWmGcocgSWdtmj4vzex0/5+Vmuk
6TcB+rX7uVo84KsHlCeIdfpo6n5ovO4uBjoy7HVbYbZ+qwvn9Q5lBNTq8/4GP0qct5hNG72BNsqB
X2FR1bgGlz+r3wLvtCd1GSJzMnnkc3V0jc5mEIWX5rA+j3TboKH5JzKOUa2F2+yfkQKsI4XqNsg/
RZKoazB9UdHffdUNVIu9Sx86XJoPB2qEV/IWM7bYXkQWo8YAMZRSpaqtEn+bURZnLFV0MqawWye2
D28Yfr4YEfLadUK9ob27+OhiV1OdkUvIGgcYmodHphdSqbAJSBuxUIUcjem42p6aBCYEyA0EZQme
8wcyOVBcqW+JNdmKbQQAPCJB+AiXwFdD6lVv/LSMDdNsjxslj9AtV0t1IUgGgFzIW+frp5xh+M9B
pjc5Cn5xz94/yWuygn+edZ2nM0eXIg6WjXbqSiQ88gCoXi3BiWvHSp+njELkTX14OCDNfqWJ61NG
f8FkprwyyU0Nk5d0dQqg0S8D2So6dkNPq3m1RsVwffMzRvDysSAiffLs4qpW8YkyRyaVJJKxvSA9
PnX0tiZxlbVcJBiIbwrby49Qvpxzmrm+1o1XThCCc8fphwJw8+a7+0OZGdq/K0tjoTZCIqQUUctO
IgH8MAlVl5WM7Gc31evheCjUkndfHWYPiH//F+U+zLKDQcKlSKXkOkVYd61Az0kV5c6bFsqyRDG0
EQcs5OoHW5C5dKd7eZ2BrkHeRzE7mQEih2LDq1c3cVfvZIvU78Vzua/JzKs67lzYqqNXaDKwHfmf
JVzkguaTcJTYco+/1Goth03kZZ2gZN9N2SzDKvqQbuiOyJ08Qbfobj1n14VIQjhtIdHtCPo0YgHT
2RU/5yZuvrFh2iqMR1E1pZaukfF+HRLZWdY3e+gjAD8zCH1EnKNp1bLawj8FHrfbEMDhHTkmU2od
iUDUm/AVgSZbI/XvRDoR4KjajtX/mE+rhkLK//eZ0x9QOR3Ai4u0YyUVmY7s60MA/8b1evlCRf2j
aY3haHbmAkeIrx7pyqXjNShVk4Xij4IDBIK7sVwcpFmYxuWmJS85OiT4zRlXtNahY1UuhHIbQGO7
usK6s0WP3yYw3LVN/ol/0mJearTZDvfDeq5OPVXzHyDZP1no+5gLkFGdF0dKqJ4C3egwWvT3I9wV
841815EEPwIxrAPNFyAAzpwD638339PecogziZ5BPxOSkSdTc92ZiKGwEzVyaugkYbXVe6H8Bx6G
VDCpZQ+kt5MziZtP8+ZUvcndJ0T9kvg7JhGEOZQ/+pPnLjeGnt/ELU32E6jAd/sjUwWR3oCiPHfj
e+jCzJJbucn25MXeBl1POWLcdS2g2mi8m1M/36u4oIuoto9tLje0qFDnzb1KLMmuMg9yEj0x6F3N
MRGz9p21DVJY3gzqZxhr7eZIWrD5cKKV0q0m4qEzj07kPv8sJeHa+rLKdN0+0zzY2YUcc1o6pBQE
/Hn90+CDbCHxmZgXWsJtbSsKK9/rEmL9NQYzgQHeOo5XBCYIL0CPU/O0KNrL1Epj2pdsq62PkQut
duH6ObMTDhegWX+tO4wJc1yxJo5yqwRqSnOzaIG74joUtESzmJQU8N8ETShQC/J5FARW2QScOCnJ
AAz14DJDgLQTcwm2zNpElswN2YKRG34D8DLTIaxQBdRSxreM+nxREDxOcbuPalyK9+1wonil4Yo1
9WD32yMUsC79NHHvc//8dK2D9c4D2cc9TeIz2p+dnbGZ1tVWcRVVRy2MCfP66fEdfGRFTdbJiXsW
G26pPAdza6qMOU1K2TOEUCE3S8jj4QiPIqmOZ+hXb6zQr8PhLOYa01ohqxkmzIk0LicC0gO0vrY1
NY6ObjSQGV7jWMls5IihUnb5K5kxFHlJfku7eE1oh82/QJRIKMDpwNcMCOFEKFXZWlxWfNRXasnF
54GzjdNw4AhrTd029Pp8JpcCs56H8I2WRl9QUoJ5WWLptEzEKspUptAqEbYreApD59OE5xw/HyrK
XOm13R1YuaLt8Z8oD84fEYHU0VHPyhWUcZM5nSSmekIdF/wunBSVcXMaoQJOo+jrqOV3jYCm3cam
Eu8hDxK2egyU47/3cjU9d9wEOsrPNEHny2OAnr18mbyNsugT7uNaQRMZqzZCzzCH28SX2AmBRzku
fy8aJMEjn/Lj+PzlG/MMUpHi44WwwxprYGXDIplyg9kGB9ULdfPVYGO0P6Ybeogmx/UU/BmxVBA5
hQRvpobAwUcbffuC1Z1GfSOu6ms3IV8s9Ef1cS3cBZ1AgO5rzBMziICNMEtysvFXBXyGAbMnlJc2
zuPQag34aa/WWx6qavk2xBdDiTzKVQvVqq3AR7UKk3v32DRs7lTSB13d8eQ8UvihC7Ie2LynCwTj
3u0LfS42SSSqBYnxiATnvRTUZP38cvuYjfyFPfocXsL+NlaICazOeJToENughvsUdLqnk3SfVyhM
1G603An5qG7ju9zypulDo90Gzb96/9opKqvboIx3B0rWnIOW5SwLFNuEk0JW56Nf9dyug8aSM9/y
+X1sP+MiJWSzT048hIdV9wZedqTGujU7qkx/tD/Qxe/mJHXANwCjZkVvfWJ4XD8hPafFpF/iZ6tG
RZjIuUPrYQrbbOHzjiGp6IH0fu7/Z9tnHK+xA7Djgmu1Mym2Hvi8rCxKLJXz4JDy1Y8m+PSGQhbB
wWx2ey6xfMY5ACf5DL5btpkJKd8ZuSim+cRk8NSM+U2s2VQppAy5Ble5/nT03IpdM/IfHVD9XHTp
Q9UhUuzXqFbx4x5ayBsmmI02wFuDsBmC2el0YxEm18jQrkiHs3V1JmG/kslSdCh9TiiwxhmRfNKb
2yjFdDxVndLblcarsAjIbc3n72FeVZCm6EaNmkOxn1pf4c0lP1x/bqHWVGnU62Yde/Gm2ZX4sHiS
HvBRbn516ZZT78Y1wegAUJie37P4x3V2ww6LfDfGyfYsFdixFaQyMhacVZO4voDyb89p6JtcIctc
zZ8SC3dvo9WGXh6r90vjveUbT3Ww3UQ+vkQNeuXqYCZaI2UIm11gPpOT+UOxWuQtdsrZnGnqH7ls
GPL4yI+YvJCwhECju7VIOQW0HlnPKbLiq0x9ZtnWX99Lnxt4qrEFKpXQF5CZIIB0Oq9kN91q9dLz
LpmTkKbrC5Or0+vR8CG+stQ+1xM81Xf4s2XIOxwuuH70veKquOhJLklQMdFr9Yl+yQpHMhQO1BfX
mFuuU0b+hNq+rGFTyc3QpCs1wL9TptUPpHjX8I644ozjpxVyBZo3H8NpeTUmzMB00XxwmMeH8EYC
umnGD4N9Wv5wYwJND8fQXDHJgV9lp9gk4GBoaYt6tJl+Ub94EV+o43E1PfKzaR8WH2TgMhquZd/p
e5UdrZ9xzm4vwr/TU82v5PhVqfcNKAYaFuTeX7ACQdt3XBLxObXBxn59T+Ytg5q84keOKK21Dzbo
kBBo7SMenOn84lVKQhA/N4M1ULgC8INLpbSjLWJk0EzH3ejfcoIeg0f9wsG19GGWAioZM4eE8Hp5
ABJ3wIix+MEpwb1HrjISaQI219+bPuLpeJhsb4hqbZs2W1ybX63SFi7BjUzknXIJdVX/4jvksS+l
nLhMlImpyReDuAeygnk0eCdc15giZ6sZY8zwygUkVEpAtE8K69g7DUJ94xCrY98FLKeWXbWjBwTp
Hxs0VB1wIoJ+WjkG25FYEP7eRSFyTuO7+ZUuOrPlzinCafp17S+3rStLfAq7lUEumzQqWwHcnEpx
taLBgw7ulqDdQUV4yr6fuT83Pp4RsKRzBzR2zlYmkMrAj1cUJgMnpZVI35f2o7ptGAIv1qDjorJI
Dg3RGNKzMA+bpuYlhxvFE1aPLL6J4Cc0JvRGp0eYhyCQrE8bnGOzbwstJm/sfWZ2244gihuOzLPa
emAQJoSdPAHybwVexudBx/oVGuma/MxKJM327lN43Ica9hrNHDXZrpW/liJ7TXF2CrR8bl/KiVEF
DHCyxbYAKMx9oxx83ZmeAcT1qXg1bcZ/GDpTBZ4zq8s4mKcVod6TaUrPPXxw1FdvIe0rxWSB5Vd2
+th8uHdL1KC5wHN+RuFWbKVJS0WXPZf2/VuTFq+F9rKPHiHstu6v+fuV832jSf9+d3QPNQ5g2bHT
MKNLqrI0PlsoUwIogOW9fz3TWqLghzxOpIRV5UmyI+3t65mVi67RU4MkYllLxf/BzdTpJj9Dx3H+
A7xsXutzMZitjdqswN4c0cYw4JaAa1B8r+NPR+lSHTYdE3rGZtUK0VU32UUSbbLA7bXbh6U9I5nl
r0V5qhWbK30ljWofyKUyxI1wdlfWIJguC88gFHJEmt5Wziqdi6VaKnt865zLuCSM1Tl9xaIscD8R
iKWdZUmKwJPOH9op3pv6MrRcEXYk6AnqtnEBXuGTt/NkHrqRi+mJ2XhZlVeNUAj6ySzA7jAoBmcl
7nYFNK8fQQZTL+x4DtIxZf1bcKi3GP7Sakmk7JYH1PCFITeJ499ohHEFEm2mr5F15CTLGp1NFEt8
5l1CsAXQSUYZ8YEk1lELMstrsnXv3GjB/iDjWbDCsTZGlCL2mBIdKNgPU15cyxGlf6TSPYMfydow
g8BDBddzYI+zel6M1w5ZF31OoG/B3TN94jlCQR+W0ZQdSLukRBlj5f/byLfz/uQEBlbz96mA/cdk
uSaptRezoIhreXpzdD73fiDrMKwy8sHSy+V02MeWwjfRaLsONvKLff2A6BymaThhfgkstTOHfGVl
fUnXOY5OQt19AU66L+cZCqk5wrqpIF8ZZkh0tXzA/823M6yNXbfqA04EdXATlbKszyQbegUoUCBm
NgC++aMzE4qqK8HYO5JuVYz4w9oxGFzkOvR6fKYPgxlhN4WTUMcJPaUPyDg5K79GjHPj9W0m/Kxc
AFHKOKTHs08TLhZbiqjiWrSWwLL21jpejMSUp4XX09esb7n2ux5KmWXGYVDpb1+XsUmeTyfKP9+r
HE5JKyrDoofH/MJPGQzD8L44bR5mZXvAyKfvtwEIJz0LUdpTq/nucUywEF3toVi0BGQEon137/q8
JkKTZu+rBlsZUp7kopI0weDNNy8lPXWFeN39a9XrA6prqa72ZdZjQAV2bwq11thylYXohnJQWjUc
J5joKFs1Sdlslv97QkRPpxq/KZR9nQOF11JFHWfQ8r171UZki87/pwdyK/SLir6BooQP1q7iyl+r
Z1vV/I1P5ZSRjxdalFVLQdk8OuXzyAJ+xLwprqJgxUppWBzh7k2X4Xcj+unpu+G9injh28i4n0NT
C/NFo0jX8SuaTcci0+AVNts/BFra8cvGXeoTw8d4mbcN3p0tUgqQzcNyjos+jGH+GOtSpnRQ7Eu1
akGSM5ay6kfP7a47yeGydT9ApJtVBVLlfG8ba1+M1uznl6aXLpeVc/EvskmLIu/SJ93Duej9fuZV
dUDCj1jnK9kuL2vUnRdXoU1SU7Yr/vDcwn5e1OPs/GtOleMiJRQbNQCwMA8W1JFTaOXdc9vBjUg3
1TgJmQ/p8eO1EpGrqZjELOMh3GRB0Lev8OdIeARIZixnL8e7x9IXkP6ijIGl7gMmKZC8yFbJHvkw
1+4/u+Pj7hCvkwC7wCcRT2EIdDPKBTRt1dZIn/cRRvlIUNXJtBBkuPYKdeFBsFDVlCMJmgG0kxV2
nzb4EwyZQMIGygUijW21sQ2CS7Wc3Cor7eh3xzvYadxnMHbSgk2z29tN6/HKm90YM++HBKaEoAqQ
2S2xlJgRWzcsSVstgtCTgqD90vqhbOTKVrJIfqtkrzqp4pZFiu+i0SOW0vzOB5rG5HaaWFokCCf9
YlT37j7aNH5b6u4IAM03HsBvVoePnqp11LdVnuzmgZ6hqgEK+esfdXh7ManefulCqgOk++071Bkz
+sMdl7lPvaro4GMDiK9llSKrXhjN6Vyi71zz7TcLL9Np+RDwhMbW57Kh3J1xyblZ6vIlCce6RAUU
fMAm61R/zqswe7OrsENPi2WKtgQlab2FaK6j2rAfvYB4NDdC8JFUTjaRpiKDHi/GwA02dc6NcnGV
vk6WsUTXugRFxpFNnyQEakEiUuRVLfx2gc9ylF/q+pOFKpJ5DOtUpISF3kBW1JjTtqz6ELCqdP6C
pWWWnoLs/UvyEnaAsDYTm9BKg4oLMVLR2NBsOAAByo7TxdrL5BieAWhULygJSjjdTM22HrSuS+4r
uss2ED3xVosVrlHwVNkZ+boUaVajDfa35FoF0Z4OtTpOmfjodAUTwqpK1BCB/MCD4w/rLGe/AYio
DLqGBxWrGk4bv3ZvZcz9Zhhz9v0oe37OZVMOWtg9ZUFFU1WlcBcFkwassU05uUwvr3hO9QFEjkMn
YBQW5VHdTXtQ+YZyFerNcR7UzSEiTwJe2yH50Xm1qc/A5lQbSTvumBtYTZyQaEWGvQoWJvEUXXQl
AN+fY5YOYQdHYBaSZDF0V4/EvH0WB7N4rkJz9skF2GygW2dZrkq0HYMBWJYqC5Z9YhbUI+cA9+Dx
MGh7dJk5AyesG2hx9fy57HHZh5bK7ZHijoWoW8aeF4tDnFtM/c+m77Dx5DWJts0qDcQzkfrriQGM
Lei7RMPMTkmqLAoE12nFZk5fVpHTy2o/3lf5giXNiPceMkLFnLIgsOMP+gQwrhH6Rsm3KSwG1z0t
iAJK5RPvy7slmTGOd2jvtY3v0IebAWasL9Un8FWQahJEX71WsuXJT1vllPkbjMWjVqHgU2+vPMXz
1OmJuqVD+TQZIIoWyDetVAGRp7xzODvOtFZBgt4W330tNFJ941IsgWugRKfyfNgFB+nG+3D1Shab
CoJkOCy1/XXEI/N5sv4zYcZkPP4xEM1T1yQAf8euPXwnovxgILfa/sStL6o2GM3n/sLgPdYO/2R0
TGvDM5JntGPTCbMahvJjbWblwtPjTyLKMfzAzWvsmQtaYuneWcxOjQnhrCkRp6+DpMyYQndCuNPt
FmG+J5B6/0NYlBwnQ/G6a8vrY1gHNUTPOPSftI5N5on0TCYMlL+KRzRlqJf97ExASlVgrXxakxpm
X+691Soklgm8bVSzlBQltp/+Hod/WQfH8Vhol5VbK8iySxL3hGXedF3dlZdjJ6LLssryw6HTg83v
aDwyMiSgAW7ps7k89/zt6BzTQ+sUDoXJRNyffxRIanhTDXM1I0vkC3YCkFZj4m95SQG891h3Rn6u
08Xv59W7oZUdBg/Rfm9cBtVZ03LShYswzXe7Jj8cpszBkiTi05RxlL/SPE0Rc8GCq7yOI62OaYQk
CWqV2IZ7fOLBgP5uFLGj0z7LaCbw3EQHxcprjz6Z3ptSP5WtvPPS2hz+C9HCSnBbgcKHC9k1kxt5
vS+AWn/AscvgBDIBa958VHbxpWVkm+qbK4MBkC+MV9pehCqR31NZre2oSyyW6sme4ud84uY50b6O
cvAReqJZZ1RQrFI4v+VB+Y6UY+cLYZDA+nwqZKI9Dh1LG31httHn1J6d0aik4BUhHP2V16+ULfBP
IJHcDJO7hqqpy4UIMoWXoc5Uo3r3c3Qi5xDvKimEvaFHTbIVVbyPK0IcuL/XszAZ5p+ZdqgdJkq5
KMwWttklxjZTR2x48Rp9j6HVIgyZwjDyP+/pkcOW4skhSkJab2oe0YUN9lCYqcu6jtpGpgb+Zi9a
pCtGl6RvGXJ+yM0FZCWDrR/zuoF9am/usn6YOd9f6ai5ci4kosEh6/fSWxqpdZIB0pbrqAT9rWVy
9b7gW5te48VKP93BLRlvWYx/k4GVwi8JYWKBJ3a3Wl54nGSBYrPM+aitl9Oe3PT1GwjIiPgjBmeH
tQcDSKVgrjmRFyPtOsxEozWBrmcOcMpWgOUJMNSN2msU2aIY/vqjuhbiNpojaQSJyZRMlKrbIZbz
MdurI9GKJHvTA7IlFao7M7bIca8cASsGE88hi8GTiLZMe84kWEmbHkag6evBn/aSEWFTH86TPgF8
gNR10zawcI5yibSf5MI4PvGGBbDrfYaCHP0bVCqhZ60ZhhgEKxjZl/EbfNBiKQV1S5Tmdu1M/LFj
l2GxhKYRlG9oVFcY8g5t6HlbkrVO5xl56SgQxZvOnCb49cqr3vHIe70gQoExJ9Duy0XeDuAIRRax
ODXRny9FSnlidw5MdaGs3iu+GAlkn7ztvKUOtHFtG85H9oydipexIAIzx68TSN8O3oRf0qKgQYJC
iQoYEDvBwANbPP1nVdXkUDY3YgiYAG/gWp5dphk+MutXNk1lKRaQJL3L5BiubgfWRZDBHmJVakwk
HYhCquti2ZXhi9DTHB2IIy95eIVqUei/RUljRnEM2O2LDw8NTo6Xis1qAmPhpfM0X3nngHnzg5tn
2POL+yVBPdMyiz4ZCImGtc54RV61NNdpnei5Gv20e6JYsaNu4ybBc328OF2ruKQTRKVdM2SlBFfY
SN2KmzViDhrYXrPI4Q27IMKpDCHGUwSyw9UMxBSYGJRaobMy/MP8J/bcWePfGNi7Syw1F7S6aZbj
gtxy/s79TCEKVxm+0aT0lVUztbn+HRmLASK00aKsnW95zNBGpwygzKlodTvPo9+MR1d0QbOLiE1G
FJNM03ZtW5fFHyQ053O9+YakelHVhla64zTQebNHkGGd9BQDovya9lYSktuEClRm+p5MrpN/SK2s
6e6AB5gk6/XyhmBBto4FnNkj2Es9IWNtvy/0vfN+qWgkNjXbekx7qdj+B+7eriL2t41LfJl6vTwA
LPiXhbqf9C1cfYlexUL4Rjt5lqNbwpsF+vpHQy9Zi9dWNePsegFvyamfn6c6bL29iCBIpu4NsR0a
Vs1vJ0oo27BbKlnJ+50d3roUdMDXMej41K8vNdeWeMDvlI5QtsNGI31uHI7BeTLqQYX1V4PVbZJ+
0hVPIUBBzuN5ytospHi1TPFPd4QYELr1c5Z8lJBQZxcZExkbdowO38/5cy+AFUH01oSAcydTCM+p
gLSZwUXJsIPjhJj7ToGD3Oq6hBdlxnioebM65w4q8Y8eaOd4jssTWIJIDcdNpT2qOum+0xlogYsK
dCf01D2mF9eN5s7FKFsUirJ3TOcAQUVjDZHMz4HOBDhpimSXmsqYUBI/zg6Cy5JxBjfCTQZJHack
kxawfK9tmk3kun2p5GC85ueKNav1AHHCTAYFqOPkb7YrMqp52ZQyIwKNQ/gN4eGS0YsYMJDbPPTN
eihDi2fYtUwsdf7WyQpvOi8F2yJ3Wyb9AfyzNuqsg/soWV3nhWs0xQVtBx5rqp8WlBuVZr3TVbKt
xRw9uibKhjHESdbqahpgYksNfrbvg77XaoIJJjo/Onyr4v9VHzp7BAmDYqNppi8RLZuc7WeZVe+V
0Yz5gbQpLc+IMVDKVYCdOZT4bk5CCkCiB/mCodw/Fe/GVb7TwhfSEtHbh4jqqlp6Z5hZDjV914js
EzVLK32p9+PTwbdkyP7e9E1LxSNNRmyJvMDEjc/JflIfynYNMP011FoY8h4MxtGNeTpSJmAAAQG0
y0/4wsDSCSrsA4HiCNaeE7dka2d8iPU+gAt5y1zo/AR4aL0v3e50yeCXjwGoY7DhIDk90oSFtoaS
SVSSkVo+YkKU7waKZxvgcR51j4UPbZspa4OF8rjuAA/g2xay1WACJwrZnvIBMqcG8aaIHvvogk/U
IGbw6o2X4RPLp1IvTFda2UZLYvLvzavPNG6X1yVPUtyvvxwS1j8a7v3562qzckdll2JUHGgTYdhX
Pa7e8UiZhYRyFnPUlSOn4uyXy4HsbU5tKT73wRjL+pcUWj02ddFQqYjk7sCU80Zx0ksY8SjVYv/W
vCUeh2MLvFrZxicJ/u9uDafYa12gBCJgd3CtLmYDem1dr8rQyfmHppI8CabGtMDYUEQiRjahzhX7
pi2kzn9zEsbqL1DdHgyKGw7Rycfb/I9mhnGHvtO7JSNM/ImJROHXABPkhSfgqfhFkG0k3aWojvzJ
tA32FW64o7zihoFYiQzfBydM7BXH5DgtuS96xnc5TjP9Nu5lCj6WYv/yGyA65aL4BENpbstwpuj0
LZwNT69qtdv5KcQSNIVYgcNjBLeYqmuwY+5AqjArD8Z+5+fkCtR6nkKvZxivO83FxR4+5Rjlg4Yi
lSG6SfoVepmmwtL68jfcFVbuQg3IzWHM+kyCHygVwteGue4IY5B+ah0dwIm86iW2ijt53qg32br9
iJoX0/3XW39nzd8hjNyHjbJbRi4/c3V6luJ6yr0HYPLwCKh90vvHEePlo0bkofQUNp3L92uiTOSB
To5BsvayYFEv9c7W4dnyhXpa6sIzTLWZwA+lUaBqquBQKOci/nt7LKfrZ728hyXsbmJRUkfyI1tb
aQUAZpI/l6NVVJGXWf8J5XWzPLWIiAfNGfwKZrl6fh0W3USNG+1HRlOnBy4qBPoR4gnIBZYjUoG1
/U1Zdd/xyE/PC3I7vWS1wdMP34dt4gLSXcFqiTrsScc09WqDB57eECnU1GQpofVU+zgxF3BEZIlY
/8d37Y8x3+BS+Sr8piw9jQyZWOafraC4cOqheLErXjzwrREVXUMaYc5j5Azjx+D7zS5nb6+qS7wH
4dxbaIg9gx/N/rcLJ5z4qGM3bLeKgW2nCDEEI3P3NoCc7tKjy+LWjaA9f9J1uruuk3ur4Gqs9NVC
3Vm1bQj4qkaCxZKc5i0ZZ5XPjdE5YEmjggUjgev3mbsngil9aIAMWlzsgoPDPW2scuzN3HlvETH0
XAPUnyDmcZS9ev3gr3yO7DO2qHKtfUIHdItLDrZFowcEw4mxD1nMCJSdtVvPiy/gTWzS+PIcQKfe
j1UnqtxwxjT1tU235xXzUrJ/Y0/CeX2xqntEzpAiXns7YnvaXSQH3hlODDn8QTmd7I3giZ/yrm3K
tiUQqnO19QrtMAk5gMc9I+f48FdjdWd9NESZs6/itR1ACmxhI00U0v7sBx76mh6z+VKYayX92ZO9
3j4HnStKKpnu2CXx2IJEMmm186UH/K1LsCLTKM99obMiEAdbFPP2jDRZrU7+1FFZSRDXmoiiUwOQ
npatrYOrl6mGF2sFVUAX7b/L1Nw9BuGR4EW8+9Q+b9qCc+ymDafACvlclEDnETQag8rS8XZTd6Yt
CdMQm0jwySMjIg1qVG/KatD68DUOFA6OH9fhCYTTJ9yjBVIXdRz6WMxNoYJNFMJ6Y1RGIMQS8CS6
E2vtzp4CkI92ClosehzsN2IdTOjpqBGV0uSprhmQXcZwZd6S10487pOG409Z9knSGRaRyFtuVVBl
/dqs+7EdGZ2k/+sOT6Emb/jkd3eV5n7PdLD5If5gmN75JodMTXrTJayLrj6aqupuktMvyFdl8B3d
IYNmGRtW/FSxcvi0yx5H6JRBxoNvD7SUkm2ck2Osn3k/ZDcnqpdXn/np43bgAnFX1CkZNP0PX5Ob
WYDERRdLWwPYjKTW4ywUinlyQqyStfXv+PBf5dVRHzgTnOp6DOJNoGK+4ZWWy2meK9dBMT7xAhJK
Xgh0YMG1ST3QymAQh+Nucm5sQj3YFO4pZV9lpUe7CDR+oTTVbYhSdwCMlc2VjsiWkKDAX5O46aYg
wSZWiX5pSIX6Fcn90SmkqQedE5+9VUNEfWUjuHIhUGPfLjCBZj45xv958pmurpxqXAyQ0kKKNNBq
gb23Xq3uXpfHaoOe/hWn1A+bg7dVffG3nqk0G5zzs51/G/nVpJDxNeEdxjTqeKjNTq3GdahY6pcd
t1ajNk3k5b+mldXCi22NC7PHHLB1uhEybIEh5B5eNgeFqofDflYTN/auoaEyfkhnegGBni8RPOlr
WDssSuuetzK4/JBl0sr0kPZVOgnPFMuMPGp3a1KP8vnHhYB9l2SuAeOFLxZK0u2MyA2eOVGAxRXD
J10jLj/W2p/GMgvVzLfLFNEIqlXe6YjMf+FM55wlZY6i7SmumiZAKbM7PxvA/fSf3DGgWFOI0RPh
jFFEddPdBUtezi4SH2Z7hLpVK3+FsPEASdYW5ZP4meRCfAUJejgMD5wonxyWWHBXV2SmrsSG8QcT
mZIZjrwv8BFr6Byt4sEEjPULCBJw5LdyFTGwYwt30eeA2WqadJZ6PVULLRpSPkU/1n893WSs9U2j
kctnG8mDWDbPoGVtQnardWGEeHRTG8BYjNtzyUzp/0PVflYAyntn9uN3gFbyM3MvAYUjcMT2Tr5I
JPUuIb3n87Jz69Zn3NvK54Jon2l2oGFKbxJbNuKJhnhLWYJmjGTDIv1wLGIp52bFOVNUeR4LoTOZ
IBwsxCNBjjPvsaovGumHg1W7tjz07TlwQGBx2WVO6OykjXTXXzmVs4l5S/vYjOrWOYnB4kPEl8in
ytP30NZP7EkZWipjVn7BGQr9gKlk/yxK/UgToVOUm1tGhPhL0S7tD2wBYnQGwRmauqDFd8G9tdk7
PyK1fHtGeODgkbzwK0LX/+GKNZrhwrSD/fT+6woOxkFcu2oE8bFyojeKhIjvsdsj+HE7kwPzCxUb
6/7vO1epeTZcChRdmdg9qIEu/PKLtgWvxAK2LVmNtR8sjyHJ7RZFmWd1QYEmlom20O4b+zxBjYoH
Lvo+Fjiht4iZ/SDefj5lPs/gdTi1cECfyLtneGi5m1cvmPCarmHb4pN6zCSfflUMEMUXN+SZgD5w
xOlXbZwqYbBGvJJXaWccV8bUCjQ4MaCod529ZUoH3xLXgM+s4/J0nBv26iiv0JeRy/DYWVlkDr7/
r4Fp0gNg6ddraf3agVLPQ3delT4XjE6ZLUU8j0NOwRxQkdqP11/ZbA6OOf1ODnSicQDsS3kCE+0x
rrU/8MIyttpHddzv2yuOK0nUwmSLui6EmMJGZ0I2EhryEJNo5jzRdJaLzISQVBexpFvPGPHvjN46
eg8FW0IddJFrTXgI8rfquD8o9yTsZ0lYyYqn2EVW7H1FUYpS91WoGQDoKocdUX5lg2vxyiqHhuFz
1rB1/O/h95g2UCyE0GJPgeQ7tJotWjXtBLnGji89+UQy+PV5oav+wm52I2V1LctRFOKDKQxi4rAr
DKmSpFX8zDe5mbsDTXJ1n3x0WtF0F7Kpjz+1Uw44omX4cvNgVbUTSjPyl1NNRd9oJ9kGw5y+/ix8
+NCzgvNnbD2nNZ0kJGGeWoSdgVEY6xIA8Aep1pdJ9zzxSTmgcqhSLyrq44MMiJ8Bm5kYY9AR0J6c
VL/jP+zhNQScp33xnJAc2IjUmZLjsxFo48ObAaBZHuquv9LhJ9IV1/BweW53vPx8jILW3OGou0AE
9vLPGcQhWCll5rjkbN9WXtBRqNV4uJYajsXD2hCIOZbMQ1iMKA2ebNrmeXKIjTiebXtkE4sBgziB
sG+dsPISZ/kQS0m9kS2kV7V2ZKii8ZTDVqecz2CzWJvVovoXoKsUFgrswTJcZ4GCIzN1D2y7xB7L
ngC9kR8E6duUo2Vh7vl8oTdjfnfwp6RrX5+euPctgmJKze/AIdQItJbFcWtV1Q97rp9wPFsIweX1
OP+1IlWlHcLEx71xJWC2FamAQDDWHnF6WS4qURmFdxZLTGa7bb2bUdQv7+gxkBWg3hc1QwhC/2Oy
qyjuCPGmPdq+MZSJFbc0p97cjzDVgCOmfeLQJ6E1BvwnxyBg/JyTC7iK3caNdfBE5LxmSn2rD57Z
6rgxxSuoqVlR7UxWXkZW14VBf4MLGkcObyQ/fARY2TpraVLZLDxmW9A+bWePCqyBFvOnnjjUrUSZ
hShPDROQnNr9me9dp83GOCBuy9mZnNjCYmfjI7Q2qcD2JUTEvdXEvHXcNlYvglbP7nbkKgHGpJPS
7vI9uDEDN5WgiFfTUZ6i5OHcRj3/Z9Gk3S8vj0VtjXsWDVVizdYZQfe1DyLhzpBXL94Jx7sH9oVM
wpGpoitw+x269Hf3MAS+sNxgJot4azYVo3SVVK2gRsHXvNE6r9FVULXCCIR54NUIAakbBifqgccE
yvvbcLWZpQGe+z01a4HLzftjviv/TVgvxN8EIh7erEvGg5YbvMG6CEfziN+mQFxzqx0NjlbFC+SD
3zgYsvFlXu3V/QqoDY0G1VjIMnmPSk0E0Ix/gmCgPsEZHEB1AZxzVog6LbNFS2pCYqSnrhDdvotR
LDqyGx7lgdxc7JXYrDnFdWdLJGzgGWNw6tAHSO4GVrEaxWyrQP1+BcxCbam1gyba8zmfno4Ogmf4
7XPrHYn4U+UsfmtNWnUjk8B2O1y/dEecDKx7PIEWUWNNbRTYH98hp46fxU7k1R82L9nLNgE4cPKJ
YWu8kFvEvWEFmFv53Yx/NBom3eplN+K2nJO7aeQtcBjOGmRSbZo9aFJFYeRN2gKry7wkEr4ALcyw
Rm26c6t1iUAOvcFNtDEP5/+h3ICMX38OM0l2G9tfyVaMwyCc4AFFzjta+K4cJmNISzGZAKGJHQ6n
0wOcW38OkhZpDIgU/8RC4uvRX8IU8vr7kJrZyJe15BzjvWcFuG5i3WFGrBuYP39ew7CLmb9dVsak
wfnLUCvWR9kAwzI/w+6awZA89Y+ZL5N6cQ05+OI3XcZ6N+NgDWAe4fL2tuXiWbKCEJ+LNxK0dwyT
0BGreIxMBUezL7r/p6/hYV1S1HMJkDIJNNJbvgepC/BEFV693Yngl6f4EEqdja9dK0cwRKyxlwjk
nkKtMWOEpV7D+jps4s7aupm3KkBKLRfsjc1RsG0Zy243RbPY5xmYwVBZcNW5ulX54vguSyZzxGCE
OyhYvA7sBQzYPnoTF26Jyxic5MZd0s5R9D6vxBMEvaWonQ2XHWwBUQOA8Gr6c4urO3M/NB863+n+
NdquRcUFjG3UOP1r6XnYhe1sUDF/+W+vzwncncINWYmrgsx2/kQaBGDxY8Alku2HYVcwrxi06+fz
HwOdLoD+lbTFGYM6y8FxE14vBDRcQc1a67UW4/IPtGBY2uHsInZ1NEnGCeJObz+pPgkvIzKovgrw
rcYpdcDjcDpeuzGKA6HjZ4s6jSO5FIssnBbywPB05KT5Y4KTQBrAOosF/+qg9WX0zePsct1nLQQ0
UP1fng8Ilgs8dMfMTxmG67cg5RPi6bgzcIDH+cCCZHMdBPMCsHZd6I/PK3sGHzISFm0tiKlGDSfn
09lm/lEKis7ML82V3eJ7EWdnBMXG2aaPz1Tk7QItVPVDVCsZdDB6N5E/vPeTy5Ik9rsDlmFgrMws
UUCnbJ1X9eAkD61R6dnm8K4bGEP5PomXIO0ZHiUyvtVmFWXznYF3V/peZZ7fqPnmNypa6vYBX2g+
fPs/iD8pBEYCBg6NcUrlk613nTpsuTKZPVnElgNNQ1MKbGRcIKuBuxmcMpuYMRW7dVl+CxOG4MNT
Cj7By/qQzcXyoDzY7IUOOFOq5jUGkrjMvyPRsw6ldEqYQPnPCLZXLe4t8tPuoqkfDj+f6jfrwsvJ
9tughfZsnLGvL8xHG8qrW2yaZSF7pNY6LzqRQ3wtfNda8u1d3YHncvliAXVENj/QvBxcjM24SxzO
7UOF9ZhXfVDCeV8CoQLfC+y9OfGgCgO7wPNlNln5kkdL3O47Hv2QnjxZsz6Fs7W8WXkRbK76lcMR
cHKxvgWH3O28SV7MbMtziEyPOwb9JCN5W4dYTGonwOZH+F7gPR59yUvWvgz1CjpT6SemEto2JXSR
MpjRF5ysX5nywOyaVuGcdOrfWuwoyHlCcoz24Rr1wCCG8fhc48trrAE+kN/OU8n5cx32oG0z6+9/
xEF/VSFH2WoQiZlmjNTpEejnZ0vd0+G9WXXctlL7lMl+Rl+p54/b21eDqSmaZOgNB1lSLU5CvHoo
1j7sEBJIUxXScQGvTxRfqMnugif7xWvvEkHMqt4gooGHAU+/SjeCGkDV4STbnBOy6Kwu9pDw76FX
r1f9PgdmBukIqj/JktvJKQVIveZElkzDh2j56LBaqqmkDyYQkONw/lAwgmrOmrZXfGNlNqfe5Z91
s1TB0Y69W5vrC6QmGWhsOBd6Oh4h3mItr5XArXALTE5NRlBQm95kWG2XsXMnHtLAvV1HVn+Aokuo
QrvtLK3LazrjpfobxnLVx+K+Z/kLWNtCGKCiFJVZNc1SLaFNhnI/lZXcLn19AXDoiQtGXr/342ZL
Z5zjWmP2ch0CTopVEYKsguYf9pwEbDqG0EowKq6YCBW9aB+eyFKHKk0R8S96wMASVgE9+5MnhZd8
eQjF8GFo6rtq6fC2eti8HHAizdzc41+89WxV/QRsSIx8HS4sfqrsMc9SscT+cmTe75i4MFLtfjc2
VGq4Y3JSnkVVHr/Yppg1i5rrXKY0PHRQFg89DRECJJRTrEhlGEa9C+IdABm6yXhd9SwqRJ3BSP4s
ermVRJwIC0I/A4pZvIHW5otkwUrwgzPlGYUaE0wIwpqsEhgDy9pDnK4Yu//ACuPPp25SR4QtuPel
HQtKaAN5w3t1ahyYAKTgNvEGHyCgY+3TXpA2dgQLOMTfBfqJekNklszc66OWuxfyRI1sl7Dl0H8q
UKSq5jvoxXJhL1W4epElWazQJss7m1K+ToZvV42iuXlEXbl5vriHpE6bPR1QUNMF+qJg+gnSMJtW
IXkfVEqdV4Ptq1YPIkjwb8GoBYIiU2YPMzOe7/0fNkUHaxf8ij9oFc68xUoi6OO4/t50gvFlF3yc
oI9OMhVzhHMgjWn1f6VbntI5HAV3bPZ4yOcyU5sY5XqN/j3V5Emra+sLVcQJ04c2AEasZlaZRWOq
OKKd3rraQKMCPQRIzyl9v3NPrDlgPsbeNV5rLLQqb6vNwf1VC67djrC/Ozp1rKNoDs6sGo49Kfdl
DuCO20geR24sYUo/shyWJXSOV2R7wnNmY46MRT+i82kY6qxS/roOsW+Fq7UJyv5jDHWpfnOtEpAc
KcqWHgHtEh8ZYcLe/4pDpAU1zR5bQ6bflHZHLQp8RDNykR28MMZjfs0dJAQ/GAPomPtkorbBOqJu
4rrxgLx208UoTnTwrGpQuPySVUpCgMQ6+35kTMEHY70A5uOOKSk3i/c9W0QVx0qhie85M8NEDskE
Dhz5r+Lu4SMIC47opWHXnt4ltC0m1WJRYhh0NrIaOWjQNKacc02PW0j9lh6+fwUxisCGjG5Rr8OB
glK8XdGJNRUbuf21cYwtPVqKrR7GNUdxoViTZtc5zbsQn52AwVG5uXJRlZfyHQiwciBfrmoVQtiE
qsX0muF7S/uJlIQWnOIE/9f4+gutZPWqtRdiGK97jgSEGZIXgSsPDj6/F65byXA6zD1dbLqbXn5E
te5cHXg31j81flCngc9Zkh4DL4r8FBXq1m4/MlSXvpFd6XaAC4MEWDG/7Ac67x0cNzzA4nlmXmPJ
RyV0JdsYx+DUTjw53yIjRr1kb0ZDIDJuFU2qURAlWW8a/KM0S+eFas90BQLtEmi7mICzz2Ov6N3P
aR8DEptedjzf2U4/PEPgprdF9mnZX39YvX0kJ3QLby2AMTwvFA5TrGHk/C9MET01FTlp1iVz51Ki
ieO8Pxp2rMV17u/bCoYYKbGtopZFcMbIW1As1Lmu00uCUQGFxDYyllSoLMUR2ZZk55vXLIm+vUKa
RTUrwUT14Vi/AEE5bgLtzCvr6CbudDmp9KM/OCWzPqmosW3SoOIZXiU1q4OqIz3DAszCJvz4qt/T
sTiC5h/1Vf3ymx3ti+y2F8W5wnNYUycGXjaxp9cSjEX16dOBb6gQ3LIXMCCoRmFx/T+5chTQu3o8
QVFQEoMde/HUynQfAH7ZO5Z5gxm2M6DzZ2IZr9VIWU4cPWoh9pvt9PkN/dGPC6Bue6rvNy1t0pzN
T3r3ucYIv+VO+MYy25FeoVOEsgOTv82aOCM9HN5CHDYMpajOKRTlsmN6N/M02bDmK8Wc2F0YSCk6
u/mhw1SHiWO4AWADwRgkDygGTVR3y2rdP5uabbhmOWomJuEMicAwZS9uSWv+tjVSSzlKEl2JMCR1
ivpywHEAXPqHTGwEkYNhXQJKZMPxg9pWqT/vY5BupWI3oymTBO77/gJ0ow99TWZ7dUfsQSm9ZEtK
Ufj3voRifw7D3QPEg1DcWTFi+PhljNcxl34IX0S9wnzcj0FfIFwTZkSAIQpHFgA1xAYuZKex67ue
e3BiRMTsZ54QFSSA/mv+tb48Ppe75sMXZ6XOVvqzF9qETKlE0MREyufypLUh7j5fngBvf16cwQfk
eGFkuPfNHdig/YO/1F/WQIWNVtG51XaW59lHN1uypEfhuj/7iVOPiSB+8t7EvzaHzDoJxsWbxbY+
sAHr1KTOQBiPoX3kntRmUgc7KKLRuzZZoNONOXjxIrCILYOv+/nsf6HXhsoMJ0/HMjL1kMXO/4Zn
SOMa/Ur4qnQQrXOZPcFYJF9MweHeEw9M4MvWGU5DsZbNPoMYVbhHUCA6Z/WiS02H2NhU6ccECrGn
sO2PoYkdJWLCCwC7PCV9mfhf03rVyoh0QZ18lgG7IYZrSTQCp6mkJ5z7+rfPdAg6BIiHA34cKHlx
+G8bliligRhxQexAr5RH7BDFDSXD4h4VQhWIM4yiwChz5UHhYRBkTOIONuCTAj1qqkl3iu54DIoT
30BgrSRAWdjp/GSLW0d4CDlsUeVbr+8sjvJZ3rU/iOjpAD4AQ7eN2ni+OY5sdrS61XwO3g8a/8Ge
at1hGoDWYYCKNMQsB5nTDzZyyr51kWUGRDhRbXYntVHvYg8dj/ixNBtuFv80KoHz/WCuCrLWxgrz
B5cBCnrkF8pkMSiwrwKUbjo9qcyjpqA4q6GaG40MrMap/qC15o2D6IXRWG9U9Wo3xnGGfiW4E1wE
N4AbOT72YC4yIBm1u8XTTstSroRWKufR7p2eZimyw6tDnWzPGYjDmi6wCxwJbRLrUAXN5GnR8bdw
ec68rOpr2bx+C2kxP0GV6MUm9IM5ahrB05838acm1qvZlxpgKGSAdwylCsCr+Cqw+1KBzqjjEzXy
Vr9XU6NpNO0lv5MJqTLw57pLhjiuALLEtNNhDaSPWwSo4/1fp4iVDh72t/8IZFqR4zgLVUW36rq+
WzyN0U4fEWlhWim4Idupw/Q7NaoWY4g9hspwEbNm5P2kXGzjEyL30cNVk8++rex9auy8MEVOdwVl
yzeT+46u1EB48dpq5w33WxsqqxzF1OhWuJGzjvJbWh9QAsUrC/MCU28dfGnDUJt7oeEzNJX9ZPSS
cdbwBIzhQdBC2buesPh25ijQH170VGhALM8gXPrjFSilOPuAnQwzJoK7tPAgR0zl7gW4/BfOchNA
vzfPwx1DqfLFNQJ8QQaUzrsn7D9U3b10NjDd3exnQnsbobK8v+MdLmK8dkoXxHN3TjyERmoDB11Y
iNu0bz9KQhwp1kNzEfqBD89arDaHKF6ZrYXv8BOHwPVa8RvkORLP4wSoFnjF6m31ZN6K/h4yYG7N
kjZLe1e4NSvT+gbqA2f06CsvKy3oDfGQQHRucmbR6ZeQ+z/Oq+Q3w9xmdFzTMcKlcPNFYp9ZH0pO
sB0pcvs6fsaZvnseYzfYmv4lGAs/53iGyzveItvwuEzfvb6mpviTbxE7yNmLIZ7obJ+dNEJKEUiL
6VT30xUuwQrKl59kMTjKEnBt7HwCV/Qt0IxSXbx8nMtklG+M6klCzHP+ZgFJ3MA2ltzKNwStIwkb
4ww61he6MaxCnaGj9Gb2FkgiDChuUixKBi0cE5cdafgFCYSFiiqELx7O6isjfnY+lyC9xoLMjeJh
gh0ih/Lr9MsamGTZXhrFZP/MO7bfLYRaUStxqWLi8EQcki0P8rGiwzx8uRJGmkszFmGb0zCQqGwX
WwGQ61/YB2Te9bl9JjqVbkZxSgHMved8sorS36+21eKSWigxeYJZc+aWB1mJIDjb6dRSovbHyass
Wbr+ooal7nCuVrN1TRqbq70QVeMCkgs4/IX20BdxVo68w8Xb25uezxPTwRdLm95pXuMbL9/bMPzt
KA4NcsVp+M+/qSbwwOEwiIrIDg8wTb6jvBcI+LDHrkOcs8hRii63qC+e/vaPKcYW4n/3rCx6gjvR
Z/A/EQJJYZQ6Bv93BB5lMgk7RWNC/WvUEbszbTZfKhn+0761+LRq96NIwMVMWauYtA9x8H/VbeRm
VLT8mWYFPKkutu19jJaoeXuHsAVwhW0+G+5I9z0le03QzQVReA4KhHSffR7ge1Be1T+TsBS02qsM
LIQlhXBbt7VbIV1rEcpiozSCD9pUmVzVYzTBRMgZ3fXng+m6W7PXhqX4rDNuJD8i/E8+z79Hpxvm
wt4Y2cw1XhDPhUTzEe1PBwH95usSxknOA7yUlcfZv4vvMp4m2pqisBKXKoFFvE4yoq1kagLWyelT
OxG+Y7sSAdI4I6vDggTXZMeGLLtHh9zmER5Q1PbnJoV2bnrkY1EotQNEpVxa9OEkH+qOHsNEpCqb
iofrUAPcZ3C83c73HvanJuv8zv1IeojEW3YinmZKgpanuJfPjpleVPcS+SbXgqvTRhU/Z+RTI6p4
mhEoDcFAP4R/NmWNd619+hO3eqQRHfBufWzo/BoviCrlePd+fokTkkTqfcV9rWs5oM9fFOwlxaIA
HjgX5FZnE/gfgMaQ1try3+Nsb1ZRvbql7p9rM0u1QRvo50b+WEJ+UWI/Wmn62poGMrbYBX2Saj+3
NRojL6Mr0r3XgIERSgtTaw9FgHdLXj/jJaEXC0AeMSJa1zwnv5yihykJevAg2GUH4ckCbU0PwrvF
vqiuqKduBaqjbtCvGQZaEtP74QYwId2GPAY5tIUvsRCr7Ut/kAlQIKMJ8yfhzN5RKyBD4tudEqd6
6R722Pz+sgjLu58a5vYQrip89g6nC66w1XMdKJVtEfZz4CeC7Xv6iCEjmtmFODaZ/377qmd2CdBI
z/QGkNOvJZI/nYAbWTRfQxEg6TgeRW1DAOOYRNeH4ZGj1AmhuN/4S7weHiyjPTxShvvM2AJ8/OAE
44JTxb3dniV6aAl3NIl4YYvoW9Jr7/6/rGK+nIBmeK5xzzK3K7QB3Jx4tBdnw8nQlIJAQ30sdaeG
dI8KBaLmiO85Ksx+JRlVMDjLf98wg0H73FY9WaPoQKRTfhe2DSi+1VDs/9FhZKOuRDn5mnYrepY5
aJtXZqEcpD1ZnDetvKrG4Rkx2kP5sgR7CEVfj02/WaTuJbKxeT7yNXX4jFq26mG7PDJkDqecod/R
abHLoZIgZjhkvOhjFdy0wzcsKyaPPMjLKhO2hXVSMQSu2PS7I4HbOfFdmvqDgbH8ZR2gCv4MpjlP
xDPWY7gIZCNVhrS2i0SAGoG9+cTMuEpDrOtp5Rv34Gu4ZxNk1iHKeZF/HRz346BymTciBn2Io7/t
kSLACGgD5+D2DNTTPwtz83bUpn9WmL8zBWsYlg4vim7feoCfl6kKx8vxPTgFRYhgWCN/qFLmtCyC
agG+yUBiEwXfr3BLvHZsC8QhnNLr+BSWjvRi88idEea9g/GWM1iOJfWngwP0SPH62ofF+TBGGuUm
qf8YN7mX4309b3Dg961Muf5x9frZ/sYB0pv2oahHy7SXFBo90EADykPCEljs724FEq1AGrytTlEK
IqB3PkJudp9ZMeVS/D80YscL/PK0vHrW6LF8edtKbbFpvvNFFaOj1X/8kViKnzTTUTJoI0G5uwGx
Dd8NsIgFJygUu9G1cXHR+dNipDaUqo5OVXF8tmNxPURuKfNwYfGv4rxHZA64EZy5uW3UK4m+WU0N
rUQRM6/lFRhMm4Rflny1faGZmMmCN2o/wgW/fJ7/UBscvetSto4vPt7BkgI929nv6aFlaxH43/4M
iiX0serN+2J91fQNPvIlR/LbQ+RoEkadBlOjIGi/LCLJjGvPTCD8jRO8ER9Ge6xPjpM0H1Cgfu8Y
1a+uWUWj9eZ5BReNzCzfmttwGICFPbD7jcM/5ZhG+F6eQ8yUrZBS8IZS7Mwmtr72VjAGiNN2rtsb
XinfOlZtg3NCnSKUygByUB+sZcySapRy4eE5Jy0Ble7STrMjI8aTT8KyHVOcrzEB7UHWzL4fu5EX
p+yt97unjyt1oVH9NopV3paL+wLdK7B4Kg2EDWrDoMrdK0tKhK9DiWTAzHcfK/O0F+jHrej924LW
5xCkCgAoOBa3Dm7fMJ7ukXNm8jcDDCTruN5UEX47meL8eBUFj7y2z4fUasMlmRcx8L/D5X8oCBUF
ybNLL5BUw8GqxoZxfQYvJK/wpMF9WX/aLOb6ILeGd4/1caWmbhJEhAnpBZfMN5sJ4SysrbFazWek
IkkNG+0sWE+knRAtb3XkfO68juIuAP5PkuzIqN2a4WqCJgYC++tVvp1wkV1UnprPZxRBuu2Rfb1Y
4bjs974nWYEduWTrZavplEeHaNUbE8ccCLe0P6uud7+p/9lhNDRtDcV17ekvg81pZvSZI2qMRioh
z5yJcyjImnCowIroXCqn449gp2huYD/7fXntUrxrhMqOXKMEEWvGIFjKAyER+DqKv7M8WvtiKopz
BdcYbior0wxPLkEKLB2dl8w15axa47xxx/zj1kZC5Gwkplh71ua7ctmIezu05TuxTMiPGX2kJcub
achMcGDvglYZ7sf8WynTQNBhMRGpPDl1GTMprjsf0kqOTSGO7VgKMSJERHSrPKrovXVY1GtA+ixJ
5aEUKjI6q8QB/TKcJ8NvFBR5DtsMo226IFkDZAP6KagU0u41gkKL4F+j53SxCrlxtBlYzQygHwfj
Kj5hr+7Hhjp3TEaYUwzLjVnTiJJs0X44TaOy8l8nypHw39ZAaNOV3iud/o5EKCmikwY0WrUX4ZUA
W7ToN8CwC3oMSsNCwXtFOdvDboA1HT1ONgeCCsyokKnam02wKygACrIeaoI1s9loyjqNYEh0QUOk
T/XsXc6ftQysSxJvGr6lP/WztjJbnJiqMfCxeBieHpM29II9pzgojl8wAxvD8LJsC0PO2qQmL78Z
ig4Nd2dWnuFXcF3trzk/EyNsJSIsnkDVbsvTTRzA/0/Dz7UYt3M938au3p68gkeR4Bsp11aTznxl
ks5xawFgxoP+BCpkVzSd0poIy5Feg71DZ5L4sZz4AlNFV3qKQuSLDfl7zglSgphCiDyFQAXr55bP
WAnonsdJV1DAYrfAwUideUDKWaJ7Z49x6vrFX5cN+aHTYFV+SjmbQl6H0KT+j2798vDWH16PqCL6
ZHiEhkKj21WdUBp4cEC6ApKGcrfYXcEf3zcvNP39+NNNkvkKG9Bs3F1C5l8biRDfBiA0EnsqrYEG
rG+1hDddtcuvjy/jilIuEGXbFtICB38fbmd2blrTHTrDrdKC/yJHdoxSCTwBuwXXJzjsN890aGfT
v8roqsChfGod042Y+QdEO1drVn1/zMlLzNTvc/KX/EFIDBbsnX7E3Yk7q99iCwNp+NLpAwyXqJr5
K0r2jwERtWyrZUNM0V7I+kdqFZYM4dd4R/jp1ydUfUqLJO+MjMb08l0uG7MrwmO0k2AxMq9jKfNH
L2UKXjWFir3wn90SnGyIg2yqLfovobnV4lr/h6SXUdYDoYf1j8R3GTzzftsd0nzdJCDJwiAOvStH
6p2KmY0fqWLbQZcC0lu1hRR07+UkcYMS2E1mYj6t0nQusm9GWbpswFE6z1Yv//wJMhiWFX1W8fbH
YCHuBVF+S0vyFocZKYxqnBJ7daR4s/oFV+rkpZL3f6w7TfRaeOnBcgUzGb+JeVvLTgETr2QfzJw3
IRulMH/efRYdl9SI0dQRdjVtH4njVsWVXcT4mF95I1ScOuy9OPmYxm/AVqyLpp3V55+GFT/BXETZ
Qy0NavxX9KsV0y6EOUKZPIPox6BTYUytKxNGGDIedsbjdB6nee9Yr182OjhrhR0h/ioEelmB6Vf3
77fsk9q72PaYXIB1B+xDIDqJ9GyRUJcS7Osgwkljcec+ibDFgnIVQfvSb/rMomUJwUwifUuKS0xh
K2T8OVZeCJmXkSWBQtdKa5Ouj5L5c48LdGFRbThyHoTN9eD8iSljwcme4i2oIlvwWMVpUqntGxr/
FaMdpWQCtFtcdsLPfriJ60SoRQiTZKAb306yeX/Xvd2URrnJkNmewnegLP+bXkynndQrV6vqhC/R
UZXk4dS2HZ4YIYm801a6QS68onZqjbA5Lk+wnkSJlxQIkIKORvt4WEryY8kMsD15LzDl7XorUCNb
0ZoL53+2O9jOCkDrXqU+cUV+jn3YSINR0NQsOYKl+hUxpDQkMbylzQ0vlcyy/slC3KXX9bUAdDst
dHcB145yS5kkcpv9zTA05q30tYWCiJyCYOi19+4+IREGT7oKtjSi/Ue2HPQt0yiI2Ij8KPjDuBsJ
i1+HGWClXRGwXa6OXsIGqdi3yeSjCBAbjKfN7ehCfXjgiyClcfSSNTYT7wGDGTILuqD4UAa/nh7c
U8mObq8Qfn4GljBowAiwp/JYk/u8LdXS+5jf+bOoludAribc+c9Tgy2GqEySd4EqeXoXNEU6jlnn
HLNQqaiPiSKHz14VuhoRkqmn53FzEXK3YacNUvZ6RGsc8ZEQC2mlNVm1Nr5jkSVGl8R4a3apDBC3
ef7VHdn+H5LBdxYkeLjAnxab2j6Sl/AG4NK3+pM1KpMUB9rdFiZH5ZFDBch4c62Bes40BcKBBr36
aBrH2GjVuIbEX3UTVFvufK8Gz0R8EhXWzj4HFMzu3Ek9RHaBcbXt6WgVCOtJ0UsG0AtAq2+boalL
uvt/v3wvSF10lxZrGiqFAlzHJNkUyVd8243+EBGlDliPyqKOBzyx3kcJg9OVlNyW5HK2wgEu3UMJ
XV+iaR9dFrNPVNFH1LUAO2Gn0AJi2H0wkAdrsJOzTDDnYpQwGECdpkzm9wLwMtTfUeWSFHXNlRDk
xqo+17xpIBMPD8hpquDV6LzBxLh9qa4T2N+aCjFUZPOSl/O2ZbXMDazYTidecO0fnGLogpK4yc53
Kz7/azeE/kvjRdbC/GcF7m6kpfDyB2LWUfKx+HovrlsftbeJAYqwS7V3+i2crY8o28WezxVLdDNF
HB5r48PsNuzI6e3Pl8kY/lfj4cY9AwCW8hMcm/Kdip1AIpS4+1F0ZSHZ+19gZUfHLLA127kxG6QS
TnEiQSI52kG3cnQ30yo4J2eu6B32+VtJA6m/0l6Ykr4SraKlxYIum+8g33UpRIhKsO8am779+LbJ
+6sMQVqNyO8Y5/Sof6rm2Joa/hJhLWRzi1HbK0o2PCOKRZcM8EATAcfaFfZZxS4zyQumVd5OaV4U
udH/zjFCVPXKP3m/0nlf3FShK1k28kqY2PeAbfgSKruoAryKNHdoQ9yFxpMgVjBbCPOnv7NCAI6u
l9ZeauNDjUbH1aIdb0csiLz9tv9enSH7ANNiY5kwf8UZNAilmk6VCYPuYzum5ip3HanDpGa8Tjzo
0TpV39TdY4FHcpg5NQwqDzKRmkazL5qdtiRjr50iJ8UX+7jHVx6d0Y4EscamF1s/bTjpj9ln3Ggc
wuoSEavCp+51SN7xtFhaa69a76aK7RLwJUB1VrJxxlQkSny1DtMdEAPzclv05aw2ZZxUBTkFhv9n
oOy9WshhAzRxl7vsnQD/YRrMpg0CirS6Uwi9wNrumlIBk8we1q4otBwB2kw07WYkN4BysbFI4i2D
je1h+kCLy+Ic1jUniS3RBEtbzECjFIhxB88GwNOANHUhjfTO7qLxYz1OZNDuRaJxGaJ8wfIEYN1j
p5ORY+DUNH8D4QRKK5xVcsLVB916B9/xY8/wv590cJaoRY6N8+QzqwfvXGkDifgK5swol8p3jkiE
ZvIydUj/0aPrTx1WiIdNmqdxg9ttOwLMSsuNm6kNnsnaB/NP84n9kyl8MOpeIgaOE1iIns4c8DcC
0R7OI0DqTpQgwxNF4sC2km4mkzdi1VxRwBIfUM1vGM/qwo/qN5nMSv5cUwP9GruA7X4F6Z9Fd3K+
UHyNfNcav3UAasFiwzPU1y/fhiFYI5LKedF7rIDp7tTSy0xZwjMMNB1ilzEZpNXhFKISUa/oMHGH
xs88JJ5BJGba0jG+F195Ld/KVfuB7bAyT3JyR13PrTMzAbxtYRRF0gUPEb9NOhlRzPdOK309r8IX
lysnkQDP/bTRra4GS/9hYl3r7FiU2Kj1BB7HbdgodDY45OdrHYr1wS4YFeAay8q6aV6Nktb/IsFX
r/L3jD3Yzi9cvrpcn5rn9/iJUlQCUkWyGAdfxVzfu2I8zE2tMlQSXWIhQZv+MwNcyUwXWKAhFEIV
e54OvCnXzx1znHtD/D6mN2ALk10ihvEsAJJtjRbDXIDgDf5KTAWN11INSx9vVBthH5xYzGVoo8Od
GNikLHUg8qEjMh9EyELoymDejN/DEVBVPsrkJd0Aby6GvftoM6okWhYUfmPhBdEtnWVqtEChzCR4
6ZjGe7tCp963OuE+53HfkA5x9PR+NST4FEPmXzhxwo+5CGADWh6KYMxJ9IfYuGaoLKlCXrquNWaY
tSNRbTObXArBBWlsXTleLsaZe72Dhp4q8B4p4sMWfNiaCC5Yj8h226mAQxl7XpzTsN9UyFJOr0D/
xZFxnPGuFY3c/eKy7ZiTEH7P+Xr+tM1xVnafqIywmnQnKm+HNH1g2x1qRk5/sjRwvPC13EYzaHf1
Rt/FJTse1TRUaDa40usHHYh2i6R+4tQ5JtOMIHBPo8nv+B4SV2vw2tv0mr/M3CSq1WifnhCPcOGy
wJRApzBq8e/89CtesTqWhW1MW6yzEEI8BByeK+62x53SjJj7CqmjPpmsP/AWkX2YP6bqkTruHLy0
leIAnnFyYNEK7J9m0kvOJq4QP8RmeolwN4wHt7xJ+JycPo3zpNDCn+bGT3s/iAMAMNVht8wJwoEK
Ttvj7MF9A4Ty86DydjYopj//ufu0YfYi49suvU9yfAT7pB0w1fBrC0LrCPXrh6AdAOsGbMkUAYdL
rUdjryD90Kq4SbM38g+7iWqfRjoatJ7yBZP6FAL2wNJZq4C57AtZDwcf7jKs3Dcd27HwHFyFVWEH
XkjvXkEojNq3sYddwJtK3Sv3MLBSIT3mfJjub30HpYuD+oHl/2ssaE+qED7/xwtU/eObDPcVu+FN
t6MnlD2LRw8cx0owQQfM7xa2c4PJiqmUQNmc6lgSre9mtTiv5JtnVpH47BrkofvFfy9t2Tse7ImO
qUbkfQjk/UqxVtW8dqlp3rc1cTHV4ZGWOsYQssLExtJ8ZEcmMFMqg2IAxCVAejFz85F7VxvJ83bk
ev4byCTXvuco2smZGPVRk5QNKYa2NqCPe2zyNKQ1Sh3r3j+T0B+gDAB+sUVjvruK+ebAr6HAt2r3
sfBUrVi3cYtxrCYdab2gsATmyDeZVT6Z0+J1EXvGNRmrMEueA9MhTrkMrU8t/881LhoLb+FSwDuI
Bbn9HSxc3AJzBsZjvus7k3lHsJzDdVNznmnde+AXDf7CHKZ5Z6jfqC2dnkrKUl00UglQ43ZHkGYd
dj85bccWSBLgUxdraHQ/dpoyBFk1I0ZyErKeJID0wXKj8SOrpO/aJcedxNYrsyGiTrEj7imFdJl5
/0dxR9DvEWqYd5P3KwM4DcAbzV75I1LDjFUVEtq05TNWB9sCj+3SYfuWALuvUGBPrcdt7rL18De9
JoO2TymGgTMAHrk4VQPgzf+vemr2e6+eGDenxetK10oxEqioZbI7ROY26v4kKDG/XMvFQzX+SOoc
ko9FF076euzygefiqlONXSGRZQwu6Ilhl7fq5bH+gi2L5tvWKr5E+em0SNxiHOJR363VXJehtjt1
2Fw5D48ci++U+l3Hq31ti4ZzeRFSmPtKxyYAcCwaIsKeEDnngnosQaGw216jrkSVCWVsne5lHd5C
00c44kqnW2UtfJyLrRdNPVrPKwhVW00w52BhdkK/3PjZrDBXizmYjYtNkPNVsM7QPJAEqySH09kw
yIDUr2FUvqoSjFgKjwLMdMEdwEPtKt8ZiTSqL31lseBe3quz4CmHEKJ53yK8kJDiSjfOReNkMlm/
/+G/ty31AuHbwfvMeytkYtMT/hph6LJ2K/bfDQtVDCOzgq0emUlEH1E0wEgmQzVyI7f/Wf1fa38u
QHzpS9XbF5pUiIXbQBdfryJ23Bm4XWOqOJcs4ZgSx0enkzwfjxm2OXfAykTUyab8qegOxYopTVJL
6GN+NSd13yao4hObSVTZ7hOM2qV9oEI2xaqIRumz6iKFjpcueSXgr32Qmnz92wprnmUlzUN1LiZ8
ScEFALe7tAKXpK/KgQsq261biFIVh6F8nU/7hrYprx426mnf2A97bmR/yGOlq0+rCF/EM95sMksO
8FVmd0v9vxB7Yf/s+3vuZzblvcezkRpEKozgkLoNMHFMVUtFlM7VcbJgxsWqvRVqiWbvtlMwZic1
Al3K2nAbFaGKRjpuLkUhnuzYq9XH8fYWa59tZ1Yof2wVMIy3y9PY7HAJVN/RSFzoxA9KBTYxT+//
69VgFpdtcW6DumxnZxzY6yIVuqRDXaBKClXCE+XhtxAAiaLFIRjeoRJp0fPQfPeb/UnAC2iwRlQI
IDD0epmDxZ0nv44TmymwClKAbnlc6CwxzUQpj6ZKfZHaKTTQ9iInuQm0Oln/OTlXvD5cxV3ogw+i
mSk/sZ0F+xnJ1fPv6rOmkhsQsyiK/ih+4J+DKE3sv9q855G+9kEtBXmS5wAVFYSnPkKGa9fE2act
Kxbu364gkzTRK3USvFp5hPZrSaGPyNrGyZ+nuhBircOEnKinj7l1Rze11l3N7ZcQ+nEzAWtT+Yb/
pjHj4qumdHMEp8gjnnrLQk3FwuSMAatemx/6gvkd4+xIgYGSncwBaW2WyRbGoIpFbEbW6LbTmOpC
2Qkjk7A0t35GQ4A+ywHS6yQZ1fUFA2ibxPpX8NBjdaqLkZR7san8YZ6qvVhJlLnmwlDcXMMODLXL
6LpRigtQGvDE3efx9BVQHj18HNHmxTm2K78gqOyKvFIu4+spd3JQ8YAiLbwdZEErHEgVSFSFwSG3
MRYB5rQRzQLHKarO/S6ayU7uT9VJExlKoVnKsALPuBziHFDakTg8yAJs4Kv+VXj7ePEXONMVjqCt
vSUk5bZ4j66dPKm3mMenyigZOfwpsNSNKdSMZ870/b+wEvUmdjLiTTtjClmEX7viCiuwG4rVrvPw
LT71ZxP1Z/9agK0ni2py9zXIqgEuVOtU1ud/VuSeK1jsA6LxZkxjxGPMqNQtyl1lQMDHv0xCIF9D
gmBk68ufRQXyB74ZKnxbHAomJtSC9UO+gvCC71ucbTLgHk5hY+5IYOMLyKBV2pj3XboZws1y2NXO
rLI4A+HS/dqHGmMPsUFffLU0dkQyJP+EjNMk0oE/va3A+kktw24TqtpI3IWLWMyALNkJvl+3BV3s
m4XxHfb9wyrsjku8kEDOZoP/7V1CIyWmlvbrrR1MBJDCp4BHNochHQNJPonv86zfTynuaS092FRY
pAY/9rdJzKWDY3EvXvYN/+zUuIDAaWsZ3lXXtsGh0IIWGL0AYaOcvq6SFJb90vXipNzCnJ7vpwom
R/yvHkN70JQDBbAit1Rq9U8eRYIJLoStI8T6hrAQn85Vy+3G75Q9dVS+F//NrTfTnb9O8O6JkxxZ
WOyDcSK9bIXdIa3PopatRgZJwBaK4bMOg/RjCsFIfCWgA4U833LBIxOi2S65eLfSwjNraEtJ8Ce7
LHWzyuKqwoCbVl1V34geHsvht7UlSVS7122p+1d7qyz2OeIcSn+9IS5L1BFq1sd5AJ8OP5N+YQPR
T6DthKU0VOSNlM41sz/+KxUCwgWebTjPMUhIFbe4EUrNgEIKWPvWeWjfGfc3uc5F9/QgxIdJHFEY
Lj5aauMLZsnwvbXEO/YQy5BQkXOOynk46jdwLGGVWHkjo3PjeM2VrPqd7pUeASX49YwYrq9ydyml
g+Sa+MRX+27U80bKXQMbjXvWgivHEY6rkzuTMYagdQn6pOiaZ9yZI7XnI/ZrUutZF299i/MMf6I6
DwJZsir4+x9Z2Yk1P+kOZpkjE/SPJJrkh/lNjwVsxl1U7FjdWmVjACGJ0wf7ZtmHnhxu4EMNFmRM
11oEtQsOCwlvgioIWur3TX74RbLe8xjnq6fMyHCnjuSZidt6oDi1mMjVAJ00iqJR93DTDmjYOA1T
kQpzLt2SeJe5Qu+Q5ZrWQBqWMjCtG2AUt73LTxXr9V8AD/1WcbYQIYpHli2al/Ka2Ct/waM0XMIl
LMsguB+4oGH7ZjJHImFwWplGlfJ/9PXCS81B8hdr9r+AeYg30m9gg6dw1d06Xj9tQTcp+9tg2q7U
f/gu08gILqNJLgskJJmk6JBJQDYpRNaCdPKjnMgFBxMUEqGtF8Xz43HzeLKuUCmwHKyFfPQArXwd
7X6FGKfzYw1DtNQ3/hEPC9hezDA0cSe5CLWpzDOyClIflPk9NLFPlEGJlzkG9rNo9jzHzRwCN6HD
gAlnFK8CEsrrrEpH0D5fhFe2oHIIjgDFo22fliWU1gsc+wjx55NQYJm+gqAF2Vfco8YWo0TjdkQz
gUoOb8pniezIMyJfgMjIIrEkcNDSKe0AQB/0tcZX6HnPkW1iH/7vtbe5yphubYqfjJ0eYRW9pTPv
1m5PmJ58FOJ1eiXmtvJHg2uW6b/RJejcixJ/wg8Tz6VXYhs7+EI2BbW4S7ZowRqSGdhtRrXUS81p
3hBe+5ltGoFCWn8jr/jHv8KoSs1pwDrijVHPcKwMpY8IxT9vMztayXfLDOYiEMa4BRQVgYLICGcU
6XHYVkAyOlkElXFoKb5Zgxt7LYKFH8SNnITIA+F9EwG1yr4NNAdnQzeWOl5JpMPLNeP2lUMy+KuR
DVIAB9lEuwpF24vYCkrhNe7nWWpOHbvTqVlTvMO0yirUBHq4bupr3qKfHy7hrcW/fsV9zQbvep7Q
BecFENBC6i9ZtfjxzMrTneadUniil+O55R7kSZrWwvnjKH06peAGHb583NxrmLmrweMpMQG6QydG
zg1kwglpKxQ0AduUsqtYwnMco5vnR6lsADCWR3T/MIbGu+VVSpQ04HY9XfkpaSJJlmX70qKmDa5u
GOjEcwnKIwkinsusFYPjg9xL2iXAepTYFZ3kNWULf4TzpEjX+xjAAmynLFgjZRGZgoBNRFPICDO/
XbKgo12cE2M5WhHi9LA+GTxsq+Z5zLFvw9nBnrqrgvdN5o7rSPYVi/gpNh8ceIwLh8Wp3nncwWBA
t8mqIUYqHIexECSW8VSXvPs7ocf+vZQFI/jL07JkXH5l6WVbAFxSw8uZ8qgcSg9qsJ8QGHlRVdJG
RenF5TD3929UtiUFWlgPqjkoeny3pstIzirKfhe8VQkSxN6VrdPoYb+jif/jWoS0lbBAZQgPGh2c
/P4/8a6dq/q1fcwy/HIbgza+5uz+m7Em1xe5Bvi/bmKl9iRirNVM+tWDS/obj2/IFQqVi0JHLt7i
XreghVJ+5EIIAhIBR53kDAo0SwquDDj0aHEUIBYa2WrgzxkdmF+PLjhrEHgVLnB1CWgeKVcV+i46
vxtHBQ9M8u7z2Mj53FNN/lF5qtNoKL33v2PGwa238g/FLGS+m/x5ZGGCkPZmzCB32fFFMXawbSst
50hZoCTwu3tMhz54NpzH7+8XUhTWOFEbNfm7K7q03rhKgfACz4gGZrbfu/O6H5EisElKExnvqKhw
rgAWaWQytOSuiEGegentOXjlu7+8zTslK/xRAeC4KbkpZ2Ih/ftbVs3ErsgvWrlwKbh/RNgdnhfc
EQTMnpVAAhk4Yw4g4IVjp4qGwBYPv1X6+hUxNXFJYqEFXVGZ85ibfHrE4Nsm9MH/enRkxx75uP2V
8gTlQ7zBk8O+89T/GQehJocf+LmLWSYVsVlt2mQ1mXwmsHM7Lh9FPbkUiPHW/0u5wgQR69XgG2hc
t7qWuJB/STSe2GQGaXpOmuTVshdS/If/jYzb2txW+4Y888SgtPXACqOZZaTag4uqdgpUykoR/IZB
Fj1mPxvXai6bFcS0+qPc3SZLl61QzzGq3SHiKCXe6a/rslhb5IQKqrfoIvPjxrVv9DLrS8gnnUVt
cruyEDG1uN/67GKIDDmHxdNdQtHvfgg5RTgGFqILAQZGXJW/CB/fUpNlqfdIPgDqIgOQm+bam1Pn
HhAiJIsXBbW2tQH10Zz09xPAgvCjUAXwsa0cFjUVakqusSkwVt8OJURqQDXHmRj5g24JMi2TrwUB
sFZLnnLTPNI8kCKMNizIqiby/aaL5imUT6GoVLl+CLVnPj05wYduCnkSM1FE6XBhXm9asRif63ny
583OFSUsBrXE0Z2EPxkW6dBxi4hFvhcvHdHKfoB+ZPn8ff/xJ/khKEsVK830RKK7ebabIVktaPzQ
zUTY58nSv8hm+rMAoFBbvP15zKFKxfRtpKcw2c3UPTaxU5AW7OD50ZGppaJv1eu0EH6+/PlpZfxs
LliqXB1uB3S+77gPmU+NfAt6HwzffrOdz7gpV4UPBUSxIrLNCPv4f2kw6Cs1zTcDwxptbaijIuc5
NTMxTpvcuszmkYsww3RoN7Om0qGeWFZ/3jnaonIveKOzKf+PhsAsnOi4LcpUIXgJUNa+e2a2E4Ws
hf9gBQGxg3sVB7JShzgiZVp3z9xetyfGXTQFfqGfR37jZxYfMEyKu0vlglQ8wCkb2yDYFF4RASUy
cV3oN3uHaYv5uCSfRGDO+r40gKa+BTICg7LQMw1DluEFTgms0KaWiJGK4/J097nFOSCkBwNMRydZ
mj9qhMnwDZUyOZ5LzV7w8fbVY8MzrUd/yJKWkjUkuKo6UjGVD4ByNL4v4dr4z08fP+/9dUk3M+iK
xFUcaDCZzgNv7vqJg1OutOwBFY4UkMCY0lCR8fY9M4YPc/U9e31NPO2Jf+ObBYhJ3oseyrc8h8r7
tVI2xmA9dC//ISuakGnXvFxrRhT0G3r+YSA6dLPQuPZQ0kcAo0zhXlpLEhJZIf7dz82xwbc0QbnH
inDGTYRRpYEVmy844Ye01NSX/3DwRfA/TtN7logUz1prRf8FpJnyKlfqrMiDTTeglX5Rqyglvjqp
DVu3vBgNKT43zSvmKlKfajrWl2WT3puONgYkML96/oaTDb0mT4igj8l8/tszkUHdIuWt1h1cvO/Z
5E8htMXGZ12VP1/CEqabuMQpTDksEPlApMWg8D3enyJjCsHh5V/d8fqoIGRRsG32TuJKyclDf9Kg
Sym8qSuJCyyk7zVIlvADC9QNKEmUcoKYEL30LcMcVvj2GshmFhqyl5zy/aWwunBqi0165hDDnJnw
/bwvtrLMg0JiMxSs2hNpk0cAh9SPU/zE9SMQefV+y/9cucCk7k97h2U1LobO8w+BsOW3HAszI5xE
b3jSl6q4N1+Ip78TqAe1CQIU8bQcrYNgR75KbD0CHmlXYnIdcfzsFUp7g7orMd3J4SUOhfhULa7Y
GUC17ZjpPGyvrdbVlhNVP+tYfEJ7d1EuYgonAVL6/pGw9z7Jmujadt1Ev+cg4R4XAjUe/LrLECqC
Y8Ut21fZGsXyp33FPf6w+baIo/7n6A/A2diELY1TPHGjU3cBRDTl2AuYZvzWmEtXYwS4z59fJJsk
otovHuc/vFWuNk+Fe6UwG2D3r6wUHHWwSAIWcgj97wb5o3wZPWVLJuXtEoQEhtyZANQ5t/d7Oo4d
QPAdsXa2TkWKp34Iw+hwsa8bCOn+gcMGaMczraK02cV1x6EG5iMa6xs0lgkalUIVkjtusQQhi/3k
X5K5URlJQV0F6Vm0ofvA2aIKrF3RLmbPQ+BsacOEVs8Vp0KkiH6oc5sSKFHJOPs0MNoiJpPG1T20
7dH6MLopl0hq6s+WQQ/0/y5bb/MBXN/FnaQIRAc/Moyc6zW3d2mKlTDUSI9IL1DxO7ljRyG3iWMQ
4KXUjLic53u+XY4FZpMmQhsq7XHxEyYEvY/MA6G409eBpAAYH4XeOhkcFY+CKCbzxREx2uFNrGzE
9jvCMWROQuB/oVjIe+5iI/QORZL2trkwM8FVzA8wkkCOsCSy3hM+ISVXF+77oZHAvt0DSV9Dk+ah
j4cf/p0Vc5YfsjAyUj52SUwZbo3iQ49tM8HlUipGWeCPE2xbms9lZS5gn8CnDG8JwwAL2p/4CD/v
I7no5QMm0wYXSP+7Q8cNLYZKNwLSl/eomNoJ/NKFRRl4ow7ffEstzVbFpDEsFyIa3mNfXsom9+AU
N2WSnllGKbuAS7ZlJrQMmfexKTT3qc6WJC9K3Y+zPPEdmiIq+6jMQdToWltZc3p4ENEnlU+eIELn
HUQrXV55qmRROfgkZDA5spBjFP66E7IsQOWe4x/g/Ocbjj6UIYgNyulMVt9NSr3mbCEx/fTFumy3
m/41t2A2rIZyJ08LEtp6PxAhk/94vUgg+N/HEPgvSBZ9RtEQ8pmX/C6eH+Sd6WXAop200NqUxJsp
yoAKi+3YY2GFUAD3Onl/ZQJ3rxk0nxY4VGnp35i5ZuOe0+0q1Nz4wNCZ3LX2Qxv9V24tNF/PgDqE
oYXQlBtujaXYsj8SKp0wuMMfvDF9PmsgnkvhAmDAnB0vY/1hVS2m10SWEcdVKDmD/j2QhieN/A78
cWckQOU6XUUNUzuJbU29ZK6JKPsGBno499OymFIgcOTTo7g5GObW0UzW6M7to8vmkTVnouLYmlbH
WP8GLJVQ/jec+pfNJ/fK9opp+AE6FtmuZJDr72PFK8VJCmGhJay2SdvxcHl19//YDJackhWLc/P9
Wi5iNccWOCEn6Yd9QHBqpC9n5IyU0sUDpC7X/XDB+KreSIFLPo/DzlZM5IPfcan3yA2V+EwxVLLF
LJ4KdmjVXV2o12h8eoxM7c+BkhpcaEdUv4ojIHqPIsJzc+VvS7VOuRUdBQA4snDfBiKmT5A5HmBU
KDo3e374rZtojyHN3My7RQd87Vj2TqOL+REHwYaZSVnc8fooVmQybDOwci3mz0dnPm1Z27rH18F6
m4Il7asr284sIa2EBi8SvJyxm1J2m1Oy+lNZfqIshREixwmF0EIhTOAfA6P4mtGXaCcSS8pJ5OCL
ln93B8ULnljMXWE/ZS7VPO0DRMxLGbYWz2xY1UrgzL2fWScR/WcMzb6qj7ssIe3ns9sDxqldZ7xU
xrECZvd+7iSqfC1TqoEZb9NdvPIMC+SnbKsvO1B57GH0evfx59lsIYO0DTpgVgdbbWcX18viTSEA
//srHT6LjyYBeHhye/TLRw9a/da8hhsHzJ7Hrq1Ov/vIso+GnZsk7KCyxvgfN0oAy8sUSQbUBaT8
mKdA9P75Q/PYbq5erdL2YbmM7weZT/XeWTBGER4tUA8DchuNNmoV0JjuRihy3HDjdNX6TJ10TDYn
CItb319XmQs2HNNZ3yLV2ve8mIKRJiWm+GqBcFh76yLsAmOwfE0JEUlQ84EV4W3yB0rAGHkNxF9Y
e9LKRuG+UL/YBI+AXhtYjj/ezucKo32eusC7TGESi1g75y90BwE0OUI0cquw54q6uNUiSYD4r7Mf
0sVJroYg7dr8oEKLda9rl+la0/3lgosqjD05ncnArTYqCRSOaETrzT6LaojXFfv+KGEvIl4+0+PV
VGx5G7rhpTWVYwK0j6TfRTsq0/3FUQPqDRoDvrQdPM9HRZLC/qVB4c2Egb9JViTq6VxoQJctWkPs
1NOOH4dIw/fOxwQycXdh2BzwvCmFPE2axdGslCDEQfDA3pNSL2naLezcpYlbWeKeiS9gKCHTRUOU
pg3/ewpPfa5AMiGvs5by4hhOaeJ1BYRpKQV25gD8mQoNYp/tLzqy2TK5GEHtgKnrk6g42X0ARaxd
R+/uWNupEZu5+P+/f91TcfqUHTSo1eGGpJeUB8ZVxGAWb2nZI8kcXwDz434XQe55ihUB/9Gsjzw8
Ev+7lB8tW4UXnq6RBb2Z0sHluVM4z/qwQngpjLyOUr2zdJJbELzd1WNYFYh+aNBJ0QhzOWI6ByH7
MF+6dUAiiVIgQ0HfZvwSx2/4ksRc1BK1H/pKcEATsceSM9sQR8LUkaY6U+uN/iOY3qcxlpD0AkZ9
5yJCldaiNtynTWSZsYo1gooAY45daSVsltKkNDfenw7KM+lu2ocytyocEVoCmRGEawkXEspsJcAx
9Vd/lxm57DPjm1tbdg0I5YBpGcYYjDQDPwI5HJMcxLqQEJukfL+0d8wF4ACjXV38ifqpjkrHo54L
mm4fr1+7ZQj3/UT8pHR5JQh0AJXblcKoFDyWtZjjmgbazdGfrhrcBT8H2ux8uycvU936SrSvYrZi
48iM6bVldrSNs+EvvFjLvfhzAyNakZvG/Ip/hLZYJCPz/Ugr/f2DJtPZxSgZO+eaWWbV2EC0hAin
WMojZ1/JrSGUTgrRPJx1tb/yeXyToy2KzUHX3OyOcLRVVX7BMXHXrwxJvonpa1ibO0mxV+2Hld/X
anW3Capk5+jLUU/kvUXOt49ZiRsAHYS/ZQ0q3wRv1+XAGw45C2VUuxVU+1OIUoUy3sTbtKu4PeHd
Rk1h0p8qgRm7xDaO6r8VCoV2swF3xNNRpsAMPxMYS4HeAKKfbfQI+wjUTMboYgVDodo283Q6HpJ9
URG2TtbCzVbUR2zTnXDmbN+J4t6dvkkbzKWOfuyp/gbnjMiHEAPBzLpH+ycqQhUR/RhrJTtRxsCF
iuYvJeSQKnle3QoY2KwTyTMgQitUq0AhRolsJVY8o44TG9sbnvaFWYWNM4E9OrEL9tpkWlpYaUjd
fw8FPbj9mCkLELFEgudso0DvYS6EiIlXduiioTUxpT1goAJFZOJXlh93HHtLKWofd+kXfu3SDx2H
yqjgj3LY4ClaEdSbTLmi2wZb+DVyJ9zNUE1qf3Z9A0Ijb9KFTYeD031XU2Vs6Zh5nDXMtnNlDQe0
LG0gRAtBE1earC5IjPQKlvlozPXCfXQ+TuTakUR72oI72WXnJwqjT0UYf0+CFciJXcxKa1xET++N
fNJkA9kHfTnioDI0mnwsHERt0W50jROr6JF6lx/Es2R+OOf1Rx6m3WGUMsq43hSi1coRnwt8ld8w
DQBoC2NePoVTzCxdbbRsfZrfBKsgZ73KRm0+0ivIoXsPZpED3V5cOoxYcNlU6sqCL2ST6Ca05GHd
XU7LiuKWCrq29DbvRo9QpuFE4Z3SATSFCezk/Xgr0i1LTEWRPafsxRfY14p8TzrvO8EoFdfKxXba
PUI7fNdTw/fbd/2IfC+VrLWMYIXPek0MmtDW7l5aPjNUKw+kNsog/ts+FcOXeH543cP35P7m/xID
8I1cENIp5lYM65GHozV6oc2xm6560GLH8wN+gkgN2D/thjOSE/xAe/bzE+yG4IOiHz78gwNo+byg
eVdNUv1NS0agbuY/Qp3Kwi8rqFJprV+CZZpxxuHhSxbOPbqA7JG4Wn8V88ZP23oEqlUaY10hUO1r
ydAbzwHUxTN+rvNmj1o+P82QJ6S/J8+W4NCUBESDwXVuFF8mdueImuHlOqpu4mzRa1luaQQ/SQDG
eXujynHBnTeJl3rXKkpkiRwYaTc3dsp6AH/jK6K/XqsToeKlhoK+Yq+mpoDFxQY3i9g+TwaA1qzM
QtS8ZI2U4E2fbINwpwxDNTWFZIVc30qbASJVjAnS7YfpBE7npcLSH/igKx8KfTNSbqpPMt6XUwFU
WBCEviZKRCAPHVtxq4M3cNmzywN8aUKMqaGgtir4hO2E3hse4DtlSjhCWijx1l/CAeoXopmOYu0W
v6HsiW2uW1/hdKhUYwq+diGhe9dGRm/GQEFUIgDN3vljziJdv2AnsV+GOLbxCNJT+fEOTsU54iSu
JUe+/wJ1XYEfXSB8ia/inE1w2XqHaDgugENKdCUZyTzEHfppdg9kzw0P/dU1tDbNOrZtTJA6j640
ndBEaoWTh7KCASzv7obfThUvRNHxWd/eIXAlnMqHFyFzjVZsQHPH/swSUpEb5lHrop+6KxTw8O3R
C/kbXVNG6pktiTs5cerDmdC29ixPh1eV4TaVzdtckaxn4U9zTqBAXbvin2MPRlFdVtkhGAdHpxYf
KwbI5lFJFqaoABnmla1wdxrgpAdqOuPgnVYfSh+ayA6cC+41drtqbEZInQUxhNibrStrGsuB0PoL
YR4yHeq5j7AXC9NjeFD+Ezcn/EcVU9DAUntVqTsenLzZvcZiwwIGIWuvhKpLYRFSiwNvG9Hc7T+e
cFzto/MY3284TMcTMnXCIKSHBzeY8ZJitbXj6Sk7RW+Q0VlGfTPkVfAqXMFhp309IIDIQgo5JjY6
H0jcVUXIjtlaEIklo6DERA+O/SkmHo/AI6FDw67cT+e9m4X+wJfK27OFuYJSKLTMcnLTRhgxUNMe
YcT+23QZ/nqjqXd5ylGQjUoP3dLR/9X4RcpKERvKobJOmMd83eFdxvCVVQaL8xsWj4Fa4UnHPvXM
s707tSIxotY6NnDsMfgg4i9D2UOHtSkhjjBrhqL7kz+2f2iZSpF5ND/UgYs2oER4NPfCpjd0vk0T
zg9W+N3ChWFBRB0t8Nu8KtyB1kXbpWpnWPLuhvDoKj77AqXAC7L+tDBplClk4jcWTWlHhE2gcbBy
FqiNuyGo+NGaFKKOj/Ip8mGbxhYYqCOG47OdMqhu0te9Zei1tpGNqSRX2fEyQgBqM7DDn3Xv+MOa
VDcVht13Xu4oC9XaqeMN4/lhggjBGAvgT8O1t9bqFLdjqjDNw9LhA2buxpGfVtcBnehP1I2EPEWn
cP8TNeVi9FMfjMjUswVJy8X2q/7Am3iGLPS3hU9GUBl5MBX9ECr5d+bSZSK6PJT/6FuR8TYzFV93
20AVon9Mj/+ypER47+a6YuFoyYw3l7p7LDS2p9AErtJbEy/amp+xF1NSiGHh90p7BVUShbPsTSzi
0hvV6LWvtHyyldUI7gdgtWgdjFPzJlhepdGoGfpPjmSjaJCLByXrnr0sL7mlo+UuY66U/X5cVAoa
TgYlr33AwcKoofYRdkfYZ177kkz51qRpSRWL8ZfCRAfQ3SnnthBvGSeiz0vu0sCzOIGP80/k4bhc
EvPp2d4xMRws4TzGOzA6zuTbgXBy0Pw40bN1IJtpoJ+rtj6sBvXtqGEPHjrBdQrbgUsx7I3Y79D+
ELGmL+ZNfOXFEI/UQB6SRc5B5I72ZjLua2cERIVGeYUDFVL395qesZy+D+LeBBb0/ByKrsrSmyLt
KwCyxdN3WLOSrb+E6JoBLCbU93pio4c72m6hjrU4LHXbOj/sDip2TLEYamNTEwAToD1Jo9okN8Y2
KGe6cfSQikw0KhNZnO7vQOhj1Vzb57O0n3t+BXTrM4mVdYXBxcfUixWC9DoSwKp2v09MBxrH5NPq
nVuPKIAaVScpk4Ta67QOrB5i1HcPKKtkQZpFZR0z3QY/f6fWd1jjU1a/QOWU4H+qp7JlYEo+hCqb
I7izTcOcxMKo6zgt+0AjRwgDLnFW80T/M/TVy38OweMK0bW080eT1h/nTHQCEWPp2PXomIa9lQTt
CAiUeI2D0ikOlQWRLaLJRxJobtQYeyiTAy3Wn8rY4dlUyUsvHpX9UNFXSLjZkv5NGM9GuM1GeCE2
Qlppl7Jk78sJLorRbo8LBabP+9Wr4wN/Bqp9gLIhFtYOpZgxnIwi9u/WhDgV+OaQ/8bRvo5N1hBu
QJMMJAOLNNdGNyXBgd7rvTbrzc0vN20bGj4uk4WrEUKHpq4mZH7V2WG80mhAEJXOqTnYr+sMpmf3
r3yD3l5ZW7zcIt7B7WIeeVhADl+KKHAWc268fJ3NfgXczS9Q2BD50whFZsDAqH1EfVFDEIB39pXJ
End8Owj+1o6YKXz8KOWTx8QxRaa7t1445DTVNky284gXCRnkOpcfHsEp22FOs4fwJf+14GWZOVjj
ZesXaUEcIfnDeA+igPxdqhP6we5wav8gys2+pz8SvjNqZB3TA4TrhoL7rI6KN/dMGCkxt1umioaN
A9wq3uGk7p/Z4MHO6BZ7059nIcPgn3XDTq1rP6/Hfv1OWl16e80ukjaiSfl2n2IEwVdihrnGsI0P
GWWvqBsynlJ2azT0xTDEHW+G1wfsdygLzqUppdxzkGqUmqhzv59siEWbBKHN6NZQ+GB1wB00FZpZ
lgC3pkCvnxVMR71of6yqmwrxtvcO4zxQvly54D484kCEvPfth+SKnmjcW3chUa+KNElzVm3wtUZu
d5GtaEBVs3slm+PFvsGhMwg1Y+vNtwgU6xXHnilkK8Ifse/Z1siZ6lio+o2mCrNA38pwxmpkvU6c
317oLiojxoGi3DU/Xww0cdWM5QjUeLqYx4O3MvGyEtoVqs+x0rOOAvNTlgcCY46hpqELCe0u5TaQ
3t/jqMHR3ak4oe7UXZQtR19CYI/GVklZu3rP8hbrrARtkkua+HdX1Q8WkWTczlc5UCa1SScxh5dz
FN1h6Vpt7hhzMEKmyRXFtghXu/SOq69vH0/sMk7L5E+kHVk2ZIQ7LPc7sh173tv769Et98EEZHus
qI7XEnyo/Ja96o135RUnz4tPi3dzTaL01c4wZogw3Nhw8vDh3p8hVAoSrJJ+b5Dtw2Z4cnqsQaBp
ZuMWh3TcvWEOzWRqEphAc7g9Vs033GTSuU8frdG91oS8rvKqxb/0N1sAM1ObJMQkA9OnhcSXZMOW
nPiQJgIW0KLwybhNA+Sqrwh/ysUmXxRKweFb5zYwn9Y1b2vqyMVzTaJJ1nPn9LSah1tCsbdxBGjG
IK4wMGtZRHXq9b9t0FkzBDdY+t2TNEPgQHPywCwEPRLjoNwWduSRIXAwlm1hVwFciYHBEJ6kX8Fz
KMrdTrm4PqXo0knIlA7aepGsSqfOtZ2QWwQk0lMdH8z6p/KImhtwMtiUNgXp5Azbg1DRgwiOBQMW
5DCHT/PVEqBiovgiVIIk+MSXHtW4Hmh2ZzvOTLFnv4smnj6HJcxTdwcg/lUTUXX6i7nDPwQOhi/N
Hd7RqLso3zKwpnkHOQUlBDM1WXp7tsZXFujy/P/BG5vYTDtke8pe9x5UJySgPWapKIe0kYUhO23e
CpPKU2ldaq1ks43SqVXNUwJIY//0ypEqJwR9rrO7Pgnxc7owyOrZsy93V/1Agwe90NpBUgScy8xO
MGpmAinv0BD2XHmBMQMZ7ULWu6bMZDNsh3FbTGBH5h0NI/bR90eE9eNFVcKVBhZiu1hfqY+D4IJz
GGFssZQKDRYZA86YhhJmp3vkVk2rUUqHP9Q5DiUo6s4fLFkd9acbCKSG+l8ZL5ZKt5hc4MheG/nw
/eHhua6IeT5lWksMlKaEj5hexZ/bDrkD0gkJQ9NB0fnwnkem6amJ94B6himLOVMFNPyVVd+gEk1y
24ohtzOUH2opzuE/nqNiOgN7Oo/bER3cLtXljD09xlIxzUyY6C3OTWwPfzfOfavZ4Sc6MbyRMPBq
Moneifr1cO+Kak8ZOmQ7hkwjBF8LvIaVIVFP9h1v4rTjIv02b2HgpsutP5rAqt9jsMlOCEKeslvR
sTyy5iZVq99ehHaL7Bpn7a7k1rG2MqQP1+CxNxPkHl8Aonq41/4ITgdDCqj+1KviupaA8e2HhnY6
+O015NCTt0N0Oc3Xln6PsxAGO7ydQ1HqKZlAYudMMEOTjXSL88TcZbyyOzuuGnQmtVxp9BxmlLN2
xdEZT6aJu9zT9xB5nd6h7wcg2NiYFBrqfEbPDAKuTTkXQFFNmkxgLSWvl9xg2UNR9/J3DJvoxtIE
0CnfrB6pCAk5ZMrZibvV6/nhcm9cRIayHNgWaCzsa3uJrMlFAGBV8E9WweHsoUynHHiR4FwFAblX
KoojY5J2NefxMsVPYJDMen7ZPwXZhWG6AueTWYbfmhbG2tXVl5U8Ucq5K6zdiLqhWCbn+0l8uUJe
MocH9O8erArmTHwUF4V3K5hHcdzY58d6njTn9YmYI3gxv1VSv3VdE3omXXGg22qbvtJ07hix2qER
S0O2yRJEOHjGglSp/1qO9YdRO5b7gMqJCfTGfrsrFBz0Wq0WM+knk/mPyU8nRTs0Pclh1GaDdHTn
BAnceitE52a7kO50KABf2LTAfAyzHJowp+QrtoLsDWsff7f0nK5fomlWqRmYXaWInnbIdPgCxg+a
yD1D6dxkxY1Ri4xcAeVrgDWjnoh0zR9ZnW18g1ts5Bnzv3H19QWEmxH0sSCsT3n4lyd8Og9Hu42E
NseJRmcVZZIsNfqa4L7nAAkfwlwgZh0kxBG7GRT2DlNEtt7u+V1i3ACSjKqbKr7BAyRAsJHQjy0y
AjTSrNd7D60KRyaZdsEDbEOCUN8Ph1BPTrx3iF5frS5Za+04WDrDVKV7rqfbWs1XQYXIZe8Rc1zp
IpaWon2YGhBCYV1VwokoH8zxureqDRiqKa/fDmjuDA1soauCoRXWMx1wzm2P1Jg3zlCYPgE+9o20
7/K+BmmfOWJac2pnW6QA0avxq0facZaGXR69djRBLyod0+eZ4+mQLATzhMAnRVE+eHRq4hLadWhV
vwfD79KKm6sidlQfgjJVlcO8e8W7pgBuIw901ttCD6CaoziuKQZydpmgQ1XWiq4XS0iQnZ8ptp6D
qd76nd1ZuQ76BiyMMGjnIK5A7/nV73TmgWRpoHV2kiL2ulil7Krhz6/RKwR7Jp0pYlSnx4dfeiNL
xIiHjCXnVwMqdy525SBc8RiMhWdoAB0u/w4JDiaVxgSfU3f7We76QKr3atYrWAM3Q0x3kZvKdmZF
2nyDkBO2IMhwMR3jqLvAIKPxC8Dm5drsZMIZNg9J+u/+8mPp2m8zKQxFwDsBTAcgTfws+Y1Tzg/F
y//MG0q1rrrPdPBMdF6arDes9Sz3Y2n84EkjNB81/GeU8OOOwlE8JtgIfktjfekpDXszzTvciuiC
qk7haYdQWN+YEUmtxiPNSlaUPhmN22goA5thNyts9/qlrOQ94SbPZOLTgU+dg5MjIMG4hXQQ9Bwa
mx/uUFiGxNsLyRNgKciOl2001N3YrrN+BJWpQmY5/jL76RzD9lvnPWvB+JLPGbo1qO5wQG+u7Y/C
eVtLxcYIGqQGrnml8jiQLEhJpHq2m/zXMsutBEL/JeADXboevfxOE3SKxOfKJ18t5FuOLdKNnO9D
czzPaoSOFcHPFsJdWhezIiod459KEYGGmMYuzXHnGKrpqVVly+A3/0RKNwlFm/1KTL1enxR5LDvd
C9Yg4H/3cZc3zOYWSo5pHkoRqVCB0Ric3aEfNHKymdXTqeNpR8T/IMxkA8L1TMXjM+vo3XrzqhwB
VAW6wVd9I0xVlYfwqUHDgEOPnX4hoNu7CO9dlGhS+kGwBudeR7O7Rz4LPfhnKOWuaZdPdBRa9urh
W6BKdMY9+Wl6nWKMhuvSJayb0SRk3f5bBfzD60iD4kJZMSVxiYYOsvm/9BmFI4qym1pCiqT/MPdn
69nSBr0q29x32/k4HOSdjNHKag595o1j3btsahBPgKL14TLO7YIwHJrl8rCqsha9wrV4SG0682WB
MgR+/TCVWpeZEZ0ORJeC4r5l6kkAuIv2DW+0VaRwe3pFrZzQ6eey5TW4vtDhGtOdXvScukxkMEBF
NtRbnLs2LfCKyBla0iNYl5TZIaRZG8Hebt3XEyX3f3XIZfgWLWreHvYexJOiP6WOge+r67v9T5+o
Azkk2VPYgaLj4q562d2qjMA4A5Dal/a5YwQHtq/lE5sns0jzwmsl5JZl1eYu5Gk0uj37DLzUVkD0
BJluHHbt0/6jdgttXFdiYAAIiLoK28V98EseKDzgLQr2xgFaZgPZCl6lRGovOMK7i7pPzlf/R42L
oRlLj5MvlDGu9eUHxRjcXpO6eU/lVhaf/bY78ZEg48Qc8kfvdNlQX1bQRMGDyEm6YAG0a2JLKknc
Zb5G466NuojlvWeynENOBS2+O18WfJCNI3pMRuWnY94I526wFuLRy+Dh1MBbkOlX9A2qYl2t7RrS
IyoDZcmIgc+skoLyj4sgW5JAXTrahXiypLIiygyLOQz1gYj/33yA1WJxX9x1nBQAuIlvLgjoaOMu
9HLTZnTcwi1JAe2ITid1d0EDhkS1Jjs67hk7/gnRTYKeeurrUuz6VaqzHohgf3g0Y9HvCQimE//y
CXpPy3DxnzMjHx6Lo8dAQMfQ+MzaqkX4gJMZwBa3HhnMkZCBWcUwpdwDkPHilwUnJ6V9JtkAjzqZ
RRMf/QWaJoz5T0+ivvQXBzuVgamPtiPUpneru1/Y1TC3WtcXWA/bY83v82PhfxgkfZXQOJh8Krx8
QpZSxwKEB2UqlB84demToShzyJn3ZM4iGtT1ai3+CT/rLs63vz6iSFeXwrfGy04PS7N7YU7/8Jrc
YlCsPClOxuTgSsZXlxz/1k4V47bvQyGBjy34wt9hHsV1TCsoRhBLcqL7SJB7JYt6R8kGCYX3xrdO
B0jAR6PAiCNU2N37TYU1qZ1UtO+bCmBPbKR2ga76VIPlBdVEANUgcQpqpC7jqFSsCn9qS+ks6YAO
95ND/ruxwvbiD12GRmmdNNuejsCFmzQUUWCCPV0rYoXOZ93/hP+u/x2eLzeRvXs9KDfnUVgNgHVS
UryIrfFhK4Lk+yBiEnAQNX8IaPynWR7YXOyL1KT1ot9JyX0oosDp1DwxG4q1K3czlXCtbk+dopow
nvdXB61H0L0VmG92NX5yfYjxKJvK01zC6CfAKUV//ygoU0fr1OfBTrdLkBXHFRCPOCD/keiJ8NR7
UUKD8HbmlyK1Ik6qi0fquTW/yXLplU6oCrbkSMsHPgafK32iQbM+Ah9q+Pm2WBbATJw9Hl3lD8EE
lcTzFYKVPADEr58OnbeiCMJ1HLFW+LZE1eiCDBKqjlDfLCTyQSPNXxANijmFgCGZ/ijAYM9CMeiv
TE4/AR7fPUrfwPffuMDliLIUaxUIvQ311O8bqzLqq/twydpTvJls58FO3184xxczNYN5RNMTPAiX
Dg4UuDtbKFPnCDd+4P+W7onmD6L354+OQ90VZsHf/IiHOKDOfpkY7ujnTIWAGamTk61TIxvNowVl
jEoQ7kitZYa+1LFCL7gdBxOL3sY8dKFlk3bEWHbdflSMdbLYbd1hqGBRbcI2n9i/28khSDNsUjl9
XhA9aKA5MK4I04NnBGFaSTVpt7W6FcVjfa6CL1hMQTFUIyeqwwzuT2Lg+J1vEifpBEIuGBGcPqiJ
Ct2TN1SzK+Kjsbn/fK/d6EwFt9I44CjauJjwoKBCe5cMCY5suLfswRJ8qiu4lI2ws7baC5JmzOW8
755c+U25hO7AzIwfp6SuMrQyM5ouJX/otsq6df1+cX/YC+/szkJ+mbAGDkXbjjpJasUXzPA5YnXy
7RO4TtURnHUkU+KOcOWo6xKJawmBEz6oLcUMWvDEgM6MOpKHSIxK6lDZOOXFYzdaC0tPoCOVtBfJ
uomGSzQgmJ+RHEvjckky6S7u0ozVuXFeb0k/ORjF7uMh1lSuucQGwF7MQXjGqsJEvKYKMNckXOjk
Y0GxYbJtnOHi2lL7qdicCWbetpi+RY/VH3UEU1dvMeoLARC7lw4E9V0w85G2YzLpQI7N9l/jp3Yu
KHhQRNEjNG66rapW9LJOru08r9UAaoZgh/AefRGgtWRN7rCsEpcNxdBJBrq6Fem0gYffNrjcVEP8
kVVL3rszyUJ49OK4lXlkjExfRqv39PJN9bmM/gbeipc0PPaVaxOWON2CbhG15dp2qMX/c1fp+ZUf
4sldu+EyquezsS+mThWJ3E1R0Sn7Tz26yzXX7JfxwBF+oNKocPHxsMQH+CzeyOvjrXsVjt4XvmRM
niQsFjZwz/DWQfwjhkqvcaMH8yK079ke7Y/yd81uXOhrZAu/hUWVkJB3qV0abRrvmj/Tln2Z4bkm
7lzWlZHEbhNg/BM45mmhsaUCr9rOVrdnE8JSdyQ8cAhge7ixwpZtTmKh/B0Q7yHbwyMDratNQAPp
YZHJ74gCDY25y8rhR9cx9v59Dd4qhsm0EkYco17v9Dlind79f8oKImvdwEpoQa6WflvJe9jT4bbX
HJTv/Ojqr8wV5Svxkl/OZ5eW586CY4WLTeMIZRs594pnwVa4SNAJqkWV+F7QEmg3xxg1V+YlPM7/
+kbg2NpfoG2PuOKWYXwIp5+SsiaBsQvhvIBockYL4tu6Vg2x7407u9a9HWmJwjleacpvDsLbsDV5
/ZJ/HSt4vxj6s3Kp4+GSAtRl95dXEalQ1xxaDUjVNa9UcO5xW4FB64mHsK8wfLkEQ8feK0pSM9+S
3xyIoaJ/131AcMJu1cXqym7mfUFheBFWipaqM9hOz1f02ovZCJRZNQLfx5b5KfG1HD4gzi1jCDOy
8c/jPl9O89RFC1T8UJV/elCvvUu/xelEh0WWUNTxoK1w39o3a5jSYWGGtUC+hBUtHvDvJo6BJDI2
Gm7PiiKyKGHdKjQLEcYZQGoulz1lvibYg36awyqeV1NoQ6imfpnhXo3XFLYaL1GxOSqHSvhthypE
Q/NtWsUNcc/czQ+YWfMonDjdUsgFOl9u6AaaAI7evn/IpixcRQoetK8yU0T+EAP0Ndtuy1fWbZrv
1OnUUoBsaaPDi1rEytdksX5OZERONDr/wQfsqUbNwl5cCUPeWUZx0bwjOB6VyBaRb5zPe7usJxKV
meIhFmvZJbCNAVMHhrg/xegcZ/0bX0k4UuAExXG7eE29qdJzuguWsBUlMMf4ky+F8ibZqlFs5Jfs
VqoFV+Hp+4jPbqlnoYA10mtKE5s4A14rFTMkyGlRB7IkNvz+Oyjm90IHKmwsPn+rG43cD0O7oOhp
8GfkGwtGvtayBPTLQE7WJOvbWmvp0PuXwx+x1mvT8EFlmAwBXpcrN2wAB6AdOkoZUWfH011JPNb9
oLCQKMSjh56/VLdhpgWbjinB1VxCB+EdtGEaJTI3iy5Coj1hyZhs6OVtdr9dSPFki3RnZIzEBSPD
eNxI7qEQUQRXPZXsZHrWz+htJeaBGNSJfHAFUgmKhdQa5zeVwGzVbdBtyNVXqv8DUpJbtzeiEkf7
CNV7SsX8kqhetp56X829vuKqAmN0fhWoBFU57KWFOgLm8tHT7+hqAMEAg2B8GoB8UabQHzS5zgtx
b7wFYISOpLYBWLz2wiKFytuBnLBvmZzZ/T0iusz1kMPjn3WfMyY20L8VLoA0YujLw8/yfmHSf00d
9HQd2QOucM6sDvKaW5okt3Q7wx/At5ZZIg0m9ykjUxDhESNudqpGSQjdZpskQxjvLJv0wcthdKGr
LhLw17tSy0XJJulJawOVD6Z80ew2aprhHvzRVEq1HDbacHTKXYapIl2Q9u+6PcU039GCMb9ruVvv
0BXimlO1+OV3VYhbdyFz2NUs2/Ta/qioOaWxg4DS6j/DTJd6w8dMnCwNurpUTzjbdFfNDmnrhNtS
wqRgCXOhZIis/4O7fvXZSlmhNrTrcLqG2Fkr/9T/Y7uaCSds786C7tmDQw/Ru/99B3OTOMK6QzQn
i6qLcBEWN5/IzECJOBtXppc6biNq73dHkiJEohG6/OFi9bJdN13tOL9FDQrHdynTAjkeZxcLcPQ2
Nm28cJ74dJp1DGzpxNi7TVQIFKuJrbAQJ5rAteZq5McbIUJty1njrVt7wp+dsmXmm4Q+DkNQI8Gx
Hk1UF8UvUH2Z2VgBx0AZlXdrTRtMFHjjLiTCAHlnNmrEPVSdJrbSr3E1gl2IBN270AfKR96G6pM1
3+0FhDtPg2KwC3R/35v6+8tw7GrRtJ3prhi6M7ILe392+csphHZpwptNhbBkPdHVrsQK6bwwLDG1
Dlt+BRQMw3ql09O0wOwIwKfq3VSE24SQcZmsiw36Px8fvhlu7zWgi9vL6ovcfKF8u9Y6RS7PBaYK
+yQaEhzIay7hKO7q/lsJSnpCdVNLuJWEtMcVs+Pvfp4xaGuiKq3ZINxTtXmgJL9PeEIgBFcuO5BH
/oePDflfNizwa9WSeeL4SkzaG/DqfXmKoDOfapHmLh7J8U5y5O+bBDnN3nTFE35ygsTWhLDmGXr9
zIbqdeCMKA8vt/why3ACiRI7hVdtEe4l49ooQu6S4ob38PgnaR0QZQQGsW1DYCUHtgJI9AL/P8pU
WTE1WUs7sDCygbhCjRMer/ilapi56P81O3xeWR/Lg9PDAky8Uagwy7R4pE4fxIu3PLyGmA+INvwa
Jv2jXGduow4u/ca27JMN+e6m7Yn0Z6dvFDTmVQdNTdoc/AYihks4IhA1oEuUkwkBC+Lz/636XMpY
2PK4B6P/jJxpCzJdyt5BHxH1eHHwxgBvQINOfu0JUyBUm5UGZ5kEoFpK85dCQgTRXVEpUoHVy3QO
3mlW7EGPWkbwgXT5oSiQumPwwe1jK3x+VHnhb72uHRiEUz4XXTJ1jYOozEeQqVDynxW6tVOA3y4u
zQLC3XCUPCDWy8kTZPWDhqopQZgV06402xrEhGl8jQ6I/20lz3qCjudIu24xIXQoMBdELBTjJ2eW
HjhwkfF0VIoFwilRyOZBaHQu4ad+W4FZbruRqaQrXbpIMEaUehHWEkCiWyCha7zut1ORKwKtV2EY
w0YFtQ/uSmtpWwQDDtbXToQAj0+6E35HRDc70ThL9CW9spoLNhVSGNISZ6j+eL4u7aSYVMX+wxyj
wa/CkOIK2Vmi+WrovqnOD7ZqS+o8B6v/bUpEcBUNMezL0LOZ9uTzEyULoorWPExp1jCyclRCHdbw
okz8eHabFpKdWytF/K8BG/mCgML4si4KBcp4noNY6dMZV4CliwZK+GkYnwkyJoACRu+3B5pqdxj+
JSt/rEfCRNdG5DUVXJGfND8p8l2vWqSxiSsQnxNr+NN+NMBHxlWexNlpc3bejWS8Q379QYjgl8Ze
GN/EHSwlW3eu5PoyHjqqER1hmqDzYAgqCgaHJX3bsxRr1/W/bpEgnfDgjtsK1T/rcYIRCiubPyI9
FogFpaO1W4VD7UbtCB30HIZP6e9Sf2Yv3lWbYTMDci438b196hm+z+hLpJ73hYudXbXDK3HWLVxA
EyNamkrnMh13V976iOufBGo7iHS3+RKQmEboBnXrFDuRpj0tID7YfqRgXA89YxjiZc/DSWDKyjsi
/LDfRXV6eISFOYupWVh0h+zfdmxFz+RTpZZwBnzOejHUViNWlEly1eZyDjVLhrJTVM2nWtyMm14u
q4OkmC3Kq9xnHOXeiJZ77Q+zur1lGdDiBi+1fQqYpb81m4zKVaa2fzc0NxsFG8vuT/rDtJsHs+EY
qYFYHE5Rdg0GrTflsAcb2xIaNm4DgvhGaA1t84ALGhnFW8zoZA9MD2tX3YI7Je/GpYp9yjfhD/41
1tuOvp6r4vxWJAvk7VnBK2Fay4m2liuZHGuZidvUmkK8VsM6bDXQTC7PNkQyTWYySbgRi4sUFkM2
tCkIC4AdGCJNwOMjhQoZhwQykSB5PkXZ93vLzil4YzI8Ttn6/V+TKNMqcg+jUd5hP640aUgH+QQp
v/JNUlVpYrkJkNYNTypL85Slhr6PZPvndhervq5He/tFFu4CSwWiPoQToJiekrOQKHx2ixEWadu0
jQodoQ38tKe5RzDXT7K1oqqR2K4dqFli0QUgqJwjBzXbD8OK3Ra04bkkWz41jrd0GTTopNJsA1WN
RhhzSFX4ioayvkofFZjeScaIzI87aUjpshnhHBVmJWeAvTsK4Dk6VKm6yqXxE3Epmdn3smjuCkHG
zZsTIV0Wf0Ra3kXHzGsepv6b/iIhaTG2nur+DQFxD+qsDpXKh6nQRBy9tmJIZHpkeacQ6EPCLcka
7LnK7YFuxxkvBOCCcH2ffhoN1IsNTMRwh7YQGC5D7BhK4otk3YVP/xmi7skhefPoMkHzheFAimGT
/Bud0WyYiBXHVpkgG/C5xu428ozw5CfEmMTa7WZhJe54jG08Ypno0vHUzFNxIU6MbtfL09zFdgXj
z/LMw8Y7oDC3IfPnniKUcM2g5BG+aaCSsbO69sSykLfjio/e2pPSJZihEb73mosUqM8D3zAVmzh4
jeNBikuBHwTuYYGM2th7INHqPMCs42vsviKjjWgizMYLw/uYxtqt4lp6sLZNZbvgbcvJQ4edA+Tt
Jjw7UHvvt3r+q+rwdw1nfp8dhJfuWU1M3iixoKCGXtS7Z4b7K7Fiv9arkMqusVn2qekU2M91LXSm
SB/0EnjdO2j3mUT730PWsetFP0J9ZB9EKwtB4ZaukFz2v+ZYlV+ehqB/kYlGzGhfQofi9/ysDymt
AhzZVvhUPwXPdMZZxPULA5zAz8SIWLWfp34HFr3YRYGWr/ZX4TC7c8Tj8xRN7n9wFrAptPWiONB2
qkHFkOVHM4qs2wHgmklObQsr4NoU1IbXf/9djfNTdlYqquqAyWcoi6XzkD9A7GkGlFaLr+LQkCud
MamL9Wt1bd0zRRUXsroseLgTI9OC8K/ALQV2KfwYsX9dZ41G8JjGu+hoqBSRLfbSypqk04b4CKL+
osvwEVlkti8U4Zio8edcQueWu3R+YbAmVaOqy9DRMoZ2YCJQSZRCH1541eNoW4o9l7iUxKl4WTGx
uop+LfrBW5IsSXQL5z2knJhiDODFOEEK/DRUG2Lpf2gNczptil+hc10qHDPhHvmo9M9nn70+SZfu
pWp48nXncVqMrcQVz73eXOAO3sMExqFZfnQknnfw81fIFJ0+u6w+FHYTsy8wEpYp/VMp7VWg9PlG
JSTwjXSBOV81x5eFO1WNncGndfV0mmszZYvLbeiFUv9dB0vwPmROB0JxE4EnnvkmIySkbRZFBFf7
ZBSpnExlSQ5Fe51zYgLS0+yD8ilzfPnugamcgZ9IDIn1PTAiLeEHYORXZnhUR/ULQfKW3950i4tk
vZcI0d5CaxG489T+te1pA8Kft3FbL0o/9JII+SSXz6MfqGHvD8IhYzbLaKkMmeulEUJ+Y3sKBg9k
8YMNupYk8oFrV2rbr89jORY50tm6VCrq2DtRJVtpWwRZSUYl+ZDwssplNVwv+nhZNQPjnBMpqQDM
xI04wZTU6dkJjxJOdDck3xOJ7xIxIxhX0y3oIDlykDnBeR7//Py8j7FtZ1imfc8c3mfwsjVJEKvi
ftv9iITehTYAKow0QZInw6d5NpDeJPAfOa7fJCFM2uPFleDKRQ9pPOW1BVydD6QA4LL/7S3A2tQC
OlUOMD0AuaI1GRljOCdOW4gZKVPHNESzaN+xWjL9sqgZfsoJ8LGg7IV90QLsW0iUDISIGs718Rab
baXE14N0QnPkZNQy6R2m5chAiOUy2AjzQgwbCmEWkh1Puu8nB2XQVlMBPQcwcBV+62tJ2I+366Y2
fKCFQY1KQq8V8p/t0Ey8e6q2louoGyS5HHzw89NQIl2nL+WLDp7d15AGI2CuYwslck63ZygOdQwR
DhmpHHo3bqNWGyI0xTWhR9EuW/c2Y6AJBk+qn46Oc804HNxco50Pw0AlJArl+7Sfvt6SbG3JBqdD
X1qwN6G7KsQ9g6bjYMH0srV0NNXRzdxMUEWaPCKgJ/N55yiI9oCpFC0OzdG1W3mMDgdRH8amwCcn
L1D0IIIedDp6EuZZYTFJdq+SlTVSgpLvvbnVxBB1+FaoPJNQKGUA9Qw1bT2LXp/VWr6auwmyxIK0
qjezi0hqxsRQJ+xjrD1eOq7SQWNdzWXzkzKXY2l/85hpL+Jayg0mAnbnRrlu/ThtIzcHG2ot2SfP
KiLd/vvAqNORwQYok6U45eQxMaAEs4wSkTu/8UOhnNyv5TIMmqx0GfXLoDMzJVIovnGU/UHptNUv
jxBidkSjXF8A1ehvDuxXYS66uS80/FhVuDkY8xe+RirLB7iKbrkzSecEBX0AYAyMk/E4YEri5QXH
KtYGq96pUJvff2zd9tdZzASUbbnju/uipD1CMDiMUoO4E4dLM3xbGQq1CsbnxmmNOPjeKfJtNGkP
eyc5UjWVqkovSmEwRHDfQCxl8SwdOjQSQMBL6jURmJkLWiPUqyPKt3DLBZlCymq69ppJ8jr5/K/i
kQ/wMPn/3NRpi7NXvdPxLErD0hvbl4TMcNfISnmP66Dwm9klAMmFxz30hJU52sJlOB7nGWDI9KwJ
WQgo5NUi4WP4WGRdtvfe1szRSY+QpGHd55wZu1iV+aj0zYuhBEGfyvtcmjCN0KGQSQ3VGTMXypwL
fpVDeYvNQJtK/zmQ02pPzPESeOSZAP+dPCVx/6AcrYzKYlH/1ZZhSwgTjbb0q/8MANafCgyjjbO8
Tco/uXMZ8Jipev/iDV7XBJMokdkQv/PoXBdBi5wgjYbznquhOSpVa9/AoHg+UEP8abNEIvZZo676
riS1b+RcuNw1LlvZBVR3gu++Ff+u3JpoKbseJ9nlai1Vo4N5k0F9oltdWXrSP6uucmSuMAY8A6LS
GPBRrfv53VwA0hgyouBBVxSFJBTPsoDQYjpiNuCVUauSghRtTazpenDiYQ6YD2EkG5WUzSZsmmhY
u1WYerSZ8+lH7aN1p3NiWqL7VxNHhIcsIEKpDKXGho4WIE308WwXCuKeVFqY5L9DsEyYm//1E6R9
nfF3hOepAnei/imfGwyP4fOPDz8zWG0Ck9a5b5zI/Dd3tOsnHkbTAzyy1mnByqJg+Pya0n30xco1
2C1BNlF32tNDICflLBAh2esPpgtuhNlUrWWHczBe36S+C4/RDAv86wDesMnKGiEclxBamr602hJu
FE6B7Aq69yQMYv2yjdDdHXfGMHJmynwkkvZLYc+xQwey9POLoZW/kyZrU4KmTA7HKmMGp1ZbiQe4
iS7hwBgS3l+44aX0/1WXc8IW1hD/AMHkvBTJhKajEhWuXXjK/R36Rf6eoiegrVXmAgmUdTPZqWlZ
bsq3MQQSyxqMx/92dWMESDByKCJ5mBQyk+uzSRCz6gFVMbXa3ZdqJGJrsaOhoQFMiXv0lksiw3Qb
0YEWlbMg7Xz/XraUa3/tOZNYZTuBEKU9fxZwR6RsZFQ2nC9G4r6DLbMhEc2/hBYLi+fvGaLt6crW
nWaEKXqdOq3CZADV2gjTlpZlHrpjEECVVDzFpOcDgJIv3wRpndOBWVkEdOBz/35e/pLsYWBzqi1q
f4/bh3ptrWRXEWTVtW1ChDhXMrLxbMAMEeW4mccwOQ6xYPPRcOCymX1Tt3zN2/sAXy7GLbP8viNz
gzDZXUGM67SBXLAfnLlBOIgFUq9ymYYCWvwBXCYZbTAO5EVQWDRdh+cPXdkpcslx4V8tbnJEJch+
z+PLU7RiCZ4NKubakRdExCn4Lq4EbUWzpd7MeFyQj29uB/Tvw8zptPs8v7pzbtOI7M3hWKdTZSyv
7SdbY3aJgbUwjbxI1JTysBvl1pjn6hQjsYY8Gix22w8wjXZ5AGn+9TjZUUzNyDw5hFkhCwT1wzfL
IIwSfj9uX+yWAzSVjd/HrGyERaLUFV9iZdZpUEf9d8kVkdgqVAAAylmAxNXtapMRsARrvrdHahsB
UsKMfuMDw8DoXyIT+eblzAIfl9p/ZwFwgOAlHoWEouYYWOeKUWGcvSuitcwhcphoe5jPKXz+JjB+
rqC5cwyv+3em7ExL4fL2NCH8sWx8gUvhNbXIMzheAidNiXNhFPFmR42/9r2zouvlbAEc7vtLZVea
qHZfS1AP5Led1vmnj+wje9ZDswjwdn8/UBwE20Yfvy6UsZeSLaOsyhAa3w0tfKxH80KXJmOGh8jl
nQfRhpikql/NfIRfl+M/suFlF5W74rM+HKa/LBKs2aVXptwMRiMDHdz+8+i4yD5rlLmKflR7mnTm
L9zyLSpQdymgitpeOMW7XfesWTyMO0gVj8UfB6em1KRdNiOgcJUx6BH/W25b3RsnQXpb+RK1zHpR
udIwH4kSAwndjJ4m8fq6E91hxk6nlez1DJHzC8nyYpnYImuPDhmaA4/p6hbxKvHdkGO3pnTcm4pn
vvxdXsR9Pg2GZJu+OTsEwUklWTKonkptt8dkB3fMmaK9ksaEWRD/CULCNOqQ/j0qPvqlqyhmAb3a
XD8zCwvJlP23jKLKNzmluNlLdWwmtqxXI2hv5F19CPL6l6Z3TZyic2qtdNZ9t/dXW4ZafdyuvRBQ
kXzA97flpHeUaRTCegICHcciw0twi53pP07fTINK89GBJZUHWjxAFzYPVQV1FJcXewzmQCGjWFB7
8qv+Msu8/b3Vpef/IWgOnJgJZFjXlEA6kXisW/dHBV13bIxMt8z6VLKdgiPND46JblmOUDXdwHgy
//zKEwW1kEsgTy0uIwLchgyo+iZ9aye0gEGJaVZzLjSuow45Re30Rh01MpTTib63BH6A87yErCg3
QCniHtoAHj1FVvx3OAZdGzJzpUNH9gsRLIBmdVCremhew5wF28X5/sKCdkfQzEFLLVnnsvQjiU4H
AQO2EQFuNZDt6Hnx4qlI9HiWYHVTzrFvxf+rLpNmfCvCzVoQucsogHZplpaIVlhavPQo55SCCDoR
gHeCF3soo22B0heUFMx+T6hq4lwKWKhL2YEZ3bx4xOb6uQcsTHZ7iRxmu7uWiSzLpe5OMG2Ahc9C
zngZ440fUwQCPAlJMny7w5rAr5K5AQlWI1gA2xUlvzpUTL8pLnkz7JaRAG3AmaxtDK8muz1e8tDK
RNF7485dLW1uVhyMKrww2ugYZVZOX9wKYyXIo93S0aoEBfoJGJQXStvi4ePec2Hhi/rLJowCtwxu
S1uqNHziy55mns0vMpZRzEgCiV8vcsmzE6A7953noJV4tnaovHUCS4gw1N0hNWhrpLotUx9GfwRc
R4M/Usagtl+hvr7TKGQ7JouAd35seuabNztY+l2ES6khltqwqxe4Em/CC1q+xplLRw6WJWTjmPyn
/MS8VctjBcBXrt+z3yphywbTXapOBXGa3dKo046bzatrsZJaO1Mlm0b0TM7wQVuoCgVa5zg5piYI
HvQwRfiftQZXawa0nYoet0aw2iwFp2mMzureFSK0lxX29p46pwWJC+brmFC0B4w9VW0zezWCx2zv
TpTdBAg7I8FG+debjkaroNRjC7p489EN50nwbBOBAk8royIfsstgb5/7H7Jxn2vmTGP/Yp3ln+QY
y+0aTrHZ1gh/kd/P6zpWe5vis63+lZOc+dJudaA8XJXzP/dMMX4xzQo52/5sHhb8bFZdtRhDlvQI
Uhods0ICvpVGxmwH5NmTLh9IOKgi8ZItWp59rVKxW1flDDukL1ulxYGk8JJS+0nR5jE1IR7no/vr
m5Fk34R2W3N9f933AQNO35vFCfXTt3jgJEFpYaqzf/TVzyq/RkzfI7I3Im/V44e79wMihWvFFxTa
tIFImHmRyuEswPFauOBhz6BKCPwSN/tzhGYTP0F17g3Fie5uio5Mu1zCDEqCBhhxSq7didgxvyfF
vs2LOzx5Y+y4qOWVjhBRnYJLWuXuibx827hL7NgHkJRy8a5Yy6aJi7YqNYeC3ur7B/SznMdacy19
snWGcoxxrTel4Tt6D8bwqvEseYCN5K3EPkFixXHoBVHELs/FXGOIQsSQVGB0PffO9yp0YO3dHr9d
48GMjp9yeQ2qdzoFos1DIXWmkI+J66g43PiSUrXb7Mdrp97DznTeJ77PxPI6g0aTMJoJDA5DIz9r
qZBPzcf4s6/cFpLWtnKPZ24KDDIJG1OwamebZ41+OYsYq36L5zTw04YUoYKOhGzghv65mu4blFe4
cHJO9YCEmzTXfmK+HMvgJm6755Nj5NGTMyqmLHAtMk6UxY9eqM1BoJveckslxJdSLDWmCvof9muZ
vSrR65pOzW1xpjKTDMjrAvZvsdWKXyvGjD4QauIOSKs2SQfejUYx3/PG+EgrzsRnWGIPw2fafKdq
8Rabq5TPDfDKFDk6MhYQL3D2r3keY8m5F5YW3sK24/2BOJaX8KzMLWQLTKAsXp4UCMlSU9n2ve2v
oFzNA/cFxOlmjMczXUXpspaGROXGSRWAf5YGoNydNGohj29JvuOS8jbBOO/wn0Taq+OdRfagHvvZ
ESHVeKk2/ssMb4WI3YC0ebwCM8LW90cBSrZPHyFdOMkpQmEGgZN/Lw8N1H9sr8LQUDFeYh+J8Rp0
dX/2yZcgqnhWyoCb77lycApChfof47PsDRzOw27liD8/pAxUeC4ZGiqfvNSO6/3Ga45DO9AgXmNM
xFyzHGN2V3ExDJJlk2I4zkc66SC3VxogWzRKe+nrdNhkbwBtfcma5RQy8hWtcgBQyHWXdUqB7rU/
udrfIC5E3WeVgbMcCwW4+TpIzzZXQCyacG1EKBY7ehxlGb3mcQqR8wFH4HZ2LppMxztDmDI3hNXy
pAUJ/K7EL/EBhy7TX+nDhmeeCmTgy59hijm/UOvAHlJq9n0Qsrk+QgGZ0zxfDInfswZ3NOzOXsv8
yTFjgYxp5oQtOoWSEPvefQ46S5KnBuK0yPASdQ63kuAKR2XdCopcBeoVQm0s9o6BMn2nULylfgZC
X+i/bc4YbZTPxbzbgqPERK/ZYb0ov7Tt89HJfcGueVvQqHb4TtrypnCUxAPGjctqRvW4bNAx6f/H
BhJnFCkUE6KwH+qr79resLePuoBL1SSztf/S8cnPdlhjn8gmvobMj10SXN34umsfH2tw+2HJiDgw
evNuORrcAKMIv5wUG0aPF02Ifhqu7EAI5EgiJYnroFQMI3/jcA+IPTNOPrvTox0EzL69SgzlD0Zk
D71IrIBGgZPnkRs5HFfPx91sB3DzTDSO3N8GanV7arh9PvfrX4q7A5dEXeL6tKntPirYfd9zi2DF
fYGu2sJr005SHydJL3KqJb+hZ0UxbzQTtWZ3caKQvOxf82yj4eL5yOQTks9B5YDoOrGy9ZlUkvCx
TR57CiC9IEj7oNQ0kr+w1ayHC+Ih3pMybOpJm9fl41bCiGbsrUYP5uvP16aHwxbpxGxEtr+vHwDz
AqCEMwMOhf2mNCbquKm8nLHFyM6rR1Gdr/LHm7kfA0LLeHVMLToTh9ttBm3Cf7LzjaJbrHIrUYq4
S6s4J8PSlzAs8/YDjKWwCoPjc4Y5oQNN8NomqxTAANZx/4hpBuUwCa5jEkUjSN2NmF/VffZVHop0
bLYYMMGpQ4jehtlyu2Mt+w7FvRPiFYaqcLEKY9OcFEmMW6p2GYg4c5YxZ/eyJyuubhblQSGiLskw
2pVuPrpf5DqZiTLZFYwDvjlFFvdLrio0tBfKPbIHknZ1GOdxdQNwXp1KJRSkjRY4DmrnnBNLz5Ie
jBxMo/L1cwbsOWi070s9cbXIoiK6ZB+9i3IxGmak2+pqT2Cc/qbEaHYvVCruDyJATxDd3ckZFb5U
eEJu4q1odfYGhffxI6WjbPBpEgfe01JXxwZW0+LCQRhqgIoFsMSFzkAw9zaWqN/jJLe+46f/DC2I
i272aAiwaY7CcC6aOvFRSwdHb1GxnC+4qe6ui/rEhc0dRR2IAo643hqnEpq1mLZWLVcA48h4L8Zi
hus/rQfm0BZTQsnZBMFSmvylsr5piWRCd5lfsWpLHIoEYCF8IS8JUBa6F6IJFQcr2vMIQkHUoyhB
cbeckDdq5Vf1f3j8RvCHwglDt8ay6zM2dm+Et5/2CB6jxS+fKtFTniVCJ/oCxw9gShdK8Cyca/tw
vInydTt3Htc52VdD321ixFcrBirMJa46oeoV0QgPPRNZS98JwoS5H6BsOkphIBMTwZml4G9L/Kdv
NhWpF0b7axFQ3dwqzPItLMRVuMTT0LZwZaRzOz5kvcYMbVFp2EztpfE7p7z0vtnAhVWbW9luInNa
TE1PsRD6vZd9Z7bjwKUHgI/+U0mQUi1QstYc0hYe/YdOL5kQGGH7Ngi+VygAP7IH6wPrG5axYKe2
uhaxQIi8Npq811VzAGnc3OB8KUUq8AD2b/ZEboE1AcgYHJ0QTQMS9CQLbrxeQXk8JvGXQDhpqAso
YDWdd+JGbLSWdVOTWyBHUj37uKQdSCFUF/sb1hV0q0+XzK44Cy0wkAtbrT7WFZu3cdqLzDKIsYUS
fxRUAsx1Vf2PFAfeiKPVSXVNXMDpSwwL6EuV/0Kd95CMmFIkoOeh7fTxkN0SXcAShhpATnB6OKHY
JgzwtDXwUscNWjs9v29YWEABpOif99BxGYpYQFqzk1h7jUVLChJIfJNBbz3aQhRgpU0X17Pyqpys
kfsVFEf5P6pnJJRqFsHmQ0yt8mS0xVc7E86XVrvMuNK0vTX1ZmRNe2Zgy0cPhusD+pCFqUG0tYWD
BPiXhUbtMyEfTPzejz0O9vJJ5GxKV4fPow6n6HQpkKad6oDMM3pUmeuwxDhVmmGCXdnK6CMMNPkp
hQvnMKVl7DsbsDCM/eXBx5FLgDLvu97ijm1D4UaOC4aaLCq3l9eBdrQRJEpgs5GFWDHiN0UrSLlX
yuShH0Dylzr06RjsRr5ueQLqr0QvaiOvMScZp9egAsZz1beXDm8MdFix4C7S29WIJYW2JcXrsLmk
xxAIycDqeIYfan8/boeWmX0Qo8e5H2UPcjMpflcPERhuFhVq8rp772gipn/Mrb0L/sdhwAgeikdQ
VmSouWP7yFwnxcture28MqNvNC1SDPjkyHaJrfOh7nS+URQh2Zd9eK8xrt0yEInF3b79kYLwxh98
DlQKNTsd3u0oHAuzx/rcby40wxhZJkjQx37He/YEAZ/FIr6gbaTEFyugxabQcJoS2D+AcjwPJRK3
AIWpJKGPz4u8JW5s6PmlzJocE/cyoHChhbn/46L2JGxUBFlQoY2tmIgJH52dGzmhFtm9pm1PSZMM
aUcnEiFQRLZLQDt6Pmgc5w7cr8oiuHX6BGCC3aqNwrEQ9oBrdHAudEphPr2Vy/imfxfg1KRBMbCJ
rxLmQpwJ/tarBSE4/wkxDOE21iPjE9E0kXde2dZvmKeyQJPcxutIyPtBvWrL56dZ4C/PrXsNer/A
HffdT+kMZerFWfsBf/6letsnXOcW3lCjHa7h8J9pWSzD1r3/H/o85BnVQGYD1WIua/vMREKcmdH/
xvUjxovpJ1S6EU5ZYCw4ZrOmwXplQK2k1qaVYP8zRd52CnvNZj7hBJzhOGroky4MhQRri6YyEHEw
6w2DtuwmuWt/OuoKEozPD2epk1kgp8rDsu8+P0atC2uCAOstEyTwAlG0AP8KCLNBTMbgOPaeXMr+
WMnkQ0+R69kCl/UYUxkEaL7/ccJFKa7rS3SyXpBnfVf71tXdMTyOzWYw6FRzjwfcXGemTacnxkAq
XSEGWdZysWMBjn1OokUZzIoaLPlzxNYAx16jJxQ08fRSWdgPGkxtP3xc9lF/9L9ZYDqgGjUFHAzf
Qbs4X2903SE2Mq8xIoIG0EQHTan79Y8dZGMzlQF/j4eOZJo2hyxQM2AlYdlXfx8jw8XSpXbAad9k
Z6pY1SuihxpRjAFMLl6EjqhCYr7rKFJtwnRvGOQW3kEZIiMfEFxTsHUSB0mougwwqlL+pOwR97hD
88cuaX68X0WKPApAAxuvAmCzsjQrvHZJrJ6qjLpPXKO6NrxwmPoUvWvoQFyY9TXIlqQxW/JwFIuw
I5hTzo7aleLBrHGKTB8KqmQsCLOdScvaYMySRJjBSnBpv1PgvznFKh635Xf6W3Ua+46Wtt5SZ1dI
hH8LrKjCttwrOxoW3bmaAf8LFs/xw6/izV/+ZB4cfrCGe/ePM0vga2rJiIU77DD3tFYmS8Pa4JkP
4V4FaRmKd+LMUpjq3PV6d7yGuDmiLyytOBaizQfiqnOSVLKBKg0RZ/eb2+wbBM6YKtCyOJfPgCVn
6q9IDNGeahyK8ttDGKtx05tjLeqR9BgKc0sozA8azOB4Pkel17Bj2ptMwYfDoV6NTWS7l1ZLSWV4
29YdFqfcVqs8C+LUuvypTadyTL5xQX2kY3QEuwQUMXMRX5N7ptvB3yjllqMinA0FTk7O8tWTFMcl
0if+eONQRN4tWxk2q0DkDKwxDhWPTmdRx0DVj5S717UZW+aiC4Zv9utG2L/fQEQq1yYRaJILdO3t
of4HKvmolAWyLLqxW1gI0Cjrkhtht0/e/b027H7GodTF8Kxh8K9ZXYUZTkBDmiXNnlkRWjsxmOT6
dCwpfjqD/jiytvFqhXQBuncdBplOfBM8ZIhnjP5W08h/QPkQkNRiAidOMFbyUFXZTSzKbZrarscO
rx0YNWUVFL59A/1VxJtM5np+c2IYG8//NeE5tvwsb40otlQvvYNFeUPlPRcIzXfnzVP2m6f4As3g
Gz3pQUYLvGcn6Hu+7I8SiDInJiefcE8S1sgkd8IkwGf8AbMT61bQWAapMiPVvGwmrJanKx6OIP/d
RDKTpBfOu+PLICHvsgPejbf/N/YeyqKLdKHKcUD+oXf+rr0iYtS7+ksgiaWIhCewFdfq6kKTinIr
AdkiuhK6TudLIx0rLypq3OT/Hl6i5WI2P3asKzJQYEb9A/az9OOBYA+ZV3NLoO5R+VYktV9c2xKv
I6MhSAn2jcWUUfXchyTBkXAe7sV2G4jv71cbnHStUf8oEoSHqgA0HCEmpD8gT7QWBoUQkEAWs5jB
kCouZBD5ttBY4c5ziKA0+JUObweWCp1XKfrI7NRG5K9KH1kFgnV/2t3nm4PT9jHsaCSc76sd4h7R
0VkqHtDWGT4Olll4cc9AttHXvlVc3zadpk4HrbobMx2cSjvGogmYGKGMZBiek0ZlJnPvzEhSmihO
ZIDkJbjWhgixPnDeK5iWQNj5M2cmDy6k9GgLJEPZ4AF3PtDxJ8InvemRhl1Ck8WEysZYBJCX4ON0
3Ks3RxT75sPjbV5pliKWmG6qi9x+U3lMs57x/UM6ypJeqZq9D36Po73Dp4KZRdazINXh0xyoK3xH
C02wZU9OF0hWtpPinYzUAKGPMaGk1U7/WlNLpO9RoyY7SE0ddBnNz25CF6SEdCKVNe0JTfrskmkh
Y3RH1eyEd3mKfJ3zat25OJPf3FDhnMpcnJxSh92qg8AF0I6UhB5dRpjOAxZdQGU7d7dCHJRVEePR
/0K0/uDshSvqSpow/AdhhBbEN+nhEBs6oSDZsTDS1MP36pr4cIz6fvjmpP7oAZlUofTl42bZo9hI
xukULYIQz0zpAIIB1WNgmBEjriCkUBq4v7pVbIeriQAlj9kAQYv+xaUnIL4dRLoZtrHq7pVxvdGz
nXGAm5EB8JLrimY6XMrUOWkeqS0tCYZX8JNXxKxJJ+k8alaJ+6jwiI3YaUfUCWUim02b94QVvYWC
/ICJ9qZMzpqyY5jZPYQ7HUqW/w4AKqDkh+7VsacXMp84Dr0C/rbJPVHq3gTSawiqAfzUo/+WmDog
UVb5EhSXTGK39jjWo32NSnEk7XIYq3ovJz6f8a8ALo29vnzhd9g29Z5Rt1AyN3VraYgGTykM2c5Q
MTIcvqN3BE0+2Q1uiRr9Y+2ctdpIBLg3nzE3GpHE/9RZks9rmRO90kDXMHqiKF5zxGNMOSX+xf2G
vb4lC8VWJGUbmResu/HnJaV0PcprrTESL5u6/5Jz5yKZgpKk7OBQIjF9Vgl5Sxj3bcXv7nLx85f8
XTksEEVrE1EoEqxBpyE2m9xSHWTAF0+dScTVJnWQtBidcWvK5BaS0e9nOHBxGvXnD9E3xiuDk3GP
BbT2c7Zh29mvxuJsJl25go1nhth4Yc96vMr3tuuI35ga5VhCCTiiLJ3sOzaqjnTHFfheDq+y6nY4
WgkDLiOJgFCcxFvmvWrRBJ+X9ZC+VAqvjKWKuWUqkTxpZME8y3sqDGkjyFAH58VrveLDFUaQps96
kQOKiT3JeDxcHiM11Za5vJa3Z0J+rH/4H9potD1xdufefCBpYrSF1YYJ9r/BY8nwjAS/NG4MzVkz
UEa2n/hNB5f9aSgLYP7pBIHLI8KH36pMZAW/IwjUSCs9+WmxwipBw+NT8utzg4JNWNZHBU2BnDce
8S96N36JFiSjIesI4Rjfsa6bWe74fZMIDefLgK8iCMx+fKX2mpyQZErWguVS0ZWByfzb1pX20l53
h96BAXJZL2/DVht7Q3YyjOH+9hzbubhO92ak9MnreQ470qaFEMx95nIEJT5OICTi5yCc8cnF1CoJ
MfO1xl4W4BRCuWAMtUb69mRJzmw7Psl2hke5mVWYc+Ex4XRH74a3eJw4eitXkkoomHsCnk1GjIvX
2PSKH6wrKCTciz7jaaMZCbtthES//y+9Ot4KqF6DPEUOOmTpq4tf/e5rROcJQGI/OzAkSbRrDioI
JUG+CuKSJH9LSqPg3ixYMsvf//m8yod9L/nzfFWnMD2MMSwdzSGUHeahxSl2U5AuasAXgk7pldcK
yK2SBxevQqbxe5S1wYXaT7ISxUCjx2yTgsTUdY+CzYSAQIvKJ7RZfcM/jnHfCutEPPqJMe8QoHRj
K87t/jI2UYGR2ACUpXGSEgwHMPIXa96kw5h3l3UVj3pU3Cbe987PG1H+j3sOOwkAaWAy+6Nmkta5
OI5J8LntOPS0R7SaBe1ptI+XB3+GyKTeYmi2l+0vfk8OzJtdiNNhKZZSwqyufw460bOOSj+MV1nC
E+i+HcCxbh2jzPgHn/PbRKf92oXljkd0BrWRlaqZtray2AIvLFlio5bpZBLOXtiV/4gptlezJIxp
3vogGktaEqcW611P8CKQehks3w8aGwyz/vEjQvBoRAh65HWSynO5g8EHZeiByUOG2KpqAIzhySNw
CGzK7maZbrLObeIuDhFfW6xYL0vMdz7d0j2kKEeFCt3UzT4LDSfHPlXCVh5cjUM+fdqVQuYqdnDS
VNqzuvoVT+KwMZORcDF3sRLgm2ZdDaFgHjYn4On++zsK4SR4sqzEZOvypXWMi0SaMwisTlissd3o
2vD6Lnzj13I3lHDj5bkFJmZuaCCtEDkt01jMDupcgy5UP9+UTw3HkHvQlrLWE6Kj5QagV7nBeMGG
x+KUB0EbERTCVc1oKjm+D56xkT83CIZ/V16LlZ3YM9AmrLqLIOsADaS4j5AzVlXGCOoEG4Esnt+h
vxPBUfE8QYnCVWakElgJS1Rur8nXOlgRCyCKthYNruE7b6PUmQXSTQ7nEnYAAbY5al3Hs9fAcGdL
fklfZQtiW7OGJgmbTwSq/gf3f2n/uftc3KAPbW8ooioMDzjz8opiQWvYQE9ugS15waWWIhYGVpLX
X5pzTFdFe8U0iSPMb8M9U/UVRy2OxRYN4B+VDsvu68cCWvumuJE8Z63c2MGNsw0+9hnv/GpMS/li
kn+Cqx6ocBlYbLLz7EXvxw8LhyewacuH/3uGMiB+iKB0yuwaGVEWc4Mq3b/PEJdR2c4dT0zXCnhw
JhFBVCp8cohjzAx3l0t7g1+0/JZVUUch1/cht2F6z+BiXPTm+b3elvPZPRVH7EyV4OzGhE6fWoLm
ZcRl4IpPO0bfSiPgxuLujQ+IwpL/kKIp9H3KsnKv0hsr1w3Efrxh6A8TunZWFkm/XwmLeTbKlI8I
qN2LjhD8xM7T4/YEYyQmd94yI0h5cniCEf9d33HbTLVl+MktO4j3qp+65IeSAD86MY8K+KzhWe/O
93tjQ/UfxvVb2IxmtXCKFEu2YOTLaw4EG6IFejrPtb18fup8bccmRwjsGij43auNmg0jfdt/FjPY
H+tUnAuPNCEgjY1v6FC9Q3Xv1BvSTecXgnEcDoL5a0G5XnVhiB8DRYaiaKlDBe9r1kdgLcmRJKwj
zHONwE523KCr66Kc6ERTT3Cr8RrMfaae2cZVaFsRyQn59Dsy0spbt2zKXy9Ws9CD40ZxJxq2NRNy
7zAD6vJtYbphYK50zBXlIlCu47MSMB8bqoQ9hf1A5tJA2b9TTKyhKs/lfNoQ7z9J3/QIDosbtGjs
QPEreb/r8eYtJKrb+gw/g6MMhIS8NXbu2mLo0IyOHr5vYo7+QxDE90k8aFQxCKO1Yp1Fl4PKJs66
uTIdkm94FMql+Y8XZ4hmRXShlKQsFfUfmy4LgQFVaOnkDDEzZ+nJ8pGWZOYja40TJ7azbEAI6gdq
bIR1lfgiVcv+vy4RwVKB8/W5anS+eGukK/bZwyt52CtkUIlgQVYuFp5MsGkRTLG+FQPqzE7Y5LSk
cWMX3tfB51657yA7XSPZY5jFEiMxFJsPYq8Z9KPe8hKxl/dRO5zlWN3v6oaV7CfwFFYhngUVa5By
2reWIXHFoFHCTQGbG53S/QbpyCqN+GPBM6WiVSGR1YwJ8LDoZnkOIH/ojyjr8TJnloyO0sIuSBHe
s5TZlkDpJk/NZ8E6g+lnHpYDP2vF01FTTJT3EAJYItiKZLY3Ap2pP9Jer08ecI4a6glBQzH9eZpY
r78kqbLgdSuPAw8GW9eEMcK39gV0aMyFLZen55+Dhy1vujMSkyUReN6L0ykFAaRROPtm8GNCxEnX
cP8qIoATfQU5XjOrSMTZsJQZ5lwkQGg3//y/w5HtP2FYO/oYdls1jyF4h0BUuKMGPuViBlsS+D9B
bKpREKE5CQqgyKDUkrFdQTtX8yhFtwmrn2BndKZ+z1k8MWXHiyhl6rAurU1h7Wk/zWAxgfgW3YUy
jZU+RSI6dwyIhZaE3K8L7yYOc3Cl4hEOP/4ct5fMI2BpfOW/FCHqaFZq4DNPCfU7CI94/Q8xzE4b
2LQ9V7Z0yNjZg7RAgednSZLGW9Mt//GzB1lK8NM5Hzet/49gJrFVjAyDrn/3jvaTVCkfG+2Tkt4t
JZ7ePYiEz6vpqUr+rXr/vjc4n49lAWOMGW2OiymL+eCl03LUzAuuj6vAH6sxnM86DoiBd9k8whAb
f/tJFVRGO80jiztVYPJEZSzA+fr0h6eUxtIHZY84ZWhoto6fhc24OXZqkBxklyWHJhpR0bW4r9bU
p1hKPhM/k24HHstan97NqyTdY2r2PAHKpFIWwUzdmTtII1KATdRmx9Lbar1XsP6DJIW5++9xCK9h
O5F5BMDl3yIW/6+lqb8bcHKh17N7Ltg8BemIHA02ApXXOpQv+1cLXuXZtl20dOHCQl9SnOU4R1Iq
j68z/cCFLVcHrwk9tlDGAf5jk6j5++/Dx/xYZ6v7MBKGn6rH0dRbYS9qDsMRlrbhQYJY7jE9KcJn
2Q4r7MObsIttHNU6x3pA29x1vBCb18C7qoJptRRJW7gYcjWIJuX4Mgab2mlQyXnI5zHmfntj8bey
N03Ez1ZU4t5/wskhux6LxEncHtpejnOYfUESnXhXPEnlralp+9XuE+V9rZMQhoSLEBTUZ6tQUiId
cjLXQT4Wd2MJiOFrX0OP6n/97HEHTBjWsJX/m1rzxX8eFRfg/SMoxDRrefByCLds7mIKnD1REqeh
fM4HsoTf35kHb1L4DGmtLWkH1SdsWXO/l5vrtnYCcfcKdQZ9V22jzRf0Wxjd81T/u2w1leJyGFth
LEjMELmje/GcnEITgCeImh7lXROxqhlelWCQLcYct3rntpHKR2y/rE31k3FPrxlDJAcQDm9KXhRV
682Crvd7llgVhLg60Yi+YuxYAhCvjU+PkPoVTM2Qe5A1Bhjh3y5vAY2tBl8L5n3uVabkfyP9h4Qj
N6jyVFee2U3Cus+L0TLUuEL19Hwbcbeppb9O6hKjQEpjU6NH9AqCAwEzSIhfefeOhr9xPlcQQtWf
SpIhwBNP/Et1WBss8M2vAtf9Wh0YR1ezmjfwRnibfwWwb8bHmEV7PPH4KY7ZqiBw67U0iP3nv3nr
BenJgsyzt7GnB66ctTkK5WRB+Kg5ezbWQeJu5+wclxsUIaFIjBnmp8UHvEM8bcLKiGQc0mywyI08
ChtbbR7AAVq+1gfBVA5ub71OJdMi9zWbR4ZHlD6hl328wzrVMKGyLNrFXO2Xsa67/fpnJzU2aGHW
eccsNsh4emnatnur4wh+/umXoI3pcva9Kl58DfINNxhFYlYOoYmHP9ePitgGKzDkIciRoru6VvHR
IVw9hH48K/m/xdVwszYD1irFAz/gulLI79XLOkeRcznpdRfdJTHPOHsgzhtlIIRqItD+BauZ7OX2
2y2U8G8fpTLatOOiY51NdILCBiNnJ9RVI1yuA0AhDFGzJzmYIpxYy6ow3XHbowvnRFu7EASPpvcg
e1iI097mK7sZ4B4u11HdcXlujVTKEd+JF+47BvH2E2RDOYKfFvcGAJgq+6s7loPloHTjU2DIEaco
qYuqgTdDexO78BOPqVdkGG1kY499nuxhQG4NyQOtLkoPtVKymh2GWGWuECed8+dvanjlk1eRs4Jp
jNaUPwhs4YNxTwmhjIc2mhy+a3PIjybsiv/EpRqTzxKqYvmy6iyo+Oe2oKwQlNsLxnVFwtP+3lr8
MTTw9BIYIpSOijA3EA/QNi83k7HnzlEAiMIzXE4ZRsErluxdeO743/dA9LG9QijgNPFDCnE5V+76
Y+R0jWF1Mtn3A0RYVjyBb/mDhA7uU/XUdheP0s2zO66vfqHJVPii6sr4co09PD4ONoIFLrQWEgb0
i7IptpW5efzonfwsSPk2DuoI+cngC/L5Z57SmscwuGH0MRWoiT2rnrJhuX4xeibfKkgGQwuiBQkB
gyOT3KpJqkeqLGq9ZF/7J5wqGxPRSNZGF6EqxluUjrIepWiqEDb2wU9r7LHRX6diaQEC39MUqYSu
xm/f+U8+C/GvdJsnOLZxzEgAOOfiV4LZhCwsgcINaSnDmrZO+tVrCNyvbKUaTN2VDQTMX8pKYEad
TPqttuYXyyUpeyHbb7BM/okwC6ta9Ljgdid2Uo0zN/jT+TiHLYXIpUE/cPCNNDJhKctYdFNhIurQ
J6PzeDz9pWnEvO3YTnc626qlrk2x1eEk06Uq/BHLTZjc1rZcYFjaJVVtxTnZVS3tRUcJ38X+rwHI
Feg22JGSho7TGdpSjNYZ2euBWmJKmomZUtzUnEkCQOgtmy+MA9wKsewRiYEcWuGvTAdxOXuxkWHF
dTPpgRYsW6KCYUJDRgUIoiQZEgUozltoEo81CT22XB1BETEpwMTO2gntHfxMEF0O3e/0s4BC95Ae
LTWjgxGIk2jLF2kahSn9OloYLb8oKlqStAkqxFH3QRfl5oNJArCmg7QWpUR8v2VmFiXCl5moOZae
bRBDpqWOZyewT3FeDb0Qf2EsUPmZLF8MKGRCPAMlE/9DQ6+effQ5KzcyISksGclIQY5ULY2HNpfT
uxUlU4dq+000n7ie1xY2NXb0fFzP3Cl+llRrLYJjD89OL5vxvpN6oyla7QG87psCU3DAzzRM7hSw
VTihWmUTg5LFbrF7p4GO7TpBvWbJ2kX4DBJBfpgn4qsdUF2geaUXvytueSejC+bSqLsyJWMrRtph
HyZ55fuzPmWmRfrxvTyKu29fyMgsQGuS/exM5VTrqnjTg7w8r4vtB7IsmgNoi+XdnwP/yzXlnB6m
sdsJCjaC1BYUxEGwtusZwNJXKsqaeBE9e0NZUxmPgE6z1s+A7HiD8+bptrYIV1MMFCzmYTswWTd+
IEnlHlK9DSHLNUrcv0Zb/6LXH0FWU/Gac5l44MP/3mZxBFbvJO5bbRw24e4SxidctWGqqO1eC688
ZV1wvIGdcE2yexcbAkdAMIgzk5PeTA/29heG8W5vO5hAkbmUG3vjrFAl8fkNgXrdtYafo6mVKmBL
cTWEB6/uv/qRel+GouV8xjQhDjKiKGsjvNi5XuIRnL8zFvrbYi+Flej6xiIEeH5xx/A1IXnScxTr
iyhX5YybRYixHwnGEnD3dlxwdkBW8dATlD0taNUSi203Bbz2oGVUews1kMTxKBS2nDrWZQKgsEcr
tZZIn/9wcqNzCvOPPjP2Vj3raRzNUUHuAkRzllerf9SdMDBzNpOb2PrFd64s1MzN2CdNz8qvgAMQ
UFxGZVDgRpC2pnw2WbBs9u3IRAFAz08gjr04bZz7ZnmrvigRLsB+oXgiyjH4zGo8zL2DH65VpqX9
gJ9uo10nlFtn3eto7spaKV35Fte7QuVUYNXtxUFzNCKpUcw6zNwkbiC8QNSyHyilRuopQ/xQpzdU
XlZgdz3WOKKStTdWX++vyziI0kW4+Dvfbu6IVkZOk4uIDKBaxumFYf8Tt298R9BNRY3wN/KrzvMJ
9UZ+1//3LN2bjjBx9glhnJRef7zE5OtscF6NzBkNV9b3/vJYhMrtA5073Lts02oy3V+Ve+JP4GXk
c49FjyX5h4kmfW3STT9jlfClyYUJhWVMQ9Ke47thRzWEitDq+kzWLmBSxbhXu9nlrVFCkp44ydzt
BkQhWJWb0tlnr2jOB814xJ2/1iUvuePmxTYpnlkw2PqIU/fWReLynxDCk86mIC8HamNmy7Ptc02S
UL0T0j84v5GHlJvcYG003cYSk/0H9EuwsIxXHCV7ogrO+8+1q/DR3l9djMLt+uPdNFNOGuVVfKAn
Lavwt8bWyGK6zK4ZJUXqpvDe0GVC4xUaDk8xjSlXnDJR/k8Rt2lfMA6WUAh1GszmwJjTN0FKIjy+
qBPtaiRrLKMaP8UIlbR3hXvPvk4Q4rPQAuVTEFoPOBvPjsDC+eBtbCkS8StmGJSx4SzbSzg2qx9U
3/lDbD7cSdYe8HNSxguyVmnNSJfPXU6FovL6bt4IEQ+jewIz/jJsQ3XQz3++isMs71teOpEMQm2i
S+OMvrgFJAlj0ZNJnE1nNFNaOUAtdA6LKDXoq/mSry4D3GvGwrULnVu215D1j8dY8Tux+ondnKyU
BOUjLVvnBwDcF+C/eQ1jg/8BseO5192uLVy03ixOynJOKzbSYKs3mGVERlBFx26/Mq5KVrFVeFDO
2q92BQAjg+2Uugj6fn0nJ/XduUVsI99Ef6Lck/rqft4mrLSxyWa8cR7MuBASrjRL30nr8l98uEyf
k/IacVJeYaU0s/fBLM2wYrVY2hyJZuXCsZwVP8itO/kYipSNIDu/9N+IcznXqom9wbKoE0PHK23q
5DFdOp0L1ULNM4uZT7FofT8EVfpZONeiW3JuhDwoPZPNu3ntVcKfivAPx3PIV96mWgdZCwDparId
9HYaLC8rEVhjIKexT+20ZKZ62p0WaGnvFC8aQUyq4EdsrC+Xmj3KEgg/FUbqQalUKIR69WVdGnZZ
WW+gD3R6I5tzoIBMnDRz4nAX5FaUVif0TiNwcxQf1fkOs6kRcOYzqn1oMCoDIY7JEeBgSrPtUooW
1YMDxZi0G2FJE4nKG2bunNWljq7F9X/UECIEW2iG8j+XSTHKlLFcMitR1KXcXEtAMkHVUwVC1RZI
/XZTajGga7VRYG/Di/Jg0tXYc6RWagz7XRsWzTSpcN1VLjXYUtDQ90OG964EsjvcsD571QvBE8Yp
6d5tgIQ/yI3lyicQtEpDNRsRRC8/llyAUZlvodWqXJ/WWSEZ1Tq/CHEC0ByDW6nJQgBwLbf2Z528
FNu3PefNkxtsZ/87uchLYw7xO5BaM+i1PRuSdZPwaZad3hhuqlsxX8HAhg9mQdkKQwDYAZ+0TLoi
RaVOxVT9+l/Bk02gUvk52GTJaVHBKkG6x53bKgA4Z/3VB5AxKnAb07DqG72nSQ/nV5rya+NGQh8p
KFKWYTqrVBoHV5l0Fa7o0E8YZsWDbbmtdqB3n8Ko7iZi30tEYNnYUXlupGAkZgMO2NzVkGKhsFkB
DSOBhZxhBeRw3XTRwfcD0K+5gu7SteiCL96EvSgf4LIa3TIz482k47XgJLBQMUk3X6zxMoeo4LTn
txvGgC4VdeWI95noSTJn+pmJ4BJWZubFrjhGFc/l6SPJZ2aWon1I57s+6yq2zJJHH5bLyJk4nMYL
MQU672MyjW1hA4XPuRXWEy9vbVMwvD9MpZnS1lDYgKknq77l3GK9hSrT0Wc87lwgaaix47I4EEXy
EVFhH/dpL+UOwwQ3dYaiz0YFQGUzbXgAaoVZ4K4Tpww9nQwDYUOfkoD11/NXDSb2RIsQWxc4zjTy
ejTRkU3ZDw8nvMDmAQgTdZ/FJbZ+d50jIfDQe6CGyzDu48utNtdCKa9xsVu74PQavVSUCNrcZxAt
5+M2+J5CGBg+2VirgTVCGps165T+IMMiGz59xVu8oBiWkyELnQ9lYRKBmtqFy2VzgkCtjSBNINbU
lF3UCxFMw4q5fO9gYLQ7Iqz+dIy5EtWvNgVR35Rlf8etFfrdZLX1WKGIXKCUr0lXweVmiwiirpwm
9HokUp1v4/r8O+xOe96IXLzJ1Pquf+cBMUyrGY/Wj2YNWVZJjBA/Gxw1QtBz4RzPLkoq32u7wO59
4X6VhPK+HVpvPhp22jGy2TTVqJvQU8XD9HazG6SSvmu46WQu3yommstJlU5RvNGZts+gqPDB1/Bc
iVfYij3+8YNcYKxFsbAw0fcXOxbKk2yegwVhZFu6txPfq8h7Y1YmkcF4Q5ekolQftq2IqC4o6W90
26KSmV9MHqBdZGx1JZEJ/RubSZlW7UzSgBz1UodU2gEDRJXopl5/M/8DOZiePyFlBlXiVTQLtuJB
CwYRX2W0A/CpFyG4L7mxBxA+GqLXKqkFM/dvkmCWy+QP0/1P79BmoHZw1iJ5Mn1oNELQq9uQm/TG
qqZ8kPYLvsuEZALiX8RCNPrexcg5jamwStGE6ZCoAFk/Oy+wBllLwzLRR5ExV319M9YDycLBalrS
ir9QgJHWkxjDwtVZncKOXZVaaX3Kq13AFOK84dnvyycfnJVmq1xCi9PixiB/LCk5NcyOs/BE0k6+
ERl0uWfIDnPy3ikMf/rfOtZsJmUdcovHfO7qwnBc86X8MPeOm7sCaR0jN3YAyrRolGABmLXcn3Tp
bIaZujLL6camcqOgtkuup+AdT56RFWe+t8nT49DJnY7bMm8pG67jE+9cbf1r2c7MUGXZrFCL5rWF
HOFZeZNI7n5IdcQ0Zocp2dDU5zF8tVktlSw6nqDMqB9RlhoVIAEuBR7h8WrduOd9ZElmYllSZnTB
9D+xcmPFMSQVMQ7pOxwdNtOC9zVQeBIJ1Nwo7U1Av2WMgpTO6yNrOM8F4MM6c6rhVqrOGZQYrW01
7QAhCE908KUj/dpVZIQkGGPEenpcBhnE1ZFSsZZfqROzLpci72FRPXU+3FtK4Icr+IB9m8vQVOK2
mxMOwBZ+qBqLtA8vTIclYlX5v5cRdkl/kFC/ps03eV0YHkcmwk0RfrA9iSvSCXcFUhPszuRJvrWU
248kIaQi5JMnM9XEvUBlo8/+R6RvJ/8vDX2b5gI7193zYbKJKN2WFJE0OQejdMJj6bsnWiFz111f
VhoFuswHGtXyKu7JrRsrbor/IXEb2mQKHqZMTeXQhRWA66QArZXhtl01e/fNlQKMYtocldncaIuD
H3gaOFgiX4bpvd0HwkXDqqEBSUcmCjCYUuPMv5bPpNt6yB4+52u55EGdUBc0IuOL1nc7Si6XbPCl
sYCc0VStABExnJJRF7ozMcfwVXq7kwK3yGOMmWd3tFXwTimjLLtp+1Ls7dv4bVdwYeRWlQ176SuO
+il8kwp2TBb71BU5/st/Fwu1edYK7VpxEQFFtjl9qg6WUMC5+5LymDqyogqqNMR4AqYa4H+n7JcR
RdvJ/ngNfXSnGbi9YB5UkFBeeHpsbt/1uG1cyvNnACx0dg58J3p0pRqpqoQ0W4NzQqF3szF7/VYk
jOXO4S2wtmFYvIlfHhzWFZ6X/Li+OqgYgKHVMIcJJY10Wbtv+05bjDfkqFt76Cogyh3QbW06h65k
P3ljQ6BrW8KZnchpplCv62Jkxc+3zCsK7LQnPlrdvY4IFgwwwUS5fJFN6rNWduh/7uNt/UVm21o3
kQaDM2A/XiCm80lvHLG+CPaRCCErnPPJE2wCISqpHRVlJq3gM7X+OCTy5nEN/L/512buJSpYnCl5
A8ilx8NcZsp/PmpduAThQBOm4t3VTLrBtsCFEb5FV1sB2pBo9h37uwZB7xbdXjr4yJ4ZHSpt6G4m
V6LwqbHvuTGM0dIrelUGihgs+ZVi+gui1R27478rUToQ/dZRqn4zGyp5cn1rtfCW9HI67n6e1fKt
R/qHVSlIkWifJEkYYaN74ddTThuYP9Ti9YNswBhM4fcVKEyzYkla53iLtmQ1VhGINWy579wvohDX
efYcrp9eqwCCYeMiLTMyQXOpiHn7FVsN4RB//Eul54OynLf2XSwgWhdtb/9QD0dqgcAcZwTnmUYa
U/np9h6GFXgsl0AXgkk2AtK7Nt+TNMmPPCHcP67AV+SZLCHi/yCE4cBzP3gMN9g+8wEnLtohipdb
f9F5I2N9h7nwpTWezAkJRhfHl0hhWC2m6vsf66p1ARrzKNcD137biq4YRMHZ5G7PAs3N/duDUfjD
o21lgfs9RgKyl6Eja+s0yB0N4dfq4IIvyUvCq53GDVzBTPeRD4xarjqp3GNm7Fp1wURgsM3ObAL/
sWjGa9f5NZIH6Ouq1F5Y5JorIPSOE0g0jgX6A1tvOmEawN54xbBunlrQ4QjOkyIDUXYdx7+bjQOw
/BDYQTYX8ZDpQ87uZe09upyFVoPQYU/nu1RzgTZulsa/epoQvUdZqSMng1xxBJggJoY0FSQ6tlsR
FGRdKqDxpGpj8mZtFMhi73jvM0PWTddc0xNsaJd2W+Wv7voNqSdGRFplaEMaaPY8Kdqow0cYNmI8
S79Pd0St0FSBkCXS4HheEoubgWTHTNOPq8CeyTIHjG6tb/Mygv5NFZAucZjotgw66TLv0eahjFBk
YakQ+acyg1OUskndFyDx9cGYRBC8FNHgy/ai5j64mh5OihGR5lGOc81wUPCJl0jgjXqP6ncqhoA5
xMg/lnRWdHPqYHDJ/2GymD9eEKEmz1K0uYtolZNdTZx9sdfScPKkRWC1hKW+EFrOoaEeI7RxPLb5
HpuTdJmbf7o1njWKI4ix8oj7HgMG4aFcfW9Saq4EzE74EoDCnDFiJ6XHjFO0SxJM9chaxLV0vg5Y
lIT/yWhLeRC+MkmOJ/huEOkrLvRohvPWrd21FcL3I7tlHY6Cvo2H+jAJYJ94tIqdQ40nvXqnynmQ
6S4D49tlzT8EY0nPTKnp/3NA/v4ISsuIHyP/Nhkqs1i4v79B12TnNFUxrx8UJcOi5ojBPdri1YX/
B+NsSz/cSBKHR9Rwtk30KATKUaPEkTosrBTlPnhu56r1RKy0lTmckgw7sEd35L1h7vPB5qz5Hk4X
4kA+udhNH5k94WMd76l5k7xlLNo/zbqJN7WgWvA1QdBUDJsRnV1aXjmQwh4MrtT9Uj3czqMuc9Ey
STSdRSDqRTfilXYNEISiV5pqdTK2aOn+w9tEk0Iw9Znn+8YmaXuwtoGWx7AcbRU31MbxkhBug6Jc
hHbUL/Wsp4uFPSB7fOPXh45vO33Un1c0WPUH9SjTgssK19R6wWLXRYs8FnuLG/gvkvACTpe2w5gz
XDAkQ6k47SLyvKBN1LezrxSllrlTkg/Iq1xNdQCN0VRTYLc4eUfhA9JrG++RgHqq3GUMdtB6GThY
PVV3jgCbkml99Gl8a/ZGhb7uAngbFtCGxgGvG7mFGJNh/kYhxEJiKkYHHYDP8qZQXEwLKrN35AuJ
L96suZl+KAw/8tWS1cBIC7+z/9BJoMLNSjUxIXIve0jdPupjq7MrlmC8fGTt84S9rAaLBPYoFQ2p
nRMT3sY34xo2UzkKgEHjJigPNjzqyHj1DtOUG1X5R51Do7bBdpjKcr0EbU059nL6H/NZtDzTm+oF
veMQDHxVOlglnknfUo2295jo6RyVtmfeHBkW7TQdDfqgYiTjEH/PkNJDWsRIp+M4Ayrs9YjOP7Xw
6jUzLSzpnh8nubtqHcLCbsIkO4Z6csFyWRA0gkYMQvwvwBnuyvwS0lv7wKXaR6WnLqsEW7G16kLu
dvpa0vPaB0kMnTWX0rH0dC3z8NQbLMWsmV6vIXKQdVBSPmM4qn5c1D7gw4TNuO/cORJH735pFJW2
phD8JdH62GSNkZajjwY4f7ysmpmoTqVEwxJePiMcLnDEMMgAJzMVY6ZX/k86OVfKnBF+ru8RU0dg
35aZOrCqZkG56SBQKW0k74fHdnG45Qk5pItIbmvU1YM6qd5HZTSACgjk/c87uIYvAAV9/e1u4/fU
AfK6zmBF+bSemUxzy21BmiOQRCP3sftQcVI2jPshZ8ZbelOVbvPNAMhrypr6ps12nZShUbqxefiX
F/ihiLMnLkgIteR/undWyi1bRch3YQpivupune3Nr3Qp3xK5PHqa3I1UOGHpYpetdv4nKv9BczFm
aP6lhs1VyX1bkApsH/VEq2lDdY9P/Ipoh1+A+f5IcojLD3hoBIQHivOk2VzTphBwADRKRrUDMt50
OSM7CR8z5VZUgVQEKGozmTurjKy7sndTwJn4QJG5sB7Vqya+KJCHswuvE0LCOkuTGUokkM78bN9g
k1l0A6jd4SOu2YRAE6Fc0Z+stsvB0AljMvIwxJoarkh+UBEeMMCcTjezGZvy0WOfxkd+ZMjzrT/T
SU8UQyu0U3jGbFnBv69udZ31KmFQVZ/H+LAe9s2Ms0FXvQoAhBFhXXYxQP/yq2zauS0Qrvifg3D0
NFxfmkgABgE8cHYo5pEY4II50w04DLzNNKH0g+B7eqK1yo2huqlCT8LFDujJwvI9Rc7xF3wsY8eV
6qbfxW/s9ZXQfkjAdFJjdD1q+rfkHpWDD6CNPqLCGAvvAbEy3oUzvFKNBTbGReRJkk2ENfP4Iucd
NPWnzpWZfFlNUptacSjWxd48/JHnomuBAwh9xuXOBxGLvMiinEYiixH2SYxSlmW1oOoEBDmL5Jo8
f5clzacoD85vZKTscOkq72q0GiZMR6F+0mtKt05gxZEdlEVnatw98YIjVBmmffSTlXIlUl2sWiBs
qJc6TLO3fQDDRSxWXXkVBf2dL1nBdpco8s1yO4lM9a5dqwyeRh2M2EidNBuhjP0n3c9BS19WDrB3
nJJlPZtFckVkpZxlKC0L1Zr0kfhN9EqkGAi+OT43j3LRKG9pQsKEQtyj23H1W3yFV2y9fREm/q4r
V9fgoE4cubrNoab3WI5UER64EZnSfjiz4ae1gC4aaiQ9BLDEmWF0X8IRjVUFrELBOCqkaKKV4PW2
RDtSP3DG83IhldBkmiiw4aYQbLSvyrhTJO4+qZqCnlPtXSA1/NSdVsAxY9OyAG7O2vZEpAFq1Cfh
LRAXnl0b1R+KcCCQRYLZW6csWofga/Z25dEzwXffAj7bO2VKclOMZWlbuaWlLBt/q66WlZQ6Y4RR
D/UIdnTJgUfpvbAjtNO6cwqOr4PMEEVoUPEY456b59AfwUHMppcHLCV09EJ8rQ7T3F58izgxdhfr
DAC2vpJHU7uq6wbaVNv8V3QlQNT/Udmlkx9DbmKOMikjS5pDhq0/Q6JS0w5MWaQk/xACwQ1sNmHF
CG/dUmbGQQlVoQVV9s5s23IpigRQJNTkbBxsHmLKFZY/oDyBpWG0BBv8uKPrqTpqCSY7fsbaABoF
RUBwlcd7WuQ0vYwg5k9KIoI9GfSzdYNPG9EnYoqMoHGe5VfNPmBHDxo8tfk573whhWJ5DEZCOaGm
ut60nJEz+t0J6cmwEXROIglM14rA/EUwMz+Z0KuOIy3crTn/U4t/AkB8BfFUdLxcLfY6lA/aSzsE
FmaqtDTEtMg7HVVSNYCaOEA4t652ZNNpC4NeN9XikgHTb6r3FCu6eAWYcddp37O4mrH4YK8mQyQJ
qvPFkAjirXncL9Tcfp0MsQ5ZQwrzWfsJSAroU2HsGwLVDlD+1+pUOLxDL4Vaaw68zY8lgsmlCgL/
G20C+2aH9NFt2Ux3bYp3LX9X7pzwEKRWeovXz4RTKDtuYFQafLTD8E8BuI8OVaqVydrjFz11HwNF
/qpyKyLyXRcT8dRNSZI1pyaIeWwNYrc/M+6lRBqX6u41A16WHCZTdu2uQIo2voaua6OXLQJ2DDRU
2Z4PETqainS3+EOm0RM/ADM7UsYPMTIv6jv2S7ALKW0CzCDSmbpNELalDQxE44tPHLKd75OzOgtD
SVpj8OJbcs63+haDQo2b3GGeUO5LbRo7BUwiOwuORWoYy8fHWLG7yb1lZNampO05pqOEUGXissbk
VrQcyz7leCHuskTl9/t5yZcPXvd2D+xRP9ewhhFxB9PQPGXQx0lxQOlgbxdQL06sE3uPYpRZIZsg
jX33VMxA1WlhGs5yFIs1pm8qaAUMVbPF/eKg6H9JNKdqbiAKYGOfbSeLpcGHMHSTgSarf4pWrfJi
QAzZKYikFKE/l55ZlG0x8N/6w0q8L63YiK8aLZk8Xh2S2mg9xwKcbjWBK4tPJ3MCd1EzV4A8wztt
9kGpAWelygRZKk3dCC2SjkXjkOixjT9T9DEQZ1bD4pCvikSsH2WcikAcCrKd5LrmV9+vYiLJea8N
eBGE/k1iht/OkBZRTgvQkT1wI/GCg+6zaeCtv0kkAqQ9goOjNy7UvetHPr9bqnei+bDdz/1YOweD
V+sD9T8cWYsh9+Iq9v1ZrbpYKwLgU5eAaTFSN1ppwzb+gGes1WpNAJrUJyElz2jFxAo/fK7+ZA8H
T1BhNLp+UnL6m30nTwNDkNc1XoAbUZoNrVgKwJ3ACFcfiJgFj5OFslC30nklcyn/bFL/2FnK6dPf
WiI8mpD3fXe/CIvMml9ckHGQVvIQwpnL2fD5Tlj5tN0orTkfO8AVbYMpVBi0J+01QYGooq9PQtNA
6D+zpWnfcZQMoT+VsiuIuWPrQrpMBGACGcCiSLPb5P+L7OW1XFptyitQRbm3klnRg5c/BQgHPgzA
IhJ/vt0/wyyAvv92brzr07SR8P3sx4hXADlhl9WRU9sMqiLNI4KrbTyXJIT30XWwXLo4hnlx+I/H
PbOU/ZmBQt+1nwR7Jw9xKIFnXchVjYl6sUZLOo5Xko9uptzHf7RJndvYI3n3sISlItG9cU1hBFbr
Nfmm7hgs7mtpacOFv5iAHgdZHLBiiw/OjkzdgIR7n1/a/xSCbo06gZgOAldSv3rB1z36b6uasdDh
alA1l+g48aR3zrf2dsitc1ieCkXqUoJsiENg8qZpBJM8HwtSgkmb7drN0Fp/w56DZLhPP+qi1S2F
rTVGtGeG6LIzQ2olHKjfZO6LobcAJs7WJbIGArw08xO3MktK00sTrCcaZbXvxPY8ewkvH3t4iIe3
PoW6lPfM+VRqPo1R6I46Wc+Z2HpYi6TtRbuYhX9eniA+cotIKisaEeIBxp+y5M7LerI82WuTXs0w
b3cqdkSND/AsV8juJvbC5GlP9pmhx1L7rL+tfoS/kGqf6Q60GsX6Rjnu7P0AZhh5ip+1tirNzJJy
IyIm3KmVH+zRxBHq1oI0mfcr9+uWkelq5rQyuNbP849Zs4SxGb59ohF1ghjel+jWdYGNgqsSWwzK
9AQ1ySYkaRBY7cyzY20jOeThmPMefcb2L6ppXT9J814EUyPBRVhaW4KFaZSUzqu/swMIjR0o9WFy
pjKKsuxm56nav3sc8lJZkU4uVQaaySv8Dsj+bdloKt/i/Idm6gGv0a2xsDXdZH23Q5UtiPUQtBk8
fIFW+vo4LqviYDchduZm7BTGOBqOIVCN/uKOn+rIOk86kRVSRkuYRa2Ezu7/m074z6zev8hLYYzI
Rm9YYJFPIJwwJViJJKhW0xrHuWGH0polOsTgtufNsYuaz7/+SDfa7bwKHBdMJHi8OWuZlDq/w2WM
tqu5JkiGSLIdCgEB/JRrBAHLhYXGzyPVbvgU4M1OWeXrA324trE0B6hQjhs48zkZMQhLyqUe+7e9
KAoAQ249I4mFSCi1ptwI19GTSG6OR3UBW5Ru1L+G7erADDEGY2+6JO3zjBMK6XjM3jAdXkYes52I
oydxbUYykF0xQz8cChQpEhpc0XDyyoQYcQX+mMqb/WEIICzgFA/EC+CkrTj6BdL3De7xR7ZG0AQB
PNkVKz1iGEqeQKn88ldK3ZO5YcHzrDjnUzR23sgTAPQT1PTXf09HNosvW9Fd31qmTxD/mc/fScrq
1eXir3b87jHeTQLTkrdyHsH0fF3BR6fxdUk2yr4LhsGXlEix+X3ToG/9NkvlvDbsz6UkTe1ip4wm
OjyqsVT+1v96YKEznALXTgZ49W9mV2gOWDr6JzGZvNmlzm0RoVuu2GSrv4aWP47PDz6MiaBnGBQz
A0MSJbXDnTKin7ZG7erLdYhRlKgTBJ2FTbp87te2JDgvtUx21fx5pgWHaudToWJG23Y9JgqcLPyN
LtakI/BkPLqlkA8Se/Cp2wy0OpJTkl65Bp3u4siwb3C6KVMAnP7hXh/h0+6PpO1TVgNkGume82b/
oC87QCp5EgdYHH7tsJKhvGXxStYYLlGRNH2J2dPQ0AuyqxWvpf7UsyakvBrrBtjIQYUiOocEC58n
RKLlav/8C2tsrj/+cxbqnGgJlRUcVpC1t34g5fXmDwjw2Z3XBtH9WJvDVnXjs6/l5t6ETKfgNyxW
blt8eZFJm+ct4Hfu4sSZwZEsHvgBjq4ZgUjOy8WjQxXcpXT3AvCbkdmqf1USWqmmPOOKWEJdo09A
ldH5NBJUwLU08jfGzGlI0C/2OR55czFa4Yu3eEp+lKa4nmpB8tIIvKkFupOZOPIEgH0JASRFTCe4
I2QcF3fHzQAzhnSX65GoQdbHE5pIHOxKRk0NfVVsO3Unq+WWy60pHo8B05kx/iPoCSaCSvz5AsZs
xwnnQPAmq+PwC/3fwmnaYCCysUBPfDoNLJCIDtYBiAHtTjvH66svmSn7qLv1wiQV/IcFDd42s4Z4
tHUEPbd6csHgZYYTmKNj01gdgE4jn+lZeqvo7m2cBLOFpU4zeuUdxih16saezCyXTGDwVQctFuRv
HapAeDuqvnfCn2dG7dwvz2hVGxdZHiJeeEyRNj/cGsXjeBtOhhze9kFoC48/VaiQ5fWHjF3chQ72
yLEEQr++dfOxnguZrvmBdsqYFSA+cTN0QUcmvxGfCALXmRVQKRqJfn/NQFK5hq9O8OSb4AW0wWfi
HLE3Q2gqIcv93i1XUlU4EkUI0fBI3GFAfO9o8840WuTe5cV3Gfqal/cQn/ax7WgHgdVoMUh3XRqE
1+sbC5/AIixPZg18/tqL7YRdV0aGs08SmC0/N5h5K1ey4xmc582BbANLTt/9M4ghunmit+CJBC7B
UCxhW17uV8DRY+JaNz8FrVBAff9XMEAEy8DqdOvJvskzeyAP743LxNfbBM42YIz8GGKOMEBzmmLB
z3HYu4e8BQdHdBHdQTqlPPDaiIkH6pEVPEfOAyQbCouxhrDVcv3Rh9uK7o8FJaOCgcd3Y4CEi40q
V2p5iw/M9yrl9t4RE3cFHinzb512Ta81Eqmb9yqe8Wid1OPiHtp8su0Y4+j+xYUzDp1VbKdh0+EA
H2krE/k4LoPxiPjeWqpzbUXmQF8gI3+Vj1U17ME8GZgewzTX3kY9P/swzVKbm9aqp69kKtv3DEYb
mwINp29j6nwxQJ2D3NGKnI9ycyRkswPYlVd35EA5FVDYZpp/jBUnBLXs11ykdrJV7hYcXTIo2UGj
XNsydCyypQrV4JRF7kexnanDXk/tYeO06UyKBgsXS8clG7NlkXlDFSkAig43HEFrPfyduI8GIQoh
0jiz2lI9fz4qQliT/x8LW/E2q53+Rl2j3UwumojiS3DzZ2dUAVr+NxgdItZ61ClK6lAQkS57cqMW
HyalO25Zjz7O2Rcka9ENcHfId8EonQmD27WPEs02orJF4gGKAKDkXanlMFlmToWK6hdpazaaPW2H
u8LP6/cZVKWe+dwjek9+aJK8x+LsYJuPiADep25mAuOgK1N/CrnGZhO+oKaIp2h/IB6ys9XmUj21
66YnBXpNE+IHGBThkBUpUFPfUZB18yjzb0B5sPqK7BZ5IBAqU2KrQZCWif9urJcwe0Z+suXXIBfd
MrwKzrPyXXMUVva1oOcfRic0/tN3L5MqRHTk4eWfroAO+Z2Z6j1RY1CM8oMyJx2IDtT3WMv1izN3
absf4xNf+D3u3YkesTkaDgpwMjudcou0RbW0s8EFALbknK2h8EqHOJ8Itlpshwv33tGTurLqHq3J
C9QYA3O8XmJ2N9/5HiWUBE04oufN5MF7yKPUxR5hz51qN/nA3vOr9rCyS1Eyq1pxvjRLXsigPIdC
Vyf8/V8XE4OyVOgNnQ7DOoQigSUJMmB7hC79Ab2ZPQW7xBq5YqKucZxdsPWnVh3R570DLYU7mkQM
ucNrQQiic6+gBqWDSdx1FJ7dvs21rElbfJ2M8acppwZxccGxGvnMgDmB8EVW8nhpRmg/dKtaGpEy
dGDn++Gn3CS5WF9CP7PzM4I0axR2QjEUJAGrVK6vvlTXO8aLsLlRvasOi7/0qiDEiqBeuWHclWhw
rn7F29m3Y4QKG9P0iqEmF68d9ufPQp4R1gjTK0urAW+CEaUnZEUPQ1om71yogZKrVmvfGjLqVbF2
o4yHszP/GUCkcWABMO9R1E8pGCjetqg2+tflltUEHIOoQagoGQA++w2EbQ7tnyW8BzrB1GVFy3X0
Yc5ME7dmulNe4kg1KA6KeMf0pViS6w3pXb1smn7rsFb/kE942jg9aYjBPzG1hVGDqZgUoUwYBomW
yu90rvWzirsX8+RyPPcWisMUbCp9bBVVPnu+l/FWlZObQYeaDTaFjYYBRKz96pyMU86yUnO/DNuc
lc0II7KKHMqEJ3ZJRmmVhgQinOq0W4hRpKRPb1QUEN4e7UDVmJ2xLeVQITV9B0pJAD9e26QlQwDW
tJkjanBlRU4Jgzj7U5f2eC63xWuUR/2Wm/kOxHC1F5IPY2ROydOWCtiXOU8jqq7TzTKah98ts45H
qqMF1+A1xqyOzXjJJ7hJ91jsajF+9pw2E81zx1sBhubffeaEkS5Bc696DzxI6/LXGO5fDmvggK07
GGLvsFPefleW3G9R5zWomz8PPZl5N4agOmDpfCC8WmLYiXdTPgZarSnMRubUn1jNg9fVMGrSn3NS
qt/SzKzswPUIu7AkuKsPEid8ekKX6IHLQYI5Ucddqh6ZXCn5SRFMOsTZmAAYEqmgk641nFXGHxyX
d1lohxW2SO13kig8MKT70IBxDSSFEBF1/XfaJMM/7+0E3wMiyV72iT9CgzMfN9LjQ72UDOm0u+t2
gwVstkI8VMVQfvysKo6Luz6W7NGc5z1WbqomfRs2QGhlsAJonvf/iCa653C31uYnow4VVzofuyvD
tKVE3heULMvNICkmCJXDz/rgMi8duz8wKqiTkQ1Ru00K2UmbfxRrOahlI9DP79zJeou5quopjRys
Ek1+V/zIbxVP4L9xyagYbSN0hxzQsGXnryEAUgo484SxXlOQKGHmAsKsq2HvqpUTPV+Jny7V2m3H
0Cm+gRdmXnSbkux5Z09IO4gAHZWSfFZy29hy5N80znbpFEHdsr3MBeYccIlaP29H9vqZ8BbWbtuE
4JAn2wEB4Pl0zxeIWnFO9qhtzVFtKYru/TZJ02GpyAAC2muGvRYnO10M4XDjYxUNZFjd/qiTlsD1
Xe2QOKlNg+e1cXwAG1wHsAwQVM8yl/IsP44PFbSmmvLnC2X15mgJiQyV82TtKtBW0qQfemTRlTwz
8jZpJyyivwkdEfJZdvtD1OwIVh2HIaeEPevjc0kMIIqAUIruYuC3LlPctYidrBsdUCjS/ry76y8L
uMTODB9cNODPs7KQ4IPZV1TyTl3ZjSM/h6cN8C1EVgeP2ctV1tn75NaU3gQZc0I5kPxjIt49jGxM
sk6RdIuo71Ol7tMbHSGZYgE161qvgi7u2xYdtGeMusfvlEmJarKoiZ5Bv3Mg62c+loyWnT4+r49Y
X9TguxISRuNU02c4av5bI6kK009KxNwtgpU0MYICbOIHhc6ZjLPXdiS/ZMn2ubsPt8bubq32Wlj4
bePR4m3Q1LfEAEeUWe1V4hhCRjo4Wthbybd8KQ0xNx4tPWvpHuSyoh9k1F2ZrIdAezIu1s0Cfh45
k/UMilO7d5NuQAzQo+lYgP9Fn3uETKt14P7ovkJRYaQoPPMr/SeXi6R3ofPR8kmJbW80V7DWHL0i
zt7VqqErbG+irx1EcbcnEV3NYEx1x+CYgsf07elSKshAz2NraKla8m2ijEZxVID3fICCgiIJ40A9
K+q7gHaOZX4cSTWpByJDn3WXmQwpSpLjU/yZCgu07BHrEoXoKnp6IdW0oLaw3em5Mkww9QCBW4Ia
vFfpT8982StG2Rx4YrR/aZGFj8x9a+n03HWT9mVu+y+etrGqKuFpVb7TE0Cru20qSbKzMDLuBofH
RBPA2SDV3Ecj64Db2EH0XY09SDdSvvU5uWz/tXa4tTeOzotat21LOdclnmQMvPVffh3qVC/UWnIq
FUtgZpXvmHGRb+5z6qMGAktMzpv6xdmkLddBlXxLo0Aw4s1/b9tK0vRbU26HFInJtIiAdHUMmJC4
XIvQHT6bEoe5oVMamt47DbuD7QehJwn+7CfijCJ/ao60oJ6T89SykPSVJJff7qA5BrYNARXovsiH
BTsM5Oor7a6vrrozvCemi0asC5PvjNHRYO4L+/yqPma6gsvJQ/oFVm+df7wIHm3Mbb6BLezWqQo2
M8KkI8/aF+81z1XAbr3Qeg9vLDKIrYeID37Vw2+6JKNEaUBnKp4+rocPzLdDbmDFTYcjGlUZLqTT
ExugAuAKOYFv1Krw6fL3wBk3D9ElsYMrbbC8BiBt1LXLxvP9B3011UIIvsTfm6XcdO2LIX90ThJm
V7IUPOhUm0uxc/EfMfTReHLOM2ApG4Lp3f8kctD6o+GA1wmsygZpp3+yUN7UlK6tGaB+oaLRalZN
vf5nptRiqB54iYPJfBA6s+IIfIJqbRcmmFtmaTqKA8v7aegrh6aYTseSU/Z5eTTQwG2ijvDZSt4D
aFCzhLV3fRWJnmz8zpm2nNcg1c+9eCI/rY9BcmAOOOsP5fO2OZuegLgAm+6cVsPJxwO2OydI1068
xoU5axCK/iPmpN+bUzpkFxFQwKl/mYr1fXEmk6i3jZ+QET9GXsYi2m+Ve7zl8G1lzwaywCdU+V8H
UCa7aaSQ3Bg4cfuRF/6jPkvLfuE1vyMV+Tcz/yaR0QUURjIV5ZJl3q0LkUJ1ES82ZeqSFuFygnGU
toQUmubTmi9URuw/J93HPedRlnyXPII6qwL7/6qZUjicCV3n+jefLJhWmcQv6zLL71mPonXwGjip
apimUX/TzGINuOJ592l9zG0uVBF5yAxPHmEAgwILH5F6L62C4BxrDa+6dW4N+1XJwYJDcWYwvebv
Bq6pWnoO3eR1yXFaR/W8H9A9qJLuBYTaGJQoTAe3EYYZ2yRxwjoqRhtHYCtGOm91k7+6avraaMdL
ZhpPaSlV9ffCAvz6He/MVuGEw19tGE+l3a0xSEpUwYJw4t7GaoUB0Cw6t3TBpm7Gg+yzPH7LnJUv
WLidC7Aiqh0ty8kPnftD55EpWqbG3aU23O3PfXHuF8u4pORxs3YYqJpJhktnbeZ5a5empIQ60Esk
MLM8ynTbAMV1rQd5dKkIghyei77LYiMHiTsORdk7TO7hJbBrS3czc/RJfRbUueO9rpVfre4GpZ3M
51Rq6O65zrWRzt+/zEEMpT7J1/+G5uk6hKFAbyerwVU9eu7+tdh/1X8ZkvZTcgjFv62paLeUWBU+
HuuM0fSkBe6vlzFrzkQyQrApCUee7xgALTXLX8arzCdOBDIaJiwfYLeApFPCkhsrhegg24glOrj7
cOsBPPfb5O/uVJdswj2IcmSAaipfKB6hX8XLfYR7JeOB+W0bb0CoBAWoeOBrak+set4huACpr9iH
kF5MfEh/Eh46WGyc23Vmlz+c+1+MnzsDCNgrHTCRiB3cyTahEaqEMfUebVLalCvXS3rDPXm78dGw
ArYVYtNbOROcFsrxw6F0I2qqIQbdjPTEcfaeyKsQpQqn60gLeO5f0ZrWnAH2miFsvtTETATIrvYr
niz45mzpNFBe4zilqjdSi6OdOzFnG94Wmt2mQzne/925KtwiUB1PFXpmplwt/w6OszUWYv7afReP
LSXC6+BHjDtdQRzWOyRYNugOvQxT/pJCnUw3MrkFESfN0Z7tUJDj0U7Ad8LUm7eO42ACPyMGiAHs
QMS6c2wPBV2fFisiARNC5baTrrs8b2FiK/lthihz1Frt97sUkyrnmmdnuarVS8PE/7CSlB4iPSZv
6PpE87KFTIA5+ai+FAQV9hNNK/3YUcUuypBKj5xryeWuuRqcJtha4EV7aSiZQHkLXryrE2IhKB7b
B8oHsm/vfACOkjpmet9OKH+PZYmqVfvLKBciHbH+R3OCvbrbZ6r+cE5qSLw9PU82IJ5XsngpkMro
iXAJPokq7YP571QzUboCd6mSU65mzJjlbt2C9nNAbkTTwCRtglSmUxW+N+zFvmSUYAnBrfvoGBsg
WU770BtiCY5q0dMxn+PePF7l8zJG7qWDfj3Mb8ZL+QN/OgQUqwB9fIqJt94+tl/sjrGnPyrgXlEm
++wPqfehpIuIddL1vmOpfigrLni4nU7UFcLl/P3BjxdampC8f+tsHbhBaaxaW51U0+PRtTRMmBRK
+pNoSrw3OMHdTLLMeqicYSDn3dC1LFVYupM9PyI3pQFzQweD89nQw3rXJ6GFOTgp1ZWaBFae+ItR
sGD8Xz4ohemt2UsgvFy4ibt7JSgcjmGumJPQVWWLjabIwSg+KTqz5DWOfHrtUhFQsE+1T5uzyfaq
KjHsACdE/XuRYUw/IA08hC06+yc6p8zK3xazKrqnHquhxahGTndXQFD8/n011dUDltWDtFAZRBxB
mfkVj5ZSFPWKyddoGgZFeWygz2xZqiwnCoqx23OohYkNMkr9rC3oZ8hTRcOTKSH666Xj2iIWDfJ/
xTYf8aOr3tmVfvO/QydOhdTdBMv52WAi8tCvMHTU6M7tZdfngPaT370c8hONhZHFcdPFm/gOHHdk
ciRBd4FHS/agkfGEITIJLH7GQBalthcMYDXVW7azIU8l0mnE0C5hN5HoaEKiNc9RPXUZdBtTCeSC
gCExW1P12N49+qkEfztOmQTTrGnj0eMhphL2FlOLud63HzwXJPJyxWgdQ7/+djrOgqA4ovRm8NHv
HCu6nlAraHsK3S0Oo4y/sMWy6yIJsXP8fUaZq3/7LtJcLiGF/D0CGDS3J5PZOjjdYcyyno37cRoh
PdUA+rU7TMCpPikUk1dNpOZENJHTYHHwirb0ECGIwFlTYiznLr6CfGX4qMWls7BcF+znBu2ZutR6
u6W80nk3cshkuJxbA6xjkchEWAe09tTrYqijACD+30I1ugPwBXrQWFIA/LEor4VQPV+sjY9TMjon
1N8mnJWjsBi10YiGV5iI7CHq/QkjR++r8mAwGpYewMjmyK0CJZi25HJwc43rAMQimiB1Cc2xut5g
hjZ08ZXAETXe/eMCttZoKjK5gbh7OUjA+v6ghPYf6xwJUOStyjapT5v1dg/s77ZqdM6m5Z5+w78H
CjTduuxa8wOsaatC5EYMSkDdYp/iruOKH8LwdvbheWGozbFTIOSl8Rh0c/Ptg/tibzKIKNHlB9xc
WG+L4uhokNlxPbwJnpLu1dx1h36nzwfrS831kMyw1jgjXKD6KMtJ9eYXPIEOIwUNGaQnAG1KoO3w
u+YmvIJVWoCkwll/s+ELqEioLS3V8A6S0Z3ldC644sy5nBTDeoug9F4grP7kRdHtLMdeEk+dxPMj
fhTPqldmzwbtxWCb0iTZoLhuCqf74Qk8HrWxI5MTOSwMOyySV236VnDaHeqeSqhQd3KQcxt0WMnO
SaK5siCk8R13obScKARW+lBnzMrb+rYXXLPLUtnOSMnZiPs1V+RpoqIERba3qWzHP8suTEdOm2g6
pn0oDaRZ91JFbGdt/wNPEAeEFWHgzRZ9xPLOgvtP9i7JLPMRUhYQtaWlWmvaozE/4c+zBTz3v86y
jitKA4Ekf1EsZ945/WH/9HmWAuQU2nRchEfie1lwg0yse8t+hwxIIPVP9QtB1KL5gk/uiq4PkrFl
9LoX7VZf3C+Ip4uAQzi+dIspxiJ73TgeszmqN00ln7wa1+UA5pZI1uyc9lT5TfYfpmFRQf5H0Un6
1uIQK0NWQ/Ts/UcHHpHrdg9jpzJxCwQQ5YHzJrIKrekPdhjTHB/uhvrCIsPSrqjrKIN/x/1eGxdz
DrhQAPC4SCqKWSVcgnWVnc2t2hC/HGc/9BCfcVfS0o+dvDsfIjythqk7N1FHqtJy1ttRxC9bR/Xg
jIj5stt8yKoueS3jduqzyXg6sCovOnf0akbNRxNCzt/1qW+kHDDYTR776tO+MrNOoc4L1QWpcH5v
ielTtuwu/tT7ZINejnojMw2qQZ0oRNrILU3uteiF+97CrL+TEo4LLeplDOnZnx88pBFaQIuf9Ogr
/sc32qkXbCMaGBj5J9SUHxGctRaoiF3m37sm4dfi/Tgm3K4DVyda7nVZkmcTUedLUirt9tjdaFDJ
2Gviv/E1sspt9H/YjWKtuwFMuzQizVHco76UOM5KTo6240ApxeJ1o4K5/zm9hLgNeGYN9QBIReLA
J7Fzk1Sr0vXN4AB3xoWE2RF6DdhuvU8+1dZBBcSt73Pp7XOddrbjOl7H/5C2xw3S60RpWUPeAtGh
bhQzLL3t4c2OpcY6qR4QK6ZZShvDNHgRrqOslv7nPyfGDBfP0Jf/e3dDuO7QVEFSHc0naDE3b90b
LwphlQ3wFNixZMeZtzo+258REFnuei9VlbtvGmzU/hL4JKmrEEWl8I9piYBocpweoTuz6+9+UBJO
rt8I5s+8Dm4IgLP51H5oZP6OhWZOcXR7b9gswVJa+s1gx8Sa4ju84m8VioCyr0taf2yWS8ysfwre
bXncjbPCPmy4Rt54UZDCrCieWhFNys/8bcH9NhnUyEtYc0EDFzr9vZMn/ffyyPxNVTWSwt51rt7Q
i3yOXTrX23hpzAusN60sIZgutNKzjANN+VAUG2lXyOB5Qiwt6i9L4vSoo4C41u+8PpLm3m9iYNCK
395q6PO9gtbrLspaEJPt9nHgeNTW5LDEwUa+JUnu15iXN8P14bDGJmeAZATHaGQDzQQdC9B3kqAl
lYsXyUbw/fscmdw7Zg+nWnXuj9ZxqN4RgeMANP467u8S8LFsCtsWGtegD6xeT+N6Hm9SW4DOMfOK
S+bArjh+ivTPDatoSZtRXq12pOOxr9ic5y+zknVDUNB5cRN5T02q0+cxisXUh2oLI+PbiRPik4C7
tFz7n5ojsFLTTZg6+h1k6vtHV7gqxIGh8h8p4vQpxYb/oEaXKPSSjSrtG6MLIOQaJ3mODNixXCnj
7oyrgGy9+1kxZnmpcPUegFFuS2+HJWMSTBmWmjd2rS62EWZDJs574tPfZErW4jK0cpSJe1sE59kv
rGDtIp6BI8iKFmqOlhzEmHYr101tiAxDvhmH2eCp3fTeC8awkTGtgAW1t87l0dtzLI9yB5EIrfY0
j5cXAVgm+mO9FTTywnIs2NBTt0tdnX+KJz5/bifcpfjaSn487tAvHempGfb4upbUcYBOzKCAI8MU
CVPsGmKEEGnyZueVozvrokUWWuSdBW72bNsfboRxNvCMnyA2uloe7KpMm/dfVJ0PYqpjCfHVwD7A
2TIvvyxNyNdcFgHlEgO4aw1dVgKjmMvKVRjb1FABFHE2MqetlTffZjRMAEao76Sg33Mme6Itd8Yi
EejO9IX/HmGEQYme/laG0PayZ3hi9jYiHOOQgxUOHHyWHcmuumI6kC447XIxtVkZUVYBnTMhe6HU
UVbwXhW3JCgV1QkIUwo3VoiT8xoPd/B/1mH+JFeWUjtrGcwWPeA2NmpzAq7KSZehhmE5bpG9gOPg
TtQNIdz5H+u1QlbIM7bz0s5nWsh7SF7p79oEZ6C90zHGb46A693Oh6lGQMAV0w+BYvGwMt5ovaGN
HFWrpyP84BuJQwNxKUU3Y+ChfaiMx7TQ4cYNH/2LsFOLuL/SQDCsQ1s0YMsy4KbHDMuwTzdvbIBh
mDjNNaGAJQfj92iAcvHkgWR9f5umHW+SexRpAJ37YnoFD+UndT3yZ3JHcOMrTV2zk5qN1+iNSa4h
TyWO1NH1U4/2ZZ4hzH9/t8ltnmNCqnN92eOtQQS5TdX12eYHvn1WZmU2xT+B3mFI+MHWt5owrhjR
oujyQZ4KjxhxUGYbjDwYCWSF7YuRzhzrUAG+O/0Gu1zSJCZoRsYx7h4A7J5n6GsnqAd1Y6K92MvA
7i5G/xLXF5l08xfBXhcwXklfpVKu0LdAp9tesPmmCtSFqQ35j7injU9enA+2YF8gZOvJGob3mHmJ
BUoavtFsDhjTHBNCwR8l9k2PlefhEhzgavB4l04xQuMZLOJRW9Og7pMyklpvz2pmRzOcXBWdAPeg
gL88wEW8g9TTx+kHuLqtlEIu/N4FrdLhojSc6OsGqG65aKy1SYaOyvEGcSQcWE04Yy7LuA/X/GCO
3jg7urYcY6st7wx8jUlAibxRc/ky18ZdqxCG7biskEpox9IT3rmhT6OyisXhlCJSS3O4e5hcfWkX
wr7S9jkJwWa3rjK5+npKJ6mlWB75kFrPtyqJAbkXwhgoUxwarRZ4pR3G+ABPL/kStjcWcTOokVSd
5AVQHYaSpb4TwNtK2gmZAOlLpPR4v8SUxqUfTwA2oZ4FHhjJcnzK/uPLHHFqHBi0yCR5Wa1q+SyC
kSJqPCWxr5ts2UEugFLTb0QflWZDjY7VhBggIDtSkURkRQOunbSGm4kSYoNNeziLU8DJy9zF2kFU
tysS3VSTHLonGgA6Dr4YdonFd5bRLQCIHqY8PtIeDWw6VNhzURD/We8vnWcLvTI0Id561yZaLBS/
yRp8kdYuiU0YjihmNK2PqHgJ+fCafiodtqoo6/LFJSHru9BgNJGE+YJ3R3QtLqqpdG5D6CuIcmnj
aVju/mW2iB2KISWERK9vQqP6lWyj0Jg7L0vQ+YhbCtiyJrKS6hsOd+BLlBbPIE2b0x9kYTcWH3qH
cKCsvGE/BMUwkRRdllnMMAJo4cH1wrGjOWoLXWub+brKTMkowTPuSRC8iL+bU4gTqs9F57i7zLtR
LcW0ZJ233kl1Lav4H2ztX0L8h7lBA6Z6eQ3f5j5oSviZup95LWrm/E+OMi/pycR1DkynYoSq4EEM
dy3BL1IZUjk2OP+MIQznyufgztLbdi3ZzyHlgku53/dGD1FF3UBXn0FE868CS0i+ZFdqjUDLaAD2
0S4HLzu9wfxr+1KDDI8LGT+IXVGmr/flf1Fzkd19jL9B5YOna/+t5Mh3BVRlGLaepHUiDceoveOa
QKlrZSsSGrwfaMB/0lndn62bKtCmIHSUtcSnUOLL0vbQkFqqArAp0/vcI+tl7HF9HVrOGh9Kz1VU
EEt3Lpr9jq/6GqLQyJ2jRBoi9gHuJ6XXz/q6ozF1x29oH69pL74hJ/SzgG9tTYZVMMw/Dz8KN7HT
XMXdwp2V4LK7Q4wKSXDQXQODILCfFp0Ns0Nul7B395KAqqq2TEEIHykLtIRlrS65wZsm3mA21D2a
cv7ZicXqQqBIGau2vixFLSShOYtWibSjCeZ2vMN/DZ6drmKZe/EU4Fdu1aVaNkNW0OKjr25S0FX0
sqdAEA7QjMGw2eL2PhDrOMUOxAf3A4+59+8qQHypjo7296xwAOH1fVVb8yJbp9Sd0nkuNh5mBeMZ
vkqTwYIP+RKjJP7D62jAPlAiPs5Z7hhxNV7gG8bzGHPpHaPPBWKVsohHkPIO9pcBZb6z76wG1jH1
7dZJ2OJ7roqjKJIqOgyxuX2LIE0AOP6VHnbOqwcGiL1kVxjd/odub7xfVLp8SXH/gaNbOZMDpMmk
PjR0H9D0oxeSdLVo/snjr2PriUxs7Cm2xytb/OQStPHDkpHKZ6JOXljkZg1QJfkRrD5w3MnCr5y3
y8qOYt59UROJr2lQBImxatZWSqCpwEUrSZG7BwvRyg0SZa5728Cho2gA3FI+SmW+Oaos7/nAceSH
0Ceqexa7nXUWnHhE94cqSMA7Vum3+WkN86LMOo3mv+DP+v6DJdq4IH+MeGzbiGHXSh3lQTOFglNr
ifWrjmQf0lzWmXbCaSinPUj9FzJcaSAdIlSlYC63FG/lf4fWqF9iVSsYSPFFk2VhrIE9bmluQlbL
WiO5FVoEoUJlrRd07llzxac2Ons6iIM2F8k/oeiES44X/YImpz8O6rvUIA5z+zpSAT5tHu1hk/x2
1G3ds24RoxrJmnDoJsHqWzUZckgVgRT4sFavxOSQNoGTPAoYgyBPCmZ+YZQmzMCYa9CJQgAAsMYs
VXqEz5CS4iAyXSl+PJc3V/zjw37IOjUmSg134+GlrG4hMzO/tAPefVS4lwR4RzWZ0d0o4qJaQogr
ZYWbE9meoS8xLrVV6tAwlb4LiumLF4XCPkLSXewVPwibuvOiI3CPPfLUxdRSEpb8TD90I0n+Aong
bPqlj2d9A0qf0xeCEJAkguKAUPQhjZhm9OLtKvzzr9KHMT0FF2P3FcrW4uRQX5/04hErferG4Szw
G8w/+EDcWj80ckn93RTsemcqlaaicJgbYpI92SNrRitE9Y2Cl8VUg1x4HaQjmte7GAKH7uurT6tG
ppCNLaSW0PAAGm3UCsRqq5p10Mv4ab/HIsLiqzAZttovtluLg8k5RvzHAuKj9IxGLUf7agQZoMg0
O+5tgBcHqpy4uy4kQs2a7F3mzQynd4KH85jynVR9zgcSPHI1z3Mrq1RQoQqVAEMcTQKsG3B7z/sG
3Mi3ZilrMQT9AgZBREDPoOVYFQg56Z+I2fulYpE/KGUNi4JhwCrrLZhH85IQ+99J616754xJiEKM
oJ0TBs4XzZWfxApWNOywgnLs/bjAk10eh5RmdFCTNx2/MKA1z6hUoOwXGAHCUy5ESBHeosPXF6qE
7qhOl2ALeAferQMfFwuqbNABv8H02l/252wmVB/3aHeUd+0mzL764CyQ8hJIkiOFBwKVoSAR6tEI
gjBDsc/ANqpUbVg5EvPlxDpBehp8l/+2EXX3ADqpZbBKpB8aYi1UQIVNxav+sejRElpEmznscDLN
p+tm9+4cVBeFyX5TVIc0+2JufrpgiBGnGVMbzRO1tpxyhRq2uqWO5aYdVWZadpDukoysEJvKAh50
Wp1Xj9TPPf0RLXgjeTxhp+65wpWBd6X24RJC9E5JGmI/XVAtO2/1eiJUJoM7Ay/4JyUtGwKL7rxZ
m8IFOZyvKLx4l0aAyCXYlJul0TZqOHolPO+K45AQF8/BbJ9MyDZ0FfAMeA7osjg9BS4WoQOC4CYH
vnQi6vQbGtVh83SSGLD0r+fl/IPLXYXh7fyOiQtNkUlOwVaHlVkhM02HzV74R9L6v2BOV2nMIfp4
kKwUNLHlpCKXIfKKrb8HauEACYydAndGDuSHfx4uxpQCw2FOdTeFzmKQRI/rP+3BUvsucEaf3+99
E++YLkuFqdlZunJgJ6ZvYez72+frYUpKtx0AcmlEVzM34e9VV/aAyxbZmwWWqadtOmBvsY59pJLd
NjsnsfEy5Nn3CE8m2ph7vau+y4IIIlgyHWxD5C6kbT51GAPx3Umq0Ac1W29fxeQXIME9J4tDF3Ez
/BPnnyADJzzf1vx8beR2QDVQytfJlMx8S/mBZ4slKprpEQvWmcp1Garj7BlwT1PBSpFV54RjmDIP
9Q0UyJ5xRIao4IwZzAry0RoIyx4aPvS/8gl4YA8MpgAxODz/5UB+xrD3feSx3aRsw3UslbJgWwex
SIfT+Kcw3M1naLFDcPaJ/q/FjKakdyT/TVLP0vlcY0ijXWExKdwwQ21AvNZ2lfxgMYS2Vw7JLlqq
ZZf1pDfu17gazXYC5gvPwtUPZr8kQv+SKvXUEzMxW9oJ1legc+BRDtOHYEtogzMfiuqQgp7AlIkI
w47Lyl0q9dFUmy8R5LHJq3Ki6n8Dk1X4ALgYVTcqzeJaiGq3gBCWoHHr496+AyZoHCc0iFWMx1Cv
gu1A3kJZzSPwGAaR8MnLC5JZh1yAiPivw0nywo83sr2S1sAbuKEfUb+MHz/OGERZnujWcBcIkMfK
XnyjVJYDz8gMZwAX9StGHJmF4lDUCEE0RnvhGFJG1Ep40t6EeJ0NhSyiNUlAH4vWVx74vd0dK6wt
Py1vqO2nYfOM+0nSr4ChlWM1RRxRPBfrKNtIEnlE8RO1M3ycpJ9GLoJcnOfXeKGdT+VDTwPWmw0S
VeLNCc1DvTOSdvrEDuD6ApKMo4/A5JnytE87Elz2YwMii6rntRl7a+exqHQ944SLFdCShAOi8fXb
ndMTFyljsO1MEeFOt5h1aW3pXneo1N+VFG3KsE2pfB/0xZteLJ/91Tfskdd2zWpK1+7zL7M6BV9i
+l3SgHjLRiTjzVrfvAZgN33rvjYe5mVVNfhIWaNwYhzVnFGFnXENGoFNftzwAmu82aXcSMjlYm8t
QphVYh+5twEMlTFV66qEcyQVtikZR7bc+urz7nn7Y0FRKHT1b4UDrme9cBByVn0muZYtD3Vr7F8B
PcXtE/P2uYGcwmVvyH/gX469TQdlwQQcTgMiRtzB1vIq8zTf8LB+aYCIAtPRY3BVXpmZc0dnrDbm
m5N2aTsH109QG+4PqE42mvZHt2JgiC0eAXCNxjTI/OqWmQmEgE+Y4htDyOXGoIGk22bsHQdYq8Z4
5oPHnmrl9gtjneFuIjrzc/q1zpzkJD77bNXhUchxcdG5bD5W4huFW7GCKVlTIEfQ9VQ7jSMrQsgU
DgV4KArR03qMaVyEJRPCFxI1vTwGUqzch7SBjx2Iwz7DcLL9xoStnDgAoqoGTUFRoZsGxoU98g/N
cmAYklQUd0iAK2iF8Z5Xgs2C+zYrnAUwAMpZ+786Aahplauoa2ncy1MRNUsvLYSutnQlqxT9Gc9j
ezLpp3IyGEFacAJ2U+i7Qe03aYnRLwcZYp1JtFk50rvfP/llujCfTDmcIs5aSj6zjXehrjGd4Ger
ZX4pybEnoMe9IsALYfNQziQBDKuOOrMeY40gTA5s3H0Xz81kH1Jf0R0ndCsC52+rZ8DNSFvxIDx5
i0+HXxtO9GthgAZ66MqK4CaE3ntrrTSfC0d+p21BbRv0MbQRRz/+i4Jz6bR+GQjrI5gS8Utrj+RL
8WCutUUHygOSb6IngX2IxtByi38qG+K617w+sm2VBCEJi3a1MvhSD5po0i21fT9pZ5TZNsNmSoMz
ZFgMCu1Dual0w7v7y4l6xIXy7zPRirA4oPgnWOilTq8NZwkQ0p5K0WcYNW2Iy3H7gTizDy2/vOKl
kbpvOHccuKTtTVO8G0VlL9bMMakUCewdxYePMB224mzeBzbPi35E4idN8v5gPJpemiL+vxeqD3C3
z0Zaf06P+VI5Dz4soez4bMmtHzX8cv/nKfsSRvmyM7r78S7SlLU082nNTFQwO0Q3D7HA20HKexIz
eG3uY9mRXndBvL9zfFuZcaclckx4AJE/4sMguE9Lb0kyE2WydhOflRg4R29Gg3dvhx3qocU02yZl
YGshsgybWqaKQk+ARAhdvTJY4lDXn4Ix9yWpT/vo7g7WR+pf1HHMLWl/FqZAKA4fOVXxyGFhgZ0g
xEnxPGO1CP7mRiq6DKAx5n1128xvnjxxzIFPyRhyBn8YnUJ+pK3r/6U2T7Vct8kfKOQWPAuVSn6h
h2xlrfQFrSvk7T70VR0+bn7+WdF+8tEpFYJqZvReUIc9RqFR3hyWaH/TwS8tNVkJbINuiHUPgobv
6disDF+9CWGTaZ0SYhkDqkXxvePW6N5erFlIX2ry15+SkSSb9oYbyHkVKpJxwn/r0xh9ZoBB7aka
21ceRkyBhDaWJa2vfIsW6Hy+lSNlIdaYGkdWhi3vkzae7fhEnBj3bxDC+ozvn7vUjAM3Om+Wvgfp
GrZloUn/Ygcm3rtgZuoqqTVdoiEiQWfF12SnT3b22tDHLvEv9poniVhHBWhi8Vp/Jwp7XK8K6yPx
LxyEkZb/hcO/SgJ+liVGuVUf2eFS97026mWN9fTVINboPK6tSe6nBeLyt04aUjK+9gEGuSZw7FvX
xAJ83TLdy1X9AQFActvQZIiBu53QJkDYXQHMEbVxmQ9wmRufTQK2vWYGSlVvpguz5OinvRaMGFRM
Q4GwKHq5XoNc9/VbFNolRBii1OHn3+TqOy6p7yA8GEu14q8BfbZ07KKFcdfb4vT5rfkW5pjE51Pk
MFd+DG/oE+V3Mv7NX6TwwhJhejYEBOOuETVywYxze6FYPtzOyuZ840pyC7rJt/2DE+hj7mMm9rJ5
tvZwHYCBUK1k8vL8x72a49wzTmlvPehnA0Tijt7Hwr20syqbZozCKgnZoc/IAqNCnI4UGWb/yKqG
3Giby1PxFEe6rFDZ4CZKRfTlyHTNh90Yl79gPSKwlsK4DjAdeXDgVtwBKGbGt4gZIOYbRgxHAAEn
3kMr7LwqIqL3xmOmdPTAfM8APKmQK0mvKfrtI65BGkI5nQaDwXdQ+RSMPMDQtFkuimoFilgyfAh1
sRd1Ow8gs15ZQvg8GxU1U+4l1XSxhM3Vnwg9z6uY1x2d+FbTDlzdzth+gj6a6Z+ktllp1UnU5wuf
79AtEomTQe+5/uq9BBzQMVF8lSi2eIcBVmUPS9iqQxHGfKCVhcnPj9NUb0vGK3J/0wBPevQYvPnl
8vcFAiaucCmVU+rrPvhQTeI61hRkMXuM1/xzJfLq93kv2iDLLkqhm+Rf5JRgj8e7nKTPocwMx7lV
LByhV7fyScZI5GundG7Nfo2AcXzugQovvgn5NoWeM/Fu0DUKKAEblL55WMU+cdSmZ7ZYU6q7eUQi
ByiWmTko/Of85JYCuMUaG7DTv3Lht7FspYEt2YKogmwbANTEZ4NKrI18IYKaiisMNWpr+ylqjEeX
FLI/9U1ItBuQ6PC1GLNmQYBCDggUN1GByp+eync9T2LSpbotw+EgCCJydDyQhObA7E8jLkG7a3NZ
CLEB9VUUtZaBWGwwwJGXWtiLcjVcy/gFjz8FSKv47UGHDhogHc9DmU/Z8tAFQLqQCzbAqNeQp4bl
gVLmJ3lr+ZqcpG0EQgCB1apokajPE4lcTIeVP6ghf/al6LmrfmEU1AlVre/AivwHPjJog4piS27y
uQG1uuHdLz5rM4xn6sybCGxTatWvqgIDZiowgI9hq6dTGNo4v/nHSbnOtmLlQTHfYU2cqd1Q/I68
5Sj0yh/M35Z2laFYOUYEChJX1dOAHdTU2qF5wsn3IFRKgXts5YvSdbLiapWIIl7+0w3bnoJRS8BC
mJTN+W7gmFgEkL9E+dw3lHHU5Yt6V5w2JKP14vGmQBTqNUAevvpLdxaehHZPe53MecNp9g7ylHNO
cYTx9z6M6F8YC6aOFElSb4iysQ7dR8LpBkCKJkbV0v7S6W/HDLcizqvUnRLeMzPThngtgoSNl37h
yrwxXSTCMb8Pu7M+d8yoGBrGrRSGYQTbR8ywyVzUXPRSYD7KXA1Kj3iBDXFFemhCNr1vziOKYes1
uFPNzHxCOTmK0puKWAB2f/y+fTT7VPSpWWUIZH/Wc5XgNpO8CBoFamephoYdLrbSIzvegD1XvBh5
TTcHh2YvNcAebdHbCA4MB/byiRfEXg+E8Cwgh/iitI3NJupA6if4pTeaDKJ5yzCAQgQ3xGiPpGve
wLpfWOZ/ZYkXEuwBjSGHKuiRSdKVDn/zPoMUyTK444EQdZ19qksX4RUmVw8Rpdo1Q3cmzZs1AmCz
MIKe0ovR8+lFGOtuCzbTCLxRpyEuIrc9zIEoXPMuy3jGGhRyb7W/VEpT+wSteEpiDmcNDIXIiX/F
qZeSW3HCrRoE6VyvEzFMlKmuMBmhrDELQgyL9l4qYja10eRZo8ott3PJz20pEpnvfEREIfGkksuh
AaraxFy8c3EUt/BLCKu5hLMOEHIMAoIfRdUE19TKcAMASeiFX2uXzV3Xi7gIVBuPcVXJo9aOWRpj
y7psl2DkuDZfSKmS9b8OYXXYUP1Vce+Vbo51VBOv8c1mK37f2bWJ7mTTlVi3R1IwoQJRFk3ox8ho
1FxJujfEWO/l/tncXrvgwaF8MFDYgLGFdCqfOLxMJ5h1R/CtLl5hD2XVQqMBI56NoVoNpwTJ8fUY
PIwfEfNPTyHY81vawu8Z9GTuGkwOhtHqP0GeQGdRf2mQC8oOrxK01gqmcV/ixsnmH9+WrmtEjbcs
Ou5faUAwD9+wKUBCNyNG7Hm8NMWuKg+sFLp8z16Lkxay5Riq8emZ4YJvoT+DpY2hRbIp/fqoXzG6
cTnfouEBXx1j55ZMt0y7PfPDhNu4NsCFn8VCjanwT/iEVvI9w28ieiAc0ned2e7xd1144KV/jHb5
RvJ8xi9sogBTRi0R8vVAeSxPkeX6rwiz4ROp4WYiCZN759MjfAEIw7zDffmdniAt2p2DRwr2pQfh
Ui5zERBKu46XXX8TDKf5PMGQ6sRWhdz4Q0YXxgKMXc8ZyKdez0NgIk09Hy15NQjZnJzDl4G19z27
95hCSIufdMjzGSJ3dVAO5IrWxZkNBJ9uo6GtXotwet1s0oRGPGOFD/e5p5oLSp68DM7D3okuacap
mr3vU+qZ7GW/2Mp4RV+iJQ7nZfxVYKwrBAwjrraazwsOpNcGFqZkYe9gskaUNv9w15ONNIz+Zrwh
/2qlmAtuov2/CJJHG7leTD6eHN53W692R2M25lYPwgCSvrK57uwNNni9YjeMsVCS/37KkBbrRFke
BCRj6rtZW9qrqEJhSLu5hfVGmQ49wRKM7gJ8JJol4eNNjFEwF4JyrR/uwz7U5+fFQzBpAsdpmfNf
zs8SHJSxxLJnoT4TOB1kHLflhRQ+vXaVkKRkrbpYSjo7nLr57ExQKgYL4Vb54vrgHTdkLqNdzslJ
JN/2qbZA8YWOxBkq7uQJrdRhr1cqXjiz6QrPxDIYO4XPBMmTMC7NgCNxSUdiJX6UddcjDqKQNx2R
TeN9dBES5GiT9Zb23gr05p3uaR3GQjykcutuw7N6y7Bczq3ntUGI6RlQHf1HMnvey0nGg0Vc9tN5
CxO5DfeJqQ7Kd1HGRBNsd1ux+Xq1o/1LvoE+B+KPVW4YwOwPAaQxQp79pEHKNuPt5g9A1cgBq/Sp
baj350btBJkzV8m0HlWjxls4NhTdiXwW59M7cclURTQosdBwqHz9GsC6FhIVpt2zhkpv+g+b3yic
yfkQ+BuE0ab/kqy9X+npcfwlELp6YWPq4iZiGpP85CnrrPQk3FHDX2eJNa9DiojOKdoNCbEooSys
DXfUh/hsyBSVO4L8ksxGUbp642LwUxTbgCcBSLoP9v34ZC7o6dAPjQj1/T96RFa4BQXuNIWz1xz+
njNJtZVV3GGv77AsNwXQ9psrn9VN9Wh8e3BjlS+3nwq6CbsTXPs+2EJX0BUKN/hvv+3bCRnfxrq0
/F/yLe0km4sGXsZD0WkYX0fwkgj/51AZxDj/Gm+TupWDIkHtqXI4Nf6LsNL2eSeAEhqDEgudDk1n
FqnsJQV/E4k9PLc4RlF2G1lb07NnFhHc0G/yxglLXJX5VbeHSGSnfRoC+iOjI8+FX9hirN/qpKrI
hhG2VG0K0RaYk1Y/5MRuPgtOoHJI2/rHRZFMAZ8adl/VYb7q0AqshplOO6IE0kWzz2MpoJqyrgxP
P+2Ug5ck4KqVzJTvgup5DAVvRWSy5hZ+WxIRlEgKebA7/1etOYt/5vqYDmxipYYJPgKKAsfgnOmL
VpCXhLN7l6r2EK9rJTN/IWAlB+kYDcNGERrOwniBHwd+YSMb6HFNH4KcTpejnrZcNQq+e0I3NoUc
RmwHwpJzQkP7PZLDfovYd58aD8f3Mk+xxscPV/6b2h9Ng14bs7RynIi01ozTipRUPmGParfndGYS
Fk7/qAKhrtHLsjr9F3GRcsGxKAQqdH9ifReR8NLVBJpLLS+TYylErcc+uSg9gQ02e47d26PtYT4b
1OgjxBUZgUjJ4zwqbW597/clePkDIWLK8ke57cyGW96Qnbc/omRwnBycI5Y86NVHt8xwCKz80bCl
KB7N3dpJU/xnBAe4ye7j9zZZ9NzvRDEUSxq1ENNAmkquww6t39sguTwIsPoiJVhTiXePKsexBnE6
6QV0nfuZ/oJmnBLnC2BZn4AzmlVwMxvFjDX8Jd6j4NQmOZa7+amaZ/vvQZ7WU7UEw1Osr33wzBZO
UO3pzcgLYtU7VcisRuGFOfyH/BcUzAlmv0pxImX2s2dK4BzRxzr2awPt6QISZlV3zaOLsHDOOv0d
NplAaNTCuDcWpX/JhZTSUsYzAnJ5GXyMN1BLG0Ngw2YHFFmkHoDO0f6wkKt9DNkb85u64UYw8e1K
BGJwa+QHOVP76+Deh6WsPhn7pO0lZoPD4Fd8DxBL2rvuttpPrMka8jy/um0X4wzz8c4Qxlo8LGu6
OjHUaVcJXvOUP6xiGNC9G+6UlhBclx4yEq2TwDC7I3GJDnOWXgE5XUCkKl5JPJyBCtD7CIfBYg8X
0xZVUc+EWqAAF5+cO5BFkJbN1WQs9pCTeY+AqFJ54buhS7f9Pf8/qVNZ1wWRIplf/MXk7czWOGUS
+VE6dPFM8tEDOMtdkLozctXx7OePQzq0qTcY+SWBQTnlIP1wv2karuOghxS44xOj/expfZ8DZUmg
T9gYIAoXt1ktc+zifSzccZWmDAG7UoOvBxQs1igl0R1IUDt8GCYYYfAw0Aqo+t/L/NwVGBltPeHV
Ya/gTyJyW5rcCNEEbrwD05JvTZFzaSYx77eJWdrpGTUYnGca+JcyWPXhwkkb8Z+8Rs9x0mEAQQbn
LO0p6Xf9L1I/qu6DfkHRdZqQHDCELu+51ZnIs40s/9scd0yLMpP2ivEP8VNmekRgEKheXVFfivxy
tPCD9vEsTdbx4mpB/8/zARoPSLIK8hC5FZUpyMJ4opiMzHb+g0ba6O1WHKN5pkTItrtjqB8AoHgf
2hJEtAiS6xAJJnRvXVEfov8WlebRtFha8QKFI791tnbiD/dgual8woOhjWS2mXhe65lNXZpDaLge
K/q6VxpA3GOEPOsFyCPsHh7cK2iqgfZFlI5nmGZEYVwrXV2NkFN7tu/kQS8DuBXbIIjaWPo+FPV9
c1bLh/u3kpubzJdDbPPQI8SSX/Q2oANd1DwEr/wIIYTCwbJCnBAToJcRJuokvmkgWOo7mhRyeyei
ZKxE+gR/EeWYFEOXJT/MH3O7OMj+iPm335I5XtGZjli9j2RnIP6gA9gQmwQuUDF81HDQi4cgAWkE
i4FB2lcUiyWHAlkCIVlY6YGlieu9nOjsNhr7oKiKJJwCkII+2pf9/K3mw47vqzThf9rcQD8UC48y
eh77SU32Q0A9ij063mgE72spopjDpbmL9R4dHHOXGmShGm0jGkuxEGAqyX6jLckTIX+Us8x83LX/
vrdbibZLwzdVEXthBDxR8Qn2Fsf+GfYlEKRjzCbQqpUHQCcjQGZ4hhTyonKWGhOnMym+rsdXO18I
8d0U77FMg30M6ecqC94v1Hogq1cgwjJici92cNMMWbWEXUdeMtU3+bQMeBfMA1zAyLrysWCmc7WM
awDi7qqdJFzDcdl8UAoP8kSeDjVgRq7ACqq8zAg0azeaPSv506Zjrv3bQpFs3Tt+IPSlesuQM1Ng
vcbFi8gOpSAH4j/VQhLUtTVBxNGh5SwrTGhLIi566Tc65/VS5z9pfOHA3beOet5xg2NDgqeMdolj
z6gGfEiFQdLV0j81KNl0ETcksz+zyj/1J0Wx7gTvv5hKOephOeo2jO8p6RvicksP/ZqZkNxuu2Cd
Cmlf5mRbiTxQeh0A30xvpk9xvEBlvhewYQs5elilq0HRJAo9vvC+sQAOG3oRBT5bYdOZqBJlXwoa
lYqtZ2C5bFt3m2ncwnF0tNoQBQjM96mtyjDPGBoObrPYy5tRD2L2pPuJnBCb2mci9MvDU/2yidJr
392gtNY6yhnOPhUBHN8qDiC5tQrEope2/tmwQir3KwWadMJBqpIbvbQowjkbwWP9ZhM2hbs/2TxJ
+5L8Mo5f7/Ip++2uCRkKo5Eb8B5LwFTuu74zxZosYQOtSkcnO9Zq8pI2dxgjBPY759XyTru/QiNM
zTBlKKCLWokv8PJRS+Xl1MqXLaFEwiw6cPnaVWthynyzCSdXky0Lzf9wFFy3D01SV3tYadJfhDYk
BnlGPrULfSUnzrVukoa7uHjcqxPSBrZlfUHeXDVDRqIdyQ/ngxR6GW54VX/FF2CN4YySQl5wzxZ9
Y/RJnpqZHJIxvv+ytIFjkrqlBx8cjb8TrCnJVqXqRpBfUgCpIZN222DxAQzW44N3n+nt9/s2ESGD
WbxvZLcn3X2s8m+gYBbqMJyitZdC4ca1teTAW0vzoOwNFumP82UYc+Xp9uP61Y2XwvQZr1iTB8Vm
dUz3WK+jKwExTxuu71mOGiXDWRMH/inwm3EF71CpIts9IMSXwDQInfRpuRh67OWRnMWr66rpV6ll
5FjGl5xVpDdsL8fJSlK/80SVUs/kAU2DxZ8car57unl45+6rB+eju8Q9t1La6+6KIJYNxsm5hL48
Wm02zxP44aeFvHQTKPWs5hR5djCoegTfPxRWd9M3/M+1BnH8Fv5su/g8Oiz1CGBvO5x5Sbh6DGQe
cYVgwytUq+48zAbzjyFyVNYXHZQQKYuzfWnTIFankHtKxIU3FiEort+0u1dOXF7bGEkQmvEexkjJ
6M1H4pPldqStKHhVRWAqGygYkE7dW9Vlh3wpCY5YCEA4b5YcwzXNTRl7sUuD8kHsntFVRZnWtRf1
o4YZ+LcG6E3VyWVvGUYKOMnEQDMW+LcvcVXdCAFw4O+Pq+9yrrbkKS9EDFsVhVtEyo5XdXQ/uixa
EJDdBpyfMT1mi8amHmfLz2ws8FySjXfynuHrf2DB3KKcXlxn9038d2wtMaAWrXj8Kz+4Vx3Q2QFa
vhMQNSrGLSbHjPNbTGMgc4p5JOfVZbyjBo8G3LPxkbH9DCubNDE3tQaiG/ItBuN5dtAETPTZa3Ig
fubvJO4PBn6KzdfT7CkwiIHSi8gPSsoWZ8BPqrWdXF6j+Cu1wGl22RGj527dczuEywFs9L1TY1Xi
UVkRWh4HabEdJWMDKe6Z+BduPrqemIpcf+ROtvn5ECCEXHe12a6W/aC9ngqZdZA5ZpLWzKE0Ct4C
Q4FIskC+27z8o4pVSGJAKX4AMUUJhllEJwd3Hs/oyVXLrhCN/Y+eyU42kKWyzuM5eSvaWsw7deuA
uhCZXUasOhMzPQpPSh0bSgPFah73PIkt8BeaRSTXJuB+XO7jqeNRtWO+pd/OL7yFifaXH3bRgh6c
IocGCHt2kRsMBdZZhYmNaHyTLAdCxBnohT+bx9DucJOF8dwQnDdh8LzCw7qfwJTq36E6V1fIiAyy
0ar3u96AwXO1tD/VfeQgV8e3QMVBbLZpYNLAHHObFOdO+GmIGXh/tA1Wm+Xri3PrdcBABTlxZT2f
H0AhiOFfrLXkfok1jEpE5YErqUIPsv1eWH85jhn5ZxWoM/8yewctYx3oUoGeLc+QnV4mHVLab8QE
eryxBrhxT8TNSKpmUMJuL/gHPay/8k3tfg0eU2JL0kOLYQUiX5T2vUXZxTcbJN4qmTMstaLPNwp3
i7076IPg8Z6DzjpKvKLwLJ36R2SYADlCKKlxXYpvMRcVdFQfOb0kH6niRMQd6Lb9DO9Z2vsqQc0L
s0oHG16W+1AcBn4fl04gVhQ8asVrFr7KIQBQPoR3g2lsIgCZrRjylk3DC/iD+JJPBoonQHHcA80j
UTpxZPVq4PHrTJWZZzcXz5VbuWhNSQ0++HRUmlUBBamJ0FsZGegd96MFo6P9CuVgn4fZhNkegDtg
jpsNzG15axYhEY6IYkuICqLQU7h9Mr3zJBI8hvZAsONGzJFNLaVVBMUj2q8XrKlia2n8FDO22KcW
atIXYl6kzipnJNk6QtYL5PJ7T1vxGC8GMI1E0GtrmF+Uzhc/7X9IqQ4z9A3Xz8BpSBlDRmdRgI/r
1Tdbd2bxqtFJZ5aY6kFqMR74h8wAze7aRr4qVTbAru4hClgSUAznXbLyKW+l5h8HPgbZg7aiDikj
2XAGNGpbNd95SLHs6IBjs3yd0bPQMS73fFaXcELKi7StfgOZMAoZX/gdgoubYZl3i1jJUeZ9lAEQ
gFt2d5H5old4bskBs0VbE7oReqv5ny32dfXGfdeAJ8gKmMdo1q7PkLD4ZeMpm9eKN35Ltqgv5t0p
OhHDWjDDy1AZu5JPMeFAEzWpVxh8TQoHOQ6QyXU9YIixHdwREXzgWIpE6Rus8O8/e8BykhMSi/k6
kwltUJbHzfi+p8Y5QGobvv8YlUYPxvfeWpER+Pv9L4MN/xB+RFhC5x43RavGrWMj63KPThBRRGsO
N2TPpw0uTvGfearU88Pmp+RompYEJop7n8u1saP9URcza4s6lCnfKn2dtAd6NvcMNw1e34lWE6H8
PJKwz2HPmE+aAv0ZwphabXs6grS/13TqdnzRB3XytlLSOAM1Xx4Hxv6slZf5cqvq53WvJEymTlJ8
+LEt35VsTu/o4vCMiHohqfroJ836w177CcjExtQ9fs0QCb8ncj+BiSP0s4Xb4wbRxYXzqXq3Z+pI
dOyfYZ0Jl15M6s6+bITPshePEFF22Km3Q/EdRWGkJpuV8Qkm3YvsUhoyFU6N9C7ndNQIyJhhFI4h
WSKRYBdCXCyi9p6HIcSgbbq0mp6KhsFouGP0H4mqn8dWg9Rt2UgtvRjl+VzFKM7xMKccqw+9L4pm
MdPjMTSynaY6PJilp0635mttEkKP+v8KEeF5dPIOLzMXHrNyPpL1TODx0rHgSszx48ZE0PG5Noiy
fdtVD4HTxQ7HJvh08f/xnbHkbEjTpP3KU9fhssK+gtp0FeIOZoEiqWrwqPHMzEbQkVn18qsj1eks
o98gjqWTYcOYbzpS0ab3E5odGDbCMEo+9aQmmNIw16kW2fcy0jBw4c2isyXrQdi/Vn9xO3Ozf5jr
K1H58R/r1yjgtJ0YzrMWkMT7c6KyRPz0vvli3ydYJjrMjayIH+ePCrQdrJsW/J3CEAVCUxy5Ij2W
MPMt4XBmybpQrDjMmTIVDOHWOIYvJ87SSV+CSkp+NKcTSyZp5CsR+Zud+oulG0v2ln4vhdwr/ed6
97poy/dZ0vEEDg+9wuAEl2jSnlcCpaOcIKn3zFY8IgR/UytS9Ic3QCJuO5gd/hUQrErZopCfCUox
USvXA5lQN1BXnXk26t/PyTiwcKHpk0l7oR/JijH7pODqUPyeBtStTKKTyvpZrywMBgga/pBBk/LU
+MTGkY0r8NMbn3zVsAOy/yCK9A/8J6WQk1Q+OXxzxYWf7xL80NCR0lK4sIKlT5XZgPkyCcEE3/NE
PqVdqYKLODSNcakaC+Z7A/bfDm8h8z2mmFv50TJtf+YIBXHTJ4vBQwaXNOQ2xPgaWdg+IXyaJpOM
iGCCWnCNhiRGCZEQ6szDNNkE7u5vV8wsrWbTQXUFoyeWFw/GGIoFheGiWpBbD9q3bndizPBq5DWf
z3yESiEKyfrNcYlwoRxSahF5JrnD5jVNjL7MKY/wFrbQ5sXUhYz3BjNzlE3Tn1dsdsW18oaVo7io
Vz9jStjW5ZZuG5Q2IyBeeoyuBVEx7MyM1cN8JqZ4iGKBtcT5miSXWN0YkOR2HglkF+hopmxuVtz1
MKe+6rPlp0BVwpSv7z3R2jStBAi/9e804CZEgSHp+aquxvPnVAXxTM9jg0vkMUidE48+pSgGNWEi
HgXHwVb+xjnYACCvMFdFctRbUjUVKST4NGgy27dC248ElKiDEpFo+QnWeHSw0Qjo+WntzMqbcSNU
fsnAZUFEeOJc/2Cw+P5eJeWlZHTlLodQDyx6li99LciuTq13wttZyUWj01RDFwPhQmFlG6ku4sbV
BqPLTC+lwZlMUgyrYORudrUQS5H2/dv02r6/TZHidV5g59L8bq+3udGwo/HIq7Pg8R+EuMMS/5qw
PfiJr2Nq7L2UMvIZbczArF60wUBbkvJKsVe7mOyDWONlkp9Qf3MM4213+HcOeBprVotpNDBFAPQ2
ZZ9sySdaKz6tTWznqfFUeODEH3+fOauM1S2yQteNVM/WtuW3dpZgLcsbQAb4Cxj8zMirx4wIxtF4
SoqljiIPKYif1esdqv/W7tnmnyhPP+PKSEoxkYgNwYIEN2ndranXDjyDklmKvMmhJLmZ4lv2ot7g
BqXQ18Qnop/ieQeMSsoXUT8IWUa3OsNkl9VO0rjJw3mRjFd5r/OoK4N1Zc7REGfh1atd52zE7SS8
Z9QOGQAuV1LA6CZnlVIdo3zfZY4H4/4+6rb9x3Bklf+gMnzNgSjN4iWufIb31MO1oTkeb4lMVG14
0CjmXeBNDGUlakJSJ9VYr6YExCHMxPVRtx7QG4NQ7/7xHFpPtZLaiAkgx1PSm/GK0RViETRouI8T
FCg17w9x/UX4JpEnFi/N3FUgMydxjSwUn/CF/rWn+6Eq1t7PTW3v8W2y4faoMZENDjfDjyeM3kNV
cx5pZRSEZOjscooSGRoj8PYm54DRnegp85POW+dQ36Z8tljI2qjcYRCQzboJdy1A3Y+OYUsjoYR4
GQUlqEAOAerRUhwQmWJnqxrjJFA6RR2Ww8AiVFxUOXOp2B4FNC8H2wfP74w8Y3JMseHeOgCMkmFh
B9A6/NWxZs9Z0iJ7QjA7J0PGN1nJZHe3bNO9DQ2lbrwAZh0L712XbTouwPGLVnPJYtSrF649LoQu
tif3XgYb7IWfeDPCxE9FBjjvvwzyeEw24JlsEiaRED/SViMcMo90K7lS47TTJjcdkJvBsWOfIi3r
ZfSmSTtrgkB+TL7tiMi1afBAzwiM3XP2OAky+aS1Et/dcQyR5yUososIXFqkvDmXxdNYE6/4u9xt
2DNurjk0c1EPkYWcbgrEZWzvN4+UVw5xdRlVN9ASQa1wyCfPlSfewCqx086uRUVFJ1NBEGrJXbD6
TLR7JOJXCQPC1JB0WZQ5yRoFVciSJ3vhiiTgunoDnuVjSLhIhlSBPjSlq0TQRsyP21vuc0iYCz1M
tvmmr/xh74M2w4PrLO0fBQB8SA/jQ2R2GjV2ldecXm8tSJeryHdSdFM0AMmzvq3Zua9CCbRLr9d1
eBCtLvQZNPVQNX0A+JRf8GIoAwGEEk+3S35cy0N+Z69kFRZV+Xl2hJl5pZKGFFFYKJ9hnbX/eBdq
fsu2zQn+Po5g7/TugZjtFZprBtN2zbmehzzs7g4cuC6cdzj71R3LDJL1/5DzRuzhtbK55w5/5gHP
ZhRItS5SOkhWIpZbKssNfq97C9aaXLtKynymmI6q34TPZwfrJnx3H65rhcwIrWTQ88xK+wG8CG/E
NVDLFH4mQfkrqaM8Yf87SScRawTisRzc6URhG3WeP1tk5h8ldodvNwm5GrAsEtUPSb2ceSqlrCy/
Q4HsZSc6g96M9CSt/yiclnic4vbOqCi6OBnJj8a6UN/8uBHfaTrN9Zj7D9qcpSpYwGyzJjo62XFc
YftI69c3XAqiJWGUxu01o2/jU4O5NMWCl+oMW10/05u94JeNXOQIyeybvLyaggqC+SVLnr34lOBq
cXZh93NvvwBOPbWUTjD0XmHGSO7q6znF5emZnWDoRQU6/j5YI5hNtV4RaD4WhN0aG4FmRK+tE0SG
ggBuPUhjaZXoF69QammBv9LW+gLSNDiD+p73b2bEiD/r73JN/YOuZwQ0M6UfYFbF0wxYePG8hB6v
sQYDeOyrZayIuFCs9f/+ghi/mJSW0Vy+Kq+zZqQuTBm6SLfgrhMPsca2q3LChSs7wbr2i1CmKr4H
0GRRz3rDqrdbs7BD1rLntsX7CtK60URIO7M/JrR2eJszS3wQLobiptcnBqwATQ6KaGTwKoP+KgzC
x6HpbGyOSEbrw029tJF09UZPtTJmpgGJZ0UwZNN975Wwg2Gb+81oHkptuXy2c3hvA4tlfHJju0ms
iUrxmTjm2W08Jwg0TGED7HG6iy3Y8UiTnwT91CIZR/mwg0l666ixIcSWnSCjYS0qyzLAEV1Q61Eq
OCAL0bKgolJhWzG4LblgeaLLQZKugl0oLEeZOVP6RUALka5k3pE8AdOce37aMhQEp81mJ9y0Gapq
MRZ7hKoRU2UCZbi62lY4giCpfrISgtgJtdQXWyUmzfUr1vREItTtpSjVoXVpmGNRC+zpS/9IvqZ7
YKtCn+ucsgRL2ngxxxIzLkufMPzOW9EQsUIBaFVhQRj/gI0622ijGRkeeAfDrRhwzLR7YfCG3QzZ
uSrVzce/jpps50I26E0zk9PGT7mFYQvj/6i21tT1KnlbMS0klFbZsPz0JMicfTmNo0eK5eg9hyko
6TaHrN18Fl/QHdGS17TioyXc7QH/yXnt86rTc2e3NanhLcLqusKJCQrQFEJwoLe58FdxelbeP4y3
5Mc+yw2BQkvCxQnngiFeSwEnObu+uv9W5Q1HRhDlDj9xZSFv4UoMTyKSHi6ctGT8sRBFSl0cClJG
ei6mH/HOnm74RmNvayz32Su346FPl1ILerdnkuN3G9sHUTxuN7BCMxG+Qh5ymmEhf4xvXW1iIURp
Sy0QhLUebHH5bPY5Na5Nlgpdtdd/yDoUW++3eUoOyRDvCeNHgMFxPK9U28l4hdmhPrb4cc2Z8I95
uzA5z8pPdEge5sAveFEcUwhdX9xUdvRgZQMqmpGv7pvQuqwoi1cK0WfXwXLOUcZs19zqFfMHKuXl
iy0HGOVRsiniWq+xkz6cdSwEtWFLljf5oR7kbVIwMPikf04BnEr4nyIdT43gkvJFWJRxAmaEXET3
gyqEYIddjZC+WQ/O8/nTM1um/ToX5dQHrQ2da4hCCP9yqKBvPt+UOh9RLKaHxgHHcBJyVpmZp0t3
pm6SZPirjZCypFijIy/v6nhhER4oSYuMC3SSJIxwmMAcKIkxc81xww93nQUqP0SUMvMdLq3LZEQT
Fc1k3NLGqsYCz1d3D82JO9vexRDncR/uMOV3bYPkFns6GETlSGuT8VXOuStiRBE+7imvh8eaRCja
Lq9kk9xMHrv/4qHtnUY3pgDEA+k+iWpJxuge1DlNju3NMuCSnlj6pIB/qOjRLBrz5ut8yRDDC898
kdLtfHl3JJvU6A14qOlEOuRoR9vlgRI7+lo2UWmDs019cVlia8gOYgoctSzwdr3kS3OGfo9lv954
KYzZgc9b3TWbIycK4YJzK0NI4Izd1u8UYmv6nBOtxIuIe/5TQAkYkC8wwXzsec7EGRxzAvrutSDf
fcv0riOiGprLKWy1cJacHW5TscbudcyGiWyalil3+m8ykYNK4MistU8AA0b35HlYiweF+SGJzZ5f
oLpdLYPGgbsEew7axkAaETXnH7kJVg+oV4R2GTKSebqWqv/OV4/FMRD+jo9qJxxP9AmNlpuNRG5y
NIQeGnNEXwHtBU2Uo8Z+rp+7GuRtslbec+8X3zFarZvahqjqvG7DlFxOgfpb3rs4DgXOb+NKVZ6u
6hrtSc7sewAqbUqFLAXkymHZva56tLNjjgy21wQK7GLtL2QAupjEaVsh+xqF+/IdMkaMI2fVl19H
OWV8j4Emh4ig8kQtfUzbllP5hwMqiH2CDIJB3a6M/bncak3uUn7I3z2pu7FkRZmc7NSl5X6BUrg4
hqiAjyCp/s+mx3RPuQmDYT+qPa//SHwyZkEu98epsZdE0FZ1bflZzfAz0OvTiiwCGLlfMM5xqz1y
NY/J9T0eXxfqbSqZtmJEtsKrZ/WnTrrqksY3nDPsZNEHGHITKgquGnVvpVztwFztmw7+4/X/F4bd
ULVenZOeD6KzRU22yiuI1mDy77u+Oh8I7a5MX7B4yKEo0/JBYxTJP/OmaeMcIXpBbfpjuQNvqlL7
naAT0oL0/JeONaEBWQnsswECFiR6QWCwCfKrDNm0DfCspWcRpToBFzrABJitnup/yAVpIQt9yM0S
+14Dd7tviwSQ2NiQZMQyuCSvDUnIG1PEU8E0RMDQB4ZZU5DPJBsbzenGAUYDNnRlh8Jdp2WUBrd2
Xxlg0hUqC3x3T3Mc19LWvZ1ad+7XRQS5l3dOhVPz43zgMrZtgyhpuhnkrgNCf3WOH6RPQZVzwlau
P+38WSHG8BbN8AKt/QjIKrZyoswLft7eCLNVcZOiTWN5i2NEWJvKl5ze9RRg4t7h5CCT6784Iuib
2BIvFTdqEPxHDs9HtPTJzsww0MqqVkddNTtJ3HHRbLszbwkK/+ZAlPkq/NEXIW625gB08kxHfzE0
Ut+9MD6TEAXZRJd8ATb4K06xdBtiK8fEh/NRWaf8S0FRTPos/PcHnLjyr8n+PoLEpttUMWUNucQ/
7WAxpNyV7ShWKZSoqMMyArRNosO50Vbo94crEtnJ492vq2DW8RS79MVUy1JSeIuDoAH1h+Pi3do5
UcgTKyR3tL5BIsol53vhcEVQ0sRdwwN7ZXWvBX9WPe3lhk0FGd1MxYcjWxD6ozv2FxkvYA8XrGDP
uDu/IL+DkJ/7VUo1f0I/g4jmuQc6hM5l9x1R463/vSxVbtz5tkhcMHV8f8YNUFrifvGWPFxJG5RZ
bve4/k8KXQ1pLml17inuhw9uE5de6n4seu55gMyzHZtcNL8JMChgxKIS8i9MVM1SAdduC9o33yJ9
03dbjYHvSEK2w20xCYrerg8+hCM8aO9+4UZ18niRGHhO9aSjgFqIsNuMuOuJKajFNobXRhHkwVsN
4OKB2GWST884pAoPATK/5gzm5O4djisJGuZg2ZH5WpGEUqKzQEwQDvTzDaPa5a7N1KJQVscm8s4p
ka9kt236gyZxDdoQ0BePaekgIHJlWERd1sCfhpK8B3lhwlTf9awpXp9mejD9RyVaZF2khNdimARs
p8n4NeRs7uUabqDtjDz8Vgv9CeYFu1xTOZX4XJAsiW0XNFCN1svBdZVyJmPquKWazus08hf/RPs+
K3urkktLQnKgfmdvYNP4GDcsceA0FxkF9k/DsuuuBNHZEIDTNo1g8E5zaU994cuV51+u9mw8RO+F
yk6dYQV157jRVNDQUuThEqX/LDwG9GzNA4qcmRm19xy2rRFt5rrN3351sHAvGlTVjjRs2nFnno6N
D6gy/S7xrYyIIwpdZIoU+UCJ9sIcQsJ7zj0pj/YMCVDEZoctZ2DzzP6njuYl4hFUpAjABJ1DAxq2
zvj+ryBhOFRiRr5Ic3JTt9zZJKv8SKpv9XaJXOyXrOy++ALJqJiLRuRZPVHBdulO83ZNT6e4q+0+
9IaG5QtiN81ZuF7UI4syIlHFmOn5YSCywyKxhR/rNoqZ3K2dLCDufEcDlD04NyJ+wE1lZWVuQyXR
Iu1ggVe+n6I2NWOYGqPi7lJpEwiRdcnyWqxRNxGjIpuraMfGxaOzcykbB7xyzAqqMasDM6CPyu36
yN0/bcFo3Ee3Xrm4ABRsJgPgupCykbxs+qPPIew2GttIUqzwHVKOJC92hNhPSEB/55Vgt1B5ioVZ
phxhWm80Uqci3lfGc8fUer1AkN7CGtOJJn77wd1SFISCdstaImRRHr4vNd9EW3MslzVwwNDOeJxR
4tDt9gyxKxWTxl+gHXV4STWBAZgHYSdrzFQwd9wDhhA1eNZnCeP3oHtRExutiTxz+dVHmDoJk9V6
i6Q01u3twI/V5S3xuPb6Rv9saTRCh4iravuSNmvWfa7d1GcFHbQN0K9afudpSisIWLHQa1jO4Nf2
USHB5v8z/YikJttGqohsGSAlAvfUi1Wfm5j4BsjHf1+Q9H83y2DqW25spPoukKBCZbS/FMQMHak3
m4OcA1ycbocWqb8OBuOxXzyshGhog5xE41Dix03XHwQbvrLjkIU+Q15fiMyVbLHBhnOXhUl5RmR/
ooLEWL9K+nvaPD0j2XW7Ijm39ZWDqb0w2zBEe4S2tjRs5tJjTaeBk7zsi6pSgsot6Am9rvO1jbmp
WxapGnMBeWgrqU1vBSCgILcyzTeZsTAk7yp/A+xbkS10nUUqB+PNP/L8QGakgJsd2JIj/hauMOCX
gtwsP+Fnh9ZxcZDMSYkGmaN317RYzaNa9QfjuRtsivUE2pEcUu1Z5KB9MJpZy8iId+b+ae35pAJv
a0WyedsyQsNP6bkCPyWEEh5bBTh6AI+IhMp3UM5kxv0l2xxdNIyjYUn1rmJiDVAL+FcJH5kkraDn
pMOEGr1pdMgqw7uAfctJAkaYHsjHeAu3pi1+GNhm4LpqTDSxtkyeN929+dczb7m3jB6nPZG7zzK3
gPHM0wr2a/IyK7skc9GhmITtUWYkh1WPGVouLsqIgVksjzuG82K5fMZGI5bdpertLToUpEm2cEGj
IIacrIfWa34gcygOZ7nuad2oZkHoWq8WPdk4daVmak/SObwn966Ygkr++iFUWpMgUcwLSdPJU9K/
O+R3Iu6LWJQiKMmPazm/LLRCkUyBeJmH9rmuCxCyk1TuEE+6xC7ynZu6tP/NyWvA64UsbeEJaekZ
N86VXixbx01L6Oor7OHlZuiV6XzdehPkHC/gtDNUnmaKNZi0xLxJ1HrD0QrHZT3zTzKdU+ZzHQFd
HX4P3g4kGS9W1XsvyLe4xaICPhjt0IVcvO2z/7H59XNE5wuBpbpu+z8Sf8Sdlj+2UO1kfZzwZrIC
Tj0NT+12OcfqIGO/XYosue1+GmpJFoPffX0JQpzVfPhSgDM0V03Ih83UC40ASIh33JF8b0+kDnFD
GaWY2hNoiwUPW5KDp2YDikNXIuXn34AQjOfZPBzAoxwdKaNhS01jeYoCuPMBd2HNBQ18SzG3bzss
C45Tr+I/DdFi2Ihjr9hSPG72NhzQ7m4QdDpLZ3BCrO7Vft8zr3CgAKBgdBHcyKMRLd0imUWDIH3O
WxeWrvo6KfLbD2Lu53BoQePSUdm8XhX9DQOu504GW7o81nMt8q74mqk8sUBaVi4iZT6vXIBXIArc
RDz/4R61E5canZffwIwBkD4ZkA4Tw0yQNZNCiDQDtUwy12TMRG73EtMHTh6wnncaaXWzoWKIbz0C
VetB4H/Q+AMknJGpcsBy7HzkHYtwE86mqruAtyjRQM8C4ns/N+qhE7B08K3hG8B4DTD3yNE1QAC9
r21Xtckzm7TpdyRf28KCO9arq1/bYaDt85w9kL5nehUUacotbBbs4MNTtYtY6ocotvuqe+FJyUdV
2Ayb1hXoVQRKE7e8OXVQeDpH1OxO5UY6oWzI5niDHsrSdLRQWbGBq9R36mGxZ7uTU5FChDbchohx
1htZsil83ENBJXp3gmaiTWaOIsZuAX4WM2PSsQBXnBe94EOoLhIJ5AgxUXs5ofe556/7ec1CWQE1
pmmoPEJ7TG1YA5sPgpwXonH4Jg68pe0BiGXNANFKzQMrSTPLLQPjXnoSeDsmrG3NaRmkJbCa7RVE
O1bg8mzrZv5EfXOooCh0ngESKT+mGz653e+nihvE1GNM5fZQBV+Ot3s7sgRO+jSDcxT8eZ2Gn5V+
wxHjgcxALMLBCFqrkSNbhVuHqLJP7QvS0u7jMzfE4hcOmKcEAuy/kyNN7drHWOGL3rddFdR2fBQl
fNeT8vTZxuNtUzUOZqLiBNfdopSal9q359sqHBETI2239jT3zPxg4ENXE16OTLX/ZLsS7ICZbohg
UD5/ErTRAHPDC4xYMGc5Oum4RYNRVa83tN5FV414dsw9rJLh9amSv1igK6/jd341sJq6REApxu21
4BBegvZBTqxNwcgF762bUrbZ5ujVrNIx57GP0UpS+47S9s8rOXeWfSMySKPefGyBBcV3i7psLJK6
7Wf0rEogzrYT94HOOdLFzrYhqSljPqgfln0RTpI/QpPh173/ZyPol6Xx5Yq+Q34C7TJ3ejaQJ03W
BVO3jX1SNXtj9IppISLR6jZ7LpXR9Uq+/sEGbuZTu02nPusKCB6sNMrvod10x4nOSBsEZ1WhmT5H
7aiNYo4Cw/ALi1uxWqNXY6ZGCn2nnUxpdJqB1EsLk8g/5Twx3CC0j7LlWvmEe/d+HHh+Kz5Qlr65
AIJMbcXMimfj7qP9+M7WDtAVdlRyyhSONraanvKYMV5N11MwHzKMH5tVEpg+vQNqDv23SyPH/8jc
J1vw6YFcrlQiQxV4ykXA2LpKGXq6ZYoj0FN5KEsIHz7qLgPCHvKSf2TgOTmBDA1PH5OhITBWeLEN
5ateO/8vkwr31yQzOuGZAiJiMwXBJ7DsT+Nc6owOLN25+sT/hRgpxyF7sw9ysj545DgPOraIf63J
8rfgp5hrIbYz3oUV9I02KUysFcl9FOCdTeQSdEc6FnkdjQcenFJ94eIzR89c7OOAUVN5LRYnpbgd
ZZ5j5dHsvMkeGguF+RV22e5iC5LY+1mjFVGn1yd9I/qvn3/TPzHsxxY14RUDoj1spPVX/20T9zxE
ztOkI9jRgeACQiMTIT74ULqxocaSQgiSUfiLaZbpb/Fb1nmBlKvSsAHCa1KXHjXq1K7e4VbGNxQs
ESFGjCFU931SfY0v/y7YekuTrq8RFordRunUHQNYYMvI4cCdy/iR1Pk0hrbeyKSUZv53TnSuLN7a
r/4001KO5ZWGptczRtqQZyQz2Beq4jdQbRV4nPWurdHvrINL53HeyFJArjxwGy6mQBwlJAwIY/jB
GjwtjGr+a9utho/ZJSwqRcdglf4ZGl+tHl5ZN8F9r460O562b4JqGO625QmszqzUL9MjxxdXp1dc
ld8UnJ3J8ZOSIpOKsEgRbkIiQisuBtzfLpI4p7UWCrCqJlxhw8iZHQnfhCEpzMX32RwpIR/2rbbd
q7BeTe7zP1lbS5E81q4AlWhrUYPBtejqXPtUbdYjaGG8Um+XYag8gZ4R+1W19q8coU61XmGUFEZu
zapys+rJIyJHcutqD4PlumqUaG/emld8CzKsx3vry3C8beBZaQ1XxSYhjgA5SwyICjW2yUwzS0fD
7kuKhUoaBhgvLq/9qBW5p485IWiFgxH/w43avVz4/5YP7W8kRKp4RJn6IYfENnam1DdFz1Yxv2qd
GQ5Ra4+2aIAPKHpvDtHlVswIgZPkWYNUGCvv1LaQ2Phb5b/Km1eLPEJ3Rwtx9dxz7WNSpazkPlCn
Png0pE92kgAXHAd5Q06HcoYQzEWGMUhneUw+6t7hHvv3B92fBQdgaC5c4DDDHfQn8Vo+iQyOmHOd
5y82MXRFI3BB+nEfV/qaXrWswWHBCFEL3o4LGSUTaBIm1oWTjsp3DUV9qDLzktHLtvNFLZ5U1txT
v52/2cxpne0N9adZRWZAFFdmfIQ9+gTDQx5T9C4oEPIwehEBu4K4jET07ZKKdzHRkFpZ/emUMGMi
C23F9mxnqzYPBA0omwnBRGwUYsuD3tOtKfaehKyA1VlqhdSq8b5IpwhaWC/k+fdPmJWhpvDa0OSG
XbnRqrgDIFz2QcvJo8O6v0ZDweR/1s4tKmIF8LswF5lUawXpwQjpsJsHs5Y3mCPLkdXLgzWw551y
VNO2ZCLti0R9RUfXwT1Gcc7HzzBR/cwz3Mnv7a48jwWGveubBHfs66bGm459tPbCfgK6JN2HVnRq
0gALQ8PNjWp0Mcz9wbUX8aX6OYlV+eX4WG45Sfsx8nuxBbCWSeroWIXQl9XzJrj06NqW3eqGRr2d
qq2PbUYC/7OVp61Oj+gk1P+B4hqgc5CJqsFedWZD15Y4mlhRHpTUYEFUtD1Fnbc33lEv6k9o77bL
8O2Rir/uo/uYryVZu0JGYtdNrMkjGw+mRnI4YFvhwK5uwN2nAXPvC1ByKs1yXlo1drSUFWgDeRSA
XQeoluxAePyVvRpLZ7GZp9lc1Y+32FjzBIQu7HK3e2Px91V9vs6+seYaLgcYnuBQz6wcqp9AG2j4
zvuuykf8F4+o1jEnti3VXFAuT81Lkui8GQJZ9tj7EryM9ht2KuEXq+nLOLVQIz//JTJjx81+jLUQ
UKWjl/YTJynaae785f07vZ+C8/AR2P53qNKo0IvY34yLxjJ/5U+v6En4x6Ay6jCxOFTI3VeHFDIK
Z4UEM2bgdpR/d+cDfwm8LLWwaes4WJiNgyDjLyaHOkcePj699NQp+THxsKcdGAPltWaayGlIeJ7b
uom7cPE9RqBc7Gp4SrfUXUDDl7xEynh7GT5XmuFvafXqt7rOkC3TpDschEftq4HnqdJesjkeSwPc
tpnEZcfEXR9iuR+a26+LRmdUhTOsmsz02WvnIj5GO9EiGqYIrsIDMCOLdwjB0tNXZtsTICkEQPEm
MN2bwGchIpHAIGPKSDy+FggZrJ7RaSbwo2lgo2jevY++boIxQaHxqHAUxmQzLF4Yt/bjK8p/l2kA
ntcVzP/KEiLVoPUWoYo0Zd55uaV8OzaecAt7lk6qQvpoNW3boxssyF0xLNcNkdmNy3cmxYPaW/TJ
xWivJoqCk51N0FGk8Ym5FfJcfVPTMRoKs7KVMBo2naJ9fPj5XW2t2Jn4X/d5SJJ/ftRV5n9FQIdP
aDEHyE1tX9pYvj7zU+Y9Y1aY1YF437uKZB0blQKmIpCXNRF4UKYRDKRaI0by89U6MxYYpzt/Q3s9
7hY0nE2ogWn9R8qw/rSYLtYfKdOWYAKSkmmIG2lTaAlzV/TGaM3JrL536WGZQkhWtR3I0IEKgsRz
T2MPXSscRy82eOevUHpHlLHV+l4IE08smX0dANc0Xye6kvEQrcTihjmtrqbxLA8ScNdnHZgfET0z
pltd6HbewT4K1WxvmV8DbSYXYcEdcd+aV7epob4hO4CPB08/3zc+U4JrzcyzlIyl6xPjYKN8Eb44
QzBv/ZF1PmA63LMiAybMOJTTh6GqutfmdHUf7FerHxe3lKXurGrkmuMsYc6tKiumiz79FqC18qHU
uXzU3S2oB94NmM7AhmgAZ0CnqLJKYnDP5fQT1UiB3Eyy57s8FmzbUnoZP7NKQpSbOkyV7YyoLNEh
jU4J1TmDeli0tmXUps+zRAbvsmbAiqcx9wOBStq0+ntMlBeTe0oX+33YOvya5Aijp2/wcQQOt5wC
2TcoOO9eMBRBz10eLJXxLKN8mTbGefIFMyLnRWmDxTZM9RddyMQ/Om+YXeXyXUj/QiUzEvZLiadz
dWsYMG0J+pVrOWkdFacbYK9a4lM69KEqEsbFsW6WJQ1A8Lvdry5auxsaa22bzjrpwppUGNXWNDLo
U0NLCbVxhqy2NVF0fQfOrFma1knLTeclaKxaw99DSzjvl0fXIDhzJJGJG/f6aaqah64m82Bbl07Q
3yvrU9J98LK7en0hMmVQjc2b9KdJjVdfP6HI/p6QY0BVnILxzbzo4vK1dRIr+Zfyc9aZA4fpNNRI
SZN1OGhIgjDReA/1iTUUvXwjxxr9suehhZGEVBU/UhKTwmBDJ8N1VO3C8DbsySCJIPIwHIy0g8qb
dT86J+GTtqgTg1v0493f5WlMTR6AJQlNJNA4/yyXCpstSItpXjGEt8EhaAjgHf7qhHHHqFOlx3OI
bPHhftYShszMQ5r8JMYHbbNSs5RRjm0ALcIrl4jEx9Wsj4HI0k6Uc/1mebyK/L8bTgiEkRgcHiZ8
cpBhAsvl3zk9W92SkwmEWDZaqyY7xHgWGjObb8cmJmmC0qbAeAJm+jJBei5kvEMMsGW3lNoe51Fi
QGqqvZ0sd/3zEQTvwozJAosEOVvntP4+eVncRnR04ri9nLlOFF4IpExPRmO+PtI/Le5MjtdiO74O
bjVzUGmmmgwff1kDutd25/XGPNPalt4Kgt6rw3lOmurg5phuBwLlg2AQa6Q8o2dmhpiLLZSFLJFE
Muwh/KOe82CtdD1Ei8jBLLfdim119PKK5JhYRQppvt7ljTNrZrzR+xffXgfBHWHiw2Mr4mKZQYtJ
1Vhaetv+XBYO/lT6c0JXi4G1Y9SkGkLEDeRNrXVQRZkuKd8y4BAjDGhiteJxYqStX0dOHesQaoGA
P8HS3oeeez3t6hki6R6wwzPjDxTMhA4lICT5aDgkoZR7YkuCTQJJLTFCtu5FgD88EbFv96gPfwEa
EFyJ/DZor5VmpGI/Wo/t3w87OqI8q1Rr7V8LX2bSVNVYllUC+kWScQ8wUX8B+uK92VCAlZVjjiGV
Fzc1vu5jv4JhdKvGvNsP1eS2gmEwWHh87NArKS9tS+AgNEX/9yCSa+mJyfLIYVuV+RD/+dkDI9Vg
GoPODoCVjUg9ZifQ7heEGOxBIasRb+DHnWQYfW1eQWCHif/OVj354l9UUAL5rc5DWA617rcXnlJv
5vpnJGPCqiNUyEa8Et+nzbhgNLMskIjunDA9qN8Z85yFdz18rXP/CbkYS9vohqe31ZrSFu0d9ibm
shnIwGSgY7PtOjUSt49B67ztgGnvkLozGVBHEg7jQQTDkWs7z7yXHxHW8i1vTvFl4p2elQksVfaX
Yd+IdondLZoYBRGdDkPjlOmcZFMxLsv2s1d8z7aPvsXkdzRitZpbucwvNTq6S9e7FWiBlz4Gh1Cj
QMVP+DT4YILnsLQ3LbA3DTzNegi2HVNJXOrUxdXtRj0C6+8gFln1eGTOUhX1gD0+FCZA2EqcAxlY
8CCGZvyZ4rDsM3cwovp+LUy33qpwRF9VG0uv7VB0YD6eRzeRQaj7VorEZPNPIrKaFx7y5ZGxya77
lqiZ8okoV7GUVPkqN/L3MMR2tqDqjRf/VG5+KI3T+Q7t0R4kqAtnY9qiCtl6xs01xdEbIOAM8tg5
vG5mHCW7c1aeQ5qtMuYCcuJxtaMsixPcALSWcUhJCaJZsxnqDRQC9oQj3DRohpY+IHq27LqUF3dJ
LmICgXJmfoUNSJab2OQixx1O9WnmJes8HDgez6VSIohKVQl7Q7Ul1mZYWYg/Oh80UL1O2ORiQ8uJ
2t5nLdeenYRyVxHKtztr2tAYm1En+DiVvQ72ZpNy7NDEDRNW3H6P5Ex7H9gfQmYDwZrWC1fju8eS
jRMFhdxDre59yIy/qxWMWoJEUPQcfDqnoXzX5e/uGKd5e2z7otqu3c7vuSlEwIOxYl2JaMjpBp9M
Fj0cxV1zV41D36NTpUNEnyELijlv+XuQrg+FYEd8Y0jMqgMPDURdvsuedMvufOBiOgYYYb/vu5r7
ff1c+fe4DFf3SHmBgyB+TUOqXxjKFaPSIcFpxKawvCjGzzw2jAwFwpPvDA+xgC8rYEI4D/fDMkHD
r40x1izXRAUC3bjtraaWcSynkhrBk/epktWQuV/NLKvc0GkxO1Lz2ttWqksgoxmkcVGU28CKWrqb
EaoUUkv+lXJi/xo9JTeoe7i4n/op03owBz4QMSLyuzNwd18Aq6ckVYOukg8IpdjVD8qqjTzarT7M
oBgLEWV6UhyEy9dEwlwxc7LpXkVIFCM7D8zwr19n/e+Fif2Y+oUOdGC/Nz4nkP0EZa+DK6cVeS5+
PoEXtvAX7EGpyetBBspsT8a2idcW1itVx6jCxqtFZ6H88aQpTKuilgZyezmZZZ8fIcJfhUExWHE5
IZG8Wmd8kThPbmARlF93eQ6n5ba3XBwDodZRtiwZWYtUmrvoVyh0Xwsqgazoid1/l0Ke25jEzg3D
iwFNEqUIZqPefHwTLduzihZmdrzL6vh9ax88X7ms++pT1D0f4yz8f9H5EqBezjB0U9CQMFkikTHS
EyYgo3g5TCaEZrdGg9hwshr0N7JOR8bf8TyG2xIXYkM9tbe1fS/IDeb4pYLtlPsPQ8YL9tbyREEA
CrEXrdUGRI4woIAUlb3ivHFkAADA9WG3eAjc9gbicOrGUZDsUi0LcOTiGeVz6V54xZ4737hMA0Ml
Q6NuAyBp3Z9/laXvzGk063pSk/dg176ADQq4tZ1u4qLCSbgEz0fakp/kmH2Fn0EsIG99fP9WEB1r
C6wvpaWQ8XEfuztBwpYJvcSdd2v21ze44SRpDjJg6cFvxVmc12RWJdhyz75kbxh2DZYOJ9vldGg+
ExJcFQruaQYc8Q7nzs+JlWf78KnVSwdl7teWsmYq70HwRIOcb3/4DdameQNHnNkKk0XKWINA1Dp6
QW5YRdNHZO7prmagI8YcI+Fy11J3kR+6lYgSdIxW+iDZmuu2mVuTUVrB0L6XvlFxhlieuNb/VUox
B+1zwfH3A93sYfu3Hp01NwnZ2gJ7J50cdHg/0E93w+l6oW0e354tStQRqCf5CwU1ltYYtoSHu0hD
TTeR12DwmzwZYe2S1HP+fFY7GaXdfk5huauzbpjMRheHw7R5qc+siEectU9qj4LXpAH6ywlTTlsW
2fWF04pCKD/2/q5c75K5VouchOSVxfmKqZeaAplc1wyvkB8qqCEATGJdGS8Ko6r31JF3DeZ7vgkR
V0jqBMeGiwjzRx2plQBG3rDV2g3JpbWJ+qQ3LYTENTkott8ZKIWC53ySEYselN18Fkrmepk/Fua+
Eo103imyZAhwYHxydXzZSPo2u+LtEJeP+SahvC/vG3Vv0km51iZwz/1UMwNYfHHcGb3kF7zsGHzO
gXpNAbEB0RAyHsqo766wsUbIN00JgqtPwPSZ2nJWg+kJ1BwyuK02c9amhAlF0Qxbt4LWylbF+zFG
DKCxK5ckpwpXRIhCoQw6iBZznavXlmJrTWlbhzmc+y5Ml/Q67viDSJM3AFx//sSP7siDWgaFReO4
AlDrTELj16C0vKadcfZhbMTQZdKJNnhBv13oul8Twc4qYNxPmzqnHrXuNjkyUAaCdVjVAJKxCRy7
3oPVu74DDX0wGhudzpmYM0Vvmf4hJT/B5cT0tZm9XiOUd2F5xXFzfn9o6EGur3GIDTKBOjCH8vJ8
vZfqMWgPYrqb7Ygy8tYjG/f/xmbn760/83i0FRT7dbpwEC2OKfS8v6xbumATvG6b+VjaStdvnVv3
UcBCXP+/wX8EhzRzFUd7oK836Z1E14FvzNjEfdabdskSvszgOCr0If/qxevWm+X0R/8GwEhkJagf
VChg60Bsp7kCjgXVY8CeOsaZHubqxwEG5orFafTHuV2XVoCA9Wn1MzZ21CoaNKVuSEgQk6IGxlMD
Ka8MxHO1OFTDKwoU077GGlZrh1+ea9JD3sZPVSU0aKKFd+eZmVLRr0zD6oSYwtWg0bu08T7pddSu
P3p+TbVRZvwZnSH/aS2gAI2zBpSP81QRUoZatT+3U1Hw4q+N+t9fUGkNRfcb+hqDVZxF7n5sr7gR
4wUqvRVRMjUyGhfrooTUQ3PqkMWjgkO38b1bBa+xycWgYA9bFLCWDcNVk6UEXTqqy2BA/tno8YoT
z5SA99Ap0/ECquapn/63SVfcHNgHacJi/vRkbiCiyVXWyqIgTT2aJv9iAhNfAjeWcYZZxSYf+aV1
p9vzcxihqBN4MIVy+1O7ZTG7iVpsGc/OaiZ6GYWsY9o66uAJrTL+LyaMCO6BFfyoHx74aD1/jiOp
/ucDuHkwShJ0ELrLIe5VTikxJeOxOv2ODjtp5oGi2noa5c60qSYAaJxh947qpiLGjuxZaZz+kSUv
SxdfjfbqiUTAxLMW0XTmUPt5CCJZq6vrDEdy8l2cA1MXu+hNm6D5YWelmfxB3Ww1slY1QDCtrdgu
WiRE2Ckf06dE/RhPwF0q9oXYx5jEvYHOKXfsQ8kps5uUL7hBMvkXBUk/BWNkgvnYzjLwB0z/bkzN
Bs/WrH4cuFnEc5nkngHV1iv5mrstP4nIxsxBqt6j8RTS5NeYW8bJr7ZXxPdd2L7q9nNgv/PfBQFI
n4zjP6H5T3Udl2ri2NAe/dJDvxYDsQr5J7BN1JRga+QIgiSYaNW8/UJCpDuyPeSBA3wivuBVAJDA
3ZoacuAnvc1e5Bc3907uf6gvguEvVxITzmSW5AlpwN2btJHngEwr4ZIBZr/giS/IT1db6ZZNaO9g
y3S7cXuU1L0DdkEpq3NxFjv42DbbuuQtrZlt4Fj1gd+7qRvZ+5Ee3hM/Yb+AIHQy8CHBeWD0JVew
EJK6OhZ+H+5UiLmj2PJjKwxH8h9AVZH/ZFZ92qASuXmXnzpqlVzNI8+qR5h1vgpJHhRY7DV7hnrG
4ZtD4ugn+GGAU1Xa/l4IS3xfHC0ADylNOOQYKIW2srr1mII7huHfV34dSGSvhZtchC1jVDOU/+HG
1j0YsSqV0HlXnYYrSGseXV780l3KZ7qeA/VvXe55LJ4GxXJIRBJBC/canuDiZlaRq6NKh+NDkSAy
JjJSGue4tnFBLsseU1hG3R6+B0D3psbWzYL/+NUoOIg8DOroJqvhCAIhDpSaMOQiZAd0GroLR6qv
SaNtlDroAVnjNghQ6pfVfepqC+WYsdqH1sMXR5U9IB3gRA8TwftIxyII3UZ/EWGAT9BDhqXAITWI
UhfV+xmjV63n7Y9KwDJ9/X/3WSGpqR3IUiUTdrzKh8+cLPBDI123MBPKCVKNfjjviP7aHn+QKQi5
k7u0D4Lt+haJ9fJhzM0rdxMsOtgrMXfoA7jiQO5iLELFpDbGajpJOCSyWC4L4NdLL7j1Ig6+yvwP
LYXj0InGMbEld40vY3+XB2bNgNRvNM6pPQucZAfhH2vu8eYenzKDLibtvCiBV3odyt4I5+HJWext
Iuck+M0QyOEiGluqXBFn5Wcdlu0XdR2L6LeG2cPoAkQQ1J2qk8j947QfYd1p+QSkgIdFzEks1jgL
qbmx9sh5Ku9+PlJRpc885rUQAp7xgmsj1u0MxsUpESC0TnErXeOxU7o8zSB+5iSOsNWYthmc5oT0
QJvjOJsMf4un2qRq8oL4hq4fZvzo3bjOePOA/DNfZfPJefvI2RKddhwMhNXaEc71x6+KOKL/Bx4B
WSpK+D+g0DrHBi7yFbWZjzniceBd2evJY9P8iycp6kHQFtZo1t1W3dl960FWWwZ5rNrIRkhjtLaY
+oiN1+XL2W+kkT+48xToPPRz3wD2tqF/WvlYK098pHIWrFu2BNY8n7OzMc/cN9g6MDDwHhLcX10d
e6H9s4rDDmFqbqY532O6Plq26ATyAZI8iuGiz8ZxCb6/QzR3Fkbe3wHKSYLj8nah63eGOzl22hS/
c3p3tq1K3D5AIEb+M5fInfmDQ4lzdPd8rizTv6MCUpZvUPozQheCp9K5FKjnVqgQS1xQL3l3iD/C
HsbYFnXiyFQFhyb763R1psdgXn9YzR/Gdi6URITsRlvJ8UsNpOLI44OrXLrAO5dGQJLmdzuDDSYj
2tQoeciKKipqecMRNA8Y1qlDIbhbGJeXA0G+Zh4e3NU7ypxa2QgGamAjWfhrM1HQMvKDxUND5k70
byefvenkiGkgmIuRNLcB2CCjemCg6sM+Gr3r3i7gDvzH0qDN/d+3FNEvt9VI8R4Xb9JVlLpYcMSd
1LI6TIyvTzDiQCyxdEaMxnC+E/zXroAbmh/TPuw+9nfWjowkw5Kk5bsqLqfyfrbde6HKTBDMHbJI
aJ8f5xR69yp31J5tns03XYfb+YBZutFfplHNZe+rvh6h1zyp1/FxZ+Ae7OwjQ8o11VOZVjPMoNaj
kYbyPelzQKWqulhCY3EDc3dT8K5KLLRbP+yZkLs28+Y+x02vLsn792w4IzAq541evHy9UamRBp32
ght01XswqD2jRzsuQxPsPJtANEhME+Z7e6G0Cd+R6eQIKkJc1bLUtjaEEbu0UikIFuukOi3JJL9b
GtYYoA5eTU52TIDTIXXZ+gEbu/1t96IVt8wUh9NIaxIP9HyClIOvH4bKmGjfcmCTnzzDBhjJCsy+
jviiUs1X4Y+ui2huWN9YQBuizpNHxcrBAJQyOaM4Ui0sCKnPEB1tZ8yUQvCx8GDd3NDIjZXaR8ix
KH3D3ibfx77Dm6l/Q/lkp7qN2h5zTXxCA3uv/EPTDZKAq7lya26lOk9ozLvUUI+u8zjLDXWGN3nO
IZ5pVz5u5+AycLzKXwXsdSJ7nBss+ErdLgcOpCjXuSEHwX+FIQ+vpt9COBp+tD9ztDsvXvKSMFlU
mGPi46NYaKOi0ECkxauCusmXor+GFSReaAQlNmWKR3Sh61AJT22jHO46xCTNlorPA8LZf3DEjeGI
Goq4dJQxIdmw1VlWGGNbZQJFt+yjxrYmPtILcQX0AkUzylR381gdb95EuBfTaXtvrBXIo3iBi3Ky
exOU+MfL9W7CCLJy6p6fBpAxcHyx1RRLgA3OG1jJad8ucj0ESOnyv48piyixVwZ4W3jI5u+MPlT/
Z8vJNLnjhxjkCzKMMDTNamceL44C8jSFZpWgFADkTRjr6XXglIHDnx9Xh9qBNBpAvMe1AZu9BOXK
/kSGsBmygvw/YK0I/Z3aybjC70n3U/LAOkH8vOhehyUfMqd4QuYEjPDSAC71auG4FApZUgLU3noN
JKdT+qOv/9rLMZMpMg1NODXFaxzvS9ujSXHPIkDw8KR6/CpK1tykr++Z16sqWI5Z2sKStTSYpBWy
21sEO5HnyVEly3WnmDK8DoXUScEWJ0NifV540JksnXpZ1+Y2EseU72JN4c2ohA3vFEJHyXSptPRX
IVIDi9S9TAnClRGpuCnzS7L7XLCHNGsb0OlphdC5k8p8+jVfdQbVQFCunddKut8sJYGB9kEYIdpO
d0ZvDrDMMbt2Aor8fbzaoQQuF3deqc2mGnYOht6Yr3bbncew3Zaug5pcnkm0sA1h6aNRSWaFKjGK
H+MfmNluOKyMILkhVK9QjVDF7TBhel3l4csY6E0p8WpgV4vximbT4qBLN36tjZE2Ao3hi+DuC0Xi
FsFznFP21ec9IiWyyreTd2r1/ye3WOd2oDUIe9e84Ff8hi4tpSKCLkDoThHzIHKAACQs3yFNqmyY
3gEm9MU3ou8pttOD2OYqF2IzASZ2EhEaXXzzng/xaPgkxorj5UiD/pubalcwEsP/fGsugk3sDgmZ
qeBZLDUjo8NmEFmPg/HZdK0G2T0DU2Wo6iD3i3l8l1kY9Hf2/qi+mIsngb4sJEFlTyOdBeLU+Yzv
fcVrmNzbMexPNP/B2HdIXFcXuXo/AK/+0BGKn+Zw36o2+KrqrsL1x3/gN5H9bWihlrcv75E8TL9j
nOjqOGbU+/OaTxULMMZc3MBoaFrCgNa3Bu3MB69izqwXUrt+XsvscEp9vs5oTj1AefXVpkqDPpoz
w2QQhQe88Zdrg9lLoFUkEEg3DNCs0BjmaiCpvavh4rIlG7rJCCjXzNVn6Z3B4Dmq9Aj7RCApCl0t
DuM0SyD3pL7uC6mersfOISqGxuyRd9XaBot0UsXdfsFzccMN5w2JqAPXSPcHjQVl5gIkNyAtkghw
5jUTMShKlU5R/tumSmDoS5vcl7RkR688MCFsDkTan2PEqDdZJO1BOzPsIWmZxl077JcUxPt/EUVY
7Omj5M8+7drM4Z8ooded6RtEvWQ7VyQi51VysLLFCDK6AGNJ1f5SRycFZpv7+DS/MgEFah4zDpWf
sYDggoIfm12zgFdIFeNwlALJFFKjCNXRh3UlN6gPPmYIiifuCIzrYGq8ol/Q5RiAa4lA1ypHWzcI
6PVhAXGg4Ip+xaUmSUZ4R+V3u5a+Wmp6qgtOh+6oqKFgvSzk5hxDxgIzGZgXk+mKoFsKXzPJYdGq
4u0ehR0kccLhfGSZdMavG8M2FsIJfkgpVJkQNdFdneE8NT62JgUkR5ibNVDX5t4k7nUjdKB7C+aQ
Ur8P2TLTHPkpJCUrjNhUNNf6cZazDEtdYAjdNs/58PT2XVuIMuLF8gra0sTbrYxEyyV+2PwmJmmQ
jJzmXJhgRoIVXiD+ATJUVn23QUKQxQSYNjSLjpO7yzW+mm+G3YX5YFYuHv/Yer9Gyi+ATiKhMq3c
VmxQUiR97e9OcX4Z7ZIJtHZQjxyXR0BvxsZ9bXEdXFV1XRYqcq7ogAkr+CGC/raXAEl4liVQP30M
8D3TbhqDiUcrasvO0HYD/XVcyWwVd0C1U+IHUCjcFYPHGZ0lMdqW8hBSj6028Z9akzCLIaXeXjss
Fbf9m9mGOjAMl4C+6lYtdBufqh4P/RvPDkoDAlZYIr/b/CL2nxfkDwXwK6ekTiMC5CMHIcXvMzL4
fukVzXkL5nW6uoH8TimWBK9ycG2tXamLOxQ7zWCyvLsdVUoMNJz9Oq8tUkyCvCp2Aau9mrmyqf/k
JZXYJ8zRsq5yZIzgTK7yXjTSGiGyPU0VnVefic+kzyKrb4ZE7goShH2bG3ONu4b4Toa+8ccMODTN
kzSXfgukMvhYGSeGgZclyRwwsJUtKxPpXrxVIi7wIyCudU+cUiEZzNhOrWjv103pfncLrOhFDexy
8Pm7grCGhJkTvHVFCSgCM1WtxIjWlsopQ0uSbNOm3Md/LF4b3wFs2Lz35oB88/R5/1ueyrYTIyKO
dwB/AJvhf7Rsj54CUtSyg1SfHeow+mNraJnTpagHFW9PvMF2yAeiZLDCtErfe3tmrTo+rldwJNAh
x3ztVd2LCFFD26kTvJuUmW3owoST+SrIsmZbC4ig1xQtx71OZD2ECPds7LdJEYf2c/KIRCcimgM1
s1svNSThLjOTE1gyo3XkOFcRUsnrknlq1A4HckEeq+0oMv1QKRu/cbhckDV4BCGh50jaWrmLpRcM
mxWaAehmis0BERIhJQVXed4bLI1mF4CrlDo1YW+bdOoTVEj1pRg8nxHo9MRbPNiYsz7ys3XqMsw9
nicBEA2L82SXgQrqq3p0C5OpbOLPrU/tAyn5+9+GhYsAsK2KUGopkDZaqEm/bZ6imx4DGbDgcedj
lyKHgFHH96NecBuldLoQoRYh6noha57O9Qe77uKX7DX2DAkxuomZ6ru7PDLI+gOVsKHDLdI03DNB
BYflKuTwbXrO+3o1MDSKx81G+Q6LUuFdhHKlbGTknc2siMR7R2lLygsi85Ti4Y7qvXM74u49QK4k
I1/vFepFQjlgZuKcjDNvr70e7IgPANM9E6Dz/9kzYDOSDvf7rd3V1LnTKtl5Cm2dOWv5s2KBhwfd
RQrc3NFVpEciRG0XsaVKCn8lJZByiMWHXoW/mdW120KFmEa5ngriHsIq0QzsCQWPC1P3EXDD+/jH
gxDFn0bjAWGpHIcRpqlF16U4iARUJ4b5YEiBzvHGLd8ByIxiLVILQgpH0/XaoIJa0vQLX2U2s/ri
TmVo/Jn3ry7dbHjtQwBwRyHFwBFisEq8e69/uIXoIun4VngH9Hxt6jcR319dKUUdgyr1cIooVopu
EWQxlje6h/PvB7g3Gc/zchZbMM+FHE1+oGTYdAu5MSAKSylbygM/jrsezvaEKC4eMLDaweI077Jv
vHQIGioIiu6TBeRwvv9q4d6AmESFiM1f0IxFgFsAQl+/3E64tp+PNZDbJbiQITAMiXD8TX2OQ5ag
FOSZ3iGTzEtn5sCkUA0XInESSTAtje0506Ny1hJAndqDgVgJrvrmEWhmv+CXGox5clIOHFUuEiVC
FesNLXtxF+H59wh0+jHLOKBwlxUTIwFPN/VQgfN0SgccaQvBFPzgdXE+Dmh1wvAM4ExIveAIZBc/
KUO+vWDEHhFKs3Oef8iG5rog0TTQ/u6kUejEDg2py03EEMSZPHqUTiM3tpnlXvCSp/lfmj353zs1
WuZZCns75PwaG0CIocZghBH677nYTRWek39rwwiaj+pmdWYaYkTs1yaFrmcxirpFTpY6jv66BhPE
UiN+Bym9CtBWfef6m5b0l752lTJkjnIXqUwO0v4OVMh/p8zpeFInSUkspsaftaGkKRZGyIicLRsu
bVEBFJHM3jaYdOf4H2U/SUb/oJxJ/WLQsfZVf3fZUmLsZQo+3ksdo/K8shskTohNarKAwCvA99UF
p7RcFVXhe1TzCiHxdFLpta8N3zOtI6vJY6hmvvWW4cCXsaTcv5M1GRrisKxEnWvMQw6ACF2AyQhP
XMwxUUQ3f7UVMMXOqfTgXb+tariLg4nXtTqe88xaRObb+6L8uCKj14bLsrhzl0i2WJHkxLdffio+
QsOL85uXvm09jAdoHKTbQhlvI3pVRy32AcYxDmW++ZaEAGPGvvrdziY61ZDdEvX04Dj1LGwBMUvE
STxhX+vI4G+Uf+j8moGNX1SN8tEP2ECzBW+9VzHjb6EZp1CiYiefqQ1MvD5Vt9mScQd6MtTfCX7g
GW8dNy30WYJCdFtQ3bErql0CneZXRBTtFRwqlWnnoh6hRbYOfeeqwNRupGmou2Y4ZGMA3yL0c6pG
w4za/gq+FQ+NCD0PFIOf7BJXzGrs23h4PqBANYstvDBguof6dWaKG53RNXwOnuJWlmBt27gWeBgR
xCMI+7p2r9ob970AIWVUplwOzNFTn/wLXHHLxNDP6vgWvAyEnU+SvtdUnSh3RZjyjCVkMNT14GmV
G98eAj3iGjH27aumFZV99LpIcnLkseN1x8j/5YjlpsZ240cHJznodlENLBx0XvtEch5TXoZWarjO
GCQndTN8A4fRUGYE0GLlhydvsbI8yBZY/Mrqqe5o+O+qYofxGus2fyN+D3KnkvLbZUgphppYuxE6
TF2GT3rhWmKeafebKYIbrI0u0nJZZbTnQvctYel5lvNgAu+sT++ZqgKSY4ORb2/v+El4JBmvpNPR
jcGxVpW/X6+nwygvhrTxZoC/Jl9GMOrHJMdROlhWRnxHuzIEOi9Qio8JzoKhdZjaZMF2uO6n0f+q
qKnD6WQKQ5YDJXzZ7MEMhOXrZE7dZr3TCo5O3BrEG2ySTH+BUNyfz/9xMCKQ9y6iwfeaEXhaT5Ja
QsbT+Nj06geWxDmOlGSvpmrUcay6xWerQk+edQMUhz92VujZ5OB9+qgCXH2RiApov2OdrDAFOWoA
Vne4/RbnRJ9fE+mxNH0mGuuComGEeYnZ90X8NjJiNk7p/Rxma2izeFbRf0J1GU1p1q8fvP/QyKwy
8/z1QTUxEKIZ5F+I4UDjXOxVMJvmD9xWTKkouYgKUcU7BEg75RCX9ncG6zhvY/ZTsathS8Uir08x
Gcp29vaAKTkw65i54ymJySdZSZIxr0MoA6DkURp91B8qBCkePIsBk1P4jH02LUtTydBSeKJL1Me4
Lz1acxyugLq9kpA3zSNJiro3H+Lb01a/1A4aRkIUxWRGrk9ZhVYlkmhFEFiy2ZxaduA6WuTd5zCD
3NLTI7VqAqibYW1CB2KBhqK3uimF6IbSlpoNW6OZn6PARc9A8lLOwn3k0w3uaPmCkitQhVaRrFW0
UtGbkJLz+hoTbXNImL4tlb2KKxgR7o/TYi9lH/hkJ+rAPkT4/KuebFcnm1MFPlA9idL+0CWQmIsA
BQo1g46zU3eshxv5HfByIVlZlG49d5H7W4w6R5Jg3d8C2fvLE3ac/ggMx/MMGER3cfo0sK/7x+P/
GXPxXugqp91+b81oJkKzpromLL5CZppZbAbFSD7+e9kBfL6Uk+B7zpUoGaQWss9G9Msp8Ydv8PZk
fYx/BhLzZaV0UaWxZgxxDOS62nxFOZRGiigsh94gZqcLiST8OogpTBJfngYaeU99yHT9Ky5oZVjM
/+SdCVQyKfQ+Gkq4cHugvPLsTiVKQmvXtw5SHAK5qcPpxIfyK8elaf0nBc8nSBwx+7efpue7C6Cc
LV3eVXrQg8IGvpkuSQHU9Yxmshi5cMaCOz0QoXhVJdv0K5jv8pVTYZEZLcMRqdwLXYPvaYE5+GuO
L2yUU24k7b0R6FXd6Y2xtJ1fqSWVIq+GkfURsybM4FDnET9bv24qTwSRFENLgNB+2UmoOE4iNecA
VdCUg3y7vUeq4ow9aO0qGQJwzPEmAQ3CbBvvACw0rHu30yHyWXqxGZVky8uxIpdRCTxmc9xads/u
aRq8zLMmUcga+Ncewb0v4eOa7gqWwFD+RZSIUaAVjuwnNbmORDHZI+BFwFFOVJ4ulAM+/LAkUabg
AxfcnxlsnN7/9KsKIuaLx9jDe8knX6DJpNCBG6XwwrwuEqiEZkwSxUTuaQqgnU2hS6TCwhL8Op9j
GoYvYd/CB8QRSshIsCDEqkYQbkaRXCRRlMtRgADlJ+W1Y9fdnZGx55lfrXFg8ZIBSoDfFhX5ziXs
Zr77Aetey46fuwE3Ej+nFgEZrEg9L0AJptaQfCcJ/ZOSiBdG44x5a/LNd/V3eJbBjQs0tlq55wve
nJp5C//F80MAKrgLW9ybl3cXs9q6YP0DCXOyexTGotr6ST/ZT0Uy+Zg/IskLYX3XYboQhcPSGsKV
9q7+fSXwdpwxSaqthAGEUhn4zI+7Zm4yBQ2C+ZyxW+wYHcEpfP+8izGeJI1sMy0Zgdt8PIa+lBpa
p6tdGvKroNMYg0zhKlcXcJz1rQ4+ZnnIUp3q3yRykfs60otPK4lD13cp384igGEC0ANZOqq+3O2C
1l5wVe5zP5BpQZOfNVQGKSYV2HJDFJOf0bRkf6BZYzsWe43DHC28pBpMLtt8bSR0uQJ35fUXedlW
7G98TSxi0e6HezM/cvm4PwN2wXId9WVQOS+Pg0wRjLbYAIcOKx08le5OKhEv6fbN10HAPr/6ykGC
jiyHXBhXYQ8Vgt1ZtPeR8b0jPItH5Z748zrc9Mp7U8K9+y6idZOwXYzZIoUlXk2GjoJisJkccayv
MHs1mh6RfSN7lb1KluaGhZZ/W1nGTs9670O7lnaTm4/A3OGQv2BX6hSYFNvnx1yoDftP7AKK+8sd
0TILZH+sO5z2j8QjQ1QEzumMKI8uiGNKc9hJPxyb27t1FPfRAppzV3SPK5cMxCgiEtrN3YaMZQsc
TR/Va/o7dR1ATvIXw79iR9rEri6ol615j0ageQnAXPAKFJT1Ehqe/7fox8XQeIDdp6AaK7VYWW1m
eOBSQekK6fj6XavJ2ARF958mY5fJDZCQUYtc5BeTUWvyx6WEcM+PXPPhyHUsqoBGbpuk8I4QYsLw
TBxX4kPkPJyxiOW2xisK3qkRMXhNecjrsnjg9Gp4KAL5e1aV6EFtlsTxrm9itumD/09y/pVhSBse
8L0yvaTBQvvdapEQLz4wnAHyCKPvBkSHk8px+oY6fB/r2wDWdGj6wC9oDrKfAEQH3IW4xHDE6SEg
lRRvRuSInWP7ymKWiz2KsVl3Lq71P4OHLbpXueExxl5FynRioi2DP97cxUCu5VWwHKDyr4iCKBSZ
lF6Q0qkHIYOe/yCi/rnWmsMBIGSPt42UhoBhJ8jRoY+FT/Vhj61NLskHMg5KXVJ3pBZ31vP46Zpv
evBaDl3UPdgAL4zr/vGPZuWNRVnbrcXSdesebDdQVwhK07PfIELH42VnoTsv34cKNcJt5H8TCask
W3pklV2idIEuO6peQYJ/sANnh65bVTrMh5rF1vWO3/mhVecK3TYsGFEqewUJRxtaWVflDMnfqQUH
TIXW1pdTPH509MkApAd8YiNxXhiUoxOG85uKvUdmRdBd+CRvD+lBUzkX8vf/oofJX8ebGbipTSYN
Sjns3zCYWXipQMpIf9S15LP/CK+O/+WWUsb4p6Iqi5Mrr4b5NbysaVoG8j2kgdzm2D4b0tbHXpWW
OLun51oeCQxOy7Lpm8GeRR2Udmzb13DWNEuhIm50oQuWnZX2ofxTOloI/QsRML6if8tMQD5m9Tji
K93ajzCBkOCGE3vgUpPvQF9TNFB93BCJjgSdfttE/x11kUESVpNcLNdk9LPtOH0/aEG7vrubwtAV
u6XQrFLc7nAo9EMWrJ1H92UiH70gjUipk076xIcS2/BeOo+4v2aadwI/C4Tx2dXnVl2hKhv11OjW
oJg+S4ka0dpFTssizSzlqUN94ELJ0odkVpN10aNkVa7sAnYw1GYRluz3scnc7mCq4g5lNpfM2T+u
mSBUDGQajy9AYCIh9PhMlFLZxYlYn49Xf6MdhWfL8WnE/65AYjVV6KkTD2Gi0/sb37AlKpzNxjne
zL4PI5VggiNa6JVrKb5zy/vQi8jOUbPYoBXGUIJPUClTjGcoyxMthLsyMyp4yfBrtkMu1BJajrsY
5QAibiWqk4a27PbQ0qXUm9tXyGnoqEeuWRXmkC7EW7d4reF6AQbtBcqQeqiezEReYa5xcD8uPH0k
9WycmtFr7h+AieGFCEHSixfbTf2bv5qImPaNYqIgIGTZ62dGTvnmj1Px4wB3WdZChDZbav5+kIm0
K8J/msm9840ismhQwOSpcZY4zyrJYeI9XkIC8fOlDOQD7C1E/WtvwkPrdW1RnUl8tBv+A5Lz134Q
Jcau3X54cY92u8k/lD1aW/02CAk6rlEZ69dqgrfEDZplmJ02QLXqOVrirp46pKbuSG9JjJ0W7PvW
6CaJZJeUfSsVCtph9zo8c6cckB330a4H6BXkRB6/t0Hh75EYvAbQaHXIyfYlIWfWJ2Iq72xn8l5T
gAWiraSiHM7dDjFP4WbkzyewOX1lPIhIHudi/GhTXBnI2pm1SL6/BsLolo1M7MYNpFnvKCs4PZoP
pmAG+qH1sGP+q3rjZ4e6yliqTG+KJTV4+fwsLiJev1tQGRyrLXQ3MDdy351nN9tg27wimJe4gffB
KGtTF80JYoSaH+nhPdiCPL+GgfU5lmksAUHyIydj1mmsL2UfGMe/k6W7Mreurz1jdofnDV/vIVF7
uKF33Qg33lgQunr97GxWYltxX1X41GkK5e2cRTZOlf89FopPj2E9AIU40MykzmeI8MUFcnss9Rvt
BsT4qVljK/4YoV4cfDI7PNMQCek1sHbe0d2CuX2klnZ+qwdVJQGML+45ydmIHGitFDuCApzIJ6eq
lYXka/mIJaHZIItcRYHqSz8xXMb+TD5/tTlNvy0oL2OEaW3xJMkpIjlez4UOD7N3uevbdjNFJcfj
UjMkXfmoh9FIHYC1YY2sBQ38+D7Aajag5zN5u5+bY6CjBwuNRID6Wi7kw5t7Xs3NZa05BSv1vtAe
IPoo0ke3+VHovitD5wlWXNkHqzUu30z8RN+9AriGLc+0ENC6mBRVg++N6dGkEs02slTwMkJ+1Zdv
Wnl6L3AHiz92JyV6x2OJp4iHN6EMTSjyXB2ze+KFKvCFKlG8aQ/aTSQX1lTRi2ZnSDA62/3Ah9vu
DnCqMHvcFcmAIAdENrqBEM981VqLo02UR83FAP2qI90OcJUVl1PnN3BftaUs7DZg3BCV2LAuDZHn
1LtDlLv9D3E0i9bHVyIP7ESbGiqJ2YNv4N+Ye4DG2Ig4uBoCO8tOPnlMjOK0nTbe3dpqfnSLz+PW
g9bcz7mRHullrKBehwyuaJY1AI5tsixLNKjxf0OmyAr1ZjuY9QUfYmMrKij35cxVJA+C2S9K797b
1Yo9I43pKexeUE2m63rsaCXBdlAwbFBrxQcR1PzbZb36H6cTbOlqXjTBXvKq+V30W0PV1nlt3mV6
RyBd+p9z3S7Mpm3QJSdrbgn8fkps4MrIIUsseBoAPweb+47Aedc4Ub7xC1fqmhaX9jP2QILiDV4j
2t1Ht6XyBx5XvL2N+ek5U0L9RyYyfTTsl5rZxcWEsO28syMxDzELq7wlTIkIGRd5y4MZ3QKckteu
6sx8PtxZ6h14+/vpx7+jV6bw3DKiuMxW0qDx93l9qIiHNeu+iOiMq31F0rRyEeq2M8tTeXoVjfY6
8gd1QwcqIALDaPfuktSOPbTZUzsGgwZJTKS97h9OXwY6g7+nltTrejg5gpVt0T5FVXRBevWElRRf
3VD4H2QNknHh6JJjE01Nrzm6ZhD///QJoRADpZjGp2rviQG/8fNrW9NhaCvXwGFqMTyRUrHgHGjI
5FIFXrB5UWucJqV1DFG78O8Amagqpo+oN8yBTT+/LPlvLcRxL3f/jWzaVOUp8ZIinA1A8uORy9CV
cUUseSq8obUVJwbTfz4Po/eSK+wKicHuCh7cPJFC0aeac1RDqYq4RGON4Q2CsIu60Mo7I+FwGhMc
x4sSawE8z4jAdjzAyXjBDtd2LgpwTow0Uxu01dIaKVFLaqlVXllL3/TIGLrHca+4nfjU4V5t7NPh
auxRObYa7mrscENsgdhtPir/i8CMbk+FJaew/KtBkAWBe2H0QDyhCpn1wnDRo8336PtG0Z/LAaH+
Bf8zKqVhIIPg4tzjr2zvLWovQR8XPctNJjpFOSFyTU5txcAQ217/gImGFIU71DmPNXJWvWrUUH10
TFlDZPjS9n7SvsgnqH3WX9brBHgIqLhS7XSvAxDfS/ikJLfN2AIru646/+DNXPxvDb83BlOzkBeR
oAcxfxpY1lDr/+xXj5Dh5zsfOLTd3wZ6Zmr9ArT0tDD7H4dqWoJj8X+uyRNOMZ0YjTDxVbV/MiWr
0cWTD+f3NvUPAS7htM4qvsUsyG+JDH11LrhqfvBEdCM0WMmsKTiyRrOWVT5lmFvPulspC163+uqW
T/Ve/BeAI/XB8jbnoAXbIeKRzjzXetEnAepMuGJ7xVliz0+L/3Rek1O24xnNysBksbQ6HWAfrAro
MTZbjjx3tID5lnrLp8t/me2DgcMAOQWNWUckp5NJDZ4xn5WPs3Wq5pPHjIgZollGRPO+jdMXlpr6
ZZxmDuLLV3waeWFhzid82cAGFmG6G7U6ueS8rh34uP/NLbKp85EuD79ibRKWnzBU/qoFJyxvNm9R
x7TGCdPX/xj7CUs7A0MEIwGT5XQfelHBffwc3GV/khDeGHnykeBTBlTjAi+PSBgUlvWrINC62NaL
aETFFSjsmBeOemC/bEpa4K+di1ND7t32thOjviaw+soJTqcQFS0T7VX6g6ozGdFnq9pTEzzHeMMD
2ti4VIsjTO64iHjgMwVplt+khKv21Nx+tgjc8hUmK4NM4309hJ5NoHfvXoD2oztdOulxOgOHm0fG
LNsX9jqxq6sJx2UbNiMQ8T4lCZTQxwohgj+Xdfy03SCdkm0v94+uPQSlBW/GRmn0b71uNB3TmqfW
ePKw2S0MtD1kBk5O6USy/3wsbIrXPukK/1f/DySQjApiJ1lXyo6mkOt/1rZS6cqIwO75G6l94dcD
21iJZwo1y74tH+CRkwYUTSH/MYzSh1XOAafTWP001vXlf0kmqnrRwdM4Qw06asskp3HuMKdSY5E0
EkcCykERd7EoERdzoHaUq9SSh2NkTkLKs4HQYwq0ORJyMYUsIfjPoA3ydFbV8VmPFP9iUMtOWRb2
5VmmF2HouA1exXHNj9KIl4SnevuECrGccfS9O4wtihDvZbOEcP7U4opHoirXgxbGXKnu/02uzu0R
JgSSgStHXCzDqQyxG1TVuZbQETU/DbuytT8oIGiI0x484zQM4AbPYvNaHfdLAq1vOHTUtJFBaPQi
lHsMp25rEEuN5pyu611QJyL2hrkG2LGK/7RYW+aMIkeve6Z0BTx2+ZjMNosGI9XvaZ62CdtCpBaM
Ut8xUmDZ0+fDUE4mHvCiY5CemYfdmYfarah9rLcknbotugDQlOQ/Zt+UyBJaYRsRtSJb7Jkrvvj1
vIGuf2woT995T4E5yeL3B1/pAOOLi333X1WlSqR2gz5MMkPa70cUbKBNmXyvRNUsl9NJaBKSg3EK
ndsjc+OTL0q5dzUQypiiiSCNyiY7uTKDcA2ZNbveEIiMMXPF3WYz/xY5GKKplXCQxlsPgcvV+d8S
oDmK52dzz0KcAUS8QnzZTb1I3vBGP5Nwg0X3wuABY3z9x4uSsgjbe24feMBSQce2KjaOF5v6Djz7
0erEqXbvGOoAeK6gsmQlqzRfNQr79LSMk5un5YPf+pqmVmjAxRUb1HyCOHUCfzu0UJXtImroLQSP
QW1VW0bkjgY+Psw6BnvXfRcqQmeMrilZJ9LVjhzd+1mq44Ehd9BQVfVT1qR5lxBHzufcvNTWHObp
hUn8XXF5AUYlhv9shC9cKOA+CKWRJnxwKqwnkdHtyv5Cvk+tSgjtZAeUsudcLccxllP6zsTtKehQ
tQSz5rjLtSL4PE2Fq5ztvjXlpOWckW9ReOLkkDvwBA2iJl856sJH/KTppnayn3lyXZheOjTaVHaK
IFbZAvwC/4q6YiqZwVQ4GZYYTjGVI1RpdHYtly2aDLjm9e4/3rjm/V5GeolI3Ktb/61fAL/qXdZ+
PLDFyzQU2jT87KAzTI/bCNoClG9Q/LIYDvmVGjYJrybvxZo7cJm+6WzOlDpqKFlvzKSJ5bAUlsbx
r0xBmM3NAUaHykEFJUrTmQrwtz+wc0rG1ecUCv/pkBMRwA/evAyD4SG9V/iDhzvGJiiJLKnFLkgb
O5bmbJj7xIxMqLxNcB4gCCa58sRLYkAG/8gnZQ9aKT5fVllSveXIl7g+FuDS2iqzAx3YfBBMdvPF
mF1sNuhFQz5d6w8JMvVdtJJvfvDbhf5D4/c8Z3w9H1yN9vEGhDgTdeOjExoP7SuRWjKFdKgUQdo3
Ogego+8S6hOjPHLIhqcdSrS9ZwbsSkK+gbR/0jjEr9dQuznuB7edySP9FLJjGc033Lhhwsy97xZF
jEJKYRbDC+LkgKjI6gASoJcgnud+S9+CnFK8iRdapmYW7WT+68+m9aLhQLBOpk9EcrBRblY2LOUy
m1hR7TsMJW9TS95lpfLLPV2aai3vJz8tv+JnU4inwWZmZ1zEFyeiTl2+hsVafJ3XPWT3eW5PY0TO
pMDPVra4kdluHWNonIAhsJsPJJqfNKzn+ddydg0HPqi+OGg1Ux58DxDfkjIE7/tokg288Gpph8TL
p3oaw/j3t4+eahFlJI/+c6dlNInX9riK8fkdOzQiVQeR8GItIoL3h2404LmyoK/DP7ie81j6Btuy
KzKbIfdiJByehjVFIKFN3P9PZfnr3orqxEIgseqnraJLl0viD5/2IznRVQm6y9/VFlSPI3Jq1iSS
Znlm8FuNxqjPCeyybtja0WUoRWarKWR7A08CBqY64fG0maiZDWnmPKeUwkKELuC/bBoTzU4j+lCf
y1JnWZj7lwyyOlQvGh3jILzjDIAETVK02F+VHGgK0Zh7kmZoKXsYtI4tKZsJKdZQEJMJAfdPfSBH
xpFhUt+tcOqKmM0BYu5daqRMd0TDeTtJQQoC9SeeDYS7q1QaSE386fyA84iYnJOPY8HzhL1PX9cJ
S1hyJSmMuiR2z/vloKVjkFJRWzFLCJX5JITyfTLk9VukeIFBnOXCvi40L88cXlBtbH+DTE2S8zl+
XUG9epRWq89iQNCaSWUbiBaT9HG/bbvwz/N47yQjAc7bIbN7fE24+akUlIxmfQN1CzD9KR1fCw5e
Ho0dhcKKAmfTfgz1Aymgq0A00kSyYkKFca/zThPmboOrQV7+H+lDlr/AiUAxyp5tf4U325JPlBo9
0DdS0x1cXgGQckC+4pWVVdsZawDH9BMIQDPry+bNiDGMSG+gAlYlx7WBRgRv13T4ryzxUxG8HTH+
qJgyDfgBvDMo0NI/nFWFkVD+zRWIA7pB/mtPBbj9D6EEq6UOb19tG7eWLeu0XDETvMM6Des9eqEA
3z1oK7ThDaUQfkRVYNUG9fkJEU7HA798eyB0GDcC04TnqCo//BU5ep/FFmMNlLtBaSH8CBmgqCes
i32mHXbRmdU3cTcWOne32hI6SKg/hE+m9Mhf92NcS8ZkIzALxFMU3klb1Q0OdFJDw49oIHLs7z3W
k/obdmOI2rbFNUsyiPcZ1IRjTDegUDvHp1ycXxicWRIiraCGeQ3L3Zsl8Q1ZS8iJtS4m5+bTXhvs
4q1rx926AXk4uLlUu2vAU4qOn59FlQ3EUc9bXYUvqBJyPUu0TZnkD4mCPfmS3LWcfcBDEGQ/Dgeh
UIViaseuqdh7Oec3q2jNUvkfQTzyRRGMXlE2JMBDR1bbH0bPyMH5xByZSb4JmRuOEZNs7dMrqTlP
mkoYjsMf+t3WYJWIwVcWMDcQvqqyXa94QmYPV14k74oQUSWNtNCoqCUYEQCRaAaobvgttgzKjYOz
sGLPQRadYSXT5mbe5ja0xT6glF7d3tmcwWYYyTwS7rFyXAU8Lhr2aff4lEj4mubki8XjVYimC1aO
Wri/ThPUl6fFJOBx8t4DMqkjFI8+E3DLsQuVz2OFKk8xkAB4OLn8c0JV3O0V/zitI0IR0cvpcXY6
RyHc0R9ZlypuCcUPpgm2/fupZzZgVCUWcdylJfGtYVE0ea+60r2x9vVwULpWOS/gvOEKLtFlSjJH
gxZno5cIvx+ysdSOUZjN1y6+z5KA3D4177crL00sVonC+QX+meE02zVemcjjqmH9j07SroziU3/+
AAK6xs0STWjG0swof74OhFT+D3DC8We4eRoA9W9ZL4n5nCjI4kvpIJsMxTMlmIqeLcwqIUel0ILU
P8AY8pJ540q9spRDnLIPuHaOadPo3f7lhjcjFZlJYrpLsVZaVhHOG9qPRoZzzqkPIBlsIr7VHOYs
rskVuspxmfk04QQ9Igl5/18Mmw0godHrmbDMkyvnwrdzc6Eo8hf+M3CxDmiekA1o1vaxC/T7irXd
cEQwkbr+mkg0SQC7BtkVeVi/8yYj5jLmyC8hsKtwm7bC25gcdz7o66s+D5/jty8RohbqULBOEaym
fGL+j/G+sI1HwzGqL5GPvtMtCVZdzRd1dbWjlDfo/znMECKD7o3RAAiK2Ry4ZeyasLTeY/XWOZZS
NfKP827Zt7Za8J1I7q56GnfqWFWS30QBO05TIA/lUGvgurImWX6zbR+moTl8wwmJF+2861NaJVC3
0Irr1TKvcoCF32r+IGBAlqgpPBuHZHDMz3Ltg17UpPL9/gFBa4yM2Mga2asQn5WfI3H0xYzKYYYK
mDru/+Q2IRiNhYZx6CzUI6IvyQ0TZJKwC+Tdb6aPBKBaWDzvZ9EsGiQd+ixRlsrVzxdom6ze21nS
mT3bYkR1hSH+B/meHw3pMxqUHAHGn/Bb4wwUu5JicwuBRq4s4Y2OP/izp3GUSfcjMqNATHTvls9b
6tjocEYxoFa75csB38mxGuanwH2mC7nksoGte47+fjON/cc7SjX88KpLu3AQKo5bY+Z3QSMNT2Xc
ozVHrnbUt7QcARFTLHGpJsui4DgQev3ykQI7J7ayaRn4k90emtMHj7dI8J+IYKRZhgLi5X3JGV0p
BsFh+GMhBjEIhNwe1jiEIi71SUk+RluX1cTlCsBkx8dK89zp8E5UJKf9buT/WBkSs6vIoTsFWkLz
P14kH0eTzKuThtoW9eEqokiT1BHd0ANBgIzAhfwDZl4ZRnEK2C/B1+uDlrzPikZDJ+0QMXC5bFDo
Jmb0j5FgGXUAig8EFpO+q2I6XNtT7Mii7fzhgRoSDSSp7L7nQiIR14L/nYcxbF3T9vNWFb5hOAWQ
r9yLKR0cFuGAgHdBensQUqJijVBGqtUlYBDBCLzRo5Oa0q32zzZ+O1HCPQCZhSqvaPoyzQ5ETOHU
1Yhsrv0gYyTDrfdWeojo9Snf1djMbQDg9Ayb+dZscyDmVE0SMXFELLDZYs8XabxFqtCMX7lsCAJz
mRCefUT27JH7zPSP4JMDQVzPtg9BA7bFyljb4kQSkLBu+KhNXwWqgnIFnRh0ZDgwQSggck22TbvA
A6eDOr6F0BCIEuV5bKvzy+pdR9OECvpTY3adTClc7OkkuztfhckAvANoAReuz+87P4h4CfcvZImA
P1W6PH+RtulQZze1ey/HY9lJMWKJiaWqWOXiQ1a2j+vcik0NCCuNYvEbgx6UGEZu2pTvEKMsBM8r
yzdffMLkICXig04Zw4/kmJM+7XI/XTBYv1AwSDROtJgM4G99FUpmLMEW6OCzEea8qgQbNoJrWgYt
DWe1EENbOhE3vhDEudj80fH2kahnrkxMHwL5FypgvMb0/8kAwoQd4QT2ES/78IWQMd++3BOELJlr
qDb0aTfyGBX5wmLkXb2ycsxoVSqFJJLgfgyyAFzX6l0YzFMlzINIIXzXaUKBehVpRFWheUphZ1ft
G2yp9NNP2VTwPUj8s6JwvpDKp4IE/UXkngMati4Nkd0VjHlmPZo5vWe/ZsJ4h/vTue6HXDDeBKdA
h19R7IJEpYIANwhEin/vTObq2JpJv5l5rN0R8LEUA/CyPE4cQTq/qHN7PP+jsMbtG6RsMdAXLfy9
MCabLUruFof56eu8PZ8aqkeP7AH8uTppS6n1goxR/V6yTcHfS7vBk1THEmVZqtQUzt5E+0rX9XJa
2CxtOXO4g8liqq1eM16trxpBcLQfSlbhaeIPDR6bkc5S5/79J7XrCf2QrTnYskhsqcbOgeKCx/oU
aL9dQfIor36ZH5ncMEUuCscP3+8p9XMqO7Sl3UOenMRn2TpJAnuqjXhsN/+sY6HspBlwwnRo5EH7
SfPHiulHLzg41sSgQ3Qv4t7CAQOi8o6nqQBrCwI7GIKc9QC6esKI02sBfrzwSOqu3N8xlfPIfDkM
cwi4F2w/ZOqXx5uN7AbXtmWNvHEff7fVV4tzeWM17CfGKhv0msjzlG6nLhaLgmi0ZE6nxWH/YDKJ
eoDn7AfT8dlCeQHaA/1/Gf0UcJQuji4zkBvXBZYEghx7yOHIA60TbO6FXFbzOEbpUlcO7YxttHDy
/PNtkSZhv0qQVNrkYxlt9uUHTFw6ntxCoQyi18Ls1iO7n4tyLLpiXVn1R24Yw0qgN7YnBkGeipLO
q4b9P0vD72dBJKCLZJeGORmAX/pE5CVKL6BeOL7HU41V/eNpXeJAGkiET7B0OkTxXB1wM+fxmM2j
od9VT7JPrhwmkt16gIpTYMXbjoeJw75OYeXpdqoZvLXeEAI8Ecf3u4ad9YqKWosMo5ZpX8rXbsie
I34Pzm4Qm7xW2WNJNOWUZwUt8sOwCbjAf9/ttMVIMBYwS2PZmYo0R8sP+OB4gQ73Gh6UiBFXAatW
NZ2Uq9fXmmQqqWoN8dfTCLeG5HXfuMy3hGTOCzX3k0yoFGUVDkYUDh5DAcY9mk8lLx1FMAyptQuT
/E+gdmlJxPUevaLa6wjia48CDLXfqJQx/sQvi9m52jVQ8T9H7kru+qAI+ROthGj47xTmDOp/IauK
6TUyBz7hOL6JJ7haDyP/yo6ZIb7iB5VGHh6veWpX8nuOxr8gOHuyrMvopOHHmm8IJuCQZcgX6anb
OsTKVC25iqcv5eUoeawpVOHfslomu8mp1350bdCXMGleRitayHW5a6fEG0OrExfnmF5m+Tlyn5/o
UUXoCU7Zg5fD07bSJ5/T8K1ys+03FRPgtN6UttrfZexUBkjFO6KgKaQU09Ktf4RmmrAhblNkfiVp
ayzZbFbcmkU9fHcIenRiIX9UWtolCfyjPZ1lWdArhmIRHEG/v6QnOzOuukjo2KZW8gkF56Bu4nVl
HUY0HGfigeCHETkI3aWgYsFyNlgABtzvLlRS7/Be00XGzNyCTh+XHVqbxT2UhEHD78iN8WkUrBez
IY5AjK0rpxc2dz7gR8yPU/GAP3Nyh8DIniYyhrGF+a38J1f7OPaa9ETYo5d93a/67o/zglTm2CpB
1aNOQOD6lh73gqEDlcmvtIMeP5HB1D9JMr3cxf8YAP76LBPUrD7ks32h9PfrZqQ502itknhuTLC3
Z8UDVSR5AZpS30afS29a/kc8joUiBJKR2UA8Xx0Ap4pxaPuv7mO6i0RmdMIjPr5Vi+u1aAZpiZSo
IjOCplryz28n1MEUekZKbTgHrtRmQRi0xDZJ2ty6w5kJ60hEodeD+6eiuzFkzQ2WWMJyYKklyLCc
Hf1+2CcBWRsluf5GbTOPHLRl8IZxFz01vh1brz2aggdsaH0RG7dXd08pCUZjEjeZIcByoD/PgiG+
2z9+shZYosEbmETHbAdyjyjuvjG67GPf9L/SPQklh9qKYPOU07i0OQVOF1Yv/ZmiXdJNHPP8Unzx
yQsfN8FORJAUbhT+wVr/VUysPX+QBnoWjihorM2TTnel05YGtEoERmFKF0gRT8YE43WRocwsYqc+
24iobKDmX5+xlgcZ5CIyu24dtyTSONuHraVPEKuf4Rywdr1va9ZUpVyFYzi2PoiLWEOGSK0p7mJ8
bJRn3KgKVlYgJiZUPUoXoa7etjyzehmyhz2nM0Ao41jV/2EVboOyf++xCEg0czD2Lb9TmwACGhRp
e7GQbknvCTEDWRDP/5bNApd84z1eME0XbwFXnxqeG/V9Gz3AiDnKfsCZCSDu6Jc6Y9CoYtTq03NX
Ia0ZHIw2Pph0jt3cyjk30xJ14E6Psi+fgfZEbGQiVOCWQ/ijJzGC/TttiCgUopIKZ4jdWFu0hfgk
GuymL8hxwmtcjRFOkStowvxF1kXNTTW5b/m6+ln0f4rrTVVX9BtwVKGv+1ZRozVGC9u5QDKcmrfN
v8/+2bWadG3kJCQ2W07pgEwbFQ3sOFYOlmea3bfeV4tNYUyjzVk2kkY2LhAbBALhORIMIbexGyVz
alFIlA0VMdT479iuf0WCbite14KhDv9vaE7st0NUaxvc9YRWIYYWEzpjF68qxHCFqEwNykFIvpbS
BcePV1lCG1Mm7zGJH809/bhSJeddqW6/KFTZdMuBhj+jmAape15E2liGAFs0AkjfmPM8dQd8eqzZ
IhU27dCfuz+iu7OJbSbSP42BuJRPrIe6zY+h4dHvD4AuZCSr0B0DpW37p5nKKD1tlRTWPWHTfKJG
KbeXiVwHV8tvDAf0f6ar1ZxtuuXuzKMVpD1RP9eSWjxTBkJzoPCOjq0vig6iQgkKwPPGhsutL+xX
+M5fIWeRc06z2cp4Im6CrBf8MjRNK7m4CCVaUNyNoO+meGOxyw+EpBvR1/HpQs7jX+I0cI6alg4X
r4SPlxbN0irlmt22TWcf4CN4bgjX31dAZW1WeG3r2iBpxcNq3IghNgvphQGvvcf+fX2NR9zYwMbW
0WP2ptSW7WC02XmgZiNouBMhIjCcp8lkpKQ3QrDeBg/jMSeW3LYP3imI3jhcNy7af1b8k3ikXOC8
kvHkTDWcPZjMeWHwneAEs+AQzAHkWIxYnB5nygvNEi0UifwAYa72DhQQ53UT9AzppulmfkcWSqU0
XTzoGOhCMaRxFEKazOQWayrIl/IeHbxXEohI5r5VwkbBMNiTqDoqPudZv5u/yXtapxaZk6Rn1tOE
qoV/XZqQkWlAaaTCRe4AtcI4rvJ19rdqsz5SzDoVfqnNQ0H1p8u6b7rzHdTsa047NphwRan9F2Pw
QeWC8HCgC182dliBZFJPd489uS2T6ib8sMT35/MbOVPJCiCviYExgPEXCW8v/zKZh5aWY/i2TUu7
6vUgzx9FzhPoXvolHFa/oL6sZQ7q1nunJKVV5SW4LzPkpQMXP8YSqlFDgNs1559EeTGqe4c/9nv/
bP9tqT6WdlcXQbzG1H5kEfBf+cY31rxClutQiqD/PYZwXcFuQn5ggeu1AwZORnx80thnQTBJk10y
/49MGLDBtDo0WmV2jf+hCZYam2syilSJZyIv/iXyQWK4yQARug3OIuEuGQp1qAbMBob3G4dH8ELe
oTtX94zCmigESrZZzC1VGDhQxxuibKQzKAvKkRDr5Plv/ptOdRE1+WIf9cNfv4PDXYqtdylqOae9
eYUqM3l00YtQhSGDLh9abtPN7BvUij169xtB/UQNvlNyEstzZLSaYjG++Posyb+BDlCaXvWWjcuB
MqTGrU6jyhuVy/JOG+Vv03HGq9yvfaFX/d3qRHm+9sGvGXCbnufbVfSjbYsoPOpMLPFqPcN36DQw
Qh8qtNvmC5lBq/7JF2tLGWAIKgUSV1QAtc/24Y/P+Si3zTUTaKDKhFtL7bcFmL8RkAeWXZ/urbZi
du+er9EQvQNb+9ATXrjg0FgQIjqZXdbiEriPJLXoicWt/6vAhaHmwR0R449tgJKSgj9HqqlaJJK9
KMCV14N+4uoTAb/1fIRB/jk/qw8qQHhNS77xxwMVTCo7ECarq22BDdp8diypj17KVZPoPooeiNw5
rerMKX6Xoon0p+d54DqXN1N0jEdwjocGSNr9jAfvcGA6TlAdT/63QgT9ja86DkOwTIK0PKREwwML
cGeCZz2hCnKPTM7PWwFvurVfVZD3aBpZ87rnO+Eoybjy5wEhiMJOOknOZbfcvJrF/A+T0MMl+y7I
0rj6onboMCPUUJgos70d7kNsgxUikUmSz9AMFhySJ4n4ymA5HWZTEI5mLWJ2MMGo96A5nNxgvkMx
e2ch831JHfNNkbToJnlev3Cgs7EbtKvZGlQ/uwA1A35VoMK9B5D3hhsMB4hKR2ZKaYuXv/zIzors
rOsEbHxewDnWEuVGnkinmqZbkjmBdowjHkcGozeaLK/momeyf2wP5hhVgbUhNIU/CjCSWbMDhsbT
VGT+gIS2pSgFlPU7vbqwvPusnv3KC49Z75zB+wppZamVulQdQX9ldePRzBKxgsP38y5HO6la4AmA
/E+TFPFW7tZA41CZL8RFNuWCfzXC2A+lLt+JjvunG1N6MJFOomLIAcoanw+QRnk4PuEAuefUWzsf
kO6J1RU7HZQZiEgNl2ZSUKLH+PXa24rSlC9clVZYrnPNwOarUPNcmIvERYPwr3SHKs2cvUd5nREV
mAuXlwYcFOvaTdXeDG0nC9Vq6iYPQHgtkPoE6qV9b/TYX3XXgDMUCjRfvjGbRt+gteoeYemZHa8d
g9CzKhXH2TFtBAkQWPHqOp/65EwInkOvw8Hwt9mjCv0uFdmlyEsSX5ldiSZhCeWHGik5WYOT4DyG
aIiQcvE7y41HlyNh43EARxOW7jx4GKBDBCmjST8kyAZ2gQv0g9ziZ0ppwYrfuRoXE1DijRETLJ4p
Pyy+xLy+uNbOEQsdZULgemmUCTM+MzVorCBzwKr2UhuaAwbKEyL755d/yPETfd66NO293l5hBSi6
+hzuSeA+bJXvdhvKm5fxblXM1jQh57lp7qH0GAqiZ5PvGW/d1HymR4logeGeasYglZEoJtriwFGk
6P++h2jZA+TvTs1SgsRQ9DztyYLJVoeowRA36oSQoLBGRVcGlBd5LWVqNPJ6NdjJoawI3O//0sY/
NkegGwunMYpn2kur/IqiZTb5P11yWzztZ1DmqRE4pORrm+yl6nNheeufl01Fltm4cJILld0zkcXU
uK0kq1+LBF7HY9GLtCuUz+P+VFbluZaCAl1KDFbpK3s6pjtBKx/WB5AlvCAuBovrATETCNQSoip4
B2ayjY5OCIKp9lJp7wvOSrvAZfZRzAtXr/z9j+y+Pet3FsscyMvgQurEEm/TQCIhfR7L7nt4Uk1R
aClKfDsokKuJnhJ6SRnmi8InLhImFZiS6+Q7CHFRLrBotHxyaaQdOWYf5O4+BAlvXhZjTBnN+h4Q
TumQW5BFbR5/AHIt6mM6/E6/kTP9YjmP2od/KSWJP3OpdeCkHO6YiIsMBfOFKnDrSy6MaMUSCEoG
dM9s75MGUyILLzXqIW0nDXDtBrrjp5oA0SkbAS3UhFN+UC8n2D2TMEcINGafvO1vbmoLTnoGEQ0b
twclOlbeVUWejb2wLEbBQBKDpQMe88fsveiyHC/rJOiZOUFGu4oSJu5WgKD6FzXSIKgHqqVH3Gt6
Ylr7SgEz1roJ7plx1eRxkOGiT1w3y6K9PTpNicdts2iYUZMdmughGLZS1hWNL7Epw2kkCR5e0t8z
dOmNRx4dJfaVfvTMJMN18Wh/z2m6BqRT+ITxHzhQGig5OEoiPDGKOHHEwuOKQlU7v0TPmaQqOBi/
onvNwWjs9j338MCaGOaGLMwACNPcKD3jSYEMw7QbzZ/cPF6i0jbsGBcleejt0AiD+ZSNdgtRRmnp
ArJ0ZfiMacHmiaKVtET+QCqlbppS2jPSFtL+U4UlaNgfKxRkuz209XMaCYxXzuxXEH4Qy/rxbg5u
pXlUJHBzWHT+Awe+PE2kgccThY5ymKUC0CSnor6/csKV4wqN1H/nQZcfYTpgYQNFtZTwc8qc05Hy
BN3Hf2Grvv60ajKO9m3laz8NPyCd7pr0skAuJu4+hfksUkhaBB2xyRkQS0c9IWpTl+F7EZLSg79v
dBVuXevDPsqt41HR/FZR2PjmdmWJQFA/UsXY/pAWAQMiXKE/tWOBkm3eXx+wKDyXLF4CuvR37gQ8
+L5/3VXgeUpwehitO6dhDjgJOAcN+NHNvtlrx/09v+tTpOjkvoU2r0L+WaocJp2Lg1OkAyqqGbcZ
dqLAqulHq1I7QSN1m07jhopcfPODEfRszkaHVmB9no5k4fcEhIp8EOy6VOvnFbOr7GY/GbmGdh6g
AAqY8N+FJwThYqc5/ZA0Syo5FLMftSHRD7X6tTFC88zwtF/TwqNVtWeXB0Kyps4XytI6qEsYXM3Z
qlnd5i0gqISS0tfdtzTcJnZYfJdzATTF4Eej0ed1UxWv0hPLKRnRxW3pKiwETerTFGYEBAGVTO6o
FGtGrvP77i3s3Kkj4L1vrUI9L2HFFLlH4ZlyPxoerffwl2Fj7PHKqhVfimhEGrfWgGJbGe7LKmHp
8F4EtXjR5t9V38OQZbvr5KQhtdzU9HGxJLhyv9RVzy1ScsVwhdZQTKj7tnQyHU0Lqfv26FR/DDYh
VqkRZ3RNAlZYEOjbAAnWrclAvdM9L0cr2GWKhumIqryLRof/SjZD09qOWQEgmoUOChK7wUNSIxXv
8GMfAOvABEPCoUQk0794GfROdy9N4iTm7vbev7I8FVs0XqRU7VDJR44CWd53lhTtnFU1HXAFpQy4
aqsskA+pWqKIRhzhq/KuEDN7gqAffHwMG2lQfBsMhapCbLZ50a//CIpj2n54jGBF0RbOkkPgkJlk
ygZiSXZiHVXMMSHwPHc+luLtRy71PUfyVKRRpVcUmz7ziKr+1ccQ1917eg8l7/2d8cgq0z3RHk6q
UULnIGLSQXpdH0EiMKimvpWpvDCdDjBAYU9r5dvU7LLKKlc/chYaPa0xGMY8LhkP83j0RcxoAl9i
9IWVWtyPTiRxD2W6WEYy2YMo8YN+0tNwSzTOkXDQu5J24rSJIeNiDako6nuEA/eEfL6PuxVKHrhb
FVaPVKap/on+jVN85a6dvaVyCQFPAI+WXFfKshCDM3LyTRXFQDS8P48T4D7S4r1iLUy6M1D+WQ5T
UycDrV5luIhLsdj2YA5k4AUGnG93wi7rAuwr10rId3FFBAB5mTZqHq0u96/xoD+K3AFhYnJWATau
ICGyDamgV6ggjHPnEKK4FmR3YhoNHdud/1x+NWqEn5LnwcGIXqDKgcC3atvETFAqfmam0mxVdwTk
NmQsUnbiG+lRsd2CZnWlYMc+RWhi0rdULx/vw9+ZqLgySDH6hgCjFOimRZtTawcDW/Y0AFWhsBHX
hRoh8SaXDTcBeT38aZz2S95s8sERDZHZ5LKyie16mLXFExy5vNCmAARtkjeQYlT8LWDGFamAN8CO
TUgxglX7GmO/6XYjy5GHKE3/7pm/s3fxqYM/VrQZCt7bssCht/nFhzSwNelqWK9HZteezTvFOm2L
xkQISg7d/D9TNFlzRjUYxMy0pszBBhpg2XYj0/kGRL7t+IIzNwuP3PvTirjofXUO2vRqSav6iaPJ
byc7G2NrboJ+B5vKapKmKZcmCji9PELOpybrp5i8oHpFu4vtqgMpC8vwU5EL3CZVl1Sio/oeCtjw
SBxe7GbydTcIMtMAsF8Gt3K19h1f42ifphV0roGdbuhtYDJrrHJRPbNhvBKneYdtdA4QhPSbgRNV
4uYF/VqxY8fy4D/emne9LLYnGZ8qNTuekJZ8O7g7YWS8BZ4LriycyDL1kJFbIvrzFoUFnNreQq02
s4/TUs1XQ3ySo+5pM5s2MdVJM3b/ZbxWYuupSOy5mxV5FLZE/ytztNxCnM6ub2ekVm5/wKWgJmic
wepdzt9qzI+33N7mEC3/s6v/EUXtQSZBqnOkxhJPOZ0m3aeEWvhJ1gi9bpw8mNnmhUSD4zIrYQS7
cB/RvAU9D/hkxJfC4SEFTNawXrMomqmzTqlVF34yNnZ7h8wlTmDW50yvDPWN85lxro6cx2rUustd
6QLIvkYbfY1yDieBahCzcszQ+c6JveWnJ7L7l28r1g/q3y5MM/ndHeOrTqUiVN+7/sXgr5d4Y2Mz
iRmypYeDv4/4X+3Wd3x7goCdcf9AgQOXTMIY9EgrEI5Y4kWp7RaU2hbqQtkb5z125PApzdJBZkzn
DkqUx5kRuo3N3bokyPELnxmE7ewZe7DCalp2D37avN44mpSnETv7al7lgsqrHb0AKqMBxpIn/3Nz
2rJSJ7hEv+QKsTAb2eKg3hiXgaJplv3S3xOnLSfzvyf8BUEDKCBOCDoztRUUR7CXuZpllBLZLnQN
B8s6N+6Tub/lHcsLoObevU/arGyaK4jjczwK1a1LzZ0Z51ROq1JHoeljLlc7hvvjXw7dGQ1F5hns
Bdey4SesJ+80EUD9eQQvIQWJbnyyUCvNwi6SvIy3qGSmlGR/yK+HQz5f3yS8TdRYM5msyt6q1J8m
uiIJroWD5hJ+cXORyViv6vpiIvdq/x3nq43O9DW+unOI9cEe/c6i4T0zxWCOi6tcclvwRXKjwms6
rwVZ3pVMWuK3tFb4UAwC6dje5qSHeLhcR7DcpKQNYVhjLH/nycQTMyy+XPSdUGlW2RsEFpd+FsQt
lEV+Yzg1mOdo/1JQPZWQ1zE59ILogwyu3kuxktoPctF6uo3wPoCSzsQUP+Jn1n00ZEYubO3rFm1W
/9KlC+dLLe01bpHBHYXaCUpARYyQyXBNWtvJF64atFAD3XylzFgtVZ9vs5tJI6rO1tcWHaqEeyXr
CEjlvYRVeeM7U56npBGuHVhDU12FTdxMW0RBxQmu3+bI/orYJQJp0w0YcYcb7hSsw2Y2Sin0Szw3
G38dLYCbTISbQbx1Hq1Rz8WVn3q4FE/D88rnPkAz45LF0W4PnmSc70MRAA8EMWUSkvdl6Ygl1S/x
RVqw691/ANyPKpZZ+AZCluMsKqc85nVYppBsX+LWDuCml9+MsVrYLpjkE/EvrEi46ncbcXWHFtnA
4Ky9vhNqbT05iXyN5JUM3YOycMObqGhpbseHjtqrtfxvOxB+B5Dhggx3aTSpmU5zSKzEYbznmyTN
SYeCrM8xOVAM3zajCeZz4+Urb1scgbVPk8sat3V2IQLvqYK+gDrhncrk9FPWYXFS5Hs8+vvu7hm2
Dm3/njIfP6jbieXUoZWs2QQk8qsOR76mz0E1l5YGVe0neYU9RcO6ltiFBO1P17gSSReamuodX/25
wQdrMXb+sgaZZgVZpFFikEruLHtDs8avRCkiXsx4odTJMxJ/nPKHG3ANiGyTyQJhB8nJ2KFfM0Qm
Bsj7/+YBthwnP82ZdiZ/mtKVg6rMsbeeHUAWhR9KawUROEOl+lwen3vzuyHMmn4fOg+kTBUKSdPj
JTc81xoe++hr+BngEW02lgdsLcjZ2VvKmVIvtL3CNXaZmwJsG3Nw9FVmiCjAOOsTgXVJSbHuK8ZM
p793JWBE3FZFKOB2GOMpjJM94BhxzYB4QKImbuDHpGTxPqLXZZc6dC7f7TJgC8OhQg0EwwY0JceJ
Xx7poyI8Bj4Elma0/c/AROh3xJ8M0Z19JQT1fDvTrdFZXml9p+bm4UR8pv1+L7S84PjHpQbjq7pM
66aUlcDAgYCe1SXVxTV05spkgskI9c7lN2Uc56htisgSXo6zgZvn9LZhtX30R6586J/2pkjb19k8
QrLSKbMKDV4s4JU4RcG+AlGmyN79L1HX6CV0G2QGVPBH/V0JHxS6m2Ox0TGwaGITcSKG5LOLz8He
qKj4LcAhS9dB083IYTbCRhFOTAVYbqR8gG+6pz8UeisDvK/qiCECxUjos1dJTsTDFOOqpjadD/VD
/y3ieDenZpssWgEJvZxUYLl7FZQrE17lki83j8MoNfkkO7emC/KtdB+kCT0pTEUc1GX/KQdEEZnJ
4w7Lq3Dj6/Lq03ZS0mJ3jw5dSacoem6c7Fgrynz/kUNbJ8Eo4KUD9ZMOF3AgQ8iWtjFn3fWROvZf
xUyDH8D9Lx1cljWSyiQ+Y3DcZOCpCotQWSwrrFk3nJPtKHStFY3mByJfRWCBFu9udNbmam6iSV7V
8tcs0ACkVPnm0jsv2Zim3yqcID0tzoubqzSLiTEMvzrgqryuR2x7/wh9wFWCPBQTesyAEMUYRCVc
nW+IayiZ1s5KUoT7uUPiA0w9j0Z0vbOmsOCeCHRMsZks5xOcSiXIfTqiOQjG8P2Y3tfF5iL3nfzj
PFhMH4aAa2SaxeJBUDVLEvuhqWmoS7gnTB2DD6LeWJMecJWrP5VgFBgBx7KlbfvG6z0QFOK/4w6d
WP2qwt+ILQiN2JB/zq5IBTenaNL3FmZDID/SlByMWdwhFtvStcbcNlEr4xpjMwu061li2naK3bin
iWH7nQHdOPBmC9JzxnL98InYZ/DW5RvBAh1VsVtXq6yPHM03bvwmvR6frTSoiQRdxSpXdhotyRE6
3oTQTeVgjMRCgeflxZ+OePqaBDl+hGWMKO6VbqnpIL0ljILnyVtrORbnHXc3uedUVJcc8JEkJbrz
BuKW8WMwxa7MwwJbn16iqdDF6ihK/4jP9jYIzVR7lNR9Y3U0j14suSb8yEIMXzS5b2OIvDwjmkDh
VsHNwHx7iD5sir4CloxQL0E0ajznfv+TmocLLlWgEhRVQ+HEqWYeB67qv4E42atpPNw0nJ0WWOKc
yz/VyWEDtN6DRXxXcRb+hJRrb7af3W8Fka9c/Q204WdMZ1dimj3SCOUCKYXctL1x142i3QbjBuNk
L45SUrvAOSGrR9wdRfPqmurXPiaTA0JZl/cX8B3wTRPoY84D2+qzDj7zNX4Uf6T9kxzgsu+p2s48
365pBc6WT7PowfbRc+1XtHgCfsveRSxKJjTxq9UJQ5h2JIOCOVC/3yMallZ8cCE36b3Ou810R398
Mqgwe3uwGOxt7HFyfX5H+6E8CPZEEQnV7xAWeic5FYagJMybDyPjfS60WmQwlEDABv0LOznWWxi+
5PFS1ezTfmkERLw+xWh5c6I8ygUqNONJGkGJphPE0TB0IZ95UliumHGhwZBT/Rt0Vz3TkjdydU7T
qZt6Ux8IzE2BWScu+xVTw4wCT0FYY9/S5pNddzfUatzDhCALbmhX/TWpBsmn/EOWj2nscqUq8j6b
iQvIW9Gb75ENwZO5n14nFXaURdlRc/N9MWiWjbmiJ0jAFeG6uxAglAAqpxPACplFPI0LwNgSdcH8
cUF0mjfb4bGvlMpX6qhZn5mWZZY/7MmTgODjVyAIlv1tQgIOu2DlN9OP4eU2+vW1yrguzzoM8xxR
Ci0pgex+t1wBhXrrnRFPan2xl1gjXZIkBiv2JpKD8zaAx0l/zOtCrY/KajPpJaI6tlgsgbSCQFmS
e2Y/lEgrF94zWUUiyb8UdJMLFB5VchnG2jBfZCwLob2u17Tn27hKPf830dxabOPl4BFXmMYjtM0S
yq6irEYxxlWOsJcuiS/1d/A0mq3OUEpnj2U4TXyipuSz+MVfyiytTz0Dtv0lw8liCfX9J6A0No0p
hq3Yh4TD2W2nx2o2ZQBa8Sns4iTm0Hx8JjigUv/VgowT4AFssgCaoxwxpYnew03FouDc7UKD4tmm
gVjl1gdDL/Fal2RWc6qxHoJKyqB6HPcuImiMwdtoiUjWfbzpOM9PZJU2VRtGNyGXymZvAv5OcgyJ
YinexYP9Cr+Z++ugnBirjUCxhKLM9Ec9CDQ1ty2kR5ZeItrYqH9Za9EzQUcQyu9SszWq6fdFchiO
9JWcSYrk5LENLrJMr0SDR2oK5kNEHK+fAMTaK/x+bkcAMrNCuUCEZ0NxxbXgGL6MS5DmZ5yMq052
HCNF2y+Xc3datZ2X88yWGFuotppDOuVxLxATUbuI+YEjZXKRCNDSALfT6z3gbptlLsG1nMS6Qr5I
EWEzsOBTyXVVDsOegVsN0qTa/YITMovXHRmyOcwd0Vfapm+vPt1dZVxQhaV9tpzEaDOQTPsEVYgY
y4t98rMdFMHsmqgim0NqNmCF6iojxH5b9ZJof8nDMBjvOSEzdWscyyUvE4Vv5efT43S35bEgZASZ
hnkbsXp/aE0D+UAZue0JgD/pdRTgtFxFeon7kqlZlzCpOjrnbqPP4IejZrcKAcE0aCfEDn4axuaw
5UEckFn7qLaTgS4YOUGonA3EZQ+ycny4I0DTWm2ITj/SVwmkEsYMdXmhcdQY+7gHa8a87dElvwi0
jXM6qJ7RBeDR68DDsT54Tzi3rhoITO0JUT5bFuGOQwoCUvNVa24rTCUZ0RpC/P1OXuVYAtMbbpRt
N/6/jEN5oiOVEQuE8sLNNn41lUvr0jLiHr7XCJT6mgmU670cC08xRTR3Yw37r0EIW9/XY2y9/1tw
9mYd4SPBRbZP/71UDLXn+DgklTpLQvlpJpVAAN/IZVSH8ps6+3J4ovqdl8+bxfQFxDt7DZqYu93n
uf/cqn4wa7ZRbcj+lpCtZcN0Mr4SYy/mEWGiUTHXL1kSzPqZDybGd4zNn5YAGz5PvOx/gxETy1eo
FlfEGip8h6n2m3x9yQR5S2tyJegt+/kDnoNMXAqyDvdJPh0cDGV3uZMF6NNLWoF0OXaUZc6C3a7+
89hrTmYkKja0vtaKi8sHXzA6mJbe5xfnSyWfeRAEE8Ue+c3HJXEhnpc169IJs7FraTe/V3WBDjiV
l3OEDogRE4oaOMgG8OabU5uBWTrUb4LI1fzEriLKJlkRPNWdQpHA1Q7n1tz1wOZXlCH7d8jYwlRL
WtABim/rrkOaWhRcDC9eK//lRCUEeYuEYCN42MN9QeIgwHKYM4W+jf+QPcy7BaNke0ewqc6B6N0Q
1GYBVPz2HlRveznqvx3QrjcXO+nBf/n38A17BH1O2SzdIpf6xBp8UxOCpsJpxaIgE5BSu5VDrUfO
9YZCMJBr8oFtu+RpEu2/SnuMVCku7rRlihZuIJEOGfnN6lfxFT6/XxAUAib0goouSGZZ2x4giYNo
5QMn76HHF/vJA2xLUoaayQ4xJXZSU0KOy4pTJXKW6yHRJz0qC7OmLDVv6bJBQVS2qX4rWgzwZLx0
kx27RqC5d5PLhApidA+C65V3BzTRF28RR0xJo6+aX030n3T84jdiJuT4OFLACXYHXClhu7ny+kOr
2gejJUOgiqqt8J6b8werrHg5qWAfe9SvCeOFBjE00zET6Z0xyUzcG6dCV/R29fUqoni5NkVgsAza
t/ZRv2Y5A3V8IQ1KFg0PVIFv1OgCcWoRG3jP9Mf9Am46cqFjZpUkVPFGjCGoq8PeNtX1wp667MKQ
hWsZclmmv0WXMKietNdGlbf8fn7sgTesAGrS6+qIgpYy3F9v3d6zrGJAiUUkywOQVg10MBXvFRMU
UvB+rIjWocsuGwbArhK4rSyYt+KGRUdPvkLBoYtPI84FAm2vkWEALhiYPkB4jgFWY2SiFXxcFMCN
Y6v7lFZbeRjgrlUvaNXzblgM6/EvrVTjGwPrEf6yFxui5DFS3sNJcjvH4N04vDpFG4A8BICoOpHn
NDeXVjVNDi9wqtWcn3tzp2NiuaodNFS+EAJgdzZGDb9AFj3kTcuaFdJt4AsJ1mu4zLThQPQuUAr9
zefsLHe2mivV6DgRRk+UwIHugywquGu229KRNi9mscBsrcnKpvVgZ79wTyqCV/Ha5XpAWogVdZzI
G1+efKrekL5yY+XbJqy7UzGfRVs37YuamK9fgfd+txeqKbFHwnhdwyarXXwpyWgairxcE3W67fhY
UnNhKWvt/WSSUyVLgaDetTCiNWCvuSPK/B73YLzRH/kBkyoG9eA5u3yYis2mjnhF1RJhJGmx1YMa
eXmDtQj/aalG7OuwK/T/owyUbnEb5IuwlKBL/w+5v0gJHsqC6DwXwRDyj3TaRu//c6XZWId1NT7t
CQ+goFyFLgmNQ6KOH0b6zKF8r16opgYfdCyRacSNLZRAb+lJBAIMXz7ExLizrXNQu5UUuBkPKlB2
G4A3GeXxG5pxZjw5wE25UCJCSoQPsaqhynBRAvhcrb2z+HzVbuJhdD4AamGiHuudNdeKfHBn2v8p
C8V21dMmiQga4Id7/LRotclFj67PUUk0Nkn4CyaD3nI/YCBM65uH9eYIPoEYUNVIA+z+iESvKWBG
cqskehklHmjvlO8jfG682AYv+aDCoBcVCtPTTlCAbfvHK8p5mRYhgRUkW40dX4EA4i2JKGzICX+Z
8Q523RxFVyWnItN0IOQm0DgaDWV7VajXkxY6MG1Ace5SjYxuQMH0LWYP8gzKdn49/qnmNz0B3pdI
lgnGKhSCvBRDk9qy1H/zn5fCs87eJtS91fe2VN4OAPy3emQ1aDJ8g4sY2DM2SVbEzuGEWw2AQiZ7
/s6R49XcMryKN4JA1Hnk1P9uQZbmS8Av3wnHUaawba42vaMPQzFmj6k78qMLswhnAtld6z6VXgPE
Q5GKCOiwThBgmB5Iw4NAwgrQPmzvPc11YSC4tPuZKrhsgALlo7qinN4+g1r0AIoeQO3k/6nzdmE4
476BhYuihsLTCSesDoqLK5kS+7Y5fu1TeeZqcGiWmTmcGQIbJDdrE7npF8Ejr6HgpFEajmxkR/UW
V6/3q0TF1iA+HZRTAvbOP8gqeriVTlBGqPYI2MjI5rphZbtP6Amn67DXllN24V1W56DZQPLWm5NZ
uWFZbqWMzd9mSsz7U/UYSbFQ7kOvebPNuhcGI/fkxUsquJ7LgbUSPymLL8NyhGH92zsvB6Dpnp+N
BAXABYiyYg3S25jyiOASRO8OT2hQsprg4E6BxzuC+nAzWpyxQcbvtgb0mhqSWPjGM9ectUbrjBJg
+s/2zdt2jmL6qcP57ikDAha7WzGajvb6jKAvm1/8UcJFHQ+cHkDE92CfKR/UNeUaWbl0K6FDtrXf
5dw7R2ZysPkioWs6IRVdRUNPAFxwfPwVkf0Kb1nv/f2KSgLRhlxFi1gKRvpmF5Uv9vUoeXT0ka5z
OjqU1wW59uzfr9nsCC/bowY2242bSPwmsaegHPp0u2pJYaa2IPFkBcScpQnxTZPiGFuJ7+I2Mzu2
KBPOEW3wrauL+MrM5Azv8y6+f9Pgkxt+0ME9fa0aN1yUUIUC81f/CN8mEhLyQ2DdNqfcdArXSuDk
+8K/yyr9deoinw7Pr2XQ+GWtvFi9feuKzgeWeoMuS+qE3D6Q9v5Ilnjpc9RnrXFCtKTRBO4QMclW
WBcYHVC1tncFMeVWjJjqubZ+n7PPHn3CFKFrweZ+TYZ5xjRFiiGTENn5Qcvut4PjOKX7RtiNwcDi
blUzxVYWX4r7imSPukNT6o+5lv7F3rDpldEl3Y0R7vzALtW5CN+m2KrIUXqY+R88irWT6sxsQpW4
ZOFwj9V4XJWW0E6b2rIXo1cYQH7vm4fIXNtshcE+zEtO1mb82jR36paFkqKrNpV6NKXsz9NG4ajz
IkIjEPcK2p+UzXzVSNaC9Rk8fgD2gK8ak12uYWA1HaOZrsofNN6mxAaqoDt4kQVvbzrM6Mvg7f7J
rnv7Jd016Koekivha5eYwc9KCMgWEstTpZwM6KH87n5cQQRgzKBsR4FDN13OeAD0UJVWlE/vlTxB
QC8teQsoXXsk795hlCFwlo7nUs7pykXqUPPXuw5pwXVRWa3GOpUoDSB/5U8ldft6k5kAAlck/XU4
Bu9dlzQToknvT2n45HS62n/yk37KRcqUQiKdrrveRVxXN2V82m1+p8Dli/+tbvnIrF2Jzec6LTSS
/00+ycxdMIHvcxqBWqMIEQvlhTV/+Id+ShnqEowDjb5iBZNzXh1VHrUpK/oaPfSapDFjHzBqAv1S
YYaVaaqyqPeJjQKiPElziuew2bED/Z4zN6jilnmFHqboJwvWVawHqq2mRz79728APAnF5NoJeh37
6HUlPSfjVFgAjMuw25flAG5oYIZPvIwB/3wFBC9po2MlwrrkIYXilzV1OiZW6qq9nY32rWTmOakH
IIHo3McD9L0Ym/hrqK33JKqwV4PYlUbKw8T4d49rIMRv/HxbiJ+6A4z8UQPjapkc71VYSOGvbT5D
WLj+/Q5y/tJoJSrUEYevTW8NnMqVCNxmkr6Ohov4UmxmfKENMpLVB4eOd8uFFEpCvoBem+JZtZri
pwOeUqWuhTD2k9wk1oVdbK4gBNkuWWHzWOD48u2TNED1g1dIjL8zYV/lcxexSxpacFaME97/1dkK
p0RoXfY+lU8LZS+23NjwiJOQizR4F9vlZGR/T598Khm8/rsacSZoZkW8/IJolFVoqK2Gfp/fhDoy
0kvAs2V0eYhG/PiXgtoOyvfZh82as2hZ6l0HAQwF3DuSV4Kas5DFnXzZ68tAgmmYbpDoRZ3rm9D9
eEaYEvkr9VUHlh9XlizTIOejKefzYFF0hRdNp7fUO5EKEMx44MKKqaDJ0UnUVZwzFYhL5DPcJuTs
ToYXRzAWnZ/QRlMWuqa8qpUe2BEiynu9joxqxL3aA0UJj6dK1dbFkihobLtbZl37o5iId2tlJOPU
6i/SQVeuGp0WOV1ZllCxDYuzLFcHFZ5KtIgJlZSXDALOxqYR6KfEg9JPRmMiGO/uwvOb/Ut43xbO
4/9/u7Qs+CYPMyqqHRhK61xALb2gqmaV7zMsf4kYSoB/l0C01yVJYEe+05bH5zYDm8ZIbK5CtXlj
zk9UQhktJddjV/9sY1cyPJjoI9E1Hu8XAuHoKOHmbk/mXCgzFo3KyKhef9B9gL7Y2AuJAHvqA2c5
TDwS60qxyEe67KY722cXLn3TsizoTy0AIoL56PYcW1vwTD7EOHv0Yp1qWrAHydWcGttt6x4pJ55f
Ziv2P0o56nSjkGNErwHCi0CSVJ73DEGdPxBR8imqpK9Nbdk85fCMJEKvOwPMFDrA3md0sR4dcPMU
se92Jn1MmmYcJmJHfgy1uGAVnARFS07i5uCny6yRGUnPCg/VjTXUHulVYUVY4G1Rr+YqXw5BfiFQ
1J5y9GcTrOGnzeUc8/Wh6KO7UuGgrk9SdoVpyqBZ2EcjvcIoxGdVtIowKPkGVTvfcktxT/Q7IvlJ
9yenOdit6UBDWCMO1PpV3LMR3gAsxARXMACLGIrpyufSqerkT1kD5Gem5AKGFxMfsRKzJ2UYBnUU
n+8UUmFuYC/TJlx8q39zebb283UIdVhhadxfp6c8+jNaC/pN2OD9cGI6b745VJcgpn8Snu7KYq3J
0aLjLaT/rn8Y3wQD/hkNLS3246tNIRrP4xdfxxO8libHm9B4fobOxnmO7pVsvxLtUJhBSI1uBfEq
7yncI0YGiebvl7iJtg+9YEbVOs7ebSlfRqBBCmDgSVO9FRs3FzgHBnom0gW7mdNg+hjYhtd208qW
33P/NI2FG2QAlPZKk0TPMeJwi594Wotdc3tZvADNXPZ8eRoBZGBuWfeWxcxlBcIoHz1CyCzUSkCO
mxyHp2rdev1DWwEZFP2QAHaLn/YpIeHMMgwEBqm1GxNuxzBJ5g+50YWJG9UGLi4sUTO9tIKFmXtG
yx2SHXx6F9KChJyZg497+Ym0vA0Q7Ni6Jlg5Jmy+x7jD7S31DtGBTKtorFYS8O25wcaQnGhcD9j2
VonQuncw8OkGZ52DWg5gw4z3rxWCZXrmm7HSOlnk/xVoQhWMJzBBOjUREw4s4oYD08lq4iRrNnCw
N80xLdNa+YXURRpAD6WQHeGKAmpNgGKKF2ZEppA7Xtuh1vpkrlCvZqR2sE8EmL0iXBHsaJhcLcQ0
idrmRkATj9OC2aGhk+HCfWxRvsVM34/9//KoReIrfbPYmSsLuSgGDjIEVZQaHP7G76dQ+QSesce1
ek0lZHvGMVnScQScowQzQGOVeM7odxqzhvbhBFL1iKXyMMalg1xtsbEnf0z2Eem2lYXTuPcoCXTF
Os+Op83fbHYAFAi1AA7CiF8cu84cVj4lpCg7qLBgFDeK+QxxtRUdI1CbvmORi6/xZz7p34qBeew5
llJoeF1ZXLG+UfV9SlOM7a/7+oxkmvLtFOxl4le4VAWZekrqUbp5KB39YcopOg097KoIlD2GUIrO
gNnzyyKJzlh6UQ26QCe1E6Ub3FcbkJ32fCGvnwdWj6rP6PU2KopHxl/PyfCn8z6LIGb7EvvOffcj
Xv9MtkqJ7WkNJ4YRnsqD1YZ4qUQTrM8ASwbgEHkJbw7DEy2MSCeOB6ds36aPlZUOD/RE6qMwebUg
aloIH5CYyYhoM/7Rfxh3sMp31eMxW56GuGEOriNyFMnVde+yAijX4gs0fxGrW9bzrQ3Vs8nCakZB
NZy60e1yAzJXmy4UI4ncDkbPtTspjv0WzVPEja3UAX6MQ4bLW+d9QZ4K52VzTahf/hzPD8K335U8
HFM/ZSFqON8/sx3rjMnxsL5L+xpHaj33bz9n73o2Xc8B6jR7DvVla9coUvaDMgDJKNyki83+rdvR
hrRuk1rlUHAvCcKT6Xmk6si3DdEEy8K0dvzDrAffjhUDlYnmtags8oticM4ivoMMEj9xa26bzDqr
1Cdp31KUZSaEbD9maYknpjUPi7NURgNPId3PidJdwW8IM7faO9LmjfUZsLvDkxe7e+nm036y+9fO
nfwnEH2xu0fo+rLOSmj92aH7OFFPNec7ZVzpkqYv1Ol2mrtASvad0bXXLT+WfZJiBaU1pfWf+S3H
4z//NKIhJaTSQwIVvMwULc5qPDi7O6lxzXW5f/0Wd6ccgEd7plV/VTyewqhYU09b50Hu9zl+hOH/
qxgrS7jbATH+4gKoOUFFGLXvWqAMGKRDgHV5B5gvHDDe/ykEKwNwj5Xa+zNVDW3OJKsz6EHOvVuv
/vKeZP0SD0nb7E4zBd6dq/UVZBcQLz5nsi1x+8Tp9zfgGR7TQhTLMcaePrJVnJD4MEAC1PiJGawu
6s/zaA6Vpv4qqV5dJlmEYRLh08DFZNM8QztytM9xmV0g2ivsDhnYIgkbpu6RBXHBa75b456ZiRrR
eN+b9MQYHYVrwIiwBHI4ajOFWRd+jPFFCAlwT32Pw/Cbl3J0unrvYOc9CAQJQRUeYCA/sVGcAtlU
nakQkCrBah6PcxyZoU7IVNQJqEoeL45UJB6mIIcy6lg7hfCmA5rbcStzUIkEnkACZmxXDHnoQtAX
HTNuoKhUJrEvPPPsWsx5CGWJxv3wgHa2kNjhvbwBg49yonLQTNuRaeqwj514Z2WbSelDgIycAkOZ
exNe1sdb70zL5thx5yt89B3odz35V5fOPNFqRILErzGUjP6zykJWGn7rWnzoefxUBOwFtCnFOQ40
3rKGg1d2jy+nXWbQa7G8hy6nu3LGuC/vPxWnMVz31RrceEmSoc9zKRzZEYxpGXhQ6rfELMBUul7V
+2MeB2opPVdmXi7jlXCsFSWralruWBZb300rqClHtojaegKGzx+3hAGeP/lC8qpoae3jzv34PK9B
KHgIisNDi7EcQkNUCBHrTVZULmAIQWkBNqdkAxCPnH4hO6PE78oqN2akZxfg8RVdHDisxCW1e7c2
pop/aBqX4U8HkHRgEHwzeJtm/DHm3KSRUPm+27FCyJ7CIijpDWyu7ARXrRlROB6/mklmpc95cVBS
d5f0C6Eq8UowV7OGg9t3FSzPu458SqFou0EuHAb6SHTJ2vBIVog+WusrhIQkC8kbNk83Pt1vw7BW
Y2rOhL1n0YGbjD6BImgggxVUpw/pKz0jq2tEOq4VD56pAGAojy1B80o41OSqwPzHbSenIWYwD3h3
8aDs9xKeYYsyWoSi+MXP3fGkjbA7gAbo1P29cQV6xobXOgAf8DuJhm7KBIXzOZAwZ9lZCMRFRy0I
YkmCnzf+iTg2FHhpMuwyy2KP3x95x96tXtQ5JUJNwzR4lCqLPDXd9DVjWQnrnXZM0iXzUzuFkI92
Mu4hYbrrahUDLAX6WbnZSooTEP0X7iTBrre1Dcvm5A0A4EYWFFNdZqBKw1E2TVB7L6QsBQPOnZKn
Q9KhsP9MsNnUhRIMS8q55hjGOrkKhRhJVVce9Za/Cmyb40R9H8YX+9ej3NUEN9b2nyOfG1mKQPal
e3mC+h7AUfJqqTPtmTFHFkOf4E3DA3JSK8xTXXByW8J33BcRjBbaX7z2XdKvfwQnfZ7Erabigqe8
LTbNyCrnU5a94seHjtssGAfiIO6IX1k8RiA7E+FrNSamPNteGuG4bh7ZprQWiKIS6RLR9PBOMqRE
suikEpO0/bIcrHlX/IX0SRha46TvaWxMEew8AkDBeWAnRyj4lWPzwKFWgDbfF+rD4vrbBq8dsB6f
jRN20LPR1xlcNyhS+cPM3LvdHIktZu4dE5g+kzG8R7ZAJSYnjZma9JTE10TDtXJY+YrsR+eM/nkW
fpWCWxmpUUrKwJmcc2ZDfpDeOGU2/cSQZK1C9wdO3yXkY2DXecvLCthWQzchMO5KGnkKeg649aeE
F5WUCJ1Z7KWr5zPfTgRf+z3iVU3G+kJ0N28YIsVs7wSODLGrE9muEqBf2qww2/uxHjvHM8bOWCAR
1ZKv7n6vq8K1NLKvVRW8xTffq32xSnFDFDsqOC5A0XoJ8+yerOb170VRTCSHCnI7bM8nJqVDHTw4
fOhyTsFWz6UjMugRisB7O27s3w6OtUg8rGgZhR7VuAMPHPU/4uxpTxXZXGtA1DBQ3G3cQZl/j/sy
grsd4opKveTO9RkDQ2ZoCKUst89Cg8wxfX7ESDO/TDHa4PjeZHYyCNhQXdqhb4HdciItJRBq96f6
gZjbNJ71ykKtdX1klA0fTdZhcmseQlIxw4Fzoh25qZoHkXwP2JFEm6XfXHOoL6+YLA4d+/NVOZOZ
PUXJmUXltoeyROwQj3wmP6zcUNfNyWVivldUtI0MuL5/226LGtTZhWQjw0bpBNvTid7275aD/Osd
lwBxsr1wDhOangZIIWegEcbE0RIpHq8Z8Ja3qqFfL6/ojXGr+0c96L9g/LNQiZTFUN4vh/9wzBWX
UCZALySkpdRcwiTriSnL1+LhIuCrAEIRz77He8cXu6HO1lkUWYlXz8qKWuC53PCAh//DQ+xyA35j
1XvqLsqmmFyCaPBPy24PlFp+QZ4N3QgDVAXMOld52qOH/onc7EnD6majYuzm9riG8cbmz1MwEnvw
QdeHzn7OkjlAq4eH2HG1azkJ936T44F2Hk5WuFUL9IzIQtEElFb7fLWD1AmSkIZeveQxrP+LLFmO
u5y2uPYKGnLeA7cs220MnNXRQ4BDntSylQfKbQmvlepqKO8IgruifogyZmYOihZzmjrAowki4s9I
1oA3DQzIhbt5YrEvdOTGSntSAm5+XMmo6bwpT+6PQPqXh++tVH7mgilmPpP3TFraEQoCThQILKYL
jLbtTcsfbOaRMp2CE8eRX1jbNtfRITeBENaDdO+n3PF0nRe1ijk/WFWnNs4PdasQJj5+py/9F7X3
MRZV8FlYfa1JpR/caFzz0w2FkdTHBHXTYwbX/dccvoQctpPUTntz4YbGHLdi915XgN5GVFfajRHP
HWmabfbQ1BeA0A7LVPA05wZQN5HLimqZ6y6LBQn+xM2JW/qH5NQUvgIycqx1GgswpY6eCc2KJmTC
0Yo01LpfvmIVddd93YXcBx5Wp3vwZvr/JsIpQuSAD7zZHbhvkze/tQr26+XjBXrKjOllS22Mh02U
jDH0OO6kEBgmMxcH0vsHVex+wdVCQH2ZG6nH5oniejRB7NdxtMdRumRB6WpbDBgeB7IGxeOYKxoB
r0D3nSOJzQ4OwOE29B3ockGR5VYH2DxQWDYjYUxBjytAVqzZTfE9A+9Qy8MdNtM13hyXgjVmhAdI
1egKeSMZz1kkSJIMUEhelWwtggd8VxlexeaME9PGQaJASsyP9owp35t2qnHch+U2fPMGfEHjRKDZ
8T7ILKEOgrZKpdGFBptG/DFjn996aF/zl+uBdRQX0I9LFAm/9NLPZOtyToUPkSmdlscxcF3nbklS
lghJpfbmSu9tqR2HnpJMbqsiYA3B/qsuRVVSMeRXQBLZC0ZdGUbsdFGxH7L1ot4p3plNRij2y55f
PuKAYSjVuum0Rl4PfgEYxTJnKC9qNTDVwDk5/AmWJo++M/4S4b4n2GR4xTaDFw2G2oBuV/pTr5W0
taN/WpEAGPfN+bzBUrB8mCpKoc6mfph/Jng5s3Uq574HQZ59H4zz0zY3VxKMXwraSXNGZY5ej5In
knQg2YOO95uyyALr2I7GYswJmmUh9DTubMNI6kDbDtkpGjZEOJ+osM4QW6HnHSuKMEEjnCo2f/TG
J2510wX/4ZJlYxG7kMYQblb7a+xsjIPVBKUNAqdsTb6V1R6+QzA0RkUVGu9syqurkyvSe088baIl
GZrOL2dzpxP29mTG9tbOlNUtPk7R8r203qqGvi9Fughsuz7Hy+jYd3WwhlQPMMDCk7Qqc3GvvsDa
36yt/sjTQnL/bLG4+I4KczN6c5mr43mjUf55diyMGbyXOHe+a+RFcvLrYmDVnpkzpvqKPpyb3wwl
N2+wNMTNO+BxBDiegKnStu3uVKE1vStIbjKD96S10EA7GTHUDpruA7+iO2Z+b809vMRWioBgN0JN
TbOKb2dfCPX8PplMgE9n7mhA1lRFdODEXE9+bp/jZEoyze3Qb28EgTojXwmyPk9yrLeepFR1kw4o
8aMtmMrm/GWRXwkTK+kUcDNFHxSEY2wg/UFy5KKkNQ4YVZZtmX1hyQ/CYLSwH8PSecylJCoWstPb
wQ+NNq7iz0/RB9PKFnOvDp6d2ZEQGsoEQXFJdRCGsYQSZxYqVcI+/pMUZEtWLyFXcRHUP6TZCev3
NiVQeOj/xsSEqUopXChzYT8Ir687IqbRxK5FyJdxz2zGEZ85qEJHLxCqzzwWkd7IAeM6tuvcF/v9
MaYoe3x7cYWnGIUTJG+EJkj51vtnXWC221hAKI73J+INDKGH9D50GRxR9AyVWJ9bpfEcdDYb83VO
3osG+XdBQyYPNuyNBbDzwItodmG2J3xxwW9DYFCP4/wGPyXs0q3655UYOf4fETd6/QydUr3vyHVM
rH+R+72tuRy5qkTVOv0DemlvbuUIILPmvk8STG8seIiz9GKDkqx1XNXIdNulZWBmrvyXgRMThW0/
wq7ijV2bO0prz3wz50LjcmUDWFf0rCsD8xrC5sH61VdiYv6wfc24voZf4UJwfu+h8YjOFGIZYYjD
eJDA3MPRtBTTSGXtTvZUXFQBiV6sjdemI1I30n2rrlUYprQtjOFMg0kx0n7aCTezX6tKcnzXJY9z
Nnw+CQvjE/f5mhBL0+VDK2Wc0k2VkcD6q6c71GayWeBMpxyIDp/8JbUssCLFzlMjcJyMzUDnjRSg
l2OAcBv2yfLX/UvbSaJGXQIRC1sGqdunjlgb+K4ZsQdIAZxpLKDVVWIQpsJbUq8K0DwJvy+nEE4H
by6wiJhF9ISepg+SQbnkXzvLojVxLgG1DgBZ7mho4Ec8PhgdPyqdwJzAuIyU+EU7fzJbYriyUptL
almOos9IOI3yKnWGxzxSX2Sk/KeN+lI1gl4JxJUgtpFEtnmB2L+GsmsIHdBM3hJHVPYkaYkUxUgY
hKoHJnXeg9Rzozc9+t5j6Hs3/E64r9160RmKc2SVknFQ67rUWPnjsxaKplwvsWA9Om5lJiIp/bwa
bkCJJZYRIlREr8zdk0UphAplEZWKYHYDar2ME1UELlUSxolhnPYjpWLkNVE9s9ReRhXR+cc0VNzw
rouyQpteX1pvlqjhVGHtbjthxgC14r9RYsvFE8scu1+qX2UrT5i7Ho67LUVhJ/LXoZ8ZgSlSk5FJ
RAyCTKbuRrVQMdXlhoOWovlUXmLs0ZsYjfKxPNj0JZ/I0PkIVNxH3cKGEZ8nwPVRkskIqacR4ckX
bZ4FNclLjU7GXqkE2ORyZgLg987tuiR954ldRxzUvmjNq37lVQZX+WSzpmbqQParDYLh39UEM2d9
bnd9mMwms4ZLG9+Y320Zbo4ZPHd3NVBaAV3Wp3shsh+SJlecr9TjGsKvZXsEdeUh6GhFopOzzWBb
gZSH3IbvVoNk86eTsdV7XbSevmkqp8hVcSGenTfrOk/69rKd+ZxC9t3Vjp5rrv8TxLw/milNSddc
eEtt93WE48U/o7dxsqLyR3lGiWKXORilS0OZtZGr6ZNOA7NxpuXLoGEgwmORWI5iVNr3svYnJfBU
lMuJQM9PwsFqoXXvdtrmPb8m64P+a0UxT+McSoWJf7o5frZcxj4uaimsFqekivPmYqkbZPr2sbCz
sjdZ7AeGq6jMWSpyvUYkWAEpJI0CzeJy0S+XcXHriqUVwE6ecBZ6hCC+uJlXg5qqH5Wu0TVzZknH
bmOwmUp00/o1tq1Fl9XuvKvpTIxpbiyavtM6N5fknwa5Zp36YAcqTZXxrZ/ApJl5DWIMcX7etbm6
ULGb+OJEhS0Ww61VqH6HbdSNwJvC9A/2JbK+rKLYgJaduwfd/EtjT0UmbhMWDo9AfdjDJ6/pw6Yx
niJCjuJFxzehXSgTt0lsr1AEkQZLLre6RZPEdmkdIJcHqS6j563vMiBYJY/2Fo83qJNHkv4NkIws
lpe4Gtp4BXBZnMi91Dm05X5ejFdcDu2hUxD7DTcAzH1AXxwsfnAPplw3BlCrkVv88pcu0YnuodmS
qA8Gssz28YzV6E3O+jIpZFrBhELfTfNMGy7hJ/qeF2NW9JDbIbxWLteRTXlTLYSkNO9NYBG279Z5
4dIjMXH1xXEThaAk0TPw4XpJbSxq5wpEo99sLL8i/mVOXcuPsXiKPEUsvc6i26nFqPiUT2jjYBB/
pcJRp0p/ppPClRP+EVoe+YP8lBNkzkIncYoCSz2ugBetfDlNV4YjT7D/ZZqiFjZt0AeNArkYQOvk
FN5U1Zu5y9wsPFzKt34gTBw/xymjFdYRDH4Eo6lOt8WwQQBWIPO7LUg4d9fFBo7iGIKqOSBv/Zag
yTZsIDg5m2A+qPYMWuUQKO3WZxzLfKgAk4DpWxcREwttmQru/exWAOtyY+eQ5Yku+FBfuRt56YcY
TLrlh61IT99MpgoAqyezhwizgXEW+9v8bMasxX4H66YqBdfO9POR+vmbHSs6VDsDZmQPfMeIrnr1
LMqvpaLu/zuYTfUQM7EmEYqjIsItfzTDTyA3/nzKz/Dj+nR8eJCPX1tisF/12CODPcSNPb4Fg7bK
t/+XgNdVLUQuL6csmIlp26ZdZQ34mSil/FJJg+lIMMhnS2iD9NKVhrGq8pNzfwLdWVp8IN9fCXKv
OsydxX9fS43KxKq5gYSLY8nXwSRHLPG1rV+5n17GRijFFJMunkOTC3acOIH6FT5feamk1TVmKY//
pI6dujkq+gCnuQj6h9zsTlmIZFkUlAHgaB1FYyzwtpH86/Hlk5XlbCpZWvX8eCiNFpQhY+xLOIRt
t+L0IacgB9Ngdj/zgRq7KUwoJic/d0LTzFtn4hSwlYIcNqDjve5m6OZdEru2/e25ukpnA7NI0DPe
SdYqrSz+W/f2SbsyntSnyabVMSVghKpez7n2OLM7H7c0BqvOPPk0ZZM9cLwSvlH1ENWKXq+WDJoN
GKhSQO+Op0z8SsA9l4rKuZf+QtB9y4DX6m0D/grBen+GhiO42dq5+nBqdoKummMYKnDCIPxfU8lg
03jNqbpWDqCMSQdYf6Lal3kUOYe2+Nb3ifFlbpuOrqckbKOB8/2j8ypBT3wuGE898wqSr9pKqmnq
WcVN/3wfG/Qzsi96HywLVo349I5bGzbixjTjSx3PFLdABOXC7OkJz0RIqcOoTvDDCDnEt3oNFOl7
PZFb9Ukp7mESK8wfcbCVjWDPS16tYaXb7LioND7xFKUvKYTIZUK9hW7lOucLsTFJ1usUTmR1vuaH
zRSJfyI2PtD/o497jfAkpOD2kPvgJMPZyLoJu8vXmQy50dsseuan3jGZfx/CareWHy6RnGE6lXcx
cckm/mkLN15PxsgXd9+tyPyLwActbCOsP3+5XRqrUKDUlkOVaDfggx+FXRpkXQGM8+tHvbtQhNFQ
7jzs1QXXCWuwetG/Ay8gpccsJUDj6CwJkwPwTzOefo/HBuNvqfwKk9r4dyVbUSWnz8lI3c4UyDrs
YmPWM7vstg9LqXvkyK8XvXPAG1VrCiaPRZBMrRXMKT8lHeyoCA5HxrV37560uLFPkLKlSqBlVbv5
R2w6HKHvP0lst1/OLCvqqURrvZTQFlPosuSAUbVmU2c/YuZXmRB/ZVSdbtfPalfcr4RkhptRF1kQ
KLN8YRQf83Jb/ARUXrpCOB49AwREmkIg/+DsnIYBPZQ2htGrgNtfc1Rm0JL83/gFAkr3Ehdk3X/6
E6f3XzOttDvu9KE9ecG6NWq1GjA5yROYk6pWI5Pujk/MSB0RYLZROou7Dtcn5lolWGv6IjHogneY
DNyeEnCl2XJT8NSFs9EdHAVJUoQNTkqAIXXT9Vkbd8WI0l+hfFgXMlG0XMSF/uCHmNuchnJ7mbEH
KwZ0Lj94s7c6vnqvZduFxBacHzkCZpdc+zL+lCoIUdFi8eduzvLhZHSCXY7n1+NBrQVlrOxcsjrC
0bfaZkPkPLWU2Pmxso/mUkf7gnDC/mWJfnPSejpRyFfPkGHH4kWz/yO2AWDmtRk2xxGXmX1OnKOh
P3GGMaJJlxTLS/g7K2XcU4GnFcrjpXRkWoiC/cf6C5tQE0uAOhZ4imgh84xjkJBwK2EbgzE0pb+h
UiHBhgE36i6f4eHwoJyXhASMhmsH/ZXRj7c1UUf5RsEiLDHv3umn6kTsMtHAE3eIRwIlk9z8tZAX
Ng09/LJAwrokGEDMaxxOsP61B1UnMh8DOOvTimH5AZr+S5wh23Q/DATRC//lbcbkG0/4fCxzStEM
gBevsgZUBP4xU/F4A7HkQvx//aMrJJXvC+2h6oW7EBWXb6R9fiwYS3rJ6zlhWn7U8rZOg5NOGoTa
gjn9h9GuDx5tcIuFcbaoOj6RZHfrWFWhJPlx2GJbkngImPT0wgVkemXSMhgFJV8XYJmmNL76srkx
w5Ri4oHwy22dHY6EP2BB5k0VOs0oFtcGWuHN73B1IB5R2doAXftvjiCZISPtDIK2hhbspBqIYtyh
z8AG0cW30C92SdEXTjBqvDbelT6WGTUOxRW4Zd1J/SwmOQTjxL3rvGDDUNcBDZCgrENZ4RvlpPT3
3OutPaslQmhD1ivvOFGi1J7t+mLkep6CUKxa5h9ruTOsLIni8m2r4K3reNLAEIMDSRZnZY5pHzpY
ZRaOuMlJ0Cdevn/MPmykd5C6t0s8nJH1eGwJsiJ8LcvrShAx/8jr4YOoil6FRozh6bVB7B84K5fU
CkoIvU1TCM1v0mJZ42WSHQgC/N0lDWXAxqFTcomk0Q27qUrs/fX/mc55bM0srV/43hjo8jEeJtXT
fFcXZ4nqU1Aa0ecbpFNqTBGO80RNEOzX5QWIuOCHzuQdZvU8OIjmyEu+aioJnU7PENaUCr3U8dl+
wluZ2dgCouOFCpvtxJMN+uP4jpVbNwEij7sf8JtuRVTQ9v5NCSxRJKddnUZGRvWbqjfPdbeq3tB2
CrzbdkXEtNZpWyMFfNJuUjiISCUOcwob2EGhF1FBYTLDsrmK0/Yl93xVWx4Rha9Hs9rTisfql053
qSmrTbxTKG0buSeKvrW15bo9IxMESDs5dRe69964wYd+IbxSsRzF6R05GMAOREE71phqB9PUs80N
pKxGut8yRner5jkFhwd1F83IcMU1rVV+Wy2vMmH/7veY2u9aHym9pqUBCMK+nT/ZdHTZnxGhfw6q
e/On9R1FZfXgMGBa/O3w+Rfn54oKJtfpj31Ov80IDIwUpDDPNPYYkB4RVjE15RUO9LNCijNCJTwn
r0zCJ/GFpUAkoTcQRfBIj+eVCDystikMK/Bo2qyY5T7qT3as0ZamlpR0tabYPpBcwbcXDqOLNdbQ
AuECnenNcDWFO26K54HVpAXK+jFIDoFTw9LhEgCocu3hBlg1ccVUnTgDtqapKtpfkLGEDAl1dDwq
p5YPuzHUtzMTAfoG089Rn7fLlurj3W5GwpWyBxOFeiDqShnOrOdDbocMdud4fw+ps/GWJBNJT4PM
2UONm+A5DHAbiHYnuOzX4Js+PCccLlEAJUSNrtXHdl5IrjxhT5eWKuG8eZdJg2d8mg7j20c2IY/F
EgtBG4MyPHmaVOXUmK6U95F0hg7QraAy/IZ0ySg1yl6qCxV0KAxR0VzQ/m7vB1Kqx8g35rOAg1Oe
h4OjyZ1j/YzQLCbxa+cBO5tM302lAJ1hTpW+gx+ReYHSPXpIB1qzT8b0hx0jHspGBPejfhRvopyP
MR5jI1REQC8OcFRt9sxgId6KHL3XqSU1jgofYPQyCJRGtvHbcPdpsWcGWasVsEr+65qTClNd07LS
TY2RB1iFol1ZOkA5H7LmsnIFiCEbXfdvoZSQdUHRxoXgnLzz3E4GTvF0UkP8t+/5SvUqe5EV35Pt
+BmmtghlJmAZ1SOpuOT7GYdmzDtrz7pb+8LgmwUOg8fGoncypzkiLz1bYe7gvSPv/Z4VzVe689zP
h8z4e7LSyHtjHucWo1OH5uHI/sX80l3adu+sTxJLmdcnO5EE9q7wqRII0BJflRyXULn0HzBzIjg+
hD/jqHHIRwtCpmjjXFPyvnJRCugc/yjs5omcoUu6XbcJMqGovECk3T4Wn/H2lY6MksxADvHZ5cC2
u0Wq/cTM6TnCOo0wX3opDIwXh4D6w85zdlmNE6v0foHOV2Umdj7zAeO/cE+H0epmKEZQC7KRz9fG
vieS8luVr34UvDPloyH9KwnNauCmkZ3tlBVJaXSGuj9elmJOBW/emcOly5oim4qo/IVl2a6yKLkm
o+8sFqaAFQ1LaNjSi8nKCXv1H3ljDR3ualWO4IfhxKqRdlJosV9w2Fkj0uhjxndrde1A2Gxu00vu
7N9vAsxilxdyLXV7H/DO5ugTXohWzijJ5ujh7cjYWWvHzgf8c9cSdWJO39qAoQcQvoTEbXpg7ive
v6jiQbzsdKhpjBLq+L4O4PfqAMEc8uzBR+3txC8evhSSr1xoEF74Pe+1rHYZQi/lEpRbnkZtLGnU
MJfDfQntdgHkXakxBrOKDns1BY7b/JX+AWjLWEmEvy3a2hDHCY6RMMXsN9gl9mF5AKStEzUClkcw
EW2ShmuDzBNIocV6MyUX3GWeYjETlA3qAP+aNLlQtpEAy5Nry688Yv+cwTSn1f2uK/UbfRPpQZCm
bbfrtTp5EEYElRq9ykJ0hCtm2c/kwWsO4RlMvZnNzmRHdhoeIMwMNaYwyah3NNvn8CUthEQCFsPs
eOJaZ+yaQiWZyduDl9Ts/Ks0IUimcpaK+3xTmmLW4aNbRCGkVgZ40L2UhhPFtRZJ24RQehITygCm
NBJay+27d1GOMaQpGLmq9wVo3WnW8cIASV3urhPgc5qP3dt411oABC5Ey8Tm8Ue+hMtdL1x8TDab
gJtP+p6jqKZQIkZxauwxWx2lq/hFVQw2/uUMwdNp6+sP2P6zv1d3kD778UJokwX5LGOvDcWaIIUP
m7IhgCsnhkLlyP9ZWZSMDU4e1/H3weRPgjNSoa94Y1rXXuZMPJKxmFVKoB2XlbpVkcF62Nsa7wut
WnKh/EvKRMRcDIHBD0uIM1dLstKZpP9OACbNLGMqR5q4MTPozuTJltvuoPgPBtJo1M0ZBbKK6t/L
6qRTmFA2OfyJ90bIOukFNGmKGUmNapCJTBdbk+lSC/OP+g1NbWLagoo8ha42iUozUgUqhMG47MFD
SeASYX3Sl6v92N2px1vBJF/DDN+BmQHXk2ErnRl6C4VXeYFwiyv3NfToFFjPAXP21EKKKOLVyGyH
QMiSnQqQB3U0sHb1ILrTKG+uwlwR94a4yaOVyGWx1NonVlF7JuTvpM/NM837toeIoNLNsI98IdY1
paGD4XyTCQSYwKOGcCBJSitNJ4c7acbUo9pYnRiXlwS3ChBI1acaKHP8FHozRYtGzgYjrcOWqj2r
inGDJ8XlrcxjRQCXVqTWplEWbKTywMMQU6fMf71lbINmuNmDIup4U6b+ZqgoHYDY+nm5IT/J7NIa
+sge3HpJ0xuTwpvnahsjPpWHk4DwGVeGKYm5rqVJ5KMsP+fnrxDGeDbeZKfjN2Cv3m5a60gRoAvg
5Z3/v5Vh8idjXGO6ZuW0p2e1kCyNq1lWyRqvUrF6KQRr/eDfxRhoUIZ5Qz4Dv6uO5WW2tMu6D94T
0O7MResmc1VXkSfYfvmnDHm/q30ZfWyYyfK9gzfbhhIBptWp6QCA2w90w0/nZDtPgXwTtGZUm1CF
XyOI1Df70EF/rMT5M3X1XLVKrHmYVZ6TYP10PiKVUF3tMoMJzDjeMnl0xSufTQ7CSf8kZXjHRk3h
CUkK0jK96QQRlu1LgM83GXKQWNmAFzcg/VejLs+x7yXkQfMrT7Akj+pcG139VvJvS4XLqcASW5K+
uJ5YP7KiE8MfMOO3R2ELg936D344VX55ebywwsD5t6/lvf1vniLqbetZc0/ZzwLFRTnJQIhOEE6U
t3Fs0uujctjTxyCUMISNAHHYb/662pLb2v15QkROt6f9WHQ2ThtA3PKr1bmGOvi0qXwih+Dmks3d
m1diV1Rmti4ooWyFxVxA5MCKWe/BuAGBFSvR03AMUK6FMTHAF/yEC6qjQ+R/oaS1qCfprh4PNl/z
UzleICVVH2jl4ea1Cu4m36Tt7AT+LJ1bsI6CzcM9W0wpBSOCVgvTzVwBagNiwbDm0vZnmTp3Pn7D
krAG0uDI4AeQOj0B5RHcBTrpUBF7h2t+ZQNaLp95CnEhoEQyXVmaEKszhZB7IKkYlDxcJZYlv36v
fBP+4PIACTZkDcjD7UQIA40GooOKW1IsUy51E4ZgIFiGBlbf8YDXjDS/xc8Vm3XVmKGXyRIqWGaM
vwjdFe5xfEKl014wbZH6l91vWJCxepvKhPlDl5nJiQyS41WNehLDe8CHvzTlGgu8SK9anPTSZ+Pw
iu/3hKV1kH0Io2Gn4VWhb4DeN9a5Vue5wO3Fl744zzBmWyOzcXHGF55gJ6gyt3hbgYaVk8uisiks
p6eg85aASnUow2ScVxWJg3qeM40t4NP8RhhJ83y/98f1KU1c1ktsuYWoJen4tEJYbK+yPihjyQK8
nZ/Sm2QBRl1Fn7LchlpzFjLXtyZ2axcYd6OECyqUxsGP9kvNUrGrp+NIo1S/KyCLjfTdKWR9NHq4
/bToB9DkT9tvWvws5DcXaUp6nyp/kCkOuwykM8JJIbTUBxyQ+YehpN4Cye0YmqYHPVmlhSMS/Pg5
b5I5W3q1qZ3Sh5hl19WSotRGGZmX160NQAScvEDsKtwOaOHqnb5nATxwOstg1P1s4kWbOPjUElx1
PNsviCQEilVVJEh/NekDG9ZwyjkFJnyqzsFUpnC0J7hZ+/D8SIVKp5GQrKZfn9syvwWnlfVzWlTw
RiSQlBSdZyJ1xTdnlIDTkheHpRihXSrrHBlJV3B99QFX6c8deogDpQh/LnNzKIA8bXYtwI1m9RuR
1EpJXEH7cG3leRxtFTmAaC8dTEnLbXaaADmvf71NKKlr/APCW7GfglN9VmfC4oiBbdtH7fGcPs4C
pnOWGTzwzdzVNKflTn+njGYB/ZbDmxR0QO/yT+BtOjIvB+ywcAUjF2XlV7wfYKX/hzFauQiZOser
JctZ76z6M5QsFSI4VaRXEu16qu8bJg5W5zXMAJX4+dfa68T4hipSS1xxX3TjuAUTnhmLpqf23ePc
un9AKqibKncm/sOHSX083hUwie1nlls610qjS0AI7OFJalhLtSHz0fNvG/yly+zaD2UMX88J/Iur
zDYaW7ix1MUbdJ1z9MKrHnnZP681oAWH+DPqM7ufRnPBN3x9lfhApsNlrsYR/XuslpSptHvb9J/9
NSNa1cwLagZG0hYFFlQkqyQe3rwvn2e4P/ZFfOuziOdfGJStyDH+raLLIZq3fWePbYr5AnxuquAE
30sMUx8aZzC6JpLlHO/e/NAi9k9HA4sUtn4kQi4+z+BD0sPUGqUxbi843ZK1NRxU4SlUUMUYBFOf
v/etMF4df8S2L68J0ikegLW0yJKYP7jt/02zwbCddF2PJxHELiwXaQLCdv0ZmAl0qvKmgCgYKxWY
zC1PLJaMBdjuYJtQpDuWUtG70Jgv7PxgEdL0xrZ3Jb9/lA0M7nFcUpHYWfR+wL780e0DV8AMFPoL
WsMnjyiOXci7MWB7CZRCDA65J+M/PFRxsDNv4o7+9SKZJLLZnCJvB7epCBsHx/Cs/hZP61+LvhHS
g9ENy+3y415Hq9TIGQcCK0cIBDaLb5A9y6WjX9zJc19sNaKwTniCbU61xbEIURR5tscTzSoGISLH
PchOEoPxj8C6P6XThdTvLjYmjLeXzrlq7LzGXCy/rcVxoa2pF0H1VlDD5//Qz1OR3WdxA2CS0ym4
eq9wCCRE1bstYwKInHL0BprG7p/5OQxmP448KJ/BZY26qh3a88/HgBzc6Q/52V7Po3nYOrOcGkYn
xQoCRTxppXYMqbkmTHOuSafLG7GH9rPhC57rgb2HQncfNnFWST9acKtNXFteA4vrQggHBP+rkJ/a
9uKPolAqQgLBhmsAqUiuqZFD8LzAsHMvfyDH5NQy4A7xhnOs+ong9WCNnbE6yTK4S1qZI65q1xS2
jzS8xdoUbXCJBH+nCffgEL8ZIiYkF7CeSo6VJmHHtxIiM85zKSTuAkWkLVW5IIhx8Xh54zZRcOm1
H+K9pmrb2vEsV9Nt9fROm7KS75sxqdZmaTdDcay3eaUR+vwufHkb7zloYM/nfE013OByU4o6USri
SMLSRZcN/MQBladnCiWw/e6RmU/UYhjPu+x7rwKfuEJmdWT14XN/D/QZzHK4uljsZhjJ8thmOL7D
h3D79V7nhNRtprhd7tWGKR/o34aDmoP5GZsi2lZAQdHlcLmmHuPR4Ldu4BW5eX6U78XDPfyyJYkS
TIn+sLYrZQANkmcrwOneDUiUI7b4VSMNsTiZFu8rFkgrMj6VN1qmJJFrr/Bb0uIiDNqUtJy2TlGx
vLbkmKE6ROZ1Tc7xxaPHqaqceImW5n5us/9p2EKHZgEtrab2K7JI9qDfbDRH2r7rvoHcHxq6eCow
l0MREtkvXKGlKAbqfduDGw8tqnua1tS9H3h2NPGIOitsLOvZYemA6PxQFKEu1qq0FgqAAhdc13wO
DwNG5jGh1rAc6H3WTsePRU98i7opzgplCNFYxsoUtwp1uuS8AhQVwUj99G7toZfFmGxr9gcorPeD
JiJ+xpI3X8ko4jKmQDYkiQy7H6iJyMUiQozrc8L0kT2/eVDAkguVfuhFH/qSGv5/NgR69hZ8VYIz
uMi+YTzXwMQapL+7bOH/MTyWBiqEo/dDJrhgVZg/2ugh9A5092oyOq93reJFhSt7z74mhlepV5l1
EnLzeKakzckw7PPpRuIA0F+Ymyu/CQUccQuVG8cveoIgTEs67tjuR8cuw6ZHTOKmx/ZLVtDdvs7N
whPY47arsrkCJqOPZZSBuUMki3mRGTjnlDJvX+dP8bc6uNrqNKtwi518bnicYpM/aPi0VarZpROd
4Raw9ovoeMi+lVBqPnjZSi9LGzldJuZPrkj3xT77b0IazuDWD0m3foHh+MvQlKDcyjj0xZ2a+JQZ
AWbX59hgP1w0Qrb36F/MlOZOZNZiNghgDPlIdnk/6Y3JqzBk573oy86NNBCY/2QeOklYZ4ukhddy
pjMqdfeVUMpHI+jfUTZYD2g9SCtnAR2Rl2RmgELrMTug02hEhnv1SvtKY/7lsoJy8DT0nNJ++yLZ
uRsvmVs+XW+hRsNZFZIu68pg5VkXJ3y+KYuUWpto5nc7oV7SmXneT/9WbueX6UHlEFeWEKfBzS1h
yjULX4QjdtGZ2sHwjJW77CenBsYtqCRlJbLACMyLryEosg4BXx7aEv5RkAv86BUVCT4DmK9qyGmW
KLvC9iaXlO44uPn27YsoY2Ko4D2Rap1kyHLfcojcMcpn77LbF8vUL+qzps4EzFQLslihuWJPoRAZ
tzV2l/X1vWCj2F9mGuB+N5PXreGFCMiOuvIaoYV1MIWpZZb9Q7DFW0lEur5PdEhXNTNHNmuZBnw6
avxQIVHlzlQywMEX1puEAkvYi1xC1VbGhc4ufgA2sotmqek1pqREyTRiXLJFrdo+eFRP4U8JffxT
Ky8j6rt3ePblnwn6ksnH4bIvdH81sv7UrH/PS2t8gwYxYv+sXiMFvoXDLMqetUoGIFJUyrgjLY9I
QVFlFC4xZaGmePA/zd+GPh0DeBzuEGlFEYTev2i3rKQWKWv5iNxFMJ9x74N5frTnfnuxSYc47q/L
DGFE12AYQpGaGY5hfbMvQiPKKrOwhX+qWzw/5NGgeVa+h8YZX7lwJKNi7rd4nDoMGTfu7amOv2SG
UNdNJlZfRbMDchTbmeSYO//AU3vX69XVmJxSwDsrifj34GFwIq8TBJL6aoBGTlGIyyksN2+w72AU
J1OApgQ0fCoYkenT42DWgL4QFW60MOG/z751MYxCA7svk/hOCabFrYGiIiFpzGvdjLWG152eJthA
XNAEalsZ8cc+m/oQ9pCKg5VYBmEh+Ah6fKJASmqOx+G6lzjBsSphPcvtbPezVTXjMTqXOJCJAaZW
Xn2EAQulZjCcypD0TqniqicGLegS/MqppOFZAxYr005SEO4j0sXzFoDOVV/xg1dPgZN/EqOieLbW
2MUU0EKoy1jJ4R3mkWOuETTb4lSLlPEbPH0ZSMfZTSpT7M1pa77eBveCMt6B2NysLk7NbZSYBrPU
SV8gKHD7tYrTJIpX9pekNLfj3q5v8zLkq2ZcPFH4Nd9B/PjaVWLdmPU5t1tPcTTRB8/bPwlhSCNj
JSbk5hSRU/Z3Iu+ZUwEhylPXCpMGvGrra6jsUHX6bvaDLsLl6mj3sX7TYwqtJAh2QAT0+vffopHy
XXgfWlYl/dMQJu3LZgooT7pA119p3dT/o5vu5iu4FvYE9B5idAodMvsVNTbudX5lP/nZTTwbTmPO
S8vbSJg/8/dRTADXt1SXL466SlAR0jMmyrRNo7oFeECZZJ2myBXF7+e6smiNjPepqFptjpFE1XT1
u15iBtT99dsaF9KA9nJZAPm5hOf5X4M2JMPqClPU8lgS+ayQ9R/GpxkSbNNudu/rXSZNm1OBN9Jm
eeIPpTAWQYcFBmQikL4T300JC4Dgbhun4qaGJxgdrvo3OCUxlL7AplwLdmSJWmwFb65/DEWxMPX+
/5v75PCx+wnZHT8quERUM6qTxVH9nwGvauNKm3L7wT3WqAs/ri78NbU3cxm2L+QinFHkQWiTKT6p
kBJqRBivX9LuP/9bm0rn/UxarIQajFbsbvcgvLjh6N2ijNdV8bHhv9AyDE4LmvXYOcErfW0lfjaS
o1Y4qyhnPuYtqaO9pIDzN7seEqVk0/ANE5PJQwT8oIbjDnDN0rZG+AtIReYP7dN6GA6apUK7PMDa
oSeOtYXu0qlSX3oeDuyikZo0w6hjzpKeLuuTmitylBG+CSuh7dinHgQWCYMFKRTlq/oxm492ihq+
uOn0s3spq3u0c8CnWdDcDBGh7EStD9wvegqFz7uVTMsigeqDBpn+Bb2ggmAtHCTVzcI1fT32TdLL
UNsTCHs+vPVLT9SU6CGmxtvsUPiD8On4Wnqnlm2r4h53zkbXfmnjxDX7VEorksE/kGrO1q/XUv8P
GQIeBZhaC/mX7h5ZkHni6VbBQpy8voPDQ8FtyuCYY1unAYzExYwKtNXQYAogufu3DazCjexSOzYo
fSbBUwbM6AfBVn3c5NSrYSTZDrLV6RqdX+uZArJA3OR5NqBejH8b7eOiaEG3Aw3ENZzlbeA9Y8vo
UnbTR+BD/3ahdGb4YbI5DhPMsZ3n12juBgrzFI/Oh1u2j4J/wWO3OsdtnluOgKvkLAd4GcL4vAIl
zR2H9oNAcv5Qqx1aP/YhD+WlygDA3xkthQjrhBZMPdRMVl36tL0DVnpA8L8FTTPIS0+YgSHmnMX7
Jy7nUqIpiEpDKH9CdtqmxfraHMOZPYumX2eapSM1slIR95NKI5qqBTSY9cH5HDSr7U8n2KO+Iedc
GPR2kdL5Hj952D+L0C3LkJ1/K2ONqNcQCVrxbxQAO5NEv7X69GG/eHXAqeJOCnh94f+sc9H8U2CH
YHFHTM6EKfI81LBzfrKa3XafbJzvL8Dr0gCHTsORBcZ7uH3n7K0Pge8yvxMInBaeBUGLIeEeD3Pr
udCRRH1RvtwnYOObCJbc1xqQqTbBGbDVNByYsPuc42za1UR3h+fFIh9KD7361KQnTMW7eGdmokfv
bem7l/KkdVdolWRXZUpStW/l5nF6gcFMLZQ930sA1H1a/+vD2NMQ0/QA/LCn84r+/rvhGaMNLXBi
g98yC+H+c2DhAtMPqplcrAMYCS8ok/AvT15mS3hI2+fTBRpnxYqQHFrXATcSDOXEffYQbdRqN+kB
lU7hjZckLHkr1tDB0O5eZwBvgoHQCGf/lkXvfcLZuH/dKTl0vXipK6hgbqupYa7Ow1NiPodzysu2
uGMjJ48CPebgE9AWcbyvV9c5Ez7Vbl/ppmuBFydAHgP4+8BuZodU+TCYAR0SendFnDWYjchqQ+GI
eE6xYGcCvYqLIkgODzn4FeUQTNmSoskDxJRj1EgfJBLkmTS/Sso9GOAxUg8kHIE3mEfpWtnlq89/
8xMXLxOb6O1MRse1Skjj1cVNZgHF57iipaDfeksXyT1Dzj6ZowsydkorWE0kqw+BQNALjKU6tY/F
mVoeDYHFI9ASElW+8PWumOwqNT/S8oK2O2HKDNMlTHE5Erp6BF6Upns4Uu8Zi/2B20Wb5m891mX2
2V0jEfregYPJtwnYXvUaaReiLslEQbkvOLQYtPCVsAxwrn/5NeIlNnynBbcxz/HoYL1Vm2/pipnw
742hB0MFBIMKiFbX+o4d3bpp6Jol/MvSdeSxpozILOEMSVhkF3K6Lsc2g9A4dnXmEWsxlrl0XGHS
TRlpC3s4o467ZCvP/RAkzvCJduQ2Xr5+gyd8c1mEfJQW77bj5FagLNc9t13sCoN+GFpLqGdNgpU7
NWRulC+kV/Hq8KuG9KFQO6DRkEPo8H8JHZyMnghJgDWogqDHqwYVTIFPGhMVunfvLoAq3u7XVVK8
2PP0Mup366XpNKhNF7enbBe2A6qo8ZCISZUsJ6353eMI1QsLs7lE2wedNB3VmCx+jPD5jsCNabMT
3D4LrITKFKf4c3nBh2jo1xRShxK4p72cXeU+/7RUnUFxzw25teAN+HVZPp3ob1kKN9n36acofrOx
V/gUxYSHuM4ZH7b8tPH9BfSLOHl6w9+IwzE0uFnwo0ad3nrQLcz6VgBOeuVaL6krH7XqWUChnAN+
0GCUIKEU5VRvUteaa2iC4+eiHuTXrWcNXnXP6OHquDjfAJx42IVMcZ/bZjm+ZPTnGQx35FQTLP8j
3Oanrfda5F0dqtyrbRubbmPfM7JYnnF3oyhOw3CmfJ+h/0+DjWwc+ryjX99g2vIdgCiDXntPOheH
25px2SHqAtwx+s+gMGFlQMLq2GcvJndiKMgoo5UJMj2o9ULCnB3bryElMkprmMLXG4VHBhjPzwOe
wbtlCoyHryqrOs2oJwycD0H5qgDHAoJbdjPTdxADHaTcS0DoBMPOo2tdYJeLb/kDQBDnF6kp04RH
rRdpAnSR7lbp396D+AX6x1rNfamhuYG/W+wnx0q4xnbuA46yG9W4uR78TzdPI10e/DEowzzc9a4s
ZGS9UyJ+hR9MBMjJJqXdMAfyVCZSbN7hQxGzkU6pcdenga9MOGijagzeONSxYyoZvrGuG5ZLahjs
QPNNk8NPzdJnevzxehVV7t8QAQEUk1yf1VkQl2OkSkpRdn3nNv2mewIpb4peQz0ZdMj9MNpKTSHE
qmWmMJe8vfDeZboEEWCYrl9kesWZL0ebn1d+HOsa8xUoNRr/apy7Cm22yFbjiGiJF+1GEQQ6fZyg
hma9V7JqymXKvo0MB+UW9pMPuLe+zvh33hZ6jtykoZmzuPUjvKdhlQ7419oLOY8TLtjUJZiDbW1i
U/P9aQj8Wh/llcNa4UhE0PYRK0UQo4UnMLS5unxB17VFGdSww9BCKuddW7PLWh+vVEMmcR82Zctu
WZcXV4/vhZQmq2C7VUb+Y7LvS/jAwRfF2KvfZzjNgtcaw6V2O9w7DU/LNWlFeavw+OYKUcB739Lg
y9JGlEMN17btUFE4JpjptvhmzI+HOXQHZAzwLynPFtjYKoiQ08WQjWCbjQAoA3xfRIhyCO1W/vOz
VvCDWxP8b2F5G5rr+rTx2uUMh/xfKotZ3TFpf9JtXK0gGqlZ0HEMNq4bbzBiAIEBhPgKlLVUyvG+
oKU95I5/WHSCqmIk4Gu9S7cNIxfI1FgBh8I0EacpLKN6Dymqa17fS2gf4yUlop0N+qinVUGjDECI
BNJrrjFQxy/TU91HmPICX1oVX0Pii4U8gV21W2CVNCJAG3I++Nxcf2wJEkZKSbjqXjtamkdWckF+
GaEAahgIOvth6d4/tkU/bmTG0tHvpPv9eWPyx4udplhaenS0pDE16kKUF84BSKsdcHdb2dWJZz98
eQmF4lrqJJaIBb1H22f+2wBYKypF8919b0rAYWf/RXTEvjz4jKRGi49oLCCzxxgyLix1R9qo22er
yEnczy3Mrm2FXRDu7e894SRiVnM2yVYUIdCKmFmkh8xtV0DNkItnwUfo4dhh84pUoDuwq6cD0gKp
CMHB87sixDonHV9tppxs1xPUI5mW7x36OycNgLxmZezKczb3TqLYr3KNmaw5rPW5SWwASyyQOHYl
fYlzSF9IJ3HGA+HdBg+XxA5UPyOS/V28Q6AITRENvoS/TuLh9j5bVQacOWWsOXlpsB3wdM8wiYVs
bRvDsfNtaGrIhaCJ6RYfkOl+MDCSKcXw44evuZzi/8Rt1Eda5JgzOHjOSQyVJaGZ2snoaWD5Fh0u
nCNBXmS4l7Bqlc4rM2T/gzIeP7iy9/H716u7WnxKfRKwuw9e6S16HxmpwswchxfCMwARKgZAxfeE
A51s5YjH7f16K/gfOyZvCWvp3j+f9VIPq8rDJ+k/jSc3nMxlEWAAj4ja1YhJPYiJQCDlKWZE1reB
jb7lr6mU9J4zotSvAnNRH1L3RaKXYgRakz9xfGeXP2QK3rDhbFpsGqOc+DgFqxHReDJA6B+pnM5A
LJi028X3qVeBd1z3iqYFvzIBwgHxVyRvXhCaCcX52K1/29+deP4zR4Jc+5C40mPyj5tgzKlwBXAS
vETqAv2IRM7poLSLMbt3Ca0cZb8m7+xEFYTc0e+/36DWe6Lmc8k2gAmV2AuCWMb4ZUb7RDZ17eiH
Kgd6p8xODA++qBg44GOe9T3XcsDNHc9MsAxQmbaL4HSZYS8CAlapOIVlvez+xSeYbvy1AbRdLNzf
7hH9+oFpc3AbxfoBdkRrIIiWNxSed3wL6jPedlTp0eVu5Auf4eORSCTyk/5uIHNkE+HfAKg9td7S
mOI/G5vM5LYCyVqHTDGrx+B8WagjnBkKanmgra2PA0Z35SvCUI9r7jocE6meV0/JZkHta6f3Eus9
9iUnrc9NjnBDNtHZa3+ZKGKMKGWDOoPdhKSQWSpKdDREX5W6H/2MElko+BRRMhKERZPjE1eEHZi5
C3eCn1KVXhfI96EEV48/mzYmr7Flu0Jt6g8pP64N+lHXZgQu+9BqfpbbvovhDsY0kASSC4RWog4l
mkXG42V9JErlne+yD9YbLWdjrLTKbOOQSUeSSgMNaLQjubWAUGdebfhpsXZHziQu+Lu4ualPEst3
7qjdoVKIiuMmS8ZUJ50hxqLfzCpuJRo0rSkO2sTGwS2znpIPYEZhqBW6x2B2AtE+4Gv1XeeRcbOU
oG5wT9EZVY8/gJ4Yk2pRWxQBJvs5vYzXgDV6Zyhm+RkWhrHEufvpIi1AF3Lj/zRipgRnv4PtMfII
1c1gV6dVfCbvbHbngZHjrGpw8kOhtVQfmE66CPYf2C0O+gKRIUhtddihFAKLUEUtWqt6ZjChKbOX
hnh8QzvbE0DsmrGs/G66shx1rEC6UAXvSMcTl5Sa6FQVuezm6EqRW07mK8BIc1OFwdO3gTOYWepx
jvjD2+fb7dOsrDQO8uQaW7f+F6AdfNTVS1ZYDzvf7paJ/7z0GKPzA1WhwDK6slKl4SEERcjhG69T
joUfS9vcUA+ZyfPHU+z6uj9CgsGbnByGwl8dzQGjL595EpgiabUcrBuBn9XxG1NAk/9ybBuTkztK
EImOyb8rIxY3S/YPZAMCMEFUzdr64ZVmGwVHICJcgPfjTXTVmQ9jbBv8KwydIpQYKRMj8Rq23IfT
yewxyJgKjttNgh/0GNhoVA6+N/KoxLF3il5SW3M/NYVvZIk05h9zhJM4BVSxLoYmnUOnQF1ZKjpK
Z2/gBpQQ8/1vbFqLngR6OEE1GNE+hQq+rgE79WWxp4de0f78Wiyi19xAM2ejDu1IpfksCV0LFkQl
mNHAiNi0Xxq7XY5B0fSxutEc7wkaIU/50jCtclrFoeRBCBQ/DnHmSE/drlbTfG/zzaHy+ch4JrGT
1Eix4BIXGq/OmqXsLMdF7u6VaMK64wSdQx+5oinMCc2apDsF1p5dLr/FiFnVMuUxHJmRNNrLwOV6
8LQxz9cOuAcnIZjSCb0dRpZWvKne4Jgvxry2xzZvAZ6QPlkCyy2ZgHi+QUaI81YVYBf77luLQbAg
KQGr7EvB6tQW0ZOK+CxKaTNHzbmBa5j0iCocnfsyecPXQJtuVFxmjGbdqT5FM5MXVm/wiVHB9xqu
x6cA4DH/VB3KYcbZDZPn1B9Y8SUf+8rRDZpYLiKs4nZfTQnMv5raBR6HBNX5L8WKazSDyH77dU/G
tOo/IyB5PFd69N1i3IR7Pbd9ioCNMZc6clRDxUiZOaaVJIjikATXzOENPEZCVqX16crGMnmMl0WE
6RR4JeO1P7KDLhnqB3TCoor1hyOD20STOByK1LCB+XYLhkJbNilRXMINrtZm1yrSmdFUG0valdts
hSGGg6JqdyRkfdVJUL+Uv9F3glVUxEPFi2HUAb9TSTkHaJ+WdHrs50g/t20fEVDAAdjQNQDPIGut
0Khz4b/da9qIxMtSwfd/D8bgg3qWBDBQcjOvncI0jTCskU5nvfYniBIyLZh/xB7DkxTR3+Tx2GN3
/roBG+HSPUBqECitOmipA1vJsW2EdkAuglPTkeoA6Db4IrkT3ZrTCwJhNavTKbaRAgHQ+eO0v/N4
kXfboKcFrQ9zfe445zg2vatR9o8f3ZJfdS4kvDuDux0UNphbX8q9db75wB6bmkTX+/vLWJfs8wEr
Ccxw3UtldIjYJKSanlxrOmxHiwCRMrSIQoVb1FKRVnoJw5ZtkP/ItNTUdK9LsvDBQdEileuqdqfF
7D9jjh5aGtRKUh5fh1BkCqCn+6g/y4ABVmIcjNx3/tFJPBgYjugHHTIyLutHNEukNAgYHye6yUnZ
AMIxRbxMJQ4X6cvBnegqjgT6t7zDh5Tr34q8CfnnPDc/CfwLf7FEpC8auRUoM2el+y5e5feFVQB9
Dd8GRXKWCLfZbA0ScBPRXV+iITWwu4rg1/94VYvbaUpJqUPh+E+r4SdgGoYcpIgbaAmLphI489vw
iU1HqLDSCg8jGvgFaRjepGQfp+JKoho07+Kqlup9ZNdM9RXEXdN6pUgifTPCwiVQad3zu2YzziLu
1UayjDukgze/WLtGDu6HXSbw9OkICivpdvoEfQLKOgBJllPF5UoJReDuICV7yi6FFRE4UV0oyjgQ
65WvgLIRNJELc88atZf5EogK3Jp2BIWT2t1x8/dBsqqaLnK4t3aFruMpnJcKvTJxWps4Na2XtoTO
YgDrCIWb5ltFjOsOXOox2ZGiv3C5Ux9yr4DisO+8rVqcXD8odCSxqWC+YXO76fH/jW0ZhR2MoYsO
YMplUbQNz5XGy4PSSuG9Ce96SGd+YPiLI4CI4Ye8BWbRbOstXUCjmARMEb6qPJpWY7RJHGNgXqFk
RtVT8ymFfzes6UHCNoRp0n/RAGpGKz4jK+jtqAdoEkGVDwxxt/o795yiIid8/I0ytwa0vvXO/BFJ
t5KWHmQE309bXXhj3jqUh99kK1GGA595OlXb5F8Jh3eB6K8UkfQ4bEPUJlNoJy4nMsZxX/8UOzqI
9KNbWW+pEdP7lGOQGes1L68/Nxp0nTevuszA2nwqaJ1lMfTEJ9uq7UzgRZYoEln5Z0/A5WTLDg3W
tTtaB0tMCe6Zs9JSHvIrJ7Ur/FD8Q/jUvPMO6WA0Iq/qzYO7pPbB4G4Q21FUjjaR3RRFomW9BC0O
vPAQN3PGNZNbd/or7XLQ46LOQ8UAKwwDhon/KCznwg7CZbZVyZ1vxfVvwE07qDVMs9eTOMCkkp+e
1AdM1rRAdHCnflQOSLgGyR7XcaZZhhWOIKR5CbBV7OK4dQPfpGh6hS22aYHr3mnLA0FTZR/VCPTq
bor0keID/k4blqhkosGbdNh8h4G5aRFxuRqsHhjRFM6EksSRjcE7ktNKU4cJkR2qFUEcb9ZzwUSz
AAkUdk8UAUqwLOjaVhk4puEl8xXjUpfGhXb+JvDdQqkjr2VdJ7m7ieqSc7df5qoqxfqwHAfOkMTN
KF+rn2FgpOngtD+MVUCYUQHNdwiV0mMHJ063fFhpIntUjKxalPAy27qAgySQGOA313oijj3/FHvq
ARBZ0MMU/1sd0xun5yhPO4bnf9i+loSVE8+FZUkmlA6lJk7hLl5iBZY6Cr2uqCodWJ65XnZpErzn
e4ReyJ9p8cRwAVIJ4D7WRIYu4Jj/e9ZS3/tNQOB9q7ZETxklFMCcWu5DbhzzdqrmKF+OEeMoxhLQ
FMgJCKxGSb63zqFtWAf23GAwT4lS9Se65pMjBSA3oPBO/yABpMSVaAGY31WtmaiuRVxMOIXEoFLd
LnN7XgFzsOf1ypsFs2gQDiHaWlDyuA0DFGTKPt4KjNQn+jldTG/jZgAhSpEIeVt7VoZtYExQ200k
kP5+Y0wJiRnEIR+GD3lNMz3xgHPZJksPbB2+1xjjYCBCrx7HdPh9vpMBlD5/BUIRbY/seAlR4V/h
e0pdNSpFfKr2I+u8+09udZdI9PYCm4fKQoKmrK9WujU9yLe0MW/j6rd7NNfoDuKMTJqC5Segfh6Y
ZaMnEW4P+gjRNFgqJKlry5kCHA+3+o9vKP3XQsULLLPj5/BO2M/2gOpip+uZF3DHGEPy5ZhCo9sM
pj2v9Ii0wepQ+JRmrpORI8Al9LRZZMmyKhbHRRRJYopQCIGbj7QOkn7agfd7KDBY/0csXi1pxDa6
LQoQ/jDluJL/yJbyk/ixz1Wk/jw361V2rCkfJ88i62HAcBi3yeydRaLDmPLxLXreQbffjQs2b2ye
6Hkhib/n62y1rIdlyAYEwfKjEdBCZRNppVJ9HBgot0cSGh3khNJI2uoi+hiHubrPiaeMxvP9jhHE
YcX4XnXi64AnmolhzCNDZvGgulXu8KGPx3u2p/Rhi8EkwJbCzkoc8P/6Mm53Ou4dIYjPp49miNjw
LpvMca5O7qzEbMHPDgpKIhw3xdtcQIng6KBt60b5NA/MC1yPEAYdnYkWJHQaFsPCh7zdZKoruKOy
evYXw/CfcM+MK8ABW09ow/HnrjM0PUPtmWLhFh1DLTxJOWanIggFsy6F/fab8YE25RTEL5OXHmZT
1Iv163HO6thB5Fp7IVV3GnNrfARtRCAydLeV2xa06REJCzK03zf/mnmu3hyL+TaL7oTAZdL8aCsh
I7dyAwti3UIi26LwrMA/CnZIEPFRdBpEOiSfSLhUzZ9/W/ymqqOS5JsaOwxL5QAAdLWFpfr9ZXTT
Rdb86ZMiWp79xkKPsTJ4U6Ai4M9ljS5MTO1gVe824mPp23oDBj+tS6knCtr8s/ygHS90ZdrpKeDp
rJ72RgcmDZnT4m6+fdHNyPxbNcOIZkgYDBPuijn5/HNDbFbx4gPvdPBQ8T65kLHUtZ1F+afvRzNu
JUg6d/KmJjKrMi0NHJmBwZdBD95Dq0TxAepmcwn+gnZfQNlYp4ygLhtnmAYWgwYsqTi9INHDYaQe
4bI7l6+PWjP2TYUN3KGGZK75bH/wCnXuM8GU1dhwq1cvkV6wiihY7SRBCh7Fh4Y13V/ggpWezFHM
TebLVgl0Ogt/gkWVLlMSYz5+hCe7/abQ9AdsRiywThBL+bJCkJcfW02J3vo8yFMCByjG4pqjE+zG
GAbfbsx7NJNNN7omdBUSk7EBbXfCFsQCjuCmDGeKuPfh1f3LiQFiJSr/SyAOU+ILjF+NLN05cES2
kYRzHLp1OpsAlol/ZDkv0JUwwklsuRERIdMQp6cAYzG2yH13DFlYfzz7RjLIbH2Hr4F0zO45gfrj
HjscHmNLZTeJQ3l0/1/9W2fVYS8iAvlzmxKwe1Kt6mfguYcXRUHQLZubS5a6iJvNLhtjryMVPQqr
YTXWzpxcXzTJWRqbbx9dcvQRvZBuSryv5tsP6v6M5prn9AB3PeDK96knAS/W/8yUjw+q0XjudzWA
Z3Q+NcF4eDMgHILvO2QPWu9NgymEo/omr5etkW+Z74bXQU3Jtq1iU8Tr9wiTmVSscpyfD8j5fupU
H6EvPTc4xdE7tS1PbJHYndY1eaSSrES6m7skDTOtNBJ80UZvtH/T/IOnWv8IYbIcw/vWlJHUAfrk
HiFkOlp/D6WRLWzEUAvNI73xtFnQIfkidbmZ/Uyd1P9eW4EufA7fjyLd83P39QJ/XeGYBTVM0Isf
nc/kwNXSPMevjXZ01I6TNteJqremPPRkXqUidxtAAZaYPywC3KiN9l+xIWNZDlJTW/HZoufHT68y
dnRSH1Ci17YLDQQaBSaOuiVt3GZzLoYBADp30IMej4sn4NcF+3cVt3ik12U1FiunthVKh/S/krV3
wrxCC+uwh3l0bxFIujBiGDSRqrwRIqT/Ngtm6oxJM8gdzjfvNSBx1QFsh/Vln+iQ33sMFVmr759F
5EklQXf5uslYkc2mlkm8b6Y7rcqHxR2VOXM5J3qgMP0X7ckwSFsbTMO6jVGVLvK4KBwCwqbHMVOY
uT+X9WoDg1Doucl+3e9Z+EaGXp7Il8Q2qjPO2j3qAb8jI1ye3Svu3VLALgWiX2nkGxS7owJyV7Bb
FSCAJ9vSaFKm8CbCIpYvQme3IMPWDfQ0BxDpssEntRGJrC7wy+S/EzNv8BAw35wSHaWnRsIPptji
2IHzA9KlWZrPuDGB4LrDUOeWc6b+YG6VRtblf0M8BkuCyRJwiSZxJhr9mvRUVe1bX/DmrJmYyvv4
KRl/6zydnxHSsv4Ui91ixkcJiOPQFtLbzW0iE0yGmOClMAJAJ8cBW7Rfxrr6HMBEsgljQAHK+khJ
7iN+YYKsJ65Eacbb2EkoA3N/Z7XsVtW/6nv0nc+EAFt/dqJKhFLmvEHIKOsdESwKLtE1PMwRdwbf
IrpMDqbMPRNb4pi1DF70YxGiLf3kGlUI+O+/RAd3TJBdvW2Bu1CAVYGU1+igBswCEnNxYJJX9+BE
pX/AKloLC7GU4bd8AMMIO4RCWJk0pEDcIi2cxBUllfz5xAG2K8aIt6q3xdIjsT2w3mBcL7XlpvPS
JZJJTfByLk/3iA9gq+pEiH42t37LmMH0HhuxhDF6d/iSqDUzdIaCdRoY7g55mub2n03k7CfKtzxx
uEdRjrC/NYx+Z9SRH0WMD3i+xKCN8t8Y+5zWgOXv0+fJnlzaKzJGBQmaOaz1KBN11afCDRLchnik
NUEhOp/1xW2gMKKh/jUroJTa3HYZiagMApQT/OhGmMljP2L/aagzhnLArUUfTmFunwiknm1TvSw2
tM4iqaiU+lykgMvwgre/xvqVS2i4FZyOMswaX/BW1RFC1/AJbKHLqWxgndOqKUviIwbIrBPC6fld
0PiNtda9IcwgN8p7t3wGclaprWaBrxVjxf95p+v4WXg5Nms5NioyhTl84uMEx4dcLIdzNKGkD3Fw
knfqhxBzH0EANWCX+HNiMlSIkuz+IJ5OdxIywMZ7Q7qQNoLBLZkDN3+GYQohF88MTjb+lS9aeGuq
9B5FEWYkPHkDGtgTYsfxLWlu4+oyJaXxMyGf1JNnBLwwxXhmym/LnhQEsSbqO5d2jw4Bp8ye+/0n
Vm3Rl0YBTva53O4pA1L/IN0xC036op4YCX57bzrKd9/Uh7NMfHeOkqhhYVeKMkqszMA5t60hKb0R
xF2dFPN5wesj0TrobLxb0XcqbGiKZuhhIAqs11jEwwHBOVNximIDYwMeDknTbjztHQWrlBwFkU+O
JFpHvv6IGRf1U5EAKHoq8GftsLCYWMyRo19Au08zFvgxF7uG8046NO8Y5/2531leCHM5bCg8o7r9
l0pW5yXd4WqEeQBeqzUQTWJcmLstHhw4QDzV8lYzngQDT7BGKawDJDny1J5z6OglDS3cnAINcDRQ
YWYCPP2IF6gGpmPxlbAhqVbNiq0AIMzjJpyfMgPgmyta70OCsLF1fkeHlCYLGkD9Td+gfTluYM4V
jGlcFEquuVS1JmpHHKmj3elzSdlbdlYqUoLRsseHDjo3mMzAowumYDTKdBGQK4mz0lBPQXnK/WVw
ufeEZQ3EuVAZZBntNNfBZJByIjfzONd/JwfTXAjkw94L25w/MQlsAG4Bb/1K1+aB0z6lAsyE4vOK
mmvMPDqUolx7qX0xhEbxkFkuhdyqP+X7DxSpJOXYIolM5IR9W8381U+1mcFmV2eSQkHU5xo68xQp
Td5VIUPSxnuIZ07B+nGrKrtp7m0S3NnxklSsO1DH/6PRiEjtqcKBDwvv/RoPF0dMSsBiCTorj/mM
L7CRcK4lnuWtAJVMf9ixoMS/SXvoX1KPiWNOujhP8nWZqFB6eOLrSzEWAms7PtPEBxdCccM7/vU3
66EHr2/h/IqJEQpv7N0FvJmidJrpk64tIISRkS2lwmHGMHOPcpIAfnt/vrFWJ6QKp2jkTbyzS5Rk
S1QMAaCxcDJgduhPm85tG+EK3B47IklZ/Fnvt92XmsV8K5pDdGQhh3e3HF1FqyyHHVb+PkQ1kk7B
3zWqqEaP+TxgUGy5NT6Dnvw0+9I2LombmQWC3UFa2eF094n4oVIRUIhB77+VNdyPo73pNlQzIshJ
dRUBsO4clbVBuT2ECiCEYkp6Zy8tuedJ5cZbMGw49ehx6VFGSMAar9Zrx1Aw+EZMPB9VtYJ/dhQ6
fFWzaku4FWc8NegUbCd24SrLesDB7glxc+T3V3R9OrRRxiNcmCxws+uZpasPzIh7rWUWIM/GJ46D
vNAouXezLqlz1+IDKdNMBjhRMNwf4GttHZKvxQVyFBHVTKoKTjn7vAlM8rtOQKUq5tP09enFFZ3v
su3uyyiKhJy3DyrHOVs2AJ34vMOmq9DKng5cG/y0tTf/FiNddDMFy5m46iPiZ+eq09Zq3EvpfeMT
1w5LdrVY+5BcIzrFIsitmaERMfeyYL6MOVRPU2Zo3rnh0dOkODMPgPArXwPINzrP6EaILQODK83K
0O6qsgpR9sFnnTOXNjwn3gLUnzom5c5lfbc2spaIFhPqNDmwMk7TC43akeJ9VL0Q/OHwRIktRdqM
yXX4NKAzwq7WxqBbD64YzVPBlN5tXDXftFbs1J1aIXz8dsIfYvibw0xgdF54Y9kwXZaor9nrb1FG
FJ9piirVgQJWuVP67jnwOkoOpkPuqqrsJSXlCIe+KgRLTx1KpWlDaU+vq5oj3DdKrsrY8lkoHmTy
OB8azS0hYYUaUE6JVMb51AtQV995AWlHttHHtwbYFsnOQnYpLx0rlqVWwFkUZC1BXEHvF0Gepunw
rehzNnilm86i+Qhpl1LZVgjLzCa91wlZYkAEiNLibb69yUUGA+wuXwNCPxl4dOK7TWR/MKWZS77n
Uj56KGxxjcn0S2vUUlfwbf1sjdSpH6d6y2RzEgaeoMJOdIrRLdZgIi++HaFslv7nalSWYdRE5X/L
XkIWyKcieioSzhm0MpGHB3aEXNTKDv+elfyz3TvBQIv+Mavv3xMomLopwNrcJg/U/0pemg2r2FV7
LPW5LS41eSeFmpSehvzpuEZBT8gzDsNKy+qgEvAVIIkhUqnvhNIvGEiSSHBQkzjlz72E+GbJDK3X
G7u6afeanOOw3U5azXOu1TPqugENyYf2MNzR0vkPiBJQY9F0AIwK5pFiqHCkZab/RzJy0lqTFomp
2UlCEWIwPK3bS+1NMU/oY0gwoezrhH/4nD47GPAkQ3vGsOTWk3n0sjvOlQFMuR7snfUPjrw/mNRr
Uhinhg4/+qtRFzlvyUY7CXJr2MZNtmcWNrfIalsRnpMNROAWC7FDEe++2h/9FEc2TGbd4AfD4ZBq
+/gJHdy06XMHV9D5wBdI5+di0LcO/gcWR6wDCJ4eCQWwStvkg8OVzNK+mN/BHyA68jZ6nXH2BCA+
rdLZdk9rEZck6EWo9fv/UquywygTt7diCRWUlJpO1V4oXXz3l8xV9sLZod4Bw6d3gJHq8w5VNved
RksgBV5h56WVLnhWDEqw8eNZvJsSk1vGv0rP8w7qt+QnEqHDzB2N1Vq9e1dtXN07hXZAodYrdrp2
znFcnuvuzr2zWLD0zCFusHK9QxtfBg1j+juqT0/379+QI+9NU5K0R7wkSLzrSPhfg4SEAgdqOgtz
PFy5bpgdUninRnivp4PJpHzztw/xY1tCtj5DIkgqI0V59VRc0F+x+rHNemP7uayeLmdHlYWwmlPp
O0o5zjqjE2L5Uk3VBnI2lzT23EI6XKUqjxmArgiB6975PIEAVsJ8uA74R9nEHdgWNcGvsRiFhPcq
9Jlby8mElVkxuG+NsgLJhHeQsn/1dJDD5FIQd+eXYjonn3Hvib6s4tsZFUpXoC5YD0n8SQ7Efjkn
TnC0/Ah8xulxi7gw4s5iKoFOlNEsLGgjs7OL4hAZxsfsAHjmhWUrwjtisK7ZM4Q9J/2Aa2Tsedkj
XGYKYHzY2sI7eX5dA0LwgI4g8RmmdizVHgZORuxV1WO1vdC12OKRCd52kHJVXBU+MgJ6y3nYRrJY
3Fq1VJKQdHShr0tHPJRFPtG+QZIl+ZHBQA2laNkauUcKEQuCS/knj4Ut2WwS1fW4o3IIWoqHQXgb
dSPJm+7d9INN5qdEK/TNhrxrTiUo8Yy2Aokkiz6Z7odzSfm+VBckVKHs1NwEm16oiUHvIeeI/Y32
R83SBPdsSIuS9fIMcr0QYjmyieZnh/WPBSzini39r8iRv4bK9PtjDq8X7/nGTP9P2C6JvGrPFZXk
7MWUCw7wucIsNbjOY2pgOBO6Q+PS/gng7RHsjTPXEBXmuhrTZlh5uL6peudMmLphVWZwrC0ipl3X
coq0j4lp6RMk8qTj/sGjZabclch/SYadpnf/Kul5Ui1VeivJGlmVJ8HwivZor8ROAg77DjVzdJWz
dzeFqqKLFsTFkeQOSYvPCyNbFrNvnzJRGRethgbS9+K3XLXUWd2ULkasNDYRy4r5kzEwRSw5T6kZ
TbdnFrVDteNFKUggzs8cLd/9QVEmwmnbffguax6W57zra8HOnHRo/xznYyLB1uaaqX+PZZBSSgEH
4LGX00gw/tNbuT1jx1pErRbXkSSRR7sl1cdHc+aDKgiqQPqBfa6XKZmlo19XSBXvMkredY4KWXVm
3fTADfOB1luz9YLBf7kxpp9OvTZSTkwz1TdjUPkxG8D6R4kHlLN7IHZnLK/m2V6UxvQp0aeF8Ac6
zqyOGCQ4ziw4PH5ROJ1XenYK0nb2G5vhu5ZswQ4Zpf2YCU3ugMvqXC+wxHiJiv1O1c9jPwEVrLYp
H+1JkSVGJmtg9Ybu7ZE0SQwGZjdvMCxvnw0W0BIiEepvPrxjHNaIk4VCEmdwk3DH8RcjgVrtJEUH
xxp7guCtoJpgqGMcCPTU/j3a9FiWM1yR3UGE0vBKYy7V4qWX473/imFFgZmWefQqgpLEyK6aQSdp
TE7M45x26gpiRMiPQvu6uMFNOPiGJ77oRUij7ACSBVaf1GZbSomyw3bWMIlo8eZxUrbxhYhshKuG
1Xe+sJYSGQGfduIBUrZZPT6ZGbXWyKBxCs5EBCDzVpje2+c4tAV3QQhtkkaJdvuKtHavVii1+bDj
24wk1lBKD0qmE/ddgwWzf2N3uGBAhuyE2NIPMArKFBjUn4ErTVSfoD32OwdnLJ2+HDKmoiFG2tUB
cic9PyUptVQGGQdxZTXMzJtShugTYA/kZgq1ufp3gBty3FUeOP3DkmVmsewZkN4uzshXgQIKuuKQ
Ca9UMJCCLF/r4DItaysriOf1d1WVnZqI4g3pzr6Vq0jcVk/pSwP4mcTVfkm74CsC134WHKRExTgJ
Sn5N9uK7Fl1Tgp2Tl253BvS2tnJDfNRbaFmzNkoJWvMqej+wJEgIlYLruKkBM3Ws3xnJ2eLzMI++
mMvIZ6eK8rQkefmFQAFGXZplnaXBZn+v16NotDeVQJJTOrPS4nPEGyXnBX4o3zIGvaOTwQp2w2sL
L2igGhlQ8pPcDDGhaCqldn5+opMzsGHMot0kRP5dLhotAnPvcPrPAr6IMJcjaAw5T3Xf+A11lGBO
p8jlagBNpiN79CgK9PIS8LFSsRfb8MuTq3efe0Jk49xuBDVjp2u9ithaT7QE8RshmmObNSz/rBak
eQy8KY+m9WAcSmuUaKBjASGmVCXWjpHbauVvS4W09MhJkf+IsvaaM/AMDZPqggqGoQhZjYZ0g4DT
Ss5Nc5ZH8rXZy1enFCGU2X621M9TWUfP9TZTJ1Y3jra38mndN3hKWmzwLMBaNdJl0w9ZxiSarSqe
MCVUygJn11hMAQb5f6mszwEA3ZCmJf1iZR6NHTiRMiLG8iyGwwqrKB7x3lfxYJaHgOYZhJeZ5Zmh
kbb1iCW2hPcqaPaUNuNEJusvM5B0uRIy2n6Hkl1Sx9AXM/n1fy1w0iyDH9GcGyjI3fxaQsVLuKzd
R50F+6u/6kcamV/SSf33O5yQvwjNBGeXCIYstpPt4wMIPhZM/rDhKCPF3mB6J4K5lU3MdOTUvNVs
luMGcEqsFquEd1xa+CQCTqeHbmCEXqAc+xxlDoIKofj7Fbx/KlyXvyh1VLSeo0HUvomcOG9hnGIh
QecNsMxr6CXaBs04YFANwGI6oXj4eh8gIqOOawkGqscn7W0yz3XFNZGcdKy2jLGDfOhbWcOEDzQw
xr+6140du+UfiVp7R/gPN/oC+4NBD+Gmkp55I763600V1FDDYVuGsM2r7iGUM+Ev6lxrN9ax9s78
K8N4OE4aEljWFGJACjzoE/SSelOpmEMmnhvjZYfUWkEskCDABtXh1NMVJ7CUsk7IQ6V58R7iOq6u
KJv2UcSKOTmfSrTcGINMOBsVD9FNYKmJs7P7Oqcap8i0EbNIjI/H3jpAi6gCY1YoKGOl0RU8vney
Nukd/R/h255DfyipjA/QkG4df0YOdp17j3+PjlVP0ijlKyj8S1FRkmWlyds+APwn4g8zketbI+cT
6fyvulJJeNoa2GjRia/01mW5dh1BpWd+EkHwO7g9FS2mFwbtIOujGtEq3pNinIT4YV3vUZP8ZdBd
nh5lPvygB76i7/lEbOXwbHtdSIajH6R0yoKzL5XtDwgrrUpV9ArZAobRU0d7rKzaNdaTbeNw6R4f
VIXx1IPJ+xvqVPNc6HSSew9rObQ3rVOAUGeGu49IWnqbi8w3EmAR22i1e80d8ZtcFfw9pMH1kQZf
coRJzCGtbseaufrZ3J9D+Gav1gE8jRA9bxhWPrEVu3/9/X1WHEdq7WRA2kBKfsq1hEWxAPlOrI1L
W2e/IvGeVTy9acUbGBqZzLymjr5RUxYRBCuulv77T4wv5bxfcINLyN+EvivRvF4WQyBkgbn15cio
Ng5EJq8kw40lECH+ea8Vs2dmmVDtKqdQsvbWD4zEjaczyB8W7VdEQSP8CQcEJBi0yA5k7SZcIZ77
Me+7OAVv4d3JCdJ/axc495R8wyqDAEilxyH2LoxF9Suxjl543+4uqffS2RRavbaI4Gq6VqERL25A
7EM1QRqF9Dw0cDG3Y8N9H7hgU9EnWOFyz5gIb8iqi2SOkLPH4votO5eK4MtebNKjJD63jTSQ5sEU
KZWGvMVrx5D9fTjJ5Ff8kLJyS/xuQesSKhdk0HM7BbYJ9uDL1iJ83yt93ZAqbdyIeUrwCd/kj++t
g2z0iPvmW0YOapht2SEpPb0yqxrsqoDoMG75/Xb+dc+fpv3mL1+oVh3r1UV1g9zUqif9mBPTaYcE
0UxOjdONkZX/5QS3eilXatZuKzh0/v2fDLZRnHHM726//QEU+2p4Nc5Z7rc9SwhEowKfEgXXSTOG
7hTjB9j+aBhuSgws3v4dn2ZHNbJCMxMPUi2TmIdNCFUtgjI345ZMY8cSIY3xEa/pS1vzbukRtFEg
9n1vWAymdOrFWwj2OMfqt8KAaFvRi/pUgrYDmF93LPAELOkZOZ7vvvOCi7rCYWzuQNLzaQMndnii
FQvmqS9EyyYh6LpkH6RwVYuqqXVoEhk7eBByaCW55qeYzg4frf9GYsL9sEexRZKSMWSLu7A/dE8o
77ZrxD+H5R+xqjEX1E7ESxskEja4i3uNUZgqi+mcrvEJ1Qpzs/7hVNfxxM8qRWZIUIP6vUXhBQ00
JY8qLpZr/2Yd/nuLNXeIH74PG/So3MHBTgudLLy5SFCRTPSAuUu5hheZWdZnAhK+I17otRhU8/Vh
QsgROygYRmAiwwqy7Nw2Hs/P4HABptUyyIChYhdmOh6YxwYOgDaCnWANTi/w7ezgeRxUJsuJZAs3
RlYzUf07trMD3+nKwUy8O5Ixwy7ffBj5Q8Tt07RJqw45SACXJn2FdTObwcxuUZ8Fu8joTApNQRB4
iXhEEJVD3Ic7GOzV+wjxu/WiP1fnr2HxZL63IJ4LTNpwUtoBbeUhsNmlCy7qI+WQSyyMDk+lkpI/
RleVcGC5TpMCAC83TmuK4q61h56NHh4QMH/tzNcI2bJXdR6ERZRX+vJfAsy70XFVqJrQI7CfqVT3
hvUm4ZKrPyN2DpPoPsffRs+9Fw2WL8Jjrt0gmQ+dAU/dAOw392m1obfyArj5YC5DEMpcNesHs5Z/
MBgBNbISHT9htxug1IspqusNHyJzJAGAtNfvISw94jYWBck/GydI3loq5C2I+nyQFORQRs9U/I8Q
lx3H8Lh5T0CRHrjeqefafpYVasqGL8uYghCTomNueOXj8spkHcdTARBcqbgCLa2HjkSftcsgQdj7
JrIGbetxn/pTQRKY5L1nLd5xBykJ+0HKYGUDytpskohKjwm5u5yupu8JPn1XOd5cJUHc1mj+iqas
zF1AMRL3Gxv5MSDMzU3zQQPnVWKi/DlSv39P+VHY0yc2S/VnX4kEqtD/ifKEfGjjh2PyNoK7t3Y3
+wiEecNnyTZCsrWNKKaSesvTa8e4prPtWre0B1f8+V+WLp3F+hd7JQGszZIvu+WviXhN1BoFGLUc
FtXrIF2gzNJdwwMX4uRY6ihKx2sKwTETd5GPyrQmVtgpFbZyuK8UR3sjDNJ/ZggvzigppcXAn9ty
qLhnBENFgwjKxvoSL8eRZnA0jqPlsZYg1xuyDCcaZ/T0+7LVzZKbyHYkjJH+9c/vOuHZcx0cdmqz
az4UxiXgBQBpS479LHRB/h1hIlXmfZJIb4ITqylGDewY9llZBaLQkD3BRaeuFc84KvyUxefFQhZw
IOKvi06eCl/wCMYmcCtHYTqq8fp8TMzk9s5iZHh3w6RnVh3QRjpVWb4SjAENRUjD9suzVBlpPYpv
yIhwWoGVZNkfcw6ALjBfQ/4tCA2zOC4D6VtBroxxlPt4nDw09kz/I8S7EFY0XIpUOFt6pvQxJ6d5
52AcGai7j+lEV8y9RASMk+7Q4rMs+kU4sdMJPU5xxpGmI6Of8fw8Hk7gXPbKqTgXeVnu8NmYtWbX
SQw/cEwqsHGHleWaEmQAzoRiZ0VbClmkAloeEVi2BoTVFRZihxMAu/fGYR35+aOZhVjC0PrrJTVk
Brlzbu//HFrN7ICHjIB0HDhWrraUJxTlik0lY9zwxH7P6Z828rnDiRDK5EpC++HSt4qbYGxgX8uW
bBV4yRN0G+VzKd6c0Hn8kbKwGkut2dwx0at1YALu+YTFVVYSyyPhh8JeEwtrYF7E3qc57skDdksJ
/sclbT2xZiijgHauqePOOTrkcka0oTVKjvToh4WeaHRNkf+c1vaMQqAYUoybv7V79tSzfDgwDjkN
G7AD81KDxHRSlR7gY5vUiSqJNdmaOmaC5/OLvQJDcnJQH9TXz2TvFioVvX+lBE2gb8Sm6CpL11nO
yf58RdC6sNdjeUWrXxALLhfigWXLRG7UTjBPCejKZ+ipP3Rw8kWdkwbhz9bNt9wOoEovlM7pMCH2
xQzFxySNFPPuRnIqNuk7xqmqwHiT3qYhpqlWw3YX1G7ykb4ZFpvgsbttylbPMGKGe/rwJVU2i4J5
9gFwcsgshmBcqAIFN8oFgc1e9PL2NLBPIJnjnLRt3yW3GAUSdRuFQMu56Cb0ACpEZT2f6oZDSW5G
6Y289cSt0elwjlyAhWPsUJNkHWmd8tf9mFRguhTz7rsg6NrnakcuPxXkqvOdbLR+r92EmEhRHduN
C7tcpqLZCM5cxrezN3zkJOIPmM1zD2/Upug0LplbrdYcHeu3O2yOBaOJs4AB44xWRz+nb1N0MiI/
P7bADfYOHJQg8wxSay5n/+IA4Toq5tsFf0+t0qDmsg5s+hxZsQfJTx7DRDrNsxbT8lFkLpRtNJMR
L1kKYTb04c8T5ngT1Km2XeXfs7swHsuNG4BA1d6V+Zau6kf3DCcSywmI53yT6mHXF7DirLXSAg4c
fvivMhfmbjdFkcckAEcB9YQY17stDyLUX/VpsKHixzO/BUlv+S8JOB/CGLkj7xejB+XhizFamYkc
mK2BHf/2KiQd0xHfaHTGemp7J6kqENNGEmqr2omUAqYOQezWc1mQcCIZ2sTTd9e2sVk1DYiGQhWL
yGSfrjZ908OWiC5Yu9FV+tL8JNpwJL7l9U2b0vL4ONyxrPSq6CodJFwEkexGEEblcTuR26qF+e/6
KQC3/AKdLYDReAPVVdg680vExcubvYvObPU0TEjChlCGc+jMPH46Sm8mGk7fnIS8ASn0jgrgmJ4h
cl8wD+DzhmozL7DSMANhGvJaHPHbLFN0zuosB1pWkrVYdNMSb3zreGGnVBaLhn8h0P3yCx6DJ9Hs
KmLnL8YaZqy8ZF/SrQTMNwPFIgSqXUuA+lT/p7v3TlyltH1K/qRlJYG7yS3Ru6kYHz6nntAxJmgS
szTWLO4LFeQH0iQ/0+jv6edMXWPYVsWMKCGjxWWxyxNdS/ku6Ak5Q4AghSk0n42Y84CA4OqrmPCT
qvFalpHzh12Z1TjWlAlRFOO+G2u5+z7+H5w0aMVytHqrKRLoZVrql+waJKt6z/bX725LmvEbKWOV
AJe7L725yOBPfvkUYxIHyYJovKmvYEeYwhh4MnSXM8z1Ptak6ajqw47OvjkBV5/xeBM209u6LFB3
kAXp95/WXKKPmAN37yW7vyb2PN+v0z4BKj4pmwaUwd05FphKU0XxNfpJx5HEBGAWokypcbgvDUEj
OSt2SCrXNZ/5UIpJev7VJYTlKIaeOeloDZ1EMNfT5kXzEXiJBG08h4SduC+ZZUGub2dokX6+2IbA
oJ0fOGoZtANYJR07be21LvvbdM8Pl8zkqUI+y30+1lao0xEGrAGpk17CHYwsWoJclIr2thsU2LA3
QqHex8WKKSNmsSzODjHWphoasfrTGoVflLijJVu7RH5P9IY/nYmNY9pVNTRViafiSuhmgYuSlFOz
7IssFVQjZAZhLFefzb1G7/r9pSzyFmu8XWDyRKM9EVMovKXm9+dhlW8td0O9KcWO5hwUIvjmOuCK
G/E5YiK+/XhrgwnkHXI6a9grkuppQfZWKEdfamlwDzbnI2sq9KMle7eQPuBs8XidqT+LpC5m0cYj
NeqQpXUyNd3JIAw1VIcO5ERrEpknGIJEh9LJuiQfGYy8Gep30y4fRO/NIoXgeoMTXmcaO92UkbzU
YLYQdYKApca1Sus0APylNkyBck3KTWj0lGixIuKmPCRrt+HHNmtJkoWH75OETqKVn8vsOkdeUrYB
dmTFeIy4BsVzfFN4QuCYOpZMWnvTdGcF0snKaexCZ9UQmOZbTnIC/jGWCjBJzgwHvq9jiQPBHAAM
7HWhv/HhOaRNU/IIlRD/iLcH9fz5jFWaNoFaEN4W0TrIZNpkRWA3NeDb61oy8SjeYm1duJoIFlwe
KhTHKZPmZS/VomdQloYbRP+QjRP8Pot7SyuSTIkgG1lo/aX8xThiYVS02GcIqSgN9S8veBInS81M
d7SOhFNA0lhK8jod37MyPQsAsJoQ4o/DnmFDKLUJOteTdGKxJ45K4mDtm1q5Camrnw13XBDgcZE+
NJb5LkiLhEi1Qhv/8rLXVL1KCXY3gMMLlPHQ8bLQ4G69VmYhSLcZAwQ/XcDqYaoZBarjJ5l8VbyS
T1ISKK7ypuVKOW4I7kKH7yQE1Z5zCmYUtbyT5OEtFIGr68lxFOAfn6jZy6F/tbwEldBp7qXNaviO
SwMkbYfg1DZKkTV8dm66rpfjvNJ+PFmV0twDGx9vwxlmlbz7XnaEeQsR91R2mcm8/qBVRozldPPv
4BzUibU5knlNzmXrmeW/9eOQUmJxXEhLlegdtWVRn9nXTVrgKNRx9Gfw3DgNB5rUeMoVnqXpbiQ1
HPAhIjprUa1pY+7rtVo+FupttcQkcxfJahgb4mNuz7QCU6kzlc9VjLfMyrAGSMNW8ND9sEwKKuAY
v0K+8xqCgQxPsIOc651tL20p+MpdJw+WBmJENN8qoMmdNxtvglmc72uJHHiv6FDMQABsHtCaXcnO
1kyWuGHnvXpakFlrr9K7RZl9MMLKM7SfnQY9/V+xomDrfVUk7EMHjp1DsChSJvgtAx+Y2yA4Ok9z
Q4xdUA4HyRHHiAOsK1RHrhhAIoCCgsf/eVtFyWKXbQ8dg6ORghPXBnecrwhaCkVG9+YGMTQRa5O1
2hzJ7Y0g/tvE7C44CmNcxC9oBXH/Iw3kZ3sJ+WGBHtixIjpKZi71gzvqz3qqvKRJDCFT/1nzxJVj
ECGw72w3CFs9+QYu+PQMVLPYDHdtsyX+pogiD8OKKBe8Fo65T2cRHJDRluulKmkOynhixR22S/Y5
L53jTwbOA+5xXKJRmRcY1sNnxqrufE4zdgLjRjbh9kRHHVEqJn+rizP71KW+zVlJebYgJT8DSN3S
rJRNAhdoElFW7EaAp8IAmSp41qmZ7bCVjT6U9iJG7H/8xmfmwFEIlHV7MB7cDVCfwke6O8COF1hu
x/O4xWV8MuLZYbaF8eEXHtQKVX3vhShaBMn+A4GuVEtQO3oJ+8npsZbdRtPtEhkH23YwPGxrI5CK
8n2zZitgDpyGqS7UVtJiBqN0aCPG0P3G1aivuPnk7hl/zcP3kEEoNT414Y7f319kt5Ri1Xp1SOVv
MTzxuTYBZFzzvKRkVxrEVyym0QHn1uUm/dy9gVamMpMCtFQlml33nKZmWHljuw2dPgXEUrtHee/O
lEp01G8TSpaNpIK1f12ZR62+UHNc/IMzHBRTwr1JKPGlZdzp9iNcmd7NoUIZKlmp2qoZmVTWksxF
RPYZgo/iBC/GyI/tXWePLX0lxqhF0dtaZdrqUxj2VZ1taMSlXNuYu1kMQUlj4H7Vkp2+6zkFJAWV
SGc5DheMBgfjFKTKxBxL7c9OOdadvw73BiucgXUkOY1scqvmzW1AU0ahK8pWHnLZoLub/oGpUCDj
mVKgMfrp99MeMS0yC4/7MDtOgNAKOKnNLjwaTcLUk2BZZg5sw+1IuiiG4s0cDxQU4WCHINOYTkBQ
Wha2wV6AuM8OO4z2HZG1f3pStNYFu7EHTUiaUlGY87DLC6lRl/s2162/ZodQKlapHvmS2KB+YQrJ
jc0/qzoog/kuJesynEaM6xPXul6nDFFa5HCcRtmQOHD3nQTThp8RgKgs8Zvx3abiOfealklUr86F
UkqOVFtzrbZ4vlFrLHkjvgadLdioFYiS2bFH3EKJO7FzZcOq0H8agpLc0ncI0dZt05Qd4K23JFdl
BXewFBXSyveBqKxE058jArU7QhI9kxUZjIbBP93q0YG+DcqT/KEeDwecEevuacmH3rlbfDjSmZK5
i2T7VUXTiWbx8J8DK20lpEZ60JWdTkTH6XNBwa6ROWF67IapJnPuCeGV72zUN63/jLV6tAin7wGW
aVtpqqow9KDM9yI8SRtCfp7ZudgmJmNyoNSMBju8bG4ro0vMaYw/YJCyzA8ShkzuFpn+guNv6jrG
FAgih5/BW20NTC4pafw+xJFUG+Yz/V2pfqW+MTYhgluSsFa6xpBX72JyXNiy9felrDntk8ODkJc0
U40lKNi01CQ7tl+q0RbQiIP91c46pJMGH1AWr/TsQotFh8E+RHYO9Sx5QpmSkJ+FxsaZ37fwYlPx
x0Im5OdwvZlg00UiG4ZaCEZdIY503oHxbBI5VAz1XeYRRnbE4RqEuGmvGnUO8VLM0ZYLSyjAw6P+
qfTRi3rPVLleHcdo996AuxsyoRDQj1cVlqxXMDx8wDYw1PKGuioQl94EPhbxhSv0snos6B+9SMV4
f8cFwcFiO4HqMhJdwk6zE8/pCerJ7rCj251hK7zy5g2dFwCbbE74yD1vi2MQkrfcA/rO3k+nDEuj
ZSxGvPBRjtid8Urd+yHxZTtQVFNz7iYNdIXvcrqJbFJpCPe5a+xKrTaOEHgzcTT6LKf85SV+oYyW
W9TNzi3/ir0KFgLQxY3Y18Gp9g6xeycg/exyOzYTRB3RSSOqxoKp2zX9kuA3mfXY3l3AwhxjBcG7
kBOXg/GXzXBNdCNX6LLVyMxRVaMsYei8KFw8N6+Fxw4ysy92OWnP4znOgRn9oPkWuU8EJB+eV6HX
/8MajkPlmVstJKyVsWpv4gaGZDZdVsD4C8rHDyRoClJ4QCBRtvxct59kUrsBMJTWGmqRXT4XDFRf
U2Ff2l7/x02lMFMmWu4Sb0X0ptQNyLnRaTUaW8bBmnaAl6IXTIAVmvcYwPJARybzbLAoey5A4vo9
dd+IYXEucsOt9yugcCowrpkHwVQDuF0wU/9uegDEuCBBTCcGsStcKsVYwVsTZU+KFzjaZXY3EXa2
M/odn4JjQEBd6d8kZQ/sgtCGzM2uRIXiueCPJt2gebae8LGbgE348YhmrG+ixRPJlNFRpMCUC8JF
4VJw34JoHvQvCxiyhU8osE5x+xEQmeLgqmNYYsH9MxbND0b2ZhG9G1NSwae6SNSvUQMEjc6pa56Z
demL/xa3YdkOuMAAoenc38UlU+pnpfBk7zrIHADjM3k3nzjhW6/fuiDzc7XbVMO0jtg7BKLZCm5D
12Mgkqwz5oPxi8qdtO9vLXDHylg1TCZQzoSYu3btOWIk/Qn0cdqWfidkazqlgsjNpUu9C4ffec4B
3MYktuqVyF2N1a/8YGGlcl5pY33wmnA6+iPx3uIKZw8zZOlPuQ7Y/ZnNr3qR9lAtMHKs8tjkD895
46OdrX7f1UAMHVcG71ZtJj19Pl1kehQ/Ul5PLpCcLOWge4VoueRBxLiPpuZ61fN0+tNn4SrLPwQu
U+i4LW1Eui75AyaD96psZYJNnqR4q+XfEs/W5JGDo33s//zNs5HXfkD3+YXH94buheLmC5qRT4CQ
R08cwuCuLd0Z45GrGPAON7iFW78H6CKDp3x89ttQ/O/LiIYRZ9CfCy1n8wM04jlKiNjCczbhhncd
40HDXMmg0XLhGYb8z1bRX9XJvyLQmMPY1qOcROw/SnZAPC79OS75+OEfU43e8yxpQmYTWXebm4nn
RwKffETs7AL0oqqwyk5hiBE6XG+Cv7+YWvaSOsui6VIUcBnWRbQM9ARbQmYd3v9sB2Qi9hBNsXUi
dFlMP+D3UHXUM80eNFNTLRwviooiDBIer7IEorfBKxjGIBBvTjPrKK9qAlbM8a+I9bct7LFejXhp
bBUY0iKqbTV++s4SVlwVh9C3H1B8SI7SEyTJR91kdjpFDbLX28w0+69JtYJMgHLT5zZH2AXF6Dnf
XELe/hip3IlBYkBof6M0HZwTRVvo9YhB3v+x9H75tiy6Y30ahwKA02AhtagrRAT1Bv+LIyZsbNeb
YCvxVOk5BtrkG0sGABloDSeLPD7M+fVaebKz6YESO+Fm9UtB1gEXrWit9TRMM/8qJYXMku9mUwX7
6w+CzCJ4+HaZSr1FYbfUslkJbTq1VvY31vLrVf2+AFnr7Lig8+VIrt7Fcx5+4saahDNv2MsPnwyD
01FjzmxX6uqcctj5Hff7JmUxmav7ngoSWgfpQVWY0XG9DLq2SUNrJgv/Um0Fpg8Tg0o/oggXNW9c
AXbd0TYOGDJvtHNcL5IC+5pY0x+C4D1fFgwy2D1Nxr2A6FG388p83oqB9oB07oJAo1BDT8p1JzLO
flwGMGsbNGoGWeAFppmli4CS34JEXgiSi9N/CLdCIy5xk1GTxadEXC7Z3hgL7pNjWnqaOe1VxINC
Zq9SJqQArFd9xRL/OCr5/rClw0F7E5tDdWrTMMHwllHmSgHaAREWBu+XuCCjjDzCufg61AUpcZF7
lbIaPtobPeijfZ0FYO6VTkti76CGkNsyGY9CECVlB25tvaZM1yJAPpB76J+9w9Hkiec/vgBZ/269
6UAUNw+Amd9P2ANZP7zbi9Zr4eX9h4TyB11WrVSF6HeHRoRZtqPkEGIE+bAi5r/e+Ko2jdrVWT4h
BOo6Gf8hRm8L2CN2qg6uoyRfbmuQ2IMEmK6kiusANqJPRq1GtgITJckzLDvOZDpXdN0p84VwjQfC
3Ka8sUCl7pAf2mRTdwLS9Smb5sdAj8i0xm4HEIiQQwE25S959oVZYYJsRaQ1ifxe013KPj6uTwSc
16O+Oj6XdgFj+a125NR7dJ5/cZWLWu6mjFiQ5vrQL4SaQE/xXFaHfA5Eht2iMOiHZ82UfmyxnKlX
iL0/YqVZTh2oYAfkJSXf3xwBL9mgjos9FUWTbKuCiS16K9lvF84kKsz6o/JyPXE3EYW4o8971wx9
+nltyHaCHDDNPhAK4QQoWGZK1MMKT+4TnGytSFLbq9fEiwPhFORZMJ8uTAtlYc3nDSqtWxIXXHtn
Yf+0WBjWqszAdAr+MUKSlEA37HpgZDcHUdgfSeHyTehcJFZnhZ3aH6wd5Q5mvJdlvVXVXmgNPJ4U
b1Z8TeXe8vxUieZwdsGU+6pFx3rCXymie4snuN5h1vbdA/5r3heCunYMCbNBqVlP8216VEM9vqzj
px8ab9G/JcfEaFLlRWoOTWv8YcnuPa0Relm2vH3jAZe3RlhpAvEDoh+/ARe9d6NO2lGKKX1npBNw
UHxl28TP06rxGh5HgwG6uR+2+e1hBGY0EayE3YQ6fAlWNYAR9OcIEu/RFG29mkofKjEK/yLpFlKG
qQIcLxypBi93rdg4KIqo4yZxy5KpbRHykBu5Ts8WQZeVc1/btTPlGwONdaInThfLn8207xVKtv9k
42Jyhsxo9YhOp9xNMqi2QXZxjnFC/b4gvyHL8/rBlAJEnlpP1GTL7QSojcB5+QAYSHOrBCju2nFo
1+yfvTtauh6jCjt0gmcViYTrp0lZf1ononWYQ7yrLEnRGyIGK9gl9UgfO5FSw9BnDpCwdPFpGI+F
QDV7RCacsqdYxyyENRonx+T9r+OIALe5H1N5DTTxwN40UEFxxYzcYt3AopJfCVKWDNke1zW27DUE
kZOf0T6YrIQX4crVU8xIbiCQXb6kDzjyOppTPqTrXWjNzG/wucUyM22U8Ce4CFZSP6XfEELOJgD6
fjpgw4KYBxRRQqYyoQJ0aDsKfudzvaX8tySK7zuTo7WhZHv67d85SkdbT92de/iPZqvRSu58C9Ee
OETQTR5QmtaToxpAdBo70uOu25tLbC+L6Ku3KzD09nnktABxANxouBOoYk/Cs+kbaOsZdWnUahHo
s6oeIX/FMmIQKtJJrRntEweO5jPuZfxCUm/+G2CX6MoS+xMyQ2bq9YNRupM4oMOjPIqmDzu7Nv8I
5BynU36in2KjPUgllJRSf4VEXR4q2UN6jCNzIjjLkCsjl+6w+JvEvAMM/3QpWMebN9p4tHAv2VKc
1N5jSFsRsPlB3IYyrpg6vxvpRX0TG02R6wQ0/t7fVRsDp+9tS0MS73AcCZmgnKCf84ZEL3TUfo/m
oA7SJO1yI8nz9OG19WREWcNqy9cQK+E6gNQlLuoK+sP1NM1+WVwpMJ5gv2i2TYa5mslaKM0G2B6Z
t1/JqRSH5fXf+3hof05gE5Od2qmyZiSK6yDjpgsNhjpC92kRPZnbPdmdFeI8akoL22sOyH1tIxTd
7+w/PxGfTtjZVd8/XQwHE4s3stBxpo6Swz9Pgdf4bGgPxPvvVQPZkLSCJGLU67zrCVkFUuC3R00n
vBJOj68YLFjl8YbwgIsFE9/sCElwchGnpfCuBzrZbUiK3z4isckkHlORgBRsMvODcLVuFw/UJC6a
+mGz2hYUlxJt8aPSLAeI8X5EdUy2T/84DxHcbkdXg9fB/iHX/Xnq/Zi5ybWtJE5sslYF7Ox2UuQo
xWASct6rc9NFJPeJDYu3Temq8zw+LwNSVDrck5pzkaLWxWku49OFSFxXR6iAJaNAVuG8BLhfviC1
/JyWNzECYAdhMzl+yPxkgqJfcNM3yyNkaJGXu3lu0OyAkZd/CQMSw5HcYu+vTq95X0ySh5oqR2ky
+2+eq+nCw7gxDPi0GucynMKqj8siZUPiDhFd+c7vXuz0AmudNoHkJ5D1MvQLKFi8cdqkAXo0O4y3
7aW3IWIMclVdk3pZ/R6meoozWpHsLVc+sL8G/Vl8oBICaytmpJPi0LbECDkDqfO39C3n9TdYGq/A
IDwT/dU6otifZydNQm3iMDO6uLeZzo3TXkp6jvIvf85VNyGl9ARwiUOx9bEW+Wi7XRTr/3t1fEwr
cmTeIvUanzCO5GN+ztN2xhHogKLXTDuGozrWQXrJp9E9dlHzqP634W3sqZCMVaFFcx6CHfIkItxo
PcdCLBcOodOsuFd7dSJShaKk5Upv768rtfpTKPD9zS1+tKiYIf1Wne9b6f8QMr3TFUJLjy+7z+wg
gXxT1ssPQ42uTtcdsrXUTP8sewM/ht+gxaU2vucVfH8X7wJwvzJlcllDqC9qsAvkj9BBj9Ctn6mF
RJiY0mg1lVos0JzlKmUg0qCI64DqcS1eRapUxa21WmkYLvqvF4iikadUMls+AFhFqExglVReyN9s
b/VphK0op/jjOv1+ImCW5yKP7p9jmUvWo2+DrNQD0QZncxW4qOC3ITz4rV4U3qx43rGq1DWPkZM6
r9H1rn2ugZlrTothFaT0M6/zKwYwJmFPYoDnrDWfj299+Gv9+xnlw5Bf2WlKjmnJMFp72tWnhA2O
RWBGQn7GqA+y3tOzaqN9TstMA1wglv4ldOWS8IxPK7MVHjQPSZpbYkG8h0Z1ZxVb82EP3xGbyYHK
FBrlu5p/MbI5EH93y/RROrAVgS98GRQs18CXjUm7UIbZc2BJy7zqlBFX9utynd3kebxpelwzHQTA
0TrQxUtZYgT60ow87IHTVbhDMQ3uRMCcd8Zd6LwwVvnB+LelcPidqiUnQU1x4+V3MJVyIEHVgsnf
ncsVJ5mf2eaB/eOWFTeUlxxcvRyeDimbjVrRGlvlQi97ZhzDXiCSe9UDMJQ2iQlqZiiNd+Q9jeN4
TYStzno/cUc6CAqIrbcqkE4AW9wxBxI9404Qj3HAKoGEsXv7nhS3J0QXkGCPZ+wFO7kKpgqDI5wZ
wMtHWlCrGe6sX7UxQtTAFBX+/SvRbwcd/gNIB+12+Dm14JdIshpn4B7P0ErVYCY//JX4TvSspRUL
ys+Lt8j9blfnUSs3LWHXNiUZsS3nuT//eahpv4l+y9ndUFKZ86kqDW8lVbPpxERrTy7aMXJdnFRE
f1uOBGc+a4L0np2oH4J3W03pWRlli15ErFh+Z6bObU00hvMABvmzj0SbT7xxNmkO5X8ETnmyHkcf
L0Gbg7waIj0Nvc374yoWLqaf6sFjAJn6sJv+DHSeLHCB6jbxy0L3kaGzO0bn71cjjskrCxYjXyVy
k430J01zzTDwMYS9saGQu6xhQlhaViu+dRsWp42mgjqLBk8sVwbcgFlLRbkmx+Ubn6r6wlTA+BuT
K7ZP9Cl7gt2bqw+wzJx51DJmGRi9Zr9Hit6V6S9QujJvL3z3Mzl7zO3GkOohTMkoWpnOQtZL75ht
zVflzNNLS2wQOp56kXr4O3ZYVmnNl8DkjhkkNb1jOBppIdz5QrcgFzwarYNxryl+kJM2eommfnLy
YUzpXVI9LgSnTbtzoOqB9qSKuyWElkoEhqbzMdRsqpFM4s0iquWYeZjY+RkpVA3X7vAHdlvHdt9f
rbNcHtprdPV8a3mCTiV3EaVKxokGZi8jmolx3HRSZ5RPrI0fw0+Z6Oqe/D7NchZN6Dxt0vQcFquF
mmbLWIofEQOKv+bCbR7hsb1WVmG1QlIZW4slyH5JZ38LFIUGyVDGx8DmJx48By85/LV8p8VKIuGA
azI/aMGXb9+rdWf5xKxhypvNuSYph/96pkc06LDhyMbUEp7clJGGExFAaVctO8oLQ/vyqUkZEjMQ
0+v/j42rQv1MqEtt6aRvQua3dFecMvSuUzUFCFFI6Ubv/mL/z8yC8N2JDLJXCYX4rR5Y/oso6CLN
jSc3h4yO7/3MYHbYTg5Nw2/gEIN3+72Msm9RujcyeP7gqAt7GnNo02sZCLSmYNa3ClO46beP3O0A
bm4HM/KB7Icye1XFRGU6iwWSibURm/ExVEiQlfZVQhQFzdl5ZITc4RoP6RWzQ7ygDq01cukPhy9D
mPlAsKkj4G+SQYf+rQDK+InJSiOAC4xsQjw/tZb3DeuB3T53foVikQeLkqk14XKFtaRrGkhxo4fd
Qkh5d1drfYo+1YqlE6PoZcLO6a2A8dJSnPvF5kG1c9HmZ6kPljtNc3Fx0ZVBUmD8TvRrLyRKMvse
bRoh8XGk5Qrf/3Qo2mvzAnms6EGiJcQ7OUef2wMXpL33cfWljPQgTfq1BnYQwoPT6YoZukM+561I
B74qVDUufWoo78/xeMncvRERag6woZifG32SYCYwTjkOf7mRbpOvasVvv6U8r1V+2VK5EL5ZtEho
uDNOYpHLI2KwM56U7L3QVKsQ8LRyLujdQkturVmFuQEC7bl8njiXnv5XugNGtA6+CfMVQpoz79Hj
NDE9N6+OOeuHoQ7chtaBvMZBchf21ITd0tBVFaxWqwerwq3h5c5GpDk5clBmSpfKC+xKpB7aAEnV
7Ce9rI+FOp6d1Gm5sFAPeflGE+psghC0FNag3zrjQVlQ/H40SoKEUF1xHOtQyPM3Civ+xiF0inAR
E8DeA77E1M+0az6afq+8mbwyw7lcpofNlNBE0mjIZpJU252AdDOdKOyCgTcIl+QYnl58DBwlxKbk
dUrYdTztASh9sLzJFeG7IMCRY30mw5l3EOuXDONMyn/G2ZFnno18zwgkSRuXYuQCrNjCxnvmGBm2
HWvCAqzrspFaDacBuYjOpo+PsrrCoIMdz3td5WH14xJ8tFA/K+wrGPyQtWYCgeAebvmM9P8gLM8J
NvBZK2+pRgiOzQ7xf8NGbLBGE5Ydk1Z3YEn/o0wIUW492e2ar/Z0s17DNOhI8QJCjfbUx/7SK92y
ysWT/LIyf42otj/snDis+FwkZTU+Xcw4O92D/mOduUWtvIMYNUMUlieunoEVs285dx8Ns7KG1Ng/
GDje23pNaUbE8UKsSVNBdgkfY7ewT8whxMSzSlfle477gj5VCVwAQh4DEGD7qPPJMmtyYs8+xotd
AfSRazK51lUeqsFBV+4/EKoMbza6+YYkU/4tj2ePOKEqEqqQ8i1T1uRkwFAr1/9yX5G45axfRkB2
EObgb0GwnJt9RJ4x/cb0htede+PD9IV8BWGNdCNjaw/l1RB04+Dx49KTLQj2ddeAVO4+m3CxKD8u
Wz1ksz4uiB7OLnmp5/vN0JycGrgDvZBJxUzbQE3ZVAfTfpu51tHMT7qhS+JT6YEw7yYI85GwDEue
REn4YOM8nTWs/Ib528KyhEvhKV2g0mwdtVpg15DcUArlPD4zxaRIi01mcfU7MJQxjDjKa9Qs9805
WS2yuFum2Vf4QXX2n1UokdbgZPrU5se8sm/ZG3L5p5MBfDaZ7XafiG5TWDKwGc02qk6iILABueRc
IOUDIuCAf8HCdmVjJ1rDjqSMT8pnxqgBQZ3RnQgXTiGd7wsl6tpvl7BGOXr714Sr4SzItxlr7qp0
41bSDGkJ4v1LrpA9KE3XPIqNmAwGpn7zP0IrYp4ipmVxfgj6KkgzDqliQiJYyb1S6ZqFSNSJJ7vd
8MW8gJ9XTaoDAG+mv80i9u++QgqETYU9i7BuyE0QpZMfIVQArzPoMTw+FzkklZyYR/ch3waI32Sj
760MMBohFRxd8bgTwq/G7aHYVRtx3qDeta1Qx3k8sVsAmUOFwedNmOf7Gu+jAZKCTKpdyYbIY0GY
FsZvvCMGKlkHBiTPCyK0CQVoZp7+Y59290fxTCHQOPWjVig8XbtbXQdOpJnWt6z4PEu++Jm3xb9w
FPBbt6A317UlAeYvWasEUtUlk0g/0uK6IMjgzAg2YC022jiy/zAsz6pLYPq/d+mZNnc2FJ6Ns3fU
HDtasjIJmndm4jmVO7HcVINrd96YmHfYmg/NmoKH7GgOGyloOIk3RIYhYkD24bMfn5N67kgaR9hm
R4D2P5bQhzlfk7JZNJNthbGwOFkQMR20oRuchC+r3IwgOkP8Mp8ZZ6WdaFNssrOwHtXSJMV6FEsg
XrDhi+HkK8OWgN373G45gvuxL158Rx3SA4QdfIz2twYce0wQJPhIPPWxMZsj5IllW0B0a24oDKQe
0zjwzBmU+EB5I+sU+y2gCnF7aIGbdHtAmhnZCwif07L/jNCg1E6a/CJU57grDJRS5nO4Usf0K8za
OJSpPPO47RhYQtJQqPiDSmvAydRJumLLM/zjUN5d/vhetIUb3hJ82yyySrNxxdDQ8h2As14Fcy9x
kgucABoLY6Ym3HEppLQdVpPEIDWt6QsaRi4bjyRL2fW0ntyH7Cd4XIWwBkFxW4ZJoqJxkjAdtwIc
t8wdChFnOxm/4yz4Q1aWjohzbMDU7w9pIVLd49OGrOkQA3tNK/gQR8KU1Pnbhukvm1BuZ69M2DKy
WlbXaDjQnNM6G8CyA8k4e2IIkgUa5dB/5MWBjblyKgiHaCwVNKYIxpGGfHnd0RBIu4E11wlcG1Yc
mpHsWlvtQoZ6GXAilUkxFN77S3/bkskY19ScPxrK44F3a7MmHtgwv2Agya1UZArkfCe7Z4c4Yt+n
66cfwpMsBNNYXrluV81r+4IbUTS3BNQh6d9YH7a5m4Gf+6IQo3S4wdCYS0d6BLxqXr92fnCylGgB
D3Ex/eBjEf4cyK/aQAP0pYIgv39wEkliyZ69zAy8GsgvmP4yA/Bl+9s+N7EA63xMzCvaJpOsPaLD
nsI+ZJQ0EAq89aXPGbni7o13F7xod+GSMY/GVmrkEBE5cEfqkIO+Mvo8IdCm64hwTeDj5GW5iq+2
jguUpapX1qUCGFlMoZbLGHj+6nl8D41Jx6xK7cwMJPGXYa5yM17T+uYC+njM//BcjHVDKoBnMy1d
1A+altdDedYgMQ2/t+9m4hJ75Q+MRBQqc3vYPA3MXAO2IxpbFh7BE10iBU9Ea7YzpCISnDky6qGx
xou68WqmbOrV11vLR3q4/LDFOw/h9Qf8WVnWCh48X0lAsQyXOSnTS/haN5dVBWG2CwNKTYB1w2U6
5IV60usPJUwJednf+zzawVs1h9Bb/0BJ3kC518jNo9s1dfD693vmViJZ/YcZa7gNCZSY5zafqzQP
Y55Rfai8acJ/GEjn2T64Qk0iO2XrQx04u0zdGTQ0mphoXHCvEqL33+1BrToFslq3ez5+/W/vD8OX
zFoQkv2rA4pXmf6bGgpHq2MNPi94VlNKDDpjMVkf6GYnsOAjG50HmZA5NRfP6n8OggAfJGJ9anvy
QBR9loTNCIhAQvEigYziJzeimeTg3eWE2tnB9n4p3sJ1bhWZ7JuXtr60DK4hRJdfPrexJnT6XVIG
tDXSul67d/zSTQPRRgZAchdlPtxdyfnHLIIy/bedDsD/ebFu0WQETxghMLFVwVnEAcSCOX3deApq
KtTnVrE3E5O5IguHE1PNRQpRw5L6D3DvqukVnTpOQeLBH8SOS1hFUGzWQEK5jZHVVUQJUXneYhIG
9BgZne+0YBieF9qwcZaJJLa6XcjOHZoF3GNbB6uO6TFkcoZcHk9LN1NCaSRRNcxPVNAyhkqTh06q
XDS+2mgU3M/2Q11qcMrGrcHyceK4wZaLH1a09sn1aairh+tz8ZlKL0Clgq9Je39H+aY3ZhqeKmqn
Npvoj1tPp9EhKGe0C4yXrkkoPPjo/g3kwssjZ4H+AyER8DvErFDap6Sx5wA7hstVjAyyveI3p988
+vsVJNPhJmd5Nud0Fzfbp7nuM+ylrIJrigVTWALddCtBrqfBsQS+L8MuohSdfCbrAWa5z8yzTYj4
0Vfia4F3GfYLOWp5/dk5IUk6ZMIe/4e9+FqiBJjWqDF7UHTIHLqpD9xkElJbRYaCCJzqDkrZFFYN
hqWMs5VsTjdULCXLUYi+2TsdgpCL+tMshFUwXs5uWe0nQTRskIP3SegAaVxj2M8B9SMKkz8fzkep
xMdyKwYVGGeV1vN08ieySgWou1d2KDXsRal33+eqbCXD6cWubn71mkwhqX/G89MrPMIH/ympAuKF
Cq/SRzpfHYyWcktqx9gZFSWMp26vFkLJD7ynTnM+d6yuLPrNi/ATWx7Hu+fwTx2JoDsf7gqg2Etk
u8klUfO8igT/Zgn8teYpe4UvqWGD1UfjIlgeYLs0sFCwyxkwL3QmTVol7LU3E1B5gXIxSNP5GxY9
r6M76G9f24VIB+/fyRwTEAeTnIZeJEBkfiZEGEoxK065mD6OLSHIXH+Wqelh28DMGxVHLwaSARxQ
S9u64/vcs0IVvfniDDpfGAVV/Grc9Vx/1OeCF2eew1VV+kJZXLkihdYMQi4xKyQXfJwe0FjrF6IR
1GTz/mNeu8c+YLbYvywQeDRcsk11UYqsHjPhKMuuUC1/omXbK4eSiIdCEvVPcUDv3Fx/FnuS5E4z
taqVIGJga1DzGxANfjkyZLd0vxj+CYzNbDE0bTm/Ug11g+g+H3RWZB6g+MP89LYyPINQ/DkZOmx5
CS4S2XKf6SEVeAXksLlwrEO78CoupyXu6Ezj9qf+y69sweg79OUZfxoIdyj9sybkDBjgtso75THm
vR1b7PMESaMe9apJMn7RGW2yuYYv2VH1RjH1upLcTJeaXoskrlj71HXNnLkIw2oFAG2bU+VRHQnp
UxNwQ2U4UW1EqwE8yWWgQOXoOJMCbxynmSPMNN/CKufZeFJN6DiIKKxO1spNUL9ikUAg5s7oZ2ME
d3hMXMHZZ/WOE9hddQH69tLIIOmsL+ormKuay9EgzJOy/d07ri1TkkiKfNT+zG4Rsh97Aw8IoCsD
zT3rraMfsT31QduIDDfavOn8JYGiN8axXGWimdBeYKXw64Ilv6a3NcChIgihTNm/6TVRtqhp3+IG
9Dd97ZFkaMXNf90YB6og6GL7KscVrccElpfKANmunoDeq1wRX59gIH6P9YD/J54o9bWN1c9do+wZ
d0zJtOUD/zBJwQHWghGxZpI3GGNJxJ/PA8w/moW89Ol72hzsYl7l1+V58kaRtc/ZtRHtMgfLad+/
dWf9X+zVOq9BFk51C0txsQZirsb5HJwG99RAXOftW2EDI3B8hyPN17kU7/jrjIsQL1sUGXDW6q5c
J7dBD4Je1oUzLp3UdG0XMS5Nb/fsrh6sKHdaN8Gi2HH2abvDT31tiGrGNDLvy6BDu895bA0mqsLV
tJvsoZp9ARhdXYjdzu1qMekljVkQm+aeqosSGHepRNWo5T8TTOpzBViGWA3ZJ9fao04kIjcvnPoH
FfuG/6uzBhMFBmj6n8+DrP3WsCKzS76cvIWyALm5a5BmPN8jZxrJxIIxiYzh4wFsNoCHP+oDbVLE
OBlfku5F+CzwOcpXrHZ/EEOofGjH5zTlX5pe/gJG1FS44uBZ1j4ZG0+5ooWSb39phvi6ld33jfWp
mJkEKgAddjbTXstE/0D7thZANe4wMJkSdjBmhrr1mnF/Un/5UyyYU3QCrYgaP2yMIULVSlBFeofd
2OyzenNhRiBaR5GFWANvXQxvkrss+V/lLdILnLbUBk7hbbLBoNGJuRGPyK9BH1QkTJVH3CpRfEeN
eC04Gffwu7DtBNUpEXtZ6+OrIagsvMqxRJHyUzK1+CboOA6HOtg+Ef1CKL6ObBytG6U4TZzhWyAO
tT/UJreyd07jKu36pkhVDt7d3N0jN1G6IZeciMKQMvse+ZS0ci477Xhtmle2XIoZgvSmRTORa3X0
yOIgy9ZJ7y0k2AXeA5msX1ORMytSb93c5+T53Zmm9SL3XqKEbKCmXDrmOyDBtvzVNUFipbko/OE6
Ru4yB3EucfEdT6LiQnmRkroCTmMQA4SxzFDseODLimRTqTs6xaH5kKhowvGAE6AYaBvLkGoWaBUf
Z0G8K9rlH6lbGzv9c9ryr5atDP792s6tGLmWMoXXMUv3BdcIsRUzmbd4j8sp8rztPsMbYxqM4PCP
9o49BaESvk8wWWGfKq1sQ0Q6VxbElW3xaCaaFGvffkz5Iu6PDdM6XdT/Cti9yFehXpVie/Zilf9e
T1YSB3N9jsvE+NvoHPNVcNFrgbWjSC1ZVxY8a7N6SV2vNQ64xUjQJHWQZwfv7uoPtravaP/IuLOy
bZU1/UTWI4w33NdLZkgbAiemuwgsYl4qHRdUlWN43oaF96FhqPg2r0b9mge+mgFxFejL9srheB37
glKFTfovbWpgYsI0zVL5whYUqjyBv8IJUBipNXNO69WLlLp1CLkUMFhEm77qCrb3iUDYPKNUa4Ev
IleQCSTkW7++xPTXPCUUR7YOcXO/x84UUyiPVQUPvXxMoU1U/K1woSN8snAWydYVqfETrCszfBA8
TXrzXTMiRqQcgleiLRNEaBO/lc74N+HJT2Fa3/v9zCT8n11AMZT/nE8SLQgokarD3Qg3OrLBfACy
jds/3N2GzvroBFxypBHSVj/d6NcuOKKRB4owCHbN3wH1vDzuDh+c1ba3rUHZx8Ln2jV7wRT4kUq+
LqRXCBsTB7zMR3vC2GJTj9lnm8iGJmZ9C/2dZ+2XBP7TENNRuubM3vGWlIUdH++/NfgFtVemHNXy
p0XltW4rvRGtGaQGFGwAwRcs0DPMyuPyTG8vkLHTlhTDDcxaJSxBXauWvSecCBkoAwvdzcBosb0Z
O7oiUBANbD44xqg1Me99ztkjYMKLugZU9Uh/RMM6s+EMMUbTqkwhVQ7ZktOdtsUUeDmC5v8pSEzU
uxg/H2rPZkwJnjPtyKwJky3bZYamTZN9KdV6c4lWEE90Se01BSBq7KNamu5DzL3VILhkeLJy+g4D
wPIeD0aoi1ECVG0fY15dp0mNDAGWQP7kcHYjEjRFbOV69oeMwjNaima/3n1V1envD3WDuIK1Op+9
bbw9ivnpIQem+3mXnF8N0jYHPAJf4HP1JqyrNvnHl1ivxc0u1BK6GK303PN2bZ9Mpi7OOmsQIQv5
9y4JclbRMbuRqQKCkeyap479bYdyrQeZdIuTCd46aooW+ffpCpmow8kyE1jXOBPHC6fzQTXErubR
YU/NLf95gFY4EoZFna201qwlm3zTdoeSRLCwjxVdY1YfVMT0tG5NumVyBTve++102ormauE/awuJ
v8sg/lSirTGDuDBKfvYaV6bFbfuaUJ6FPWh1i+u0KDa/QNMdHqeUcBINhx2S4+eCk4js+I30tCRX
JPq2V+LfgAVv9+6jqffHHJHqohKPex5Oh8BuHQXLznSLrmu1NAwYl2HPMuO4+vwL5pjnJIQrdJPt
DjaHcX1Xa3oeqj3r2FDDDhs4bOJ+YpxxZ26bMfF2nkl+jWbT7qdnSURR9gx8gYCpVQ3P/fzY435n
kDTHHLWXnpa+rJVbnK87fnfQVek5jjYgPZ5sPqnDjfn1svMJnJqMPf2DtoahdQ+oVO8NQV2Ej93q
8JtlWOHq8OC70lF3zMRUmmWaMiLa2OPyLhqtXjDfjXcQHu68rF2tpEq3f3JYVx8zzMPYGL2q1c/N
GfN6qbXeGE2JWi4naAEeAhylYeKks8D5O/cLwEMcnOcb8f70XmdLSyEZTiAnZPWNgUzT7z8qtnLR
phTdjehDywhYNhN8SG6Lk59ORNAcMwWwEEet5X75Jjk4CU9+oEWsC8XUdCvnjx4hhKg1r85gWxnQ
GfMRWxJ/JWUX/i7vk4XmcOnRiOXgG6wmgOCMZHHHYM9IyeaK36g325hmLxsKBgpQh3dyuH2erx4i
mWPs2ETxUSiu3fY7s0KIdHBNhEEttGWZBtvmWgdRKS5Y8RR3He/cNQLxxfqGDtPiuZ7rBxPXm+vE
wzA2+thGf5W/4saqeCr4+/8WxVXmeH+EIw8gMys76qTGBGW3KVP0sJes3wqx/Jt63i5gvvGxCnYY
NNnEsrl/C4BlXqjWjPUt0vBXy8LBWDyH23Kp/5A5bXMpmTUrE1VVcCyV7udyoSt9gg3DTeO+2VWg
tPiIwg4NJqgwTs6TGdDMdoa1K/58X2eAqquJ1hB5PPliKIm37M6NCMgP+zr6x7XNQDDHPH8+8dSm
szboHFVp8YhzUjYgHT+yUYYyavjzV+T1X2gIbZZAeN5VvyTzz+itMFv/fQSxfHAAYY6xY1txK84c
KprRIv4tERdrpCZc81agbvD5IeHwF+ACckRa/i3ALWXofkeGEDlZunOpvKFlnnMXHm4MloBb4LZU
PaAU0Opjv8coP8IoHf4QHsAjhGzBS12wgvE9fcYEjn4P4ZMD4pgMMuROpEqZfpTJvceVadF3pIkg
xr7Mz4Sfz6l4cjJ/Az+mr5Zsmlc3A3ZmdkHEIyNpjMHCbYNGNomAaZ3038gy7vTyGjl5WoQWUA+2
gPdfrUQ5f25SMpTeflcdU7xFrzgLAfUQM5P6Yb3Ajz2R2xRXKIjqDFipl/IfACao6BhUZQl6MCpF
pSC44ndST1gcrda9Ht2HynO/MBVot8yYG6hR6mvhcdAv6J6+dMc9/qBqGmjLvrTYd6JCdxurKJbE
mwggNnAaMFNHhp558PaVnpCU0twFklEKoz3Ay3bgUWb9tMe+XGPcFVZzEcV2JRTlOHF31EQ0fjnL
FbioBAy+ZC1xnWQNRMRqeVnWIru21PJxWPsZ9nXJw9/fw5Duty/sjP9LxsrTvhgqN4lLjUV7/CTG
Jsdjfe139jhDZlqdNXiJh6Vb8H5/KTkotAcsRvDbSKFuRzObWvNl05im8mCo22YF0NNf4Q8a0d8N
/ucJvu/01TI+pjx1pbeZWDDBUQaWT5sPKi0D5EC3ei5RYHtBEjdNeU2hoyzCzjPrv8+dL93Wq7Rs
BEwR9s69NU2FR/NR1EzMSVLc6H7ZeYa2kpcfa6f2tDuvt7oqpRZh3QRqX7Q45IZwp6PjF34O6GOB
74jTeFr6J002RMZhuVscqPvAnkY70gyuzWNOK9O+VVj7PBTIo9BPI11NToX9+C+/gAvVDA3Fvo7J
aQg5AaO9EDXZMFMkLelH7dID1Ow/ev1971vvAVO4V3DDlnFhLmiAtxmQgrZPClb3WpaWNGQlYRJT
1p8QI0whiZC9MsIKCjF7dia9eWdmssaSHH15z4ZmOFFoFxYciB3xZHm2aJwmLH0crpO5qy0e1ZOG
95PyPCnPVe2P3jTTizQPsBBjjNFt69EDegUUhxRaMavll+rUDe3C6Pfn4zJti39j7Q7p+vo0d8Zm
cnDBv5um/3J6BH4/fjpscMDfC3vuoWZT3gL0b14EEjahTCGqXYrNx7T/JQDk5iprWNJ6t/rMem98
AY/XRiTqDwuGMrwTEHkMWERWD3AMlUECDbyZqfDTQDRIcm3+IRwgEKP3Tp3CJfasOqVeWNWZ12ac
UTgn+fmsW6PEMvoCxVWFUGazmUmxoPeNUdpFUuNehMrPW7gT9CFiqseXaar5EuHKRNpLoPruoGeX
QsuHA3EnGRGjYPIYFUTnjPpzDdvXKHzrx1knhitK2SjMWfwgQRobu6ajF7lvdSxeXRWSk2uPSl8/
T9cB4bIARS1FeWdL1NLYCZQZlSZoOazGk+nQIbe7pbPkUIWTE9CH+TXj6srk5aEAPTvQWscKqABj
Ir2EL0LAPJkB7dcIA12otM6lNiyMMooBDOCZBRyy0m+VOWw6iwhjkEa2sKKNJsaTVijTgAT6EQSd
jfyoZv19LQN2um7cXxH4uZkwXlvJti/N/QVe+RsrphTLSdBS88a+BmUD3FiRP3LPYQOQRkGnVxpe
KRoRczhn2ENKnWJYH7T6/USGheKDx6AnZwlQdKHnT5nYkfzT4P3z4iQJIKQBHZGOq5EAjxcXsWgP
3LaURnhfWZjVm5pdt1CM10ebdKY1RUcEsDkgqvY2UADFDkHK+bpNhdnn3+9v1V9Jm8jTxzCEc/7r
2I84rFSJz56olbyy0WxhEY1qXSBOTKBpD/xx8SQAVu/Dj/g3jB/L8AOk6gl6NoYD5/8CRdq3yUke
neuA+IvrcJov7ucHUXP867dXzxjTw6AX2Dueg73/inlt64bB/WtTpO5cTnlvlT569FH8MUYHp/Yj
A4dxyVw/xTXkCAUVVIFh5CDP3nxUjcXu8j/INERVS9hDBiQy405grMecCOncO/BY4VNWVYg7eLri
vdoOPU8Rqp+d0v8jCIQneZRA6nME0CBYeOmY0DCjSIL9IWcGpv+H1N3RQJ7esW30YAWsYptQfDJ3
5Yd2Gqhtc4O0AhXj4EcYMD6S5tDH3iKCTSsWTWQTTxPlsRhHLdkQjJSumy8G9+bBgkMy5sxMnaUd
y8f2bRj44eOyPAxWmHrd9CLt6deawzw4KqJ8HnzbJ0W8aHfJRMJ5kyAe+yfRayduVbDntktrknQB
Bknfy+tdlAU+cetNkFw3ocRUg0I2EmRlYXQHn4Qh7dAm0WEgPRVOaUCdCd+G3/+m1hguvK1V/3hA
LdInwCDpsti4HMQcShDHvNGBmmyQZSEYkjCpSzg2VwrUkk7pS5SiXotF132zTC2fb/taZjQzcKHF
YANqkU/W4SVuvcGibX1qAvgYrlJS8QeTLQ0M6PXv8klAy9jQlBPVROkzSyA91skOG1DQvHj9bvUt
EprWd6Nl/0iVI3W90lg+zaX23NA2T+jEqib5CH0gCylLcJTXEG5OePt5klU7gOO4zvrdTnGc4EZg
Hc52veXhWMfyDGGKgyKl7OHONHnMwPYtcVkjbBnHGeDIdCcpYyyhf9RfP3wmuCtPztSqHI6HjUuk
Yn7a1HpOf8uNLXNq57t3zeGZcKyfVS2hpNDpvIyq3uVvZky5luS42gw/ArVBMv4h34Z0jHCLAbXR
eJHMrYhjXlRCVpKcutV+H/epT++nboLSXoib1Njj9x+P0Hz+tNX7xCV5zYS9Ljo3JmsONWVQgD0O
D6VvN/jJbTlpRISLqGvWliuJHZLJo+dYvDNBakErvLnp8JhSz9rTV5V3laOJAfxxwUenALj8rCQg
F2OogVKu90CSACCQ7j20v+ceazLZTyMtJoGVEqMXIr4ojAXVNhkUwX3vN0584w388BuedCU1PATH
f7Ez1ZezQYStqe+sDpcrwSB3YAY39Qjvz008IeAapnI4OYxh8mPuBdASG5nwV8dEUTph9PurlxJC
NzSkVdndPFl7AnrUDGZX8v+ygt+7PKgIirFP8X25RltPSJ5NBmtRhNjrHP2DejL2I2OkqM1lbNsa
gFwrEqCs/TVcbITfXWw8q/nxh27ZjHg2EolQlH5b5QXdfKCQ+sGxGQ0icGr4yupCFHIsBMHoFpaR
upI8YcEcSbig5eFtPEDHP3+jxfEAM3MVH6+twXscB1i5ptm3cOLfDbEexHkJsxXVAq2j8HlQgcv0
G1ZX/+KsuLihOqe4DTFaNEO/wM5sNqYrm/8CBhNd23v9eXqRrydpsVkLbdN7CWzNzN5WJvsbnWf7
rSr8LCe9vlPwsBxEPGMtHMyBUHMgWcnLQMf38sjg7sS97oy4mbemVIotN7dNjxNWI/5pqEpJzi3a
edZWczcCDwJ6miPgHfSKmz90+iDnsTlxhnHV9hrYXl+kpup5GH5jkGS4nWnTVtVuaxg61ZXy8wwo
8ywuXQw3GLlDV+Crf9dqaT5JdSTO2HY4HSbt+g5vheBSx8lQRx3Y+OKyIzz1KNzfgML08o1twARI
eM2R5TNanpBvXBZYx3MuXfxGFq5tSrNKUxDqASKQUXJEE4gBnTWL6N88tteOcXR0ri3xnjwC/Y5c
g8EkJ9dwxnlcLaslqXD5n4V0vG/sZ/G30+BNQRRI2yamndP/hk2Il419KFjBbbbuLLC4IYlrcPDy
5MdV+PMTu+RvE3/pFnY3zrR947pk+cDE/3ytiDkWjjq5CdlTYqA0f2sMoiwYiilV+xKB+4+iJ/me
mGsgIKkrBki26TSWe4Qup+2zqWixRu+XpYqgCnqFH9G9GVnZ2xADkRj7nZ0PfZWGrTsJCNk8o38i
lZAFsl57ullK8yGfOYq+aJCEd3bY2N4/k4FSZFFrnzvB03tsE2d+SGO9iwRWPZNXvRxW2nSA0nCa
yft3vG8//WbYn9vwkjdPUTk+BNxPoYmcbDvCJRpXeLgvD3yPefZGaVqz2SZzoOuCow1xWxS/ZbUk
kuH1gZccPiN08tD27P2HsqW8gXhYTmzVeUG+Md+viISSkmDj07namXmQ2Ijh8MM/DeCz4CnfuQpj
T4ynyF+22cGm0Jg2T6awC7sIxmyVpFWaiXXnXQOfDGfosNrXPMraYDUICf4/va1UKxoSz6EEJsEY
OSfrTEeniNiNVkNbvAI8P6qRH9PAteZVM+rqWmliPlvf9Th5D4+DU/RNLxUWq2nlXmJU8UjbJUOC
ZIEUfA+hVqPkT3CySqLo9zCxi29K87T+Bg2YV1XZh/qiCHrn/Np/kTmbDhDkXVilRfcPlt1d4jqB
LJiBvHJFc8FG86GsU1xZ9HslhmmXmmXGqXb1x3QAVF7sAxVfRFJw8eiV7ePoNjQWXVOzrZ0RP8G6
LY1KN7DRcwAJ7IaAkvlpGb8wZAZbzokboWosHlJB8Tcxh37n1DntRS0L8+LoExytY8B19GsIMKlf
ka7gSA+3KUlRYmGbEfT0bSoXJpBAynYoODuXZHLgKxkuCV3hVaY4CXG7skTCZtFaFAdcruITGsFw
QVEeymZWTYmlLYYmKwjtr8ALczip9Icv0C4+16FBUrB1/oHhBEvkLc1K9q9D4w3Usn+I2KIpSVW+
LmQKDzGDrg4JLRuOrhs3p8Dgwx/JzZzQLEXMi+V75m8Vx+jk+wbnoQxwmgAeNFJZi/fAiy2yKrV2
21+6UCh85ia/HMST+zVS7rx144HZq9ULOBsaLba50WtyNFjZw3PF6Wgq/NxIExAeN+waXXuqEd0g
38M6iUA02hFd13l3LURRY48GNskPCkwd3E4DSrXny3LglwQ1TmFXJdIvM8mdEI2+UeWKk+qFhzvb
9Ze6N66FaOZ65EsbJhtRI1iADUHgfS3hIjCr7JdbJBRBgsrWvY1XkfQVK6Vy4dj3FqXdDPkXUrYh
1W6eCkuy6gOPwkoVLhw1vBhjUsBmqbBiBzhQa0Vk4Pg4evdIr7Cytlu6BKNcXWsAQgc/Z9BOVxkU
jcF7Pfi4YCdAIgwBrY44vNu4QgIMeJeGpyeUf5qeqn6OHHsmscalutFIKovvVPqWaFQLyCUS4qyF
vCijullUvDERNQtsbxzb/8s3AB3QQ22JVlDKSjKZj6v8GSv0chPnXjWWlYTZwOOesatgxMBloBhA
qOHmfgRtF/+/pApiLT/hcwmnoKJooE6aEthkAg/hwUIdrPAo2yetIpDg6fhxmpzxwjFxefFkEflu
hZG9rI5AO37U2LzDBNzKd7DzJT++GXvzWCVtLCA3aLKPgRhAZ31qld9kixsgGe8ZPD5xbRyPLCvq
pW8wsYsg+ql7FERLPiiyEZ5uK+UT6gXsQEyPolXkGYWAoc+7dqOs2B5R7c5+ELHFtISkUi7LtsLt
+AlcTNfnTrnnxdphlPlz4YB4pObJxXf4JsB+J0pUb4RoR3pdZ5EUht9vmkluvTozKGbJwwGsRbAX
+I8uvhBe/m53m/wlkvVV/D8Mfu7zviTZwaTe+zFlJ6Fg68FODr6TaL0oF3Pp0xmeNIMA3LW4s+gO
rfxASMyKbZ6BX9csmi+d5gH+CbQUC4h6NZE5j0ulXGHLW/YdCRCfSFmK9y/L2vsj3Do8Gl2aYay1
W37QrpxfCQpx1TTUqC9GF7kkK1VyUN79Tjiv/FeD5Ikm4iE+lPgWrqGvwazFdC1vykj3APhGDQiO
gVm/OFJ65Cm6L1U+Q0K8xtxePZ4GGOTCB/sJ7qfIlvvbLX5wHHfK881yKqmwb3NcJa/A18+SkZgS
qMQiZD4ip2QohEu9RLHoBfv1GSrkvBJVOgzOh5zpg3zU6WpsaDALBQF+8tEiz+MWIe8nBY9oJC8D
+eztnXRWMK+u0RIZeSOdlNxaFe8hMuJpzymfR99w2jKbDzZq+u87WOQQ0VZbx/f00Yh9d1nE76BA
nKFaHRVnSRGzdNWmMYG94hPMLm5QlbO2XKtmMykTW7yCb3f6a75sXV1gZS+y+lLRFU261hU47FQt
2A0Ks+FzqPiPBF/V1szc4yCOoTi8iQkkpK2p210b68lrweqh6YXLjInNoaJIPQWUt9X0LxNf72oi
gYdM5SFEPrqJdgOrcsbSrYRkJ9v74fltnNx6QHOc85tG4z/GsVFFZCXxD/UCeDZ+tWlHxTdtZwec
9azx1MInG1Lu+BjV4J2IwKeiuwY7zH4wxGBZyKFmv+506gHLMLsWfu5tHPzlM+wiQ83J63LFkYT+
ZbWlzONC+bMhCga72+npcZzyYAvaYzB/X/wITjPmRQ8EpqU/qcMSWcT5n+z4zZR7cokCrxffE/9C
sptcekEVxPkNnsvVbLqF8dBO+VvBLnpnlbIxc3+ujt4LV6tf7YUSy3K6HRl6CSBXai3+cKbBFBB2
Da0MEprnwlqD2p/VasmE2xlvgIO6Tc5USv9N6uBQXehy9Ctv6kh6FQqY7Qyw4XanzTNoRug1uIn9
/upcrAsY7JI9BwxbZaIpcFD3YDa4vSJTGLnEpq+OWtjuaY2xocSLzWUcLvQIfr0MGPYCqK6g3wRX
xBLi0mGZkQGrSAvGP49DdT8ab/oyg+bxMW/AVhQ3QKn1Gkh/v/TDws0kcXn2NsamsjHh5c8wtdkm
kiZLSOPOgXwrrwYir0YBnlTUdAL9gAJdUTejhZEfvE2sYULFLL8ejcvsIyDuHbMbtYtjwUMUeJ8P
exhsc4waoyhJnkAY7/Ax05aW919vjBuCPRXZJZzfk/4M2I2DSgWUk9jowj9xIKbXGplv31I/kZ8O
S1Hw+PjyutWNkY7cwk8H8GsOw+l4+05IAhViStxIbLYah8FeFjqOiouUWxeIxr/4hkUhBkUuTT7a
RKlBabEJDQSJfLNaZgq8PYd/bPq4sCA4wpTC0PhLUNr6ChWzYE4KorNF9HoZoaO6TBExAqlSm4Kw
C2LueiuxpUgEEUckmyAMVG3c6nNm2GpCgRfjzxoGxSRSq1gyNGJmTh6fgqDXK4e6HfSlj1zelZv5
JaisXq1RIEgrmgF7UmUt3nQqku1dmrDtxKeye4lBROxV+qj0nFiju7DVP19ZjZmDylQWomNTYmTz
huSbmfZwfMgS68MNv+w64HhM0O6fvMhn7QB9i+TT2JJ0yRfXafBLuZSsWQcC36A4bVEUfZWUa58p
hZ5gFHX/yWXmKkVBv1YQnwkvceId4K60uBFOtnyHEkVhGmJ3UlIiiBkxTPqD2RMDQ27qpUzOmiv7
5LTpSzKTbeSwW1UT+qNUJRHBpSofP8kQ3Vv1Vv06H74rz3Se2jCrxgyzV5ZWVoTGe5Ptvjsp/eVQ
Ey7pd0NfIpx80f2ykNKSjrTlFXO57H07YdaJ4DmIGrCP1MvptwUvftHwuPdIFXvfjdHZ8nfDHURc
4eBxZPV1VwUStdLy47K/xos5H13sNX1YOv7c/W0DtlX4WVnJMfU8vFMjprAcqNNaSBUDBcjXoZ+Y
CN6rHe40dPrK8SjL9Z03qXTZmQ5pUcAzAgDDmFy8E4S8ehSIBMltYuIC2tOrVLxElr1IZNoHej8E
665HgFwstnAUoz6GbFw+A03V4X0poy0101+VwXQLVU/0CMca4F90jxuwgQyveJlC6y3rvvjGu9gS
VoCXXdOJVljiABQ69nb4X7LL/GR0dWs4KbkG9hrqh0FKpjD6blo0KVQfV8P4QeYqDFP3xyykldlJ
rKrdMg8pTrgbxO1zXGsrQOend6+CyK2xVObN4ze67cP4egMbRmP2IKqi6Hu6KKP/DjJKV8uSsyyl
ROIi0sWCvqRHtuGxs6GK2WGBBur54tjyeVpMdsZ7M9pFwqPKb7OfffPMAnfIktk3rcxBICuamrvj
DMNHlJP0ynV1Dt5qn0WVuij1RDAhOQ8Qn6O7w4pjn+ulAB/cdriPrxSEz+yLIvYBId9sKl3/FuBR
gDDxGSM/iAUgF+xgHbad7+C/d9aEPAfWIUWkJYyd6c+o5Fr9JhCPrmG/Jz7uR8f74FhTQoZqeZuy
wXXKl7OYyx8Y5ygTx+yAcP2pRjFory+4U6qELCRNO9LXR5pyM8602QjLD8iP9ksChuL6QheOPEGd
i4Os/ewdHFCcgL1O7nmWgHmnHGhJE/NCbCNHOMC4huFz8C2CHRXAYtGa9vGvF0oGRp26ewULnT9G
qTXIFivYHzHzv11QPpkEwTEN3JoMVYtVIwYej01tibcULeGSqTR+ZGHKrPgv5sa6cdg/cpTNxM/J
J/5zJayIWIaZA9xpESQnWI/Onse8cETP0UCv4uRaeOPR7jeviOYdJQ16kOARt42p3MBRJcDktk9D
wi/qWBB5icr9UPkoiGE2EzDo5QMhxfFqAkif+8gizPP7qbZCU3OQel7EYUMSUlhHtjeBO2y8Fbx6
Dy34s1hrba/6pg/ggQwh8l/j79ybAxoQyd7gAOVquJDYueAEy5NDDuIkp3nzItzpHY/X8vQ1x3NH
fWIALoPoQRI8CNhISnL5k7V9uYG3QDlumpDK31HV7JkLPTYta3fNAYnCDzHLccjZxgbKY0rurTGQ
bZqNDAPzTAI5XlMpG+yPUUZe6+dbIHa8yg9khftxhAAH20wl/jDvhArUXBrAxvyNb1M2oS3Vcd2C
wH1QgvZStKw188Tr5l5TYjvkn3Gdw3L8DnA+/vMVRCkCAR2gpswVCyAvnE6SvPwExj1B3AiUCmjD
s3UXQLKSUZhb2n9rK+K3rpLYhQmLzg47PEAZPs1HcwYt3GGHHmLKcHAlVAUUa2yToCtMeN7QcQRG
Qb2ttuaGahXkTnCVHvgnAGy52egN+vkIgkt6MV8kbPNJ5yimREax8SKQ3V8CUhmMNDdxahA/WQjk
Q9G+VB9FpHG2s5xnQ+EtElit65trCWLXVoUI32rm43H+oLVtA+xWhq4GSSqCKmMrnxYus9zMJDLp
y+GAxEPaXN8dTx1QG6G3w64kE9hQj3NhOTCgvwhEWPYQGt2DP1RepMerka0vdXts5JP6unQIzqx+
5S6SrXaJH/2DlAmYbNBmi9asRic6ciMvwpl2AZArJVf+Mxw0PqSyejYjHZ9fuwoknbgS9UTSzB5j
ZFlx9ChoTzvenf85ofZ7agYXkhHta815RKS5KnwKHbqbxRoBLmhcru+GgIVFBAifi5h2IHLZWHMD
kzAEdA3pGEC77jG7X4wYA/1pgXNUxbH1EHGxr8rl4MNESa3AzPwxieUJMISvDGRl/vstogKZqCYb
cjjjmb4LhnkgRwzoczppVfv9915IE+fhp+WGN8L7/NnLJAtbJ+9eabIy5boFqs8k7P3kKwb96Kj8
BDjJwgq1sxAnDEIKpZ0keN1SEn4t2gD7nGG0HQ5nBk6zkDCoWg+GGokhTup4elzOrdA3Fw75cgas
bSiPlEM1Gz6IT1ey4UibErNPkSoTgOVVG5JezL9QA1KO8zVRJn/NA77novW6RUuf7Sj0rmQcMXDH
cshpXAgY6r4orSRcaCmmZ1D3aR1L/GIF2zVEtJf8WdMX6pm2ZBnm8SJ2xVTEqJAPCt30czorTDkV
RQ367B+lnx72ASha1mquhbWnxEVizonmOfALKwgqgnKUtpSXpzSVzz2BLTFn6UMPAdjuz5mz5c4A
Fq5i276PxScAFFYqRzB5qham0NI9TpAwEDvgftDb2YLAMYMw4SyU3jpF9DVdSD9c6Udyf8Ga0uj0
R8EMkFRFtLKnfPErx9v38XaIB/AbGEn2Uf7llVQxZMIvS8vLRKhquEW5cYIcpi1gz16NDsaJ2tZV
9kLJPIP6adIT1gnTcdxkNKfVWNLg7tMrR3Lr5d8/yzGYkTG+ZtouY5u4mILr2P1pYc1DZ9HX5DdH
DY522jzLyXGhNY2GYjVYaKHd192cVUjPCTTuaH24wJjvFuGYCbZHvdCrUTBKJGv79aNLaGj+RYum
M0ukRhO4eXqXw73+dFlYJ5w210H5OzY7xTgTgzvtrYtXqRocvhIDM3RKNi1gQQXL8SHD8aITNiZW
x4TYLAgbX4Rf8Em5YuXFdxv22JqIb2OAz+w8fbxPxPMRBtg0zvNFaTim921fxsLW72aM+kSJivBn
ZcutJ8Pjqm7HnhCxA5lA4aY3c1vTJg2ri+o0acj2Gvrp7X/jri0NU+wVZH7mp9fPkUSfyZPScy3n
f9miLzMIIVO52cKWkUaQgce/IEwiDrE+wBq3x9RqailLnvieqAxXVPkIc6/2Le6QJ8f9Ir2ykLvR
t42L3BfDlRqbVh9a+AF7T+/psPmI/Ei9d470E1Wt74Ii4s+3KxZTINswGCQUJIf3g12bOxQ/8Frb
+/0hf7+hyVv08V50OSiamBQjDii0+LEiy3ZnDjVfm6vKKi5Rf1SCHGekrGSDinRUDpGh+cTRiux2
lo19g3JTcLmiAsSXITImL/J6KbPLJ+5tOMqqhEJz69OrfGuvSHXute899zrqzBDyvIyRW2MUqJTh
RCqRjac8et8dcVYSvl5gDEp0P1fwOaBsnhNl14pXsVzewIjqQpb1k0tCksc5yGJJBIDM1ybE8MmD
LEi8ONiU3rlp2gu1k8t1zG2GMm9EU+zZX84zbJroLDTK+mhiGLqcvlSp4EUy5qIjELClKrnTHscX
dHNOfWBYz2jcjXXu2FclUy+JnYbVG4AubNhtwecbyRx2aCxOENlgSRUHA6ayyGYO8BtqwcnnDWTL
1b/FWhM/HnEhx2KwJzpkrwHbsOFm2rHRGsWVXzh6EEoK1rDw9uMh/Yg8g6vyCQMSJn2KID9ruCTp
EDiDzfSfK3H3jANBffavJQ/myBN8hcXxZmQRqT+m77MbWGyVnJe/qMS4lCpBQVWj+AlZpMXqLdg5
IP9JQ1AkrM2BJje6A+9VJ3Q0Bm3DlOozapl3QKtdVmVT8c/LPTduPTFQn/LcjS7Z3DQxzoidtFq5
uSeAekNcON3NjETOExQ7Xnc79ofX+m6uxUIZ5yNK16XzJ5cIW2T0u4UnOAFfGEWrM9TGRz3Tr8Ss
+Uq6X9Vf6m1deV02VBq6Ar9ECgmE9LRcu6Lsuy534ensvfqesT6jzb0R/mB1QMi4+Qi1hS6PmRrO
Na4FnPya06jZkzAoQw8uX9ZwK0xTc3k9ACLEI5QjjDVZw0fXwpyVsb9AMI56hQhY3bB6PWdJV6Re
LAAdWn/p8xDn2s1q5f9I95G49UpzSZ+FWn3VjKBpiQ/mZcbxla7k33veKfZZN6u0txTcwf/hr6nF
djMZczDs0fsQn7/M+u/WQaus1GCnoAEVZ4nI5DushCNd5bY422u2Mn5UxAsY59l0R5ttpLvncdYp
lX0CUg1lwK2TPkBSg1Ps1eS7jrqZytZeHDpqWb8VdUgPqKzX+JCXEEU5eyXYEkDZTsb7IpF68CpX
HzZfKTBvKaVFi5Hi9A002PHylf0L+GKwiBSOWVg7uH+2I48pxjx1SHNjPLJkCycAgErtqo6tYB1D
0TLI+1iJbkbwZ8a+7lVzpgQ9407ObThDFgX1y71u9ZzO3Xz0GXNCs8LNRf3S24ZPWO9pPGxlB/xV
MHOAvLjVxzCDTm4wtSAOs5Qv9IOGjO5D5Ned/tZt//Q0Y3+VjhR5KXUyhYoXrdN4dw4LqHoGPZbB
sONrEoOMb8fGoWogc+atAqc1RY1xaWTbhIyiwgH05tnIAkHLLem+rKaHqYh19s4Bqc4O3I1Varz2
U8uPij+ZPUmBOojR83ycEQZG0EsMDK6re1FtkvKPUttk9KV9qeE1gLNi9r+TIZL+TURFx6/5Z6UK
tbzQ0WGfhqI964EaYOM9stZbEcCKm1h6Ype807lG+MXQ5aYegiyU2nFUyMKxsS6zxSdCrXd6Fl3m
iSp9769HebDzdoKCJVQ5TC8+87L/xE1Jqu3eEy4LzuMdrRox1ooSm9Llx1kKcVBJs5qL7+nDlgr5
zhxJKlYZf44TF00rE9f8KcH0bU3k8SYibOq+8cUOG2r+JjXxlh3kc0eUzyHaZ2o23XTW1RoZ2JZa
OzmiH8743TeZYQxxiPFJnwDQpNbz6Hnrlw9VEkgSgnPIQtEH7qH2+3KGxAU69yIt88HJmoWeEdua
q7/c9sCENX7SkULufbueNpSpkV268uYwnpZ4g152UX3wdnDd8sIzsd2RXoY42dehEb5098TplbEn
hZeoynw7Q1bnmCduAf8wJRNm07rH0dbbahn2Gno/SMptb8mdfaGrdtPMbjIWhZa/whlM+NKtNdZC
XdQwAQIgmK5JvuKBMXzDvUUknLcSngXV1zc4L7TEJc7jJ+jz3MT3yvBi6SOU6qOWLo4M5WbDRcmt
uMoNeaKZa67R3V3kNEik2AWElZdGND1pXtj8UazAoB6EoBuyCFaSUAtRARW1FfzgRx93FdAAdd8A
a7zadfP5XvSC0r6THTebTtMUqJCGC2QcMrmNDGGGSqTY9bf1xop1JZ5NKZL41BXFSvmM36MNv5eI
jvoL0mTGeO5wzJa7Iwi1LRsnEBCz9YpBkzbt9EtadYw0bxiy+qJgLqr6zHlxCZ8nRNAn/Mqrqb/T
RV/YYKZW/XwPc/+5f0MeITMZbLOdQECeu/WZfqMNPVMUN0tY3mc7ztjwZ6UXFLY68t2TsXuPIvBX
R3HrAGoK3iRpXhT6gXfe94OJaytRvPHaHZ0j5uLS25DSYzc1IiGTQItlXAKKs+1V/c9Fm7NoYURw
XgQn3AOmH8ugfYpBZnoPaVi7PDQhC/6c8mSx6/4kLfhmfGC3j0DzXrX9fJAOlSAy9EaWPk9Nnort
oNKaO68uV+SSFw7SyTtjRFUr3ktpERKdw8CXrNNJBVVCf7ujTHCw9H8bm/WrKkTMjV2ZqkEiGToO
mqw8HgqRO+dGsd5CgM9FupTDMJTtJJcpw9qYmXdwxfSJC8RlnCc+O2C0yqQsq+e8fhbtbfHtO9K0
gWhdqOJPwaF54SslLVcUfG6CI3QELIHVXFvi5OvzY9b1vazWE/h6wjsF3gvRNXmvclMOylzmSpE3
PkKJCeLLL9fATERpjpHq6vtnDUFHhmzSldDx/zMa2xS0kqyBc8TMCv+E0DL05Q11i5FxHgFGvIDZ
cZ0qN656NsnlH7nHtmBrTiY4pEy2Qv3RMfdM0EnsmRq+cXn4vwreNMOepLVQUCnGAFZtOu79xGda
j9yWPn9ovNMrgGDLgS8qvJviHlp5Q7wAzPPSjS0ppscosd2u7SGY+V7JsKGS54hr5nByK2MgbJd2
ce5pLDnSdfswrTFaT0gM/EBoaWmahTO8r3lK6WGurlclTpHu598JrtZAFkSp8NE1N2+2iW1jI9sm
Y4f1RhSdnQq/MpB9JQ3W9rTGIpVbqulc7GHK/MDGeqW7KuggaHSVOaheaS8RTmTK6fCjiHI4I0VI
qA2eUm9pk0qleGSH/l+YeNtDCNR9GiFCYQfHP515cVHXiONH1kiHGYtmi5ef8w8jXW6LXdZqXdBw
iRY6NMbNSsl8/B5875AykOCSECCHjy7bLoY7kiSWGj8pO/cSCZFSWShQzXFiUcytkDCDQlOm4PyD
B2Nn2xv5RCeSaVAQI/Smsho6EqZkGY9KJ9RsZyRkhJwnvBzxbga8zLIiE9CjAK/oBLdGEBKalYHJ
2DqI9dZZ5CxqBajpwIqOyUy0/RsABq9k0l8s15/PSDjQT36XQ01A9KGMpSdzqlawVNB8ce42mGTF
o/1uLpE9IV6vpQHZNp2beM8mG9Htmpcyc7/MoBpTtDzW+Sa99ZGEmUGxze3+YBfxcTTTnFrey19L
s9fRyAZJEbryTFTwq2jZku37P1KqSWtn+m82jV5hHntugMvjS4W31rxZbzrkzcFQ+SZGV7OH737l
RZ5x7moIpgmAwE6vhizDElNE6ZaVX3D3NBcpvKHyxURSRqfm0ZlRg+821Ir/+Z6LizBX8d++f9lF
w7/rFdc2rxsgPkm5GmdApeXYn4NsP7O7Y8GjfZapvhgghIPYf2/GyGb0P8IAscSvtTx2YBt10Cmf
281H1qEdUx1YIaSJPFQ8ScqNv/kPrx1MA2eQ32//pOFtKaiEoQ6M7kuuo7bMv8m4YLHGm8IMcq0T
ybKQcK4d9HD8fowCYt4Jv8/kNfPVAHYysGGXcJ7wKtxxXZ4LFph2hrFKxJEhshP/NhSaMO5/gwNu
jUp6eGLqy2N7Jq8MQ4dSFhuEcdWJWnUZqMrLzm5kLEUHfUouay6U8KLvhWczpUP6uEtr4gyBmlem
JYQR1GNtJWq8Uk99G/VC9xsjUOSPxHnEoX8m+tigTUvLVFjPKan5YiwHu9+pGEBoRhYLbJRvTRsO
+IGQSPy5hchknS8L9xGO2maKAzE3wZ9oiinabwFp+cDY/Gs08rals8oU8uQJWrJ9ijafY+tJS3Ld
tOZK8ER35KXQWMbM2n1/5vLuzB+JYMgT/aAySOXS38vKnVni6G+MRS2NMoi/Vf8OtR8FiougpkSX
oSX9nLQG14Zb1d1yrwu3mtePo/upTA1x278SRXHsOxveZeM4XC1lzL+wvwCoy3+rHPyAm1PGKRCN
yBT+ZruvFzBNortCefLnhPF9+CnykRtUiYun8HNs4DTtLsJUzZN2W25nfkyGoXTQrTaCzt8dH9hP
CJWJdk2TXzfNmwg1hWri8ZepPeHKpVO9TsFPf1njKQv49vrGnT1zrLHL1AME1UCgijZdqHSbJpzc
L1oOhiI+cwuezRShqgnlAhT3EO+VR8Ii0cOKZpM87r/s1EVczI4Jh+HPn6FPrwnCCfdRotf7Vxng
d0UBcutsfS2F5ssvWQFVTuJUcXT0iwr92OWJGglhQLGHljU8PaOrhibpJ0Xwe4szO2Tm9Tmu2IWl
Oh7Vn8vM2BM9zT/JgEqtGdvNgYa6xNd0bQb8wNRgXGeM7g1c4x8LwoTGRY1XFjVB1brJXPRcqU4m
TixEyENWzPYLlzFtSA1unPKS1PDLxs66wdyKbUrvNtr031xZWkruUQsgyweWN57ukuUgo7bdYFfm
AERSD2a+ix1WuxGMzOA88N/IpbTOovGDukTnwZ+dB3mIjYWntVgCzS1DnzAP/QQIp6GTu63b3dq8
XXXCdh53DHNUMUHSa0aaaMtoqGCAL6QQz/svXi2IjlNLifo3sixQAoYCM8JYwuCom/t6ONSuXPkq
GRR0aZ4N+4UxWQFcoBbhbVq8rOUhJCt/OQqZU+SehoYNK/q5kj16dtXWb3ELhoNUYddMgWJaAl29
sILgA2FtzjdmWbWOxkVd+0vVglJCYP35Ba5a5jO1behY1lUT88NechqBbHlifFNmm0OThrvxvWzX
LczHUEOmIqgPoeFuFawg9+2QKqfWh08pUcXPnJ0fNgIc6W1YIIM3maZIJV0G9IOn+Lzyr0t/GSka
5dJHqu4qj4r7EBXJPS3ewS/J7g6MBkyPh3jgGbqOuoxxwj5ii4y7/KRxdG4u3BoYfGSR+lS9Revl
TSOYFTohfgchNcf7wUYncZSOC0rqaiXr21b5xg9umCWCSPun+1QCbCivL3N9QhZQ1S6h6IMabrJh
0FoGnqQchFikOzaGO9my7cQPnWjc+vtkaBaeH6raRe35Ckxkn/VzGNbm1uhP+gBDTedi09Y2CJFc
qLdG7l/V9TUmP59D60rrcZLsULORhiK6yVKu+AHCZzjc6KN9/saNB3kB3rlNXdszWvswMO3i6kN5
Bn14yg198hpq9s3W7UoAF4Apcamg0rOKNjvlkG/Rz1OjA7hhPqlVlKan/RSnm7kXKITegDmQqvTL
IF1Ilu0Sxzs4t4VLTQ2TDW+mH2rTLuvwAtJ7G4fcPX88KrKlCxmVyAm8x2W3mrUDnmiyVXlY+qJu
On/+SSb6EYMZ4wRf3Si3RwYCV6W/Ei8RS48O/GJ02zmbjJiWIw7pxcgdjYVC8gbRTXvobNMqhox6
RMooigbo0zP3ZII343sHGAPz+n0Nie4v3HfQujtJBUhpTYV9nBCEI4RH4kDNhr5P5+N0T7HSgapL
EFrlTn3g9LKj5K6IZ32fsYzkCmqCw9zAQ8B6ZvU8gr6cZJo52cslJR0SsKFWQaAIm7IHbmh1/Spu
fKeiCWu3rgyD1ckpFD4RFeJasDZn7dwiJlAZyeFK0GV6UtToN6KuKq7Hulq18VSdUwi/00ppuPEF
I47NjfELt+q4rVIR01NHvDszCbPad6skcfkIKyxQlOmWMYQimu8Vw9R7C3BkbUjLEoM/S2Mg38gZ
vvWpWmw5mN4C8XUN26rOb46PAdjYP5rU+WGTwBLoOkRIA7eYbIL7sR4SNKRgWRx85OCUMKiCB2Vr
PI8LN+xEmCGE6UqNzxMCle2il6FDp21ngvkNAAjIT0OIscs7uo7/Ih0sF6NGGjLDAY4U8RVhuq+i
Nu2aoNw3F0hLqC9oVCYSUQSyvOtA7gXkcZM5a+TdhP1RKEn2erROxIPZO8TfBUENxc1hbtFabawS
6vASFFjmydj0dlq1RxZh6SQ8q9hzfFpW/zqltRhAjH0vZ/vEjHgyFBCzZqg2AYnpz/Cugx3vrVjM
rbOZMxvdcEhyj8GwBT89F+61ZHKgnF3XKBxeqgoKwfek/Y4OjZzJ54nFczRLRGa7/KrQ0tf1naeo
KmziM6/S+mGF/7ryuMCS+NPtBNJd2oJzDG0vDbaBcjPYV72A7D+Sqhd6SqFqzsZdMTUC4Ld0VbGv
KmnxhE0TW998XwmAlYXqdiOY7wsGiokVXwX0uddaN3MqFq5pSXpnOWLNlTBo0tHAqBuNGPCkE1ED
ngldMOYyDTmMyzLW+UAZx2nBQ211pKLf5baWwEWnmrh8FEtlkrNMYOnnUsnREbS2OC82EO6YztdZ
qo4EePP0B2uP77Pcjh17bj7A2HiSSV1l7SUuXVJQ4lYEOXMvORQdBVw85QXRWIbdbzHqEGtCNWW4
D6MSldg+/vrUmSY0CpXR4koDZ2WD50EWJuYnBw5Ae3nujuh+LRUrojHtzCyT6DNWkPd7UaSWlFx4
/8kSasIqOzROGNCcUaXNzqjD1/4fFnp0P7gpOnqXyGvi/+UJn4iM7hazWsrbLVYQKvCV3zPZgylB
smMBIIwutQqLO8lgpCxMXBUlp2RKYkt30xhdVSgouZ6M0qBEj0LP+oWw//WDBsKyzMfFIVNj9rCk
qoCacsEuj5YLjt8LbokDIiPqBYZrgEmJGNWTuGkM8njt3Fl4kFjDRkLcSQXKQmcgTcV5rZjxJikw
UWCKfk7Q0KbcotxxgnKdtR1s33WsgMW06esxV08ZYuRBB3psRlXwF+cXrKiSLfUOp6sU92LdfvQT
8Sdy6NBZFRxUQvOvCcN/7zfetPkxgBY16qWBscuPS/v2DRtEQmk3Rq/DBKTEuTTNgPBdAnOVy87Z
U1qTLx/lyoKS/IVYZnmEHneBFIvveFMAcvOqTs3ss8IajhbZRgtKhXxksz6hw+TGtL4iuP19OsUl
dgj0dbk/z/MWXuUDPavSAQEM2sQwADQgBwIzs7678ua1l7YK26y1B+SY2dUMyISHnuerDhsqOjBb
QSYoIGkL+BxNyfyr05BOXNjIZ99172JkJP6jlDMc8IUZ3STUkpvArjTR+6O8+sFqW72F0O38knzz
nY+EElRbzj5X7ONgktAULxFmFlcDJchVVGgeOGz3I8NjVZvKBZmdIyH+ZrUqPT1luer1pZFhWFG0
TBCD3QkVfhnDKdG4UFR467uY8IDUvHR8LpYGsBTmCr+vk2wYDA8pCawFGCBfK63ZpnAagK+I+Z57
saQWYW+lKrdEcqLvrqQ8NJmn6Zl1zjWcNNi3QSibUK1sbQVck3wFVQxtAVY3zm7XV/lJ66h6RmdY
z7YQqnFODRNeGhj5mBqL+gVPE/cR4cwnQEHmYZomp1rMCb2AMtgf0GA94DWV00O1dJQnMTPErzYC
FMBt1bsIoNaJ2DdG/XHIL8PA82ANGA1KWChAW3GE1y0sSbvlxpX/BIjS7fDc/seDAkmxGlx1qdEF
GnOXatKnZW/5Q49vUBl+mLviY7/aSTjmniHpW1G95eZJFI4Y9SHhFsXdfmY7alb3U+dM0/H8T1UO
SsvZxfh9APjwJVbYJ3LERwRpeqn0F0Qm1CpmasnSkyauf5i4iOiDx7sBsHj/4S3Svh4RAYR0/y+6
IjJWJUIKlZa2TvxhREbok1ZR5g7aL30usnMJpCVsyseOyvS2zRZbd9WyJbhn/2mIxMjp+27yBrdf
RBJnyVrvb293uVMRCHt6ane0xkEkcYDC29HU7bpcnzXlB9MpR2twUl0UXN2rm4GKRyr+2JOU0i/N
MfMQkAze/wBvb/7T2jM/9tL/wAkqEtIgn/H8V3iU/AUsIq4Sw5spFQ8JBIvUaAHIhxUYNIw844zL
6OLJbSwjLFM4wzIoYLoxxmewAEQdh4R6wGbEwWJ6nKoXZjC9sfXxMEuU6dhQuFQWUzAQOTCYBM8Z
GS2pBeIQX1L5Kp6oad2S7ZiHXOReVSzCqnXSEIyKEHaELQSaxsGIx3hNMQYYLYhxIDDYqUVLSxUM
U5WAI5ysEV3xNEzH5aAzA6uP04gWqzLAlOBjEXOf89AWqbKfmDzOrpfIHY+XSXxluiY1EJIqY3hf
k4GQUAu80Vg2nhp/FInHC0KTLeEzPPdklUlFy6lWL+ilvIbtxN88+ucrA4tk4aq7tYHuZIoI/97e
c02dR+HRcTnuEcR6sDqPJUQu5L5th837jT7rMux6Nm387WGNSRe7xXSzCnWjyHd/niRTrtT9UKVh
oyFIgunWkhO2+JSXtajTdU2NCRVHFbuIn+aFjbHc1e29EoKiotoaNr9M6nRkSppRWqzufyt6Q4ju
LNGO3tgHsvxj/+gGdrodu3EaCIyWWJquV9xFaa9zGCgVLPfjfM8VGfSG3NhXzg4juunNZ/zyeyqc
8fvF1g6yLfOJ5Ny6XZFIiWH5+a9AlUTphH2o7bZZnPci0KUAKyq3qys2lnsfn8bBTMbBQCxVI2Vk
8X2ZtZ+c1U6lUedk/7xK2SDfkP27t3Oz4ZFJX4LF3vcZTCA90Y0FLwaf1+Cp4H/xYkzlUTXxM+5y
NyE7VfJ/goMMWcjDJPxDRltWfePyf+06cmJcRenLJu/RsgJ09tyYseiP9Wxkz8Fm/z/8DwJGGFXi
hw36ycWHji3ZQTvE+B77Kl+1tRhyBFB4je1ReQ+8pkToZOEaFiqK+jt04h+21LHdNZt4MpMqrWSI
jcVMAK4jhJcLUL4TIw8cQLl/kx547xYlpCGgUOy/kI6d68ICtww+MVwN+PEPe0zVwSMd12beKYc0
Dr9ZYZWufefMhpOwc4uXHO/RwfW37Nxms0EPuRw55BFiiLef8+kVFQsFg1HFnA0z+OvnB7WMg00u
HgMEUqMhs7SfiH6L8F9T48C1odimNL8zQ2mXpVRRqTxEeWmDFn+4GUOGhnlJmZOqpWvYwaNnF5/P
XDLMBMPA+CN+hkgFwJVdu4I16yUWJXHP0pJHVqY87uqvyuaMpmU6zMXWEa2ufe7XbewrM1y+2+/R
rBmOBz+dQeFVPxVzKsRQmOKrbKbjmXGuZ2GTkJ/bTFvN8MfKcLtbldKkdCXJEL5VtHU22q9hTdwB
3VHBHnFMezfP9y5MlhXj4Qh5i86/7I3v6kuqprEOdcl3BeJgylluwFkD8Pu2gTyUk5uECi9bRkGE
6pSBWvVp2T/xyo5+5zaFOoqSl2kt/VBUF9u/rg5gB5NHh+PSSGl+IXQ7knKUoR1IJEG85OG9IFB3
dVaC7MVdqwuS7NAIMiyZE6ZYU64l6jdWsBhMWQsh21ZYJ8T+0YRnXX9JdSsXkililmCh0xyyoMra
vIX2nXr6pLxiFO4UrsKOl6Y5DPrVpC43hRrxn9zC8I09RWNPi/B9wrrOizdaWDCZFTtkF7LJ4dzq
m+ONah/PbtEPIka2hCZnH/kpXsBewP8TbgVuVFlqsy6FRgwFN3KUzBobNPOq1dApgGGxc02VQen2
/PKrc38FSlEIWzec0yAu/Jbx6eALaaIeZaWkbYsgSLnDy+yLzZ+qC+5Qllmtax7zKWJydCucJ/nB
Lg+LsikgOWpcsxPvLBYFw+Ev4xAlDHHbAlrsG79JwTtQSia4kLIwkCw2r+Ncfte3PHr+KOuHF59N
IcuXQGnmxlyUEteI4xgqHCXlOdox2kbm3SSzdxsANmLWW4kgQPzpuxXYzeYRp3DDhWxfN+Pngh7u
amaUiEs3M/jIJ18eAxA9rnUJ3VtAgFCZ558zhXUobwdbDwE5yP3aaPnpX7bwVSx8wKIehORGgMLK
YFWl7mQ2amZNHrkcYoYq91Y2bCzOJkKCAlfQuRMGRnlLaIK+CIGx5WwzJndSMAaJqoockf4cVJTE
orMDGe8id6ORBLgK9SLmHrNT5C2RmpFJdZ4UvKfZtAZNBn0CcGZuVyOgiX5yrt966qTrCONEGZa5
RuDF60IjAXjyGlJTI1P2lfyCGlu0RCw4D5QkV9+E0PyOaNPE/dqxrUGR/mt6N2tn/KrLXkd1wc7Y
aWcFSD33SZ3XFYvyM4J6GC1MJck8JshXHGbZaNkK4XyO+2jpfG5x1qlAiDl9FymH3PKzcmhHbtnw
Eqqj3tXyj6vZ6b0PqkGxJDJGI7IxajyHhZR3kFEihz6TZtreR4p0Jwo6uJ9ApUrRMjgjbZ4zA/ut
iulQhgcc1mRUk7Anyz2fT1CYWfZ3w1siBB0/mv3XsYg+tha6XJqjEhq+sfurb2jvhUiojuxuu39T
mGfB/YgyoJkQrC/KaqKDkNmELaBqDsHGUYvoOqS3t+WY/93ys2PiE6vowp7gPQEXe4u9874OuL5F
ZDs1/l1fXO0DSHlS2N1EXacJTTnq4TdAJYQwsBGilwQ3aVqmjHzXOLy20q/X2z7tCk1wp9yXS+JX
U6V9WEueDwP4oPVZnIpbXbDNdYTzd6k4UpcqiaC9SUNamL7BbSruomcdZOQzpZcLvERcg+GTtph8
rCtj9CaRh+8hJgSYz8UVoRW+BGwRislo5MMbr3imx3ul7d+z/i0i9zCfRW/UO/P5cP80HDSPb4Kv
9eYqxQsvYFOM1MPOMfO86AqEJcjvIsVGn0aajYZus3TSp/iUiDxLg77S4L315CoLVtKOw0mLu0dZ
62aZqiFsWFrf+TXZrF3hHaFBqVL2wGmhOWu5hGlWZH7L316GCGe9x/c+on/oZKWqEen341B3eb2V
gqfoEte1IJAZrd2uKrMjYu0qPhOoNcyLjkB7BQTDyZCTdxDLuhn62hjz4xVbuyiZsJ/+Q5UhjpXi
AFfVK3Da7M8M9aWi7AMAuYgt+FfD8bqyYtFKIUXJ+beBzBekIJ/DsfMGPPMXhX8lyOyb+q+7IQSm
y2mk8C4oL0j18wn544aJbVjwX2gYQH1vpzn7eVwI+1a6UwWiWS/aTZ2HfcHQi8knx5rjhrD9R96x
I3cODglht0S6Ncma9tUTXIkizh58TfgAcja1iC5uMOo2iIatFwG0ZsAGw46QGso5pmt/YCsaY9X8
hShRDGy0jC54wFYkJ+KB/Db1aIWjnPb584WKJ+BHoChXMM3ljgHKrape4T5Y8DJK+7oEpcWXr/mE
b20F0lbP/oxGvu2fY17yKHlot5p3ak+ga+UGK61xPp8B6Dagh+PIE4HKxK8lX8KaYLWcZT3Ft3wg
jRTCSNk6iRpRIu5xjDpoF2BO3eYz1cjMv6EPJc5ybKlWx/Ph+eKXF7qrWV3uPPUAQ3zTpr0akwAI
hNafunlezEcjm5CP9FWJi7zZeQ2Jh+zNGwB4IDd0Sea0LUQ3CGb6pU4RA47LBLNJshgvEFUE5KgI
IImHxEoARK1u4oaNSV6k/fVy0JyJTcV9UgR7gNxpsYqd2rECEnk2r48Suqlod4YpWfp7gVNNPA7b
TvwB7d6lQVWd7eEpc2Kv5wpq1hxpcNGOk1ySPpg5WAxT2g8pNBSfFlNXk4u5wLzSfPKxkqKaSTEL
t14i5acPfwjE4cDcddMbR2+mFZFH5pckuqHokAnpLx2suA3BniyAzBwqMtj4Urpfj7CV1x6Gu/b8
Uu2JB2P0wX2WXbSZ8Ro0xnkU1xsMxVPI3eeBlvhTbOw8lR4tnokFcOsFvdXHHHjnQxAT435nC39I
4/FExw5nfnvIw0iQKEqSOz7ViIZJLote9oWmaono2ushCHZZfQ+jT0h/UadVFctnfS9cv0H8ltto
fASukRJr8cQKDajwWA3fonOGYgD5uqiQbSXN1tWNbmjveqfJoSdrXqUm90st0XESmmhTyHV02oGs
lLVqp/dJEUF8dtYcN+osiwwtV9atXB6GC4P4tO5UXgeQdwD1srLYVM7SlAhIVCvYrjsq6coTS3HT
eD1VfE+Nbrb+51pyrSTWxOd305F7g+jegiChJenc91Xnje7V6Re/JbvvGqvxw1vvla2g4O1mer8O
66HZukO9OgrV5yUT3U2vgpdtbSGAWqAYcaC3EOr5hJEb84gQKq9TS+1dWbci5pErLbSyApihAW+s
0ji3mNir5nCuU56/LHdnSRhmvqSiTj0v4BWm0O4GxFFZWYZkjEyCr/V3dgLvSWWG/k61ooeoCUoB
SDtXbpfEIvMNF5rYqMhvc0bOaPes5Npz3bNiKyfM/WqVZpllEUEWPiz4xHu/UnAzi00g/YztBlFU
RANya2DPnT+MsmgtZfeoiaaUyxZoqSEy3YUFPlo5nrcVVN0+7WpD1i46SBU0raXFoTA5yALqP5ah
T02CwdxZOXTqThtZXp0rmCTLlhSrrA2YJl/UKiAFHT5pSSdHq4Q7wBUpUYLrRLCDsOJEqcLzpmx+
ty5V768gIDXypu8kCIL0KzPFXMaeeWBY713bMcrGh0pW9Pa7+1kEzmBeiN+dvHuaiixKPBQad5rz
kqqcGy/AKoBty20u5fb2ZyedDHFFrKR9Wp/Sm2Yy2oTEMdl9nS0XTwH2lO5+s7akmVroJc9cBDyY
oCrLbkGdGFwVZXCHJLSTdwd1kQXzYq93QpP7JAqxNirsUdJ8/svEopevXg/zIA+PLaGyjMuNzMH3
yjYKojnb30yLjUf7F4k+JNlQNEHxCtOlwtnx17K6qJBrN6twuFfdylWzPMUHClcM2Tvgi7hOeoHd
spR9Q1clNzUJflyUxUCWhhMdNANN+gxuq5pNzTTEF/3WvONp54OL/IR7n3jCcL7tFBA2XXnLD4xI
2CEKfeiXRnI26L9ZaVXIJyVUYJDWC6WkLSLTpHu3qhqYvwdIttEGIMTLd6gfcIJ+QF2RNi0K6S7R
5v9Hg/tIaUedYWuIcVGGReHoEJaFpTbr+HBqQhVu9ojakhornRiqxBkunT9wuKJ9HlsqOuXrZAGx
jYyhEWiI9GMa7OKamHk84MPapv8y5bm3hSg8MYQNqG8WyR/w/mMGjEDCxibEa9/tizMkA7PTj4AE
xj897QX34YOprEhVPOuz1dZvgdr7nhQOSWl/TadyfNgVAo9jYwS1cWfKJKGqVy5XaDzJ7y1h1hTx
5CY/AbBCP7i/4Sglz+dCz1WU1rXSQipqMvDA5PjMtdYNc8n8kvJMgEg8J5ulbXm6Me02eVXxlJ9E
mQXNmn+IZyBSq8fpFOwM3HeJbJ4IPjGuxsI8pmRn21AT0EmzcHMFmPU4OQ0zTKjU2C/d06c7civA
KJUi8ommKF/+sKDI/qBx6OfdUvmoEQuTwxnxQ1p+94yys3IESuZLYhoO5hccZW3f8sF7c4Q6EVIT
JXJpyhXAQeGC1rJQSY0w/G9PPjqJgKKPJlFQ/7tQrxsIWOEU7CbnaIicGXHqnBQXNFaDW2ahqcC4
pnt7UdRpkEJqWetz4ESqbyINlhRySUvWIQg1rfpd+OvXneRUGzn7nMy3jV4p6OMqTT96JMqBhM/y
ZSekF0g7KEpEzWuShZCt1f5rAxX8EE+A0vR/M/Q8FOCkAZuMV+BBKOq1x0PfZVYwH1YWLb7vMTKV
pJvl7GPrRv6ul07i1ck9tA+17KozWwalnb6B5fkjLP9Cfb/0MjmV1uN9w6vypz/m8fESYVOWbqVx
AdQetwepaNaDula/r2IRfkz3mgr66zkvk11exaJUSeew1fXk9uCg0Qqrj4FhDGxJeKeBIBaw/nJz
tLgHVD0HbYeXQ4iK9d3CVCA1O5nwuO8H6K+8tSHtCl4o1nbFlCuzsEXQsc3p7D4iI7BISlf8vOFJ
uQc4/wI8CXgnf/bBFZM33Avi7Iaw0/aZbC5FECNh2aLeUDPhSaC23eO64Q63NCG1OcREYG2fvrNZ
QDRmEx8XNIS2VKxz49659nANYuyHXsbjXNT3enC6pq2W+miP2goTy4sWP4Go01kwqF2WgcpIEzbT
g+jfuNDy02mMJhmm34Cxz/g3Hkt7C/F4BF2GS/idQqxOOSYcI51PnND0RgjUD9Tiy6a7VegHIGdH
5ig8i/hlqoYa+9DGlsTH+lC4iMYgXfas/X3ewpP9l/vNUL7qvw0Xgk9MGA8M0ui7bp29M6cj7p9a
KBpfZPSetw6HJS3PenXlE/tcgJn8U2JQUiMhBLGTzEWmTzWbJtWJSPttwJAFj69xJ7A7LEmg/IHp
xhtGN4O//pxM+Y6uEHYVY83or6PSKDhgyF0tUCyGvGFVGFyzFp2TmSKIWPYnuA3MlHCW8ZtH/Gu2
dsjGubyGBmjkwxYlSECvLXf2SB6v9O7VgzlDq/pTfm7b6pisuR5YZnaCzKhlnTkWvTxw8uqgNuhx
AM7nIf6Gmy35HZXWC7Xf3XgwmZU3dg/0b92Fsx5tUaLFPIsN4nl99tblFDGWGMQ1l0SQQdBuJjZt
is8HeD3CW92/cBPbPmx9xqMRr0dbmVi47lMmClRS4vGCLfh/UWzNShaUxjBt4TARs/T65r280Zf1
mn978CuNPsIKW2YG1IG4N7fnaA7OdAtSYVzN7yc3kWDqtYipkKeN8UmAs6pVwZJRuP2YXDd7aS+b
j2cEoq0ima6PxJ6Fme8tobP26FXk92/68VGOPuD87gH9Eb52NdNboZH9Vxgrg5RwX7qDffEflWdN
LqytxvWfRBed3rRQ1RfCoiuEQWR8f6GVGiOBXuu1lTJ+eEGJxphJ4zhZzfpyHVICgrljfoa68BqW
0kopp4barhA8r0InWG+1D7ftuzgNoDWffIftxNANxYTca66GhwH12nGQ2hyWCRehZOcdbS2KbFPh
XeAwMcdTn1ems6ODugoAjgBnRtZmk8qcCR8YliZVsVNz1vzSkzT0x7mTElAuL9jno1zAJU/5Xzb0
wIwK5eoMgl8kejEAkvnoRmZSmsQi0FI/ebhO0w1HuDX2B+hg57kS1smONrlOeZzDfKMCqmGial69
RtX0OXuZkP+G3OuzxoyPbyqmbIFXQT8YFw/7oX/YwfJxS5HIF51v5Odqvij6XG+I4n6di5AjFY9W
taZE9Jz36cXBXe/zDPcDiMrDMs/IVc4K7iFuVgZwE3Qr2ghs8ux2xM0ZdZwSzaDhmepxs1fatFCu
bBH+LI05j4kzt+hk7RtM8HlKJFtBtDQyclY64Et0YjBdggVVW1ucsTQk+DizNDlMVoC/HPAMMDPf
U5PM0+qDENObtA+r/vZxA2v8pSxEr0Ax2Q6/vyY5BI2NtVA9JLjY3NsPems4swqVhMt0V7BZk5P3
FCcpdBTxAzm0nJ3ilZz7aDOjFn1zDS6cGGqbrzASI6mWqdCRh7B7lDvuX7WKBN3W8+7Nl3D/zBUO
D28NcwnJRumNFXI2wek8zDhQjz+/8N6hBPVWHZQRXFOa0gl4vHgRcwH1l0diib9i2LJvf0O268/6
K1btJQ0CRpkhezSMTtwYFixmJGc93iJcUTM9iL9lcO/k+yoKyTClBuQowmZm40CBY66FgAgLQ2vV
qguZzAXwuzibKOLpCyJjgT6YsFnKEaEpXolnJJKEwE7b9iJRepWbiwaZRscid8SPVbVRoA2S778C
dZeDex7FmFNSeiJSgj3XoWDM68stVL7bsNJjg2vY7f0RPQgZanfDmGc5q7az106Fz0G6aRwmeK5c
utRAzZE3/7tdITBr/UFxl8wIeIXc/i45tok+Zd6LBUyZmwrj6JAwGL7CMk6shJ5uiBqaeb8WArwA
61mqCF1InrXdWmnJIA2A158gpqw4iiiFpEsMem7erS16J20prltVINtYWCH41yvWOfxJkvBDo40B
BuJc9sGS4YsmQc1OUquMYrV06X6iUKQNo2DBvCAr+X/4u3bySt1yym5l9zhDxmNlwW1JXTSfnq+B
5Zr+/NP3McfMs3APFbDi3mZzALq1dFtVXoWINWRp8PwItcMZwFK5W8Fya83vM/bAuxcWhDY0jUUK
Creseip0IqCPwcRQRXFxwb9oaP8wELxiEAr7ygLJIkLASfGRJtxm8dog4yshO8Pl8DDmD/EVDX/i
loKDTkeCUrA5jRhvlJBoG0/Z9z/BRrcnKgHTQ9IA0FN+yW+nYY8syXB4yUaRXO3Y8fXw3Rg6aEKe
PhlYzu05CnGn6i4VZWclnGP1tKb+QcKWAEqE6VNCsGt2lUfp4yhJ6JTBRzxhJNrOiUA7GQ8Yh97L
MVZTtdCmTvxdNJv/XRA+AS34Pasg8WOJzk+zxVvAtOSTa7p+cwOOIceHp5AiAeHUN8GJxCwGj/8P
0hCTwc6Eilg5oCs8OwgW2hRMzKnUNPfMxVuXcS/MGg1Z3Dhc67i56iMHJAgb/A14fRN1Mk746a2W
FDr18FKNT9+DRPsMFvjIIXSx87m7ZlL/YX6If/bNA+3WB1In5pRjpxHAlh1JrnA5Ba2OQF2VySL2
48N3Z/2NhIQRpzIfOdnLwNwKZrcvCw1Cl/s2yOBFx6+W74mCFStbXJj14H6c1c2bALujV7os7PPf
fkfbKm7IaqMtchYOMxIb2sft9FXm4jW9ROQCyl0newVz/22600KvCtqnoSejJBIQ1+oGfc4f7kRL
2soTeU2jxjtnxG0Waxu21ZecW1/HyAYmWStINtNQzQkhihl1ytxYIOsY+gaup2drx67LhqLS0xAm
uHH09r8axwY2HgprW28L+utuPjhNQWWRt8Y1RTVCKRTwwlk6OwPJg8HNF78V05TNmtdXSWO/+XrH
6xLS+88nTq8IRm5KToLeceQQyT0/KY7A6z6oyVTBS4J+JBkHFb3rm43Pap7MsCwBsbNNVXT/5d+Z
LtTC37W1iAKsp7VRgVWZujk0LXRAGYOWadjl8qQuRS8sc19g2u/wExdr9o0jwqoL7+AP5HZwsmIN
yNmBPbYq86BSwfgwfDGl0ZXhMeiizOHAbbbgHAtTDgFA5QcX1JpMHh7wa/R/ojEVNteb/6OoTowM
3/E43wWdOz3pybMszrBZA+SGkQtxAn0WVMF9D6ZSxVBeq0LDSx2Pz/r1WEnhHFZKN01EjXLkcYdC
jvPme8tYGEpNvyW3dBU3qEYZVEqV69hVdWXOyCQgyu0G/LeA1b3bEPm65hMquGdiV+5mZrm6eEwB
T7GQFNc9+U5f/6VAizo/0r4zCvMRVr+RW0q4Wtow7RfybK+x8PYylnMqen6pqiwnrNK2wRnKWaHs
pUCfFapSuWdb3bkAlgPOC5sZXFjyeStiHZTP5KECjUolrM5p/qCKVkxWZ7EfMAZmK+hBOUZYIHIV
2hYY7tHnNb0Zznv6/xPWHM+JbCHyn+t34UWXUOg+u/sc6TNkFeLH5G2FXSSuHotjtL2erKaJ8Zd9
3AvnYp+S16lAGqDAY1YxgAxRGjaOrchB1FymQY0tWs/iqKP9CJVnWlnhcYTadlEegfr+y7UtIsRE
qYwYX9cGVmKbczp1njRGSsjwNeMbJROAiWuk3TpWJ/8dj/U7zmkRxQK+ZbHPni7h29SQDCV1EBmw
6N+47GceyzFWuwgkk6W7rtsTs6/Ed1lCVvEd3LV6pluu/W6SHfpINlVxaJHL9S9KUWYqcxycgz51
dLjpPerCWIgCKuV6MU7mEA+y0SmsT2rK6nELW428ifNZIiQkjMYoZ8zk/DWwO734DFGyvc6sdXWn
dx1zhzEe5dv2eup1gpj6oyP+tQ4Gy5tM6zhmZB0ORfu5UOJPU2g3d1n5qkgfaAkLiTmB/AHMpiej
odDRL5lEpRSJH4v/VNLneidQodn4XkHN8z0keyS1Ua9/4l3l2Kn/yzPRaRQZBU4JmSAhzG4ghb+y
pq0DPjxv6mhyZ/4a234I9DygGea0ZaOc928x7hGBhZZO19rxoBest2E2H0G+6DPAy3+f3c275mik
IPkvmfzPuLAlYRY0ZlECgn6X2cUyBYkUYDNwwyHgdngyeoSJ500iPW2l+G2LpsWj4CAJPMOi982d
vgsa86MFv+03IEhbEGdv9pgL2mxPWGby5YEDyH9JgajQLmgraswbkBXB6JEib0PNW9J3ruMuHYe+
7lSM71MuGgyO5+7cLoXB1VjnF+OKdTYQr8v6S5/YMpqx0Kaa1+2e8BDwYRLKfY4+yUlcPFI2BD3+
ztgac/vAzUBzO2fXiJ0Q5EpUIhLmeZ/NYOu92AQENbdlZEYHjChV3T4EvYT5+TP3ZDys6NFBUkdF
QbUAGDVtFLJ1OrlEIer29vZwP3WSTqlp6j9PoPtMwdY9+M56z9KOEzmwvayrim2Bjbnta9jvOJ9O
F5Eu9jEFgAlhMmW4KOwyBw+YaU8dnnXLvUZ3lsnEDS+7smsU8CvaGO593F1Sfz8gAZeK602ejpV8
LMY6j5ZLtG7xVqptCRdgrneSnBew9Zl82wS2zVjqxnZU7peVdrIKMezJB7BYeU0ccYAI2PHq+1PP
I322HVaEdkmqU2AhDJdqsAjI4NDTXUMGHiuX8f/JzDjflWE4LL1hdiXgNQeIOHhry49qgmy76B7m
yw8QvAQXj7CQqOVjWrlv1SsM4mXthF+puaYHc/P8/r2SCv94dTQyLLTtRfcC02uO4bwAbf3GOlg9
MANMFEcHtIo4AgcFswXdiMYrdV64P9Le6X1wILzKx2JmzJrLESr0oPHANf2KS7ztpdtVOPezeFKw
Mwt86BcYe/9SgSMGDSEuCLxZiCJ94xik3UrtaM+37zRaPVvESsQ7iKgx5pduv24Wy2pfAYLIWb3D
yGTv3Gymww+o6cJJIwmYpnCkphepxzbkiWqIicoPGq5unY/UPgP3Y2fRXBfzHMkla5DQTl88R42M
7BijA968mRPRwfdtuQI4y6K1Pva40jMyfDPpJIehI1t7ibF+uzAj0sJZTUmQPCYoAOK5f+mqTHNP
r+cv5a5WSbKDLjPSkOSghgpbScBg7LxVY3KAPFITvAZMcTYSz8JU4U02jCgLE7zUqSJgv7YOT0/b
n5nVM17jsExUH1/Cg6X8DN79WW+A9vRNmkzx+bb3hrs+vDTQfDYrWc3VAqTexfQ2OvZC2ilr57rX
hvPu/8l+waA6+4Jis0/o1khbE0IMxIcXUIHyYZ0S3yVh+MyBq53L9VpK13vRYlOhCxHzK7M6nfoN
gVkC4b7ac75R//hTbTzoLtOu6+wAl8YdE8S20hiC93VfBJssliRZVg7x6VEmCfTj5qGPqzdvFGx+
BH0nZ0rePOYThBANkrfyfOMyFpCWOwIgxkGxEoa9wTnKFxTAUkD00UMH5qS09n7YWlJ5OwJpRxAH
5hunzdJHV9RBbUHbEIHaIk4V0gQRQTM4wECC05NQj0DCGrJYv3gX/XXXjtgqsQejg/A6X76NfnN8
6fGYsc4mdO3E/LdcntZjCxZCSqeRHEX4vZ5Tm0iJLT3K23rb5HnMVcvBbno4E8yGnpJ1tJUCs95j
1trRfKSpyWYvMY3ET/eobx7TOwZHZcKXLgYRhEq27lz7ksSgz63vQ0TH1d963WCi9NB06QM3pbqe
1SFKP+R0E7Z74VE9viFsq/U++ywU2rp2EPBW/351wntzzg4TyIWfOWvByf4rrRSxYdMP8N5DfYrv
L+Ld57aU2Mx0xb4Asu+4php/Isl6WNzGAaQGq8XAF+dn2J4HkWmeWAlWodJtuSNN2BnjgEejM3tq
rfUiBcr8IHbeB8RWU5G5t1vAsx83lx/YpSNulspYobVvnoZH0CxcOuD7hXo0G9Pf3yR6CIeHWb/+
7n7ikix9SX/QOs7tyZfSTvhfNDhetzYdSTHXuQzuTtYdc/G+T7/OEg0dm3HFuR5SrFxkbIxihbb+
HWaTjmLq/OxIizc+mcmtLx/XYFt6v/nMvnCnuuV6k/Dgr9lSgPq5rK4OBc+d470mTRjhnZuxtsf8
1rLqOUyqdbEHFEF95YH/Xy6B4lPFjGZF0AM1Dvrvy1LTGuigYwqNBOYhY0M84W2chRoPfVJxLBoc
CDR15U1hMNDNgKnghg4WpZ0/4OJ4rel/tJl4oDhD7X928mCJuP2wfa5I2vrCZ4D2tJfkx8jGnGwP
53jENyB6kdJF4fi5FYIL6A71qiOJT7GwBt6NRrAU+rLiXxKFFfSZzZik+oRJHrYqUNecr/9FveAq
WnQ76gvjLtlw4JnLv0735GozIKKdFev4NWRrG2xB9dZOoQRaNQkK/5xFXrzZKr9eRzbQLfTQpsYt
Xoj7QJOYOsYeZouszVDHi7R5t8pmab7hpg+tx2ZdJwgkw5jR5eB5yPjLSX4siWXgPDMotw+CKCEy
u3u/uao3lU3TtslehurCWwsK2OqpSvjDTTtDiJZ5WVA9SnI5t7bWC3teaFwsdVO4ZrZpc3dCJD93
96xtXHRaxCt9DdQNxj5egRxSt8nKR/kGKdJwFxGLQa8KyIvjgdUChcRpHnMcPddFlPMFAm5ykwMz
3aCpCptsGRKxz3OzBGm4J0mu8k0yw4LcvQnCQLAcoGoRdqGR/JjKBv49fkIFOXn/XZkjjt4Pgx8+
bKsHiuyqC27dUakcYHna1DapurxB6y52TcsazgXYt5x0o999y+/XPMSNr2nSeZwcyGtiJVqAYEZu
K4aux5bBsohfAgoMWPWCTsqUDdt0jBGw5kWD+rpkHnyKWcm5wA17LcExnqIj89tVB7aHMGMNQkkn
PKltAnaBC5ugUx5BKgjPu+JoyR9+kec7hx20bwf6W4W0iHpVpjtNky8vOp08TsO6g+Gv6+i0CvL4
DmvfyNAMm7khV1KJz1kGkFNJmGGPu1ZnF26k58NREV91LKmy/SdQvfvGAnVFiFpPtSZlaq09cbQo
ioq6b5dReaOKQ0p3d6mHMufYh9O/XfTl++bfyfr6vkUxz3JA9rHldn4Y0naqYd80xfGBUW4l5mfY
/g4f9eIYUFdCntCOzCBHKHaPIJUKJEeJckizFqfLlnpM1ZDAR15FfYz4qz2OOLdxWMNmmGGRWfRx
eJjLrB6RLnv3l9i4XMeY0YZNC/QgldiJuHISSzVUb7lfTvq4ndOurhjhUDE06jO2S2kL5q4ah90a
v+d5bLjLtidXYUhogY5v76tpEyGhkdLcBhQLzL11u2c6hroHGvwW2uB2mfg9MYX1h4LNAeIwPpwI
/+HRKDzVugkKLkWKqQONOSFF7bns7HCYU8b2OjjiTm0UZraL1+YWq0Z7pHL8Hi4VDIIuDbLQn+AJ
CPWGSN3WsiRjAXoG86w0FMMTSW5pbdqtdZttG/ovsMnB2hTqUx5fuvcDmu1mdP61BFcZdf7kxxkr
KBuANBs4eY2zkr0Kpdkrg2six9KtMOYQq6DqZlUaTDSgHl/6DXfcuV07P4V/uL0hFIHZBf92Xb3v
8XDtdGRPhPFOlkjB3wFE/rRLu+pEm1RjYdtLsLsscxrON4u3bzAMnB9pg5AEBlj8IJf5pnNhfNlM
0G4vP/PdBFOgvwvqmggkEItgX3pl5VzTC69jArnpfKOVNiX9m0CzsnvMhcy71yGe2HYzKvXc+8X2
0tQNIqXzeiwQP8J8PTr2qA80n/9cicCDhTQkFPkC0r0CortUuqHxadI2FwQV7xcSh2R7IZW4bfQv
AdQVFjZDQBLUVp/q76iolDD9eHwd6VujsEG/bFihbPL8eDZIxWhfoqGx2DpJWMK7uDvM5aJasCMF
jUSXoLINdt1eDOSo1FWdmzPqsv/9oYkTKDi4gW2NcTh5whRX1YuJfXPQJFeUkelScQ9hrg16LkaS
M1cMMUCu6pug3At0kY4eO6hwG/DKMdvoHubGF60OOk33Tvjw07xNxHrb2bALHpvm0/VqvH9pTaV4
K1gjpzmaISdh0CkBE/NoWxDIeadN89c7+L9xc5Emep110Syump59Sai9uj9G4YDMM0YqpMpiplRL
YB0vQtPqMRRGbmdLOG1uu4vhCWiIoKL+B8fzM1LdBeJGNc8oQPS8IlD91Slk7JnBaMv37Ri3yN/q
8h53+22w06QBkiri2uT30ydX/xnHBiiT4nkmFkKd7/DfkjW0YEUaRePJewir05+A2y0VFLoILzJd
lNQVmhhnaK9Xre4JunJxI0kLXl7jK4W06lz3jq9K/+s4oGEAw5cRIZiOByjRQ8HUVb2e6qJI8CDC
Ln/bkt6IRhXC1BaL7v3Ty0jxXJ5k8texckBkgSqrzcEFjQ68teScvwB5s89iPQxj9t2D05B4lWYP
xe7nMS7I8tvEsUuyZyY9gSrj2L9dpNhuOaipq5zQMtxvoN703SIUYXAPI5vnx5D4Q4tT6RFpBowL
UoK/tKIxnlxOXFyww8YlPc1sVTGmJ0jHcZqvKmqOYBA2O6UdcWw9OkICkn1ZQJfdW0ga9jKboOBb
UboOcj7OC+T0W3UoWM2nUNmzPswWJQIqjuZfbB8Q5hYFPRRSwdjWbZKPT3r3Aneq9+mlL9vR7BVa
IlHSAA+WPNBiK8vQf73zL0YAdiQhH4vER1J6Nd7AXTmSI23AzGS1AJrl9rcNYEDjjtW4ZTfG83RY
bmXt4m5JdpcmUulvw8awIFLyPKlXgdz5kst2UmD/lNcr2WsoQ1LQ3E+MReFqYu9TCSbrKXaUvm4U
03KSL9dA0ly8cAS7icPtvnShpXhTp2OthD3HXdc8fDO6swvgn/4cbcWyb09gkGHs77dKFt/hekJS
FISN4jJKi8Xi1IvpQ4ajC7YjimRfxXtypC3cXCdv3msWTTlwpiCJPTLB4bVHwk3zzgRLCEqnRN0n
NgJ0GQ7FZO1n++JxdObYBNYnWCsEvvRFi19faFybs8e9V1WcOyhv918F26ohHKhbClzErO33vKK1
9dmvbVObJoi1sAulzporLSp8RVHey3GR63xWa9fJvqItdRc8L+m+GVhAEohhH2pUGjaORGFMhHJg
ks7omQGouYUN0E9Cz4C1+mNp4vyCyUQxIe4gr7HdEJzdGielw+T+3h+i8CU4giBuU2sZmBnNsLto
iIAdwVpb7NLXPztJnhLk5NDLxw0PV6jSpUVbjOJBJiIA8YusPlu5OoTTjA5Vc5R50ujBVLhkcAAT
gK/wVyFF4mhxsYk8WxM8TEngrryACq/WxXX2kXt0YT8D5LsCAOYv5wEvw66cftxFaAB9nx8f406+
5OoVKFSTRWtd5lvSXgyvvMbDfZatYPPPlzWz8wDAL/4/n926SU7A7ITXcB0nKg55dPYvVLN77srw
6XPIN4sZHu/d0U9xG4dYw41ktFcBHBxkpXYGMJDKifU7pQde5ooisrAWJe+xtfBeH4AoI5ab2OqD
s8TB2mxElDFFk1M5QBElErMFlN3kMlOG2fPXEc9BuXO0fvN0BuWlGYhTOGCTDb33xYY4HCl5Memt
/zqlFXxye28/rVrZtypnsWcCyqco7Z+eB5ClvHwntsL8VRfAxajHef9UWCcwM27ORW8rLNMbprv+
gSaMXc7cCouEZR765mAcc3x5dBmG2BBivto+9vay0Ga7y92rk78Sl4DBP+qzyWe1GZLo6IO0RAbq
W+AW/YX75qltxpG2qvf7r5YtZ8ADpRp6/Jk6a63C+EAn1mLUE888ckkclzQuWWJt7NloT2OE6rg+
hL04QQW52Yfq4Wseq7Bl/OFPsYcHMPDd1+WDDio8oFViWUoJEE05LdjShZ4uYHIvPloN+N782vbq
73zt2XfFf5Hm1th0VfgKZfkQbYhybYEYlACrQAtpEubjnnGMCSs0PCNLZEAurbU4FoJPwRrcrjpx
XXI1hyNfludr5YDipw1hgu90s3ndB5HMqWFoWCXqIqlqZ+C17F4RPJ3rvwhQgil2OEzMBtwhYlPP
Yj61qrFVytJNhIbdxFF65NLBTqvMWqnUlkirC6AGh0wIExJf2ZoUSedrtXjtJQDT+wRXc/rrTTdQ
y1SIMlL583LhmSar9oCNd/wzn+y9qa+ccFD5puykv9XJ3kmUTj+syLGlOrvvVdlJsC3whLFCQkLo
4CmMhAJFxU+wozL836obCBgYiCikgGyAzXo6LRaIiWRiUJF+hPEYhdgvWa5goC4ccMP+qVYKstVK
xM3Mtb0VB4yB4dQga5uZ7ABoRSgXHHfKCp+RJxAGP/IV1jSQ0gkwzULmJLt0HxNoqgmxI5vyT7Kk
Gfih9ARKgWx1PWppyg2UDzOTeJGb86AaIF5J5ihVyPnD5HHOOkDsZJt4ET8mbgquJrulH3fLxzB3
zwNma4RtwVqnTlVX9gLlbRIe6XtGcjhpFwhz5N69Cm9edGLmvkt/Vi5JX8WXL41GoOrMbqFkR2sJ
59uDGRZB85Yz/t7lkQC63+8SGvNEiG6Mfk1352Wx2hDqFwtvAuZQiU7YZ2tGFypENoagj3tC3r7Y
ViBCEf/XO/Hl3S3uOPMnBZUl8BkCcH/9zkZzr7o9jQkWoAKJYnyCWl0G2o7NgtbD71yMe+++vvay
u4gwO9AOqAqpM+XTpK10YF062XwJUurdR1OaYCREmYhBmTYkZA35UwskmSdaU4PYUvVgl/vWWY6+
9ki7L41J8qUPoV1mD2yCV6dxI1Pbiclu/Na7ai9Q2ENRRJxBAVI1qXh0VrXoWAvG/yECT5iY//ZB
9z5FN4Bxs9TKEJQvr5Fh++VODGXKCHmu4rcTmDMvd1mMirO545OaqYwZcUzIMuxVV7XTMJSmVquJ
Pu+LhQnlbHej+LfQ6WAe3vO70DRPYZuD/oKYBcnDuanlhINhIaWJTS+HtNcU7scS/xez2npeXrw+
RuC9njyCCj22xgsdZZtHWPFXAg6f6UHfnD+U+hflPzY7HfkJ1uXwSrgVGcxac6YoEkqNcZRgUcNj
bG7YXsAGzc3GOULwgFIHUKfhH3fpq5KDgyitv5HkmdsbayZIeCtqsVGzcwSbTamf8YiSv08hemBx
gy5BgUMeNI1XCcZpkp4zoHEHI7+03KHGuGqJLVxOivzc8TZj2Wb7RUrdjQZpQ3h/fInQVKQ21cYc
+EvfASHkFHJLiTJR8rIUz3Ind7dQZd8JJZMR1lOq82d5bhcBB85mvt1fp+rk9DcGHVd4Mkasrwfp
BZwqyiog6ockVU0okA1W7C/PkI/bYIdbzxHg+qLIocqtnuGV10EEKuT1i4AB31Pted3omjYa+gye
BScG5LaZoELGIAyUvLG+tIKtEoeHJ3Biuej4AstGpFZ+s2uCCEQ0LPo2GOd3o/qSj09PhPUl/vXE
k12MTj9v9otQA+vnFmIIPMUkQLVTmrrGkajDYguWTpT/wV7OWGhp7LOKO2YZU8e44l6NnCkwqTjg
jxp4MZEiEEM+lyqWSSd9/lbuPMU100zJT3JMv/+M3pvJoW0VznQ9GLzDjRsdJXyphxQk+aQXT65a
G69/bKbMd7EBuhJXkwt6uOywNcOcMXFYlVl97X2uMu62VfRPY4XXz8wBIIlwxib3i2q/YwBgOOPU
cC9zBP3E+78H0w3FYmG016UVipWuoFYThqIfW2IL+eQ5ESWYj6khbkGbTwtGFm25SLmfbeWlyvM0
NcY0KamC+4P97QYFh3jfiA0fR+hrooOXa8b/QhHLFOqk8+Sv9s6TpnL4+/rr2Gwuu8CXdQpMfO4D
Z0DhtYHtjm926LGbqNs2cNJexThuTSReOBlUxjyFifzIkaMvAlf2AYgpptRBPlIX+rQc4wX4PXkE
6je1lnCWmirdMVnmonMw/ez7XW2Tk4LDn2ugE9IDHF4bnjuuQ0m5qvRr1txoX6qcV9htKE1JK6bt
xEqIxEVHjuSF5fSSEanlW7d8Zt3J1mWKn0H2I2v5BKiJE7QRJr2ExsxkRqHxFwScpav4yqt6KA+S
vK7rbXI8ramFsdmdD8xv83T+CGwLkfaPlEbtJTQ4KbZ2rvruAmAJkjLE/J6/aFncP4oWh12/US6f
/fTTy7ESJAaygmHAvj2/A7ikHDip+lkdUTxxhJV1yPd/hibLxMQTeJL2wSFr1rk9/cdDs1vDlaAD
kPrW9dTM6QyqN+0OD+kTCm2lCx8WiRon24Srq+mL6VzDHGCMJ03JFZniGRuy1r4NRtyJQp6PV4/q
459Sg5c2FK2nqCfgesbHe+6ar30hlHa331L3SY4XWcMCEzWo7Iu/YmHBT0qOE41LyquqniCVvGOn
tuC/FSsWpd7qu17urbD3hBbXImduea2PrsZnMjWCWf1r+Hb0kA6SfOef8jh3s/ezLaANKaqUxoOG
XcRK0LNHR5nL23TNhVaYX/T8lxKRn0gf48yLQhZ2Ag5IZNQjpSa/+vYBhr9ZyZH0wW0TSk40B8ZV
xay2lsLti55vT3j+8fq5KIlj/wS80J5DDkuaObr01OiG/CmffWBM9ViRNLV3P4PwPXeSMDe9QgJl
/mRBv3XqM3qgR9ETmesz0GvuzNiGhbpRY+EfZ/KLlGql/Eho9sRihBh43/ifKsOZKmo6Ep3yeY9r
IMdEuiIvbq+2sDU66s5I+gGsfxkuxgLWuVyvZ6bSLjGwNyOVRsro1vpzHp3ovmkhAm1OzoX1FPMF
abltdWkTmhrgi5NUmZzFU1neCE1hjXfsIXtWdz2/XVaf8OdkL7+C0xSsa2UU88y9PR+qHDZFLk68
XP7fUVz4qS5HyJ2UPqhADHGRVlEMWlmgInlF0DoCnjhgPmfIpz07w+qPUWhhqgQ7ula0nXuI8xGf
PsQuHlSvcEgrNQFyY3pHANYF9zWsvtkSxXO1hK8IYyMOmdFRqeCJ1w+QO4QLzbmUYiTV7PntxYtd
Tyfky5YzFvQi6R0OYUO2gmZc5MHaxjN8pbCKXGd4X6l3kANsU0Y/2GIr3JQkN1IttJKH5RC0N9DS
V9/mqicvxKEPk9g9AJUV+TU+MGObO6ocQBf71Yd0CnnuDmSdwtl7hFwoUgTQAsZYJ64ntkOsqdAn
TvHlZlVA1fLkhT5S+a469Ac2TTeuLmPwdFNnTvQ4D9Zj3kYayF/3Pv6A2GDeNL5QA5Yl4mWQmMcR
DkVeVCUta0PGWvwJPjMqNKCg862uLWS+NTybVjfXxc1My2q0Vl8uE0xPYk6bReF4TtTwk2/aj8wV
8lO8qla7biSuVvL0mfDi+hEJIzEGR0zA1Oh2BmcV52W6o+WCzSArpv0PB56xMvytQejVGChV49dv
U7zuJjVWBmmprl6sDWTLJovm8xUUyiDVbeaYX3pTBizq2LAx7Q/zc+z9ZFg795ivTzEdfi3IEEOP
6txyAm5MHIYD3JjziDv9hsuQGRlkXllDsb2AWA7gpyIyLZWkxpGiik+kCuUqNIW9cVjyxGQ3q69p
IdSBLbsEZ32VqSbrFkqAxmCKrJDxhyi5NZyCapIXoO+wmk6vXPlMh/5maQ3ALKVPbOHPyVw7SuN5
g3sym2PGXn48RveBwhMQmRLt3GFySkA/qGvZNm0HDNq0nWV8fFonef0l/++2wHzce665H681tDo4
u0C9d9RAi3/WuODanY6WQcq2QwZxeqKB+T7CGQcTKt4OsXCWhu8z3PbD9zxdgH4xIkVtZyRAKm89
L/oL1W4ZB3iBGFv9AqHCSuPEWvFuo3G4ATpQwH906fZm4l+F238JXdbLp3FwoQ8e5DSxM7yRLPNj
pvcVJ6lDbTFmabxv3zZ0G38kp8S26t9lACq1NHqrDx9yyWYuiJehih5uSwH6UC2+uyQh7heG95t+
WWdt4QqfIfd3Lrg+neRbnNL6GvVAZhWjzYqo1RoD7HjhZM4i/Il3xnyIetW+/mxVPfF576D+MY1n
+mRV4MhqLdNVt349lgVPmB6RPpKtyVpvH+LUDEEJKifXZQ4PB8KaP/r1AyNeLBRga4x9ji1Y26ew
rFJLCTm+lbrx5shoUQwcb/7Qm8kGClx1lCThHE08a2lJAXrvM32Ogob0Tkz2AyjW1hwojSQ3uvmz
f6hjCZKDtgKisGWsj1V5jB2FARX3od5eb/wTjGjdP+OzOJrhGQUu4aqU1xWxlZvet2Zx2/e4NmGD
gw9px7uJ6VK6RyByv84xizZa5dZUO95vvqJ4MMI+Xtuvax3fSsyh1ASNwdpcbIQ2GIPrFXWFwM3F
TfFayGfd8+tNAmflBKb4uTGrPZrGpIPhXqZBkgsW99G9SEV4sS/Pvi2O3V40Uv9GPmkmxgUL43yg
8WHofNVf9T3rMUpgLE9NEr/R/a7jwKzOyybXnAojdjED78rOXMeJrgiUsQ2xdbzgFkY7CkNmGWtz
PlRdSpM1Iggb/M88NyabR0G6fpo0iL+d6sgrK/n/jAWwEO1iHcNS+Rjbn/+RGMHtBCjUlKKXL8QZ
I2jmKCeImgKqMLjmzqYr6q73yW4uCWvuuemqUaNb3wPp1g9m59x0TcI3RooOVSl6LyhUlVFpIm5d
+IjcE7BeX6sEKBtQxVptIAo9VauKLKnyW9zm5NoC64Sw6hD1Tm+uGzXKMUsufdF73bSxNmbo4qzp
HfEBPpMbtDrpyQ3GETyY9ozkJ97Xr3KBe9PLirfTC0lVruBvpGo7PfVNN7T+PrY38RH6ppGJw/JN
Y91Fl05ipKgKBxHKApg2wG5lRjHC8NFOSriwRuYIqz7h1kZ597zHvmwxbOHI5vBe9MV7zdgCsXqG
U7PuhCPzZyRpcKVs4249nKqnKkouSsuehZe4znUw1o5EanYgDXP3RZ2eiGZaJG13ge/TZOiekm92
U5jhA5T3ODJV91iX+Tgf3Gv9REZFxxFL5FrLmkbL9FHAJ4w97zvWJAyx4SdQhVdRCLEVnmNOJfd9
7jAhDJzjedW0q44aUTPfFw7tD/xgSNnHfJgIFn8YFZGHLkWQaRuIiCpLByqaEG25W/4Li9589Oou
uyR8RHfmk5gJH9CWyJhTQRP4aN0S7K9b79LHvSw+LyqnsbIueg8qDH8G2CQSAE6AG3z32830TCst
f10X92BZMOBMJamquixTAy47lwb4KdyJDpNYg/OxmTRT1ogjLgtdjH4d5irSJU2eYjWNGIgIUFOh
nueGhhiuEDcJQRGamx54fyjZpEJxVQMZLdzzawdwcTNRUznAAYLXAAQxtBklMx29+sifV0GelPau
YDUGFncwvM3H97EVwe5zJuqAANWlURk9xkyTmJiUHgWESpest6C7FpqkjJFn+gqxxya8ZLAsNJBc
b5eFGsko1FNTgNrtCfglbjefejgRiNKSFNC9VJ5Y/vAcEgdvYAPE//XjG2pC6KrQJHqOHBmvVkFB
SQNtGM7oB05pk/xaC6EshRMas32dxQCVYaCB9+B2IjJMJ4h5zuNwyUkbj2NKBXpe5MNRa823rHIu
NQzQnm1lTJNLNSe0wUFfXVN9lAwpoY/kHAn1B0A/zVFgiViS/cZafTAvYetK7nAB9Ry/fwVLBvgB
65tGRsRplunEer6SxC3sC2Lk1pO+2ft+83GaasnxFL/qiAaOD2PyYO8vi6tUxjGkXwehyjsdUq7x
syUh7417cSxfLvH/3OkfgNkeEfGzjgyNIMXsqxQuU1XCAjeBoIPlpR4IGuD3J0lHFlt5SP91/RuO
YZeyKHRJ8vWPtd0X0IB8pG/HZBSs6FLxiPwLNvhAMSOE6kxFl8Aht7kuZSFN+50GF7myGugZxOPo
E66qJY9Yc9BibcickVVzxg+gR90BC9e2KAl+ObVPxB5J/huE+bXxHPvTZu9cKUaDYokWNfmFdvrQ
ZKDxsvAzur1FwDR3aLNkbq8J6Lf2uyOsJvQKZPPTmnf+hzZRxaL1UdXGctaovdW0q5kTG4vRzPlh
3/6scM7DJoYuq8UJrC7EuC6JQl+XHcpjM6iaZeE7NAqT4pL0npI0HSeB4oqUnZVgCKLy6pWvgdfo
hnbt7GEpNYV+t1whB/sCB9wpH4KXf9jwCnStiYsb6VxIHPvyCp8IdcVG1qHnwKWIGV6o6PqbYTMb
ot7VzqWHhIwxNmyXTCrE48I2YYEo4LqODz4kpcScKln9xJhWpK8FrKuPxlKoBNE2Kc6f4YAJf4Sl
kooUlzVNICHeUum41nMGlVuVmqzdGsJOk3txFbrvc0zWXSP2XvszyWwI3G+H1NfE9qKaRJNUCqo+
nRqMU+CxxIrtGyewEEvvrhmUPFiVaCUvBSu5l5mLAznW8e9HTTmSg6R1WI5eQBGClrkNU0WWv04A
se+H4XmwYzoLejsvXhExe1yitKdNH/tKZZ2n74c04nJC166z0XkRX1s20xhPE8VtnQmu4Z6IcGFa
N3PbIpI1XnuHhqqpCgNXnhsvLFBEP1zMiaCusz9cPJUBgQeHzfCwq9peWu4cz1ghanlRIp2mSv72
iYGGvOsRygAH/JIRS5DExIs+Wf4J0nWh+2EZDaD1lk5PYzIXoF7ZF1iihV4q5/8t/pNsoKSrrjQ4
6b+dlhqU60UK/sUCuMLb057/6KOyeS9XmiEZAO8RCJMcTY9M1nf6gK6/h3B0chUo3eoUCZON8gHM
33H4vo5LSnnh2YMb8sBRYU1rV30t0UA3V5qi8d4yPr6l/UEXkHxlEuW1BATEwOvLUGfW42i8wjhE
7tTyxy3ZUftpECpdMLE5UlENI6TsrYhphyLNsb02usfi6Plv8+vO46rfxEBGGoc7hxIqAjd8NSmU
Na4U3eZZeTCf6dR3/aDE7+gonSp4EiPAMplEJdiWAwRDVsZOKRM5ulLsqoLbj3lmqwz+rSGx6hQs
qumyKBjMfc4FbPUrCvELmyZ4861X2FZ73VaHe5FY1qAe1MOnbx43TKfwKQk14PCtWUH0Cgcqjk0P
kanVTQc6YifZAhTt+7tiRF7hVdKmeIkumnOdEGni/wVzGU/KCMJrqNq+J5ayZ8mJvEew6Kon8+WA
VBlDd6/JvczJghzccC4qODNxme/r6q8fVkCcHC3yqI4oGDKvgFLqEh+buEQRmDOZlENfCUta51Y4
W9kOye3K0T8eBquOmJsXKH12HkB9fScpE3v1O6j5lIpvgs1F7ZFWza91Jm/6Y+64rLTERYNpZJwJ
Y1PcqZyLfp5kU7HeDBZfP3YfqZR0BLwg6yCWcumCD559IUouxa427TLMwOV6krDTAHa812MDaNRO
RKHK27/FhUPUh2fVv5SVfnPBgEj6ThEPkiAp1z7oNS5NxDx7Z6QoB5IZmwJnp2fd3HHCpMqnZ+L7
EVEfngJF7fCyIbgIcGSDFnJH4+mCESbLRSvKidweM4EAyz2NXMxJECDQp5veZt0XvHSfzdKjWQAF
vWItUd0qq7IhyaTHoH7KOK5+GR5qPBJ/fqXtIF6R+oDlA6lglQfAoTlyQ3zpOqMn1QMNM7SJh9jd
4Xq3NfNJEZJjDZzXwO0uCL6738S5vNrc2TLYFeJWmPoYBK143bZoUeZv9BmV0hwtP/qDuJHDUqqE
+qd2Bmc631HAb+2hsp81oAXcSui6Z001bihzpOxfsfmXGbOMcSqX1bLyxKHqbojPZYHly3Yvbm3P
f4dOYf0SAnErZ+Szn8ep2VHUWyKa94ewC3Q5CJ/1VJ5+C6+mmUJzvINPGaGDrSfj76GcAOpn/RXY
IHxn3QumlRnDYzx/43kRDG3cY9gLSGLiEn4ELZUqQmimT1Q/1Pq37sCjvMFVxSWXd8p0KXCp1ggY
yqfcslXMHEq9SC80FGrBnzydWmFhZ4GWxLCGYzzGvtLQk+nVUrf3yI8z7+7u9pKHpqnSL2tKmGEE
T3RCUY6vtEL9RHrhy3UaWGEFr4DoTCFE1iwcqfoxfOkDcL7UFM4OmNBcLosA0MI2jryifqzKqjjZ
jnmxVsh3xaxIuTtTcYeFHEqv2p643WnpCDnEYKXUDFXXZRysr310TcSgtpF+APCgKn31Re6ZxOHK
ABjM3wKZaDZ1vMS6e1cp9bMnF7zyGdncVNMGeOvf8l4MmNdry32xdoP1T/uu4/tnAotFGJZXT4wH
W4rTbdg8YL6T02h+2qX1T1VW1CfHG4FHyT7o+uGl70vw0c60VHDhPGXZlGLD+hl3a8d3LGQIKRsk
EMfpTDiVL60zpnm8wQVdNdoSItgOFvegh2o59/JgNPiUxIHpjZCmN+hMgcd9cpLhgMHd0Jh9x6h4
2V33chCnyk/rsvyMBqlPIXOrO1k3H+WBLzZzs6U/uMtynkRo+Sce3+Dq7mwvWp0nMmx9Ky6HzJ1x
LuA/RGeXz2hDe/anpH8XVPUIsGqmeq3uIJiYPT54RBBLJm6N88ZqOKMsE1D+qRx4NL9HarCoCwlH
+EOq0PKso0A7oT3bXMfMEdinqw8DHqFNkGlQ4Oov3wdX8uasZAiEdQ6rr/vQjB56uniYvdysq2sb
QSqK+Ib/Q1lNnV+BcU7GPeXY7W3WBSkxe5S//ebMX2BNmxxlzD7be66UO4apUWFziYTpzcoWc5vN
N55hvLwr+fwxaLNelUrGVIX17YboHk/URipjtKRx5OygCkuEMFTDhehAu1xBc+EzY1j3/Jsl9oHL
sgx7f+OyMeSa0cG62rxg846RKxa2XAPyuqohzauZkujqhxGMC20JeYJ26U0/Si+xiDmObe6gDT+3
LAtnS0AqfmwPjUG+3BB6cEp4B0ZiWem+OfCLyCuFj/UBAWcH3QKCkSW4HxqA8c7e03zPrjtBPQ0c
ZeZgqWVjof7Vt897H8E1GieatjDLszMdutBvaDJeOhnqkYRpQkPfv54dh0/gZVEAZnE5bV9HodAq
cKOFcYl+xjYnNtmgY3OzjFU0KQChMMKAWrLQ542GqSfUw2EcczI+omcUq9k1mkyXoSIdGWHalMTS
bkXmHbIwxLPZkSjqo3WVlQ6Yg6ra8+kTIirjnVNK+EawukYKbjSnc4XfZw2ny7s6XY6y2UvtnoFA
ME6xNhZ3ExGv/CRkSbQantMJ8P3d4h3s6xqsKOf6m58S9qXR0ihhiJiVKzZYJuNybmCV+4oetUz+
0PcSFwKjHmAKH8O1cC8sFk84P3del8LeY7mgzO5lPViMXe2t83A0Z7V5njIzGOobxadsHU4MkyqK
4+oo4v0KCzGNTMA6T1R7Z169yk05qZsx1lyvIZfpZrySDMG7UsVC54ZOzb8l7LVNcqXITrfGJH7w
zUJsLQE0oQWtazDzWsX51KcoLkg/bbo5kKEl/mQbG+V480xXHnBFc9OlMzDwF+mj9f3QSxbPyfB9
heIsO6G5eNI/63RArqgALC6rQrORlFEUkvJcuiE3zJqXAExz4605nncluvB6cUs1zRmYbCOaZnIx
iGyez1JvPiaQ2DBBeAh6KMgFiDaSzqmGaER7T1g7jHbjM4MLCpECWNQD/hJ5faZHtkMRSJRCAyUV
+DXoiZ9stTtyg0MrC15XaNkno8e3szqR2JjasaTCVq61CCNlurTxoO2HC56mQ7Ux9BjTNdDjAiT1
GyqU5bwxL1DoOjDjWUK87JZy3YTnkl2J4IyU5a1ImqlWGNguajhxfzCuQpdGdIz4BADYh0JZlgj/
H7IxJJrheFSYvxlK6/5ZELcsNgCvdL0PE6kVbG3rMLoWuOIfQiY01aBVy2oxvoEubm11VsYdK/Uv
ZmBoE+Rsj1wbXJRZBxECodfC4TwDTfhxmxjXnZzEVuQF7S7M4JHDdNWcOYfEtoU582io1/4H1ogf
BNdk8WfPBP+gcijeYI+WxWs9r3ZTpTcVm6m8rDLTUbIVVRxRZ1+JSEi9pRBu5o0f/fEpVvokGIuf
KNTxfVBlGgKpKvizgyZ5T6WrOd4pvuPuw7ZRrDyJ0MOCIetDLPPBuusKnz3cXJDnw+S0tgJMpfs0
IdiEMDLv0xEGJeIwZxvCrsb0Sk3kBhasYiGH+Wb7neFq/Jfw5x+t9nzCfCu6BOM5/I63S164BZDF
6fApAOPUhczfnCPwD8QwBslvcGbbrI3JELgv5RaVMUxTdOEGPoOiILW/zzzpQ7bm7qe+Hp+z9yA9
AKmJvtN190xBl30IXj/zctDMdECvNe3YULy58BssGuuLFwIhsMlmqwQCTPyJU6xEQzNd/fTZFJ02
I4Q6hET5cOEpSBn5PAoJh3+SmySSrv37jF/239Qmo4wzYO+TzM0lXS1soQH1ENqEKb0IlJvmAFkS
RJ7caj3LnTEkI8xRLbzNohreLx+9DTYmXxFUI4iGYxHqzs08iM6AfD/kTWWwkCa94s750jUem75r
E1g5LefW/NMitTr6JQ5dvnY0Qgx9EQ6SPVvj9a5ZeiLOiHGHkO+CbbbG7fUE1BbZeE6KFGzmq/f5
gV+uwtB/LCcHj5mofnX33Iz5a/TcvBG5GhXFgyjTibFdkqwD3WYSh/iwKnjrK+Kt3hLTl192NZTX
ETRu2WjjNvX4w5LOM+Rnw5jUHzNv+6tZDYIvBXbspuenWC+33eeZxFA3nXQlDYw+v4Ivjm0N0uDp
4t5eLa5jB8B5TZH16yglU+p/e73ShpHBVnBfiCCdpnaivo6bdtTtXQU7ZkqXIKc8vKlnu4mQjpns
JOwChtPzd2o82bn//jO8z/tMesywxx80QMvg6l8fQ1XLAPKu4PUYk8Cu3jLXCsU2i5fM6Xbvmbco
BYJ9lDKFZ0SP+TN4JPJvEINzEzWv72lKgdwo2hAZkXYIWrQjyPno+Y7Nj52DxdLefOYkEM33bxXA
PEjeXzFicVZDJEi1ZiQVf2GigrtTZZSKT3Uz3Sbl4/9IpwELRCyV6VkrG98YoKBKiwR0jP/xvD/v
Wgyf5pJ3u8YudAv9pHh8Jsaf2n1ETZF1Gio7YjFGBRkMTANLNli4gWMkFgGsUR0IsUIS7Sf4zCtr
qomOfzFK037dt78Fpf7JjeYwt/jEMOEA3w+WiyDLzjb4rRubvfswYXAIUxuRtyGfcmiCn3+SsCAT
rXP3ddAOrUklHzat8OHrkGd5cdElLL3FyUTPAbzF37GuM+9enbM45kJ86FJNPn4MRjrAaB6UeseF
MDaT2e0aZb/3SJdwnu0kOUo9bA2F9/7nuykplhgiqNrw8hlE+M9TRogPiAimTnJlR/DRDSQm455Q
XyhfoypMzR14GsC203yZXqYZ4rmIV4oupVoI1dkkLaxEBf0TCRsXYhTX3X3SvZb1XhX3jymb/dEO
O3dyqhZLpdJMmiS+xPZXDa4zo+xyhzDozgqMveKyJDRefkVOJ3YhWYjfxs5nryo/SV5M0qyuZ7iH
WCLI1AaZexXEZFM0nsLLD1EZL1S9aRgV0rpYsGE8dK1/lUlqZvN4dkFJYU8lMtXiaNtb5DCy84Ty
o5Hija8l/imCH1yTje3vcE72tDMUtIsv/Inic7OHaMF2dJtm74Af0TqrSiYLnI8lnBcABJmLR1d1
+NXmG1bcqmttaodN7ODzlXc20hcGaQnmfZlieXD/aiUizJUDtWmM46wBdICL8EmqDyyHavSNDuN2
seZd3YyQXrS3J9glsoghgLaE7hW4aTT1GNh9B4TtNEM5netV5Li1ngmA7P9OhBvHAvdKb+ljBPDA
/gebZdrVFI1aWk/n8L7UYR98kIp5rykCuaxp+BREshWoV57o2naMWvA77Gkv6NWY046vAQwaSMUi
6/tTTlNSutLCNY6Q81bTBafeiaI1urHRQ3IGojzMDs8b5ko8kihAYHvcRzFX1xmd3JDXUaAQEe86
un7Nxe0S6jXjr0adjgtmXEkvMZ4yV6k7dRrY6B0HtEwv8IcXtsl126JWBLRSS2B3/0DzbhaSZ0lC
bBeSGpCBfLc2vWc/0EvTEwCMOEdRN/fkxlRXKumwlugAXqclaYRb9/ZOrJJOiwgU45+ihYMhF6Nv
t6qqY82nPyORs3P6ohvq1ny/RUT0zSn86xohRmSSu7pOfWBTlEaKDeg2H9HZnR0Fif070Gbm6MBg
5G9j31/nSpj8qHmYUfh0K901ukb7au4WiMK3RFgKFiLSajRKDUGspRw1BdoTIV85O6s78nn5G/jx
COPcfNuWDKCzB5JToFvL5tMEzeildL24THnPlTQinQ1+3GOUibBvhjz4Fnu2Z40dZwt5XIV+JqRD
sEdTVV3fYRuPtXk9qqfEHow0o9+oz6mtiZS97LPAbvLRyD83qSBzri++wAacOFG+lHOUHhwEvP3Y
EIDn1Je2tGVA6vhXzZXBrK3NqPO1c3gIcgXd6XXvNpmIcI0uZl1V1hiRed0tlwjPN3fG59+XepK7
GR+IMZNzjeH2tTw+u1norrWYwZXYqR36vlrElNLutu5qdemqYkNwlQRQ0VfezZtMmAEfmHLk2G3O
+lbKP+drh0r7lXzrUQOGiWH6M/XkU9+BESs4hCMAWDdALHrgKrJyi4zhgW2++YBTTklUI6GHfYJF
Vnj44qu6VZnVfmrugyWudOF8V8PlKxBk0N7wSFdbltuA2CHVxJ1t7UcwnILarna/kGBEXB9lSKnA
QOOfxxjcR+wkA1WLGMX8groH2tyGfQajkzisdpxogHm9ttSgnbNoVrbUkcarZZbrbWmBiTpDiTkX
zTD+wrp6Ip7gHGSJ7h0aMLLthV0KuARSL8Y21VCuxhR/sH91wH08274QgusdyJ069Dw9LzxT0L7w
tm8QrZBzdqc5b8XvDoYsebQI/WORSxLXtBhZaD8VTi+jUs0nsDcw3t+ya5pvYo4FV5klOKesX23A
WDTSflRAhXJpnNTuHxIRbwKDT3q4S9ROojFt/r6KyLBDxa1ZsQVXekklS2YuhvcTE6lfjtaZ1Jnv
5UThTAE+j42qWX+zQJuf6g72ToJDN9xqIyXy7bYXiUoAaktjBGEIs2rogs7fAiAwFn0xpK+YxZ2v
YjWgeQLs3yS3rb5iXyRwRTkUphntjTTen1vDCpioOjVquXWnolXyvE7CNKsBm3miv+qAY31mzyaM
uKqWXlGIjpRi3yGh4pApJJ65JYOAUckrqxV6iReU+Xg0nXHWeptB35qNGoUiM0zsGMlN7fNp+RXz
d/TFJHv1xT3hW5HVSSEKg7nSfrkrVv4VIo8lvoG1DpRMPrduo2uOgmY3yYlyW2XwCICfD1DJNSdt
pWSrTE/pVneej69F+lKLhsuxnE9Y2CR0Fpo7cTC7rWVekmp6cn1tviXK1e6hm/llRxfM5ClWTwNF
pTXDVmzxWw0kP2H/Swfqspvezih5Xf/zmqVzUsbnhkoTP1DKPLwdTSw/UVKTSElmG2URunza/A7L
SxQdGOe4C5AfC/nZUWH51Fg2KURG6udm5HZ2/FawPMvbo05Cqw2otWkFdiHCwuKkloqHc8zE3jDq
6CqebWZ1tyCL/fn4R4uZawYsLMMHBXqMqhiaI+qs7fBE39SpLzDVeKZDQpAg2cRttNYrfIyYzhlu
QjItQaSj3oAntYIie+GIkqQUqf9CA7MxUZadCZWF0XJ2ndFU9JiM0xbf/v674xOBq8ZQkKVDlZ4F
Wt95m/7JG1uv3Vr/w48cc/mTdhFr88GazvWWJ9Jhj1/VHsNVrEJfr/WZcWNc2ITrYJJJKxE5Cqn/
o6hFrPH5HzQvXua4UecRoGLqEfcXyvYE3yTjVnSy1z75d8UC14i7lfXAhBJfYfPv+jS370lh+MH9
O2MxHsVQ9i+h5wUqvYh6Sy5eZ1N2ygQI4D1tfr88Q1zRmW1zpHXXy461IQtq+1d6EBFlcAnLADHv
i6MqrLDTdFeHZvzoX8NJb0VHsCphLFIrjaloxoqjrxyszqNNd3OfP6zuYwP9EzshJrMh6rDoWYFn
YxxUEIuoKIG4tM2zgO/VMz5GbEsEEQ99kLVZC8fmR9tLurP30hfG4LV4YcI24BbiyNOMk21dhpUb
g0nzR3Cmf6tzN5pLrXQC0ofkHfBd2GK8NlqZoisBF2eoqtJOrOsDkUtNIqBRwYS8PHNgNUi4Bm91
a7BrTe0jlG71fCrvVkFxDlvXKqvcFMWF6AemIbx4CGznj/CMWI2Uwm0+Gm8DHwxxh0knlDrsB4C/
KNDrxiDvxiLpV/Slm5z0T5NV1NAWSTOwxNBHGc5Y+PblXPVG9/2yTEVXtsWNeZE9SC2no+LdqH45
4bzdpfVw0ChMTHsno+wyR3A3sghUEpV45fglxCEaLnopz7jN0dAPudcONPqWN6yGnrLgcGOMnYRb
ddJjhDpiqHCwi1Vhwn311fwuuncZ/ICftmmbUSKsaxoFu/+UGlp2bFs+ppxAFAgWO+Y9V488Wr25
KWiG3s+A+drjGf1rTcze8tv1xeXE+FrIn+F9lRk/BvxGWsLsqj63sZK4MantsvWYbuaeaE0lfPSU
QFrfNaP/OyayLUnfR18lkvQi+BuGTtLfk8ZfY3186Zbr33lS3Uft8CzslBJwy8Juc5Rgxmj5yDDV
7ndIDl/G6qoBCSIjRTVbJDj1HwGeGBMxfHCu0Pz4fca5DLe3GOv3q3l8KpR0MSNEQbxqto/emLA3
Lgbzk+SCiCKrjeARIKl/D6EmhC23NX6JA3FCS0NsrFHtiK12AE0MasXaF6GfAIIQZhQkieZFlpjo
Flfxyq5rkX56bTO6xdgaiGEg3zyd8IeBlfpuYWNRkZqU5+zR8jadA+UYhpT5ZaBSsHsnbkZFF1vS
TrT8q9tOClvvLm6DzKgJO0I/LACfGm1fm/+rdy4KQdIimjA9v3afRQsvEcQCAZn1dxiAgN1XZE8R
SQxhC4xbTdYZC5N1LlReg4dN4f7H83yziU5R7W0oMj3MplSVyimEmgkopdR65G2ePBRBaD3JOGtM
UGQP01kvllyxKMT4joRjgaPoG3fXweKCpatuor4XIRPK/pHw4jDHUaZDXCWqFemVUuArb6RefM3/
kgpRUYuzzwRok4ZL7j4x/McJwBrMMwnE2QKJeKsylNGPWqxD9kHcApfdEQkTS4VXmvhlZTBNqR3j
sw5OtwhxZqeAAM5zjfub8fxCCHFBQByH60cKRYzK0v9G8vKaBVh7Y/bjGSXqgR5hLnE7Kxtm1fTw
ZyHCZn4MdWi3fGe7Z1tWyCnBl4wuXIN3YUKoy99p2ov3D6/3/WwHGIHjuP8W7hSgD4G74LtIvQ6y
bAucoNMZt504FaF/2Z14CC901IZNCIhwr0o+AFoE3qI5GGJiM/G/OpY0zHCBYNaZblzi7+N4YXI/
KVTxIzD7WhyOLTSm2Kn7ZPELdcmt5AJJVPNwpx2idwdKPoYCAxhZWuDAf9ge7d4v60qyJpptIUxq
quU5GY5xsK8RIZTS37EnHBZa8kV10RR9znYgYD6BuP9xpLGcgBfS6Fc1qlJf6k8TquqhrXxKXbSr
8BibY3qYXttV1GF8kPStuKhB/2MmXjrLnM8Fn+wu9ivz0vYb0SbhboCVC1M1CSsHyieLjF6ji/b9
jp3wMdHe+DIaCI+SAF72fihKtXrBtUNVzW7yi4myxJt0vtOKpZKVZXH9iN3wfSudSO15OMoS78Dp
mDpVHwdXiFrDGYe5ZSzdJoBfyc5uHm7ylrnf8dSQmHMJCRdHi+5TAjqximRrphrNOLew+sShNY87
6Fujd7CoFdfLWrr09w9Gtdb2gS1DTnjU6iY6YW2bZHcq4ArsLa8H9kdRsPSonkLHw8fEGX7ynqPD
YQO7lLiuSLccelzdEgLbCDjJAImnkPwBnV4x2vWTRa1wLHpW1aGaA5D8InlTpdnJC2JOoU/O+1TA
4nTaZS27QrZ0t/QsdOrYhXSIleThru9VGZaML2nQrJ/N4UrZbzBLJ+gUy4gn4yMT+7JGqdupASMe
vN5URmCSsaW86egfKFSlL0ywn0QjoKsLQ74yUdZ8dUb7KjJcqEoXQ2d5O44c0TnjU3jrTl5/0SSz
QgB2wojbCIaViKLaL+bi6hvjY+yOuAfbHWJAGmeqfHGPXexF0XO7NMXoBk49Nk7VjWAkPbHatXMv
1B75gpkHbUBmWcPtk5x4CPfvJO3WvOJ00nA3qleVpvzIxw9uRnvKAp7C+lrWAy2EYxzQYwmO8naK
eSo9F/+Wd0hyWa5QKHpiWqm7nNlZidxwxQa4T0qTN301Adv41Vu4aMat2U/P98sWdmbor52jZK5a
FBKop1Rz0VhN7mu/GE+41sKFG8CQZ7rtzb2nl80C68fUC3wti8w3255kZiLU7BcTYs9thxR1TeOM
kMDoQcWePKctGbPn/WTGxx9QwZgyvdTJ8XnWjMKmODFAMKGQ37eKh8wK28YO5GzZPltncRIP5n5K
KTea4CJ2LY1XLAiA66gppvq47EXDWwUWf5JZCRe8YB6p9SYzN0BQOhWI4pq/TE7MSdOZKbYUYhCO
4D9vIPJSQrixF2kFNDxiQP46Nue9yBitvGPvVFzBRaZu+54SPeCMGp9wvuwb7crGLDNHCTd4sb6t
3tviCxRKj78/KgSAZ0kawZ+dWAsezaxzi7aOqlwS9OnQ9iH7BcipulBiHvjfQW+Kdxm9812HLfkn
v09GdjDFtONrYc9cvD+7BKBsKpxkk7PcMPgqPL2p5If0gTMIdDTd8nw7tMEx/7yTCn94I1LmHBeU
KMGB9Cd3RyAsSTHpXiEBJGQGHp2qy0/1hSqo3ftoqcL/jjxW9AJPL/C4dDKNgYY0uG9l2FCgxko3
8zmrJiBdysgfvfGDyoqbZdWCrEPoOSpued3xFvXJQEWI8cjXknE5BwKplhF/hyL26wprAGFC0M//
holcveGbanfBRTkS1UDnrrOI/YS0FPbLIBpwZjqZvv3udjJzSxrqVbkJkafYq1lKiaykcyPpySUO
xNokCZqbPwE0T2L6UQOHMHbWNNAEqMJPxAkjS50mjrmp0dMiBP/QtOQZxWuMS2Lb7aO0OVmM9BP3
uec+MOWydRWc4EerWodD8lsBPKsm2FA2ZNYDhlCPLNYdotWznWLTV8Wab/M/7K+ElVzP7JqOWz4D
Uq0cvcyOAWkb5VvL8BcRbLKYKvfr5ZgnxmyW3qQRWjZm96NXJUxbKR+xlRnbCi7akAMbk9mkHrI0
qU6lDYmrjv0EX3l7NrEaH/vssFjONf0zRpQAnQldtoTly6L7pXRngjdiBenRrmfI6WlqkiFZ+PKY
cyW5yIsJLPOtTuTIJ0nprgWA1y6OjdPl45EfuG6IaUmu1es+581kele4p1M/0ykcA9KRS6LIbl2p
svqd1uFebvss2Kp5Ki/pLSpBvvuzadNG/t5Y+Lu4F61LYoAzzM+sairbS8Ek/71xOQeZi8FClMQj
Y1U34JqVbiTm4rd19A5/yV/X9PNL943rqwZWfYx7Q2d88faR5JxFCctYbNzHN5WnyhvI74XCC99/
Jf3n7TDWy8BMCPM4mWLc6Jpwh1IQTzjNHJU8v6msGmY0KttbZIdu5Grj/x21Z9kbDVPExSLy/er5
6v6URlmSK6yWW1osBu+Toy7soXnoyf4Le1DrfEEtzvPnzOEKiubnNK6LoKv1gDiWoxV0Rb8e1x1T
vpvY6osERU2gcmMTAeqUA4fbE3sfNH8YD018rPvzgYVjnoFaYl1hLwpHxofo1hj9g0m0KpdgYyze
P6DcESV2GyDan4IJcBB675ZslBSejWF45JCPtJ57dGAg6J2t+URcRA+MBOqhVBVm4mxWBThlDDHU
1GbCTcvftLdg8yWw7UH1luI50HuebPJnQ1kh2xXRAHPRfGDY/i6SJ/exxP0RoyWXU6meNoH6mozx
W8CrsvU4GjlxKvVzHbtC8NKtvLitFvXszqhPNKyexXDQIiqKlkBLjTs3Ft6pr93d9ud71SsH43sV
fzAwZOiXJV9ZkPeyekhrMYbkF/PpHB4G7ouFCCyGM+TnsXKPb4XNdPwDr7KMwiPYC/3hLjtbhNp1
Kz50S8EF9ViOhnUtP8KMQLtI6YZJw+yIUSEWVX2kz7VZ/TR6U8hUSpcMLwlsHbjQsseTRyZ8EhSu
Qd7Z449lLBVt2BL800Iuhs3aOKwdWf7olFS6NgYXfnL4GFsE6ao0ZfMPJjT9CIc/Wb86hx/hQNBl
cuc1HH+nin5LmYltW97y8IJK5NjKLQ2DPq1WufeH5u5yCXxYlzvYmqOBFjO4H9TsPjnzpZEk4gj8
xfxd55hZCoIkiJC3+aZXss8KGooKVBpIfFau3mF43PdmGe6+ucIZ6ZSNok+XBYuhXZQX5TmpRpo5
ns3n/zFPyqw7Kx+vBQw9HQaimZQQdHJ8tVvrgC8+1/Q8ZBhisqq0MyWhr6W57O/lwJ99JjSFSDYW
s8850dJYxvR3wk4zIC/e2/9r9Y8m5W32N0tIRs2Rkh9tyunjk0lJiXO5NuK9MU1m+ymxe4rLPXkK
Jzhg9/HsJpaSxYtFznYoKIt/HYM+VVvcUM6RrsHZHt88VIk98xKlICaK2ilzKufwVMmU1+MR99Y3
YaF040bCkkx0KdipJ9RcCxAcZQPyGnoYzVGj9DvwKvUbCgWBmv6taL4jlyzETPZl2bB/eis/rwIy
ULykA5suSwFIwVNpfmngZdQ6j+rfZS6pElEQLEZoxDgsFG8ip8utdJR0TX04fnGe3JSZppDl5M/x
4pqdhj/JLZfoo0MhJMAvv2XZcZrCAOCX+2q3zHIldEJg3YretNWH2IK+JCHqBKiwHURFgAEBLNOS
wLY/A3e1LMgiCoDPx48F/zGHBC+Kv81TYDTJBE/GS9hwPQog29m0q9RYFuyJfE6ALotNZVL7LDFy
Vjq0O4pJOSf/1AuedXfgrAdb1elyCxgBW6aAsShP4wljVA+KiLhEUJeSfCmr+C9MkUC3RDw5y1xs
TbSYxWf2TeWVEP39nxHB9oS89zeu6HfwnAe89yn036OLFf8DIrORzlbEeZK8dZgj+0MxUsLELlOq
la8cEOBc4XArXxO8pPLPTp3vZYoRcAWabtS++LLWGU0qe2fahMurN5MmwjeJrIkJtMdoBKHbrMD8
tH4Rk+rAI4qUrRamhpmvFmhVjezZV2vD3OkOh8EIz0JibD1dwmoGS8rBzHeZHRD9+lDumA4NINeF
HC+yKBMPoVi2YBW/SyxsHm6dVGDzXbT3L3RW333CntxnGjSt+h6Xws1zh6uzl0EIDPU5ETESOobY
sz2w+izS6k0Ev2M2l5duEOOYiXHn/Fy7rR8KNYOO2SgFa0RYV+5ZllL7E8h0M+r3ffMb4MSkJrEZ
JJVd8HmvYsBheuGGgeqXZtaLjfRGx1HrDfYKfoDCZFCljhKg/2847zItTLqSfF9SGmjOC/SRV4vq
0niwBe/lzNpKxgvBjZ6H6jix63TUT4rlRYu/IN3LuhLjdJHfJBO2xIP1AD5zxT/hSo7yMB8LyDpw
vZqUy45K1/BoghH+9OwzlWPGIoZNmlPZ3pR6fkrinfVpO3dySAFmjE09leLmXK1ro2mssf/fe8L5
WdG5AiQ4t2v1JmnRiQOlmiUfElH3iMzel1cF9AbJ1ETTs94nKKcRLCqSVMBi3p2lyPG4SyZojwlQ
dItqYpWZDrkvNLbDsHu7r5Y5mwVLNbDs/tCe1AB/nac4nGHT5bzNFRZHsifcmKCcO7x31dNJz6J+
V8Obs3zl61zEn6T3fhw63FYNmcorrLy7KDLK6M05BzmTFk5HgM5VJymA0TY5pvxEHJLGkeaPo9bL
Pyi0VmZXYQOK4bj9iEutdtHDfZdcc9Vm2AeB5yIKjq2bJ2HKcg9jCR5siBU5VK8tDcV0vJCNgfqy
BYrMF4s03UZA+n+TrEf9E+S6bx8NCxhC2BT9qmDUwpQU9RGws9CeqoJXVWD6r6bG09y3fJKzBxRy
5QL6gK6C7kn2VkO5DhkBv9OLIkxQqTy2lyVmRCfn8i28rYG3i3HBWmqRU/ytJfKoXKzk9O9NLQdH
3BXPjCJMTbOZfkmct63D2UO1ZZlRoNDpAnMnDgVBz+7UQITcmyagMeNfzTBlzWi5T5DPFh4lYVa7
FVowQB/hlXKPHM1r7EZEZIfVCI1d2T7dTMtzxxa7Z4A8nCnekoRtVQBYfGRU0vMwzFkL/ipqHsOY
1HQU8j2lgp5UWF9Hxur/H47f9dnkgFbBxAENiDYGTrIMjBUisr1njLVaHGUQSDWZ/vWREvWt1ik7
ZDHBO9YzjuW7zV+l4C2MnzGfWqytUDBTPPY1VfLZWX3AecdF49AXeSWPbwceidauQKMwGD0w21aA
7AojnKw9v0oX3i6XPPmFteGb2zkF+AWwxqurNGEtd3fxxaluV0WMyz2ccrf9FPBIP8emnsGAQJw7
eKYtvfX//vZkbXNy71fw9nFSUGyIeAMD0NFzIb3X5Zmdb/QwAIC22pcCTL1VwemkrvDQX77/LYi2
xDKRyBQIbPuWu+iDDL9qIZ6KeZQMyeYNxK7vnLF2lm4E/PVL53x9dVwDla0uyMSkg/517KyiaYiZ
AYZs26XgSqpc19kU+UBJYIJJGHhg/druMilXloh9ZdDY8u1W4cjJpwzALp38izb6hqm577EC27y2
aE+XZmaU6SdWSM/Ypv3K+ELOs5wOfGgp/U1aQfiu8JiGB1wmWkCFlNhQBLRbHOrDVubvLVCnWrQ3
qsKcxHLY0UvKiqJLP+OM6LCw12oWUV/ss0OVWww6C40CJyZ03Qq3oi6tNJkDPoCwQXDrkn2c7PhP
Y3M3OyNOx1q4Fow13AplTCj0Keui8y9ScxDfUhK5CcrSWUhUcLnhToSWS+S3qW+F03edw6IAOtOy
8U/fmR3mi5E+WOIV1XTuRDQO81fiYgavyB/OE75f1dGLk32+CKP9dsZg27AFKbltxXbPMu+4kqbp
bHptZOpCNCFnHga1ghmwkTlsNAHS9AxR5YHvce4Noae+Okn/B7fxwdP0bUK5njXL+3kSd957aAfO
3NKPdKb/QN7J4mHTqbtEsxQw8MNl1pWGWq+vl8cJ3t0JKexAXRo4tnH0BoWtV25ZbCh1zt57o0m4
hvcfY3nsB2QLroikF84ukPA5W1BbLkUzrGtP/l5ttDqofj//XqvRDoh6BlH9mmCKXA+RFgRAMLKx
sDw2rC/CxKQK1qurMyOp5XiyvWBSQaoV+8g3rkBaKyZ647MDOpeRE3BI8Ue8e55ZJ1mNqo4IJq8N
HWX2P33xOU7lAOctC8vqhwU/jhsupX1+WppWtJjn9ynKLvgwZapyKu7ZRKkaJnCzwYJ4RrOzOvbT
O/yDTxHVNDr52BFaXkz74woCiKeBk1xBdRB0LXBBCL4cHuQlT7DHx27MJx1P/LTl6Kuwc0BfKKui
Edygt5Ir5iR7wQUvj7EoqewMfRWBvduf5eM3nIZtmJV4m6e2uaQlRh88vtjGQdIjCdRAsSaQdR3A
mQnaDMxpcsO5aOjHKByb/ZnU07T2t56X1xb+a69QrfrkQ9rU9fCvG77s57JW9eEnx5bwIh4uU6Co
A80hxx1xAkagPrZhOzp4yiQ5fNJEjgIXtHUl0IOJfixkxB6YG8GBOGqgkVyDR76YxGXk1OZqgXsB
Hw4Nnk78IHAW+AqawFXg7PwZY3E0tMfH7rvW3biGoX+Eu57eleCBBFrWBhemBJsQqkWg0V5VZrJ8
rvyh9Hbzxgw4MkX3nGmzOULPROUpY0xnl4sx7R2Nyp8kG6++PKs61967XR+b2NvodnCxeWfp4d5s
/GWRUK7XQSVq5sBtsPVZhFbUbL5n0gDdguqdBt0rA7nIYEHDr8rD1JDg3yqy5ZAjNY+3yo4oeDag
6HmW/zv/vcvdNiSyqeHzMev09eMq/GIcZCy/Krz2KnQgtE/JcnoJ551kVvPkWC8gWRPTn/4OXU1E
a+wSHiwatJ60bN+AymBtifQl0422J6yXoDqpRFav+jovbymweOOwXVefFlepe/3+7IkEXyUOt438
u0Xb+/g5O19OGNTqyDFNswsmAO80TUuzVx3CzVdFMoME0RaR4jOXuBhapupWem5qds4pmJcAPVIX
Fu0zv7Q7QKRRip0rBKpQ0vc38HP0V4W2EBdBOqXrHmE5G9ktxuA9whr/yTJyTZZTE7NnI6/cTbPo
qNI6kWg8jOp+PTCQoD+Rp18dmdbKKslVAdqbS/dIfXDY6G+U1relyO1TIekTXKb+nDtPRObnGY+y
LJAYLw+tQBDfWrqox7B31pRzLx68niQEWYkDSpe+jO7+3tmXT5aUQDeAJSdWJBpPQxhlW3dL0Cpr
01ZigOTwP8J4uP4xODbfN+aIrdcVlr8zbMfOtbnlbh9JowZNQ+7ETVE18q4sq31yAGjhrU/Sg+Wh
MdxncZr8CJ//19iSkHX5RIqw7ytxXqPFnK+a6XfFLqs8PpUcL7Kwz4YDePN1EBgI+2yY2Wr1xWB0
X/ngmMsLnrpfk3j41Ora1L1j6QJFDvRMRGFdUawMiuqpQJBElqTyb1d5/mH9FMqi1nawjo0Of2/s
fEQ9IdD/AdgyKgMXEk7JfR0HjCwajXAQOi4pJsFRmknS2eaD6lYxqNROW7xFFa5jtom0nFL74fZe
B1adX4FpEsJxZPpJxJUMrYsKhordO4BHlILcDeI8tpg6RnS56Pd5StKIZM4ZfPw/NukT/dRwJdOy
0Qx3siuWOXLgjwa9H8MPUsGH7a2+Os12HyLVs9yHZSqU+nwjSa3Mcf9qT/Y/9LcpQNZwCjCzD+Dj
ADR9/rSyCONHUiQ8PQQowBonhoPHj+1z6lRyiaVTXF8ytcGwtGouTN7QsOkBM3y0XFSCPFBUgoQ5
Kvp9UJsefLbjQd6Zu7zPxwdeJGquEbF9t/l9KkZ07YjqkFU+XUTL0c7bE/9nz/b3Y1OnGFKsRJvR
zawOYrolM/G1U/smBT3NnuJzhXybuVb4YUAAsdXcrjDxmU6PEdNFEMDibXmprpbtv0jFAC8fFOU/
FvhqoT2OT4FvbWeDwIHBDiTtrS3KjzhNzTylAvai7AMrCzdwAfWFDWLPYA2BcJ9XoTa/ZbPiN+dq
5PBoo5lcKyRKsFqx9e63o8vzy9k99syzpmVqpB6Omab0mngSE3KWZO7TmKAAzh1et8SQXicyRkhT
aa7n0jYF424SBzdUBsOfWWjg137SOrhxi4+Oc1AVS9AHxsD9Izj9hRjMCDePN/1Hgcb9miDcKFJn
eOfLenMgCpkD5ruoST18Q7InZt1Sv6kNVPRDvHMqQAli8f5XVb3kNgvnHAhSyV8ndC0J1BK5RGTD
aoK8Dfdp0wlOtcDSd9i2kpXB3/Uvo4L42PE0ZCc3PdC3Q/C9AmPy+nHySg7/FWm1+IAvEgB91Xq9
WA8eSDYe/J++sFbJGMaNU7fRBkW9raIZy3w5TrTYP0E8OukxIYKPuDj/DTe85ypSi3PPHtV6XyUe
S4hL+SpmokLPb5LqaMHBHz511wFyL9WRtqiAEZ/hNhsiZZYZQuSAaxFE1C6JjUUH3ZdeTsOy/sxb
Gmx4cDIeph61bp++jirnOQmc69yXSDp13n+btm6vQsaQAl+EqMQRm7hvoExfguOvInBxXHaioOdD
6ax6ZlJvW88HeSKXUmSTcNJdCkuSwB/HVVjIYiO5njLBz+GrzRLiCz2KL52xhkWFjamyRuU1x6mc
XYwPLbX4Rtprw6CqZ8C2i17DoVq0IH/7PdQ2Ory+ae71IDD6UxTybKrL0imnGLHgXx3pfUXUFD1h
jKJ7l49YewgPpN1jiiXpFlXDjWiQQJpucyTcFzoWJZgthafapfuhz793tIz07Xux88z08bU1SMgJ
S2yYTCJobEvL6T+6itar0T6VVdNPfb/HtcK6mBukk7A6x7alFy6i/yg6v8dVx7UKdsxL2H3+VSe0
PKNBLQd5uD80zeN7c0Z7XKr23zNL9wRFj+2WatBo2g3HiCiqXnXiZmwzkqlaQqiSZ/PXJab0X/MO
QW9f2TmDm+E5mEPjCEkvzN2ZQLsDoSibFaAUM2C0iLbUOjRdL0Pmn1c3tMUyY6Y4AjFcr2Inn04b
47UYCu/7zHSwCYYiPbn28pIKLFfWqv6CQjPRKpDCR46XXgocvyrXgInseV8CWoiAY4TiGjEaYpfw
C6GH/6Nbgso0ZzUBjETpDmdGnQpjT9F8oeM/23jIfz3RbPFZz+iWSyYWH8Q378WNyBT2Toa74w9s
AAXskXcaZAUBkgYhpDE/I2Uc7WW2f5CTOJuYk4HLC2QFwpYJXZ34fXi499Ol81McSztSIvx81TG8
Sh3JRwUkSsaKg+5U4e9+mwuSUlD2e3Ol3lNjNIVyhe4WCIbeSfSPpZAf+8BnS40MLeBM/Hk7AJrP
fCfUcb5g/dnz/7JRCgSxTPaBjlfdoG0aQS0vhVx3pj5NPwoQZiAuVQ8dnKjOh1Z6WfHOgOVX6ETO
ScKj7dkV51+1DdJsIEEMd0nqkjl/+YLKls2wRVN5wfpqrCF49eAMdhkOxo27RNgolhZUhc41e5M9
JqEut1gyTZA29kHBC5cMRv4iOXWC/EH245/kOCu0VFqRN21x3jILDp345BII6fH3kHU1vSmjhL5w
rXoanUHkJQ/oI1nDV/bYmS5mRJdjA5HJQjxYl/jL8c5Q7efBAZG+jjWZubLkR0mNqUfRBksVTu5e
GWn+IP34bbpYtsmFpq0IOokAihVuE6sJnLq4PcV+sOH6SK8jXoRPDDYmZsooIHENdNOZ2KcCUP7b
rz3dJ76TUYfQtoA6FEXEzxSZl/yM590pAgw21WeD7zAng6IiEkY5aomU8vgcAhmU86fWOMtyZaLP
ZuLYYUjCVFOdJesTnB43w2eFQaSV0op6wjTcrR+DuLM0qlFBW6t+QilBtpIpiLIx2tcrVGV9mATD
PDPCuGYOKSWXUDFwgUqbrY4KHj+zP7zO/pZfE6k7GSbAmy3vwF0TEec28vR+FYkaLK8oSPK8KJlS
rFx1fqHg6ofP5RAidQWbBfaoE784L80g56kSUa0oPiJ2aYOw9BNSzv2R+PCYqPKYpp3b1LCndKjv
oggSjusZMVvzBL68ZGb1FcyKDXl6cjliQ99xYLEUsVm+8DzUvdagrRpdbjsXNvHKbLrHh+cSUA7v
AhYcBZ+vCTBRcx05IIcXDVbmBAKwtQNTK3Axqy2tqWd2QtiN0q8NeXK/hPSWhiIn/VcnK9LeRQRY
x2uC27U/fv5fCg1fkZJuqMjnYupJugO/eEduKdKerrBvBocqL2bsokFTbJle+0k29QuwYcpDuOrx
kryz6HMwLzYLxiWlDrp3GHAO1KRPU6cSVkeZOV2O97cH5jfBBYijQjRNxbnqJdiM4hZ/PYx98+qE
nX4bEemLIsvS8Q9jn+b98oISKxfkL27kP3+SqmwFgK0y1XN0bQcoWnEvJZxewreaVOy0G5M/O2vN
+mXzOsp8uKHrFr1BLQYMP1uOjg3OesE+leEtAo+LmnJDAbgM6c1wFGyeOeU3hm4PHMOgi/LD2pTv
2djicgPlHWEhzu8BxfKgkBZRJOcM4gfD/zcMGTiwE9fHLaRtm4ZRoQdi/OderzvO9q+sL1t9FiRN
JAo2ags86UNAwrbNHFTm2YzTVhotYJhGllBLJNj++S3XNSm4+7Xam8SugDzjda12PJ8Nc/EH9akj
SPKDWbBP5OwGY4EPxzUrP28s950BXNwJpYUeVugSaA65OAMkDiCiEyN8S78xZMxGcFaZchWfQOc/
Su+fHBp1yVJ1NGhuIOcwDVzJ9g+XGN/HHjYJymQKzUDnLNgWI7fx3oMoVo54ZAaAMxBwAf80yaYP
hVstba7+rpHmWVs9U0U4rs2+/kk7vDZkWyJv9u9q3O7/1WlSL7Wm2h97gDabcGnBG6H80c5VrhMa
HjXdl24Vj6tZ7RRK4SQBpmE/PhOzOr4thQwL5Gp3NQ8Yw0EVuiM7PSfnKvKZVpTMaxvsm9Brhy8D
xEcSajPtvs7QHBTviOX90bq7nZSDaeVJysDadRgcsX1x5IccSktWkzue7zVxP3f5Dc9XHC8uVrBA
YbY7CqM8AdqSjvVbXV3WIDfum5D6lBlRzk0ZhtHqGS3L5hGEfHyfu9PQGsuhfT/zobHjvIFcEEJx
jq3P5D57E11gPl7FU1jStoX7dZf4ZE869eaq1Dief00KLC1eSMuRFbnv45FeiihR1Wm88Q9oLOy9
qVvgN+WhqI87tmFPwuZsfQW8z+AEotUDWcjLD2vpjzqUi6K88/d/sLpEJGQ3F8d5G5vgnx5v2cyZ
t+VqBsv52irs3SbtW+NqCwKNU+EQzTlsAuR9lFRPJVEAim70KBFZ1JWvGwuNBHiXekCTwkubuVzU
wQKMi6GzXwbEpbb8XfNMWiV7pQO6Wv+qPh/JFN35eppVtytTFf1XN8HfOdiXhulNzTUaXYduiqt5
Et3Df5oMBeJEoXtEsxWgpNqWQXRwGDEtfgv05XRmdum5c5g0oaznFuYhYxEQ5BoBgvfKp6jN4cTp
vho6F37rs7yfVUJfBZEXjYnAZDnMnDVT586YGc/XiVRl0F0K+woiBF5yLFqbwu80Vhgqj3mbxdav
OZ5JEuGSu4DoeeKExn9CjPfNn0bX1cUIGwpbFJVLuUBhBc0WCXelf0rQxMINGHsXMAASbmL730Wb
/fJ9jsF/2xyKzv8YTWww141yVmJ+wr2Ln+qXaJkQ75+uv0uHV59+KQ1w0GVsbpG4pkII2+RN3Zlt
KmaoxWR1hfP5FTEtdHkXgR43a+++mv2EqHZThrnnz7FIFVdQW6dbXoa+S9Twrb6bw/E8r4jRRS7R
o27kWoISi9bTSu23dHG36Arr9iYnSFDhrcBP2Nj303SWq16FFWBcy0JwCPd0TWGZVLLx+J5DoLaP
RzMEh13nGlfrhgxAznS6K0l4YIzdCW/NKCBM9Hm8JAbmF66EZK0VdkxvthZ6h9t6os/Y3FbBrYYB
OsvtATSQWzWSbgn1l77x10mfZkfDGE9+0dA/J7yAa02PqbgpMI5jGKznqoBy9Bo01Eh7AtO9a+5f
Ngc0833aGqvpKD3JZ8o67NHHsuj41/PrD1rpBarvJmsxUJ5gQiZDx39+kCNjcLU32PqW24JxtCnQ
/A8zlphFC3qg1el02FezR6zumNR/155u6rMuuA1oiDYY/C7nObRUBJ8ex2HCuzcEJX+GDtB2/nfm
CoIvFlxRTtO6yNjHkbv7GToYgbtppFWTjyBlh+r1M+F2J+BXy7p1aV+WJUReIbN+AzzMHHpMHXtG
dIlE6dYmyn0/vt8h977wA039yPSCQ32mdnlmStHpRDwyH+/p7/isFHwI4eUnJLRh3OLqEe/hq3Kg
S4b/kFvlaB5uwd/faDQZWUVdj3tQPXrQoTUlnGRR7jfgHGRMZ0hg27DaxSUNQLhhkPIjUV15eu0v
YgOVK9vH9SyqZzJ82k5tcQ21S2CdOzBBJ0ij1wbXRhVfZlw+kjfrEkiLycbURCWjtu0XLehdah58
mTr3xZwlfGIRCfRDJ2lewuQamhd7J5yL3TDT3i0j77fWbp3hGTHP4HN4n7aKD0czYad910IwSuxd
6J4VICqonum6Z6x+w85F4vEjWxV0yAbVBuvWlg7YNxzN5Nvq8NRpm/5825k7AM0g0U1Z47aT1xE8
qwoT1zAW9Hj8dTUacXNff1xg80xTxNzbp6db1njPhaSrCRg5EJhckZPCBneUG0+zqzxLLYpn7VBk
T4gCdxtrB84vXYgcgCtmWDPltgv1bGUHZPEQSWRQmJmaL5Elsi2vPCeNOy/+Nfedunr5+CAQe21r
LkRY7RF+O9lEk1NMbIbVd7aI/k4m/SOwJNjpymka/GXBDOFucYEIh24Ir/nWDUYXoAaGFEj6J4wH
loCf7AOSjXvpjkmhtqIBSiHHWuATjSI4LKf6x7IosiocBTVmWm97yDBjGUYPyO/Fa88HhBBwajYM
yOyN5BkLdqE1IK6h7cRwQ5oOOG9GWflpWJbz1z1hmUjNZNpexVOQTpo9ph7LylwR6A+4d+546eD3
Qzgros5taelVN1v/y9wUerb1qy6OeYS3Tpn19zAmvAbf6Yr1yTTShtDp3NrOtwmnOrIV/1Ze4FG5
zleEbl2+NvHn2cBMjblGhv7hYlmmb5DErrU4/ms1kCM9tnKbOp4tUj/8Dlzg8Qq3hDnsbmWcRKRm
4QTRaTkQpFspLr/+0qSJHhNsmQGh+HamAESl9iEHXYUE2bqrj7sPOQFdjr1Q2ZHqgJMBa4HErLIF
a5PwU/Lb3zyfN2ACBTr/IkBd/xQ3RWkZcttx56Rr+TYFoHK+9XvdwAmdoJ08c1J8tloMJDaE+71u
mIS4WC/Dr6DnfSXv9T7xyCAc/QrANBbZBvDpde/TEdcazL4J65q4BJEr2pQrhj9rPmVL3rBPYuzx
XpGigzpROejGhfjQG5Gbd+39kni7A9YpGifCsGrZAuMn/6fVfjnDTKpPrZxlm5R45dP4Dk05mlM1
kweP8h1jwgstV6Hcwce+BGC33+hW2mAZ9/HWETLy+CK+1ycx5fn4MQspdl5sT6rccD6IQKJEdZKy
9jy1Y/eoo42VhdrADGnUrPmXT+HuRTHOUmxR5QNb64UPFmr7RC8ytgLwN4oOVxS6gM/xrQ44a+Ss
tRk5NlW8jM7SIwqFEojn33l4uG8kxkGo2zF5RBIa5WMG6kiYVjYksLPgZaquLVUDwjJkoyUJpHGv
k1xHTjipFX0Q2ZFodxcfJrr4zB8owBeVUe8uf1zFUkb4owZF8fICYmw8jyj4CYaM3nvoW6l7pNJ9
f8fZ3jZe8bMZ3Csa7/v568ate899QVXBtt0NPECzVHp2kU9clB8SJmDD4fWIfsrykbFAbUGhRIOS
spZDiRx7G+2S7Wfsrgqotr6va9Ym83XxNOr51PiyP4MGI0k+puF0D1aFTODFcwsywJBIOu+1OEDu
p/J+VtTmrtNRJMJso37gqLkQWsh4jK07t8VvIS7A/tFYnUdZHrrcfPnaCFA+n6oqoPMqB0aKjrQL
sOLXdcRzJbGHOVIlJMb7LZZ4BAFKEUA3mRv3IdgoMAqm+yy0apdOsw3gZ/Dzu+9igGR9A4PS83e9
wA9LKqBUISve1k3zGPIIh4i8+lkCPkYEx4ZyWKgIgDgKK1vruFVR/bOpOf6W//8/IEYHCj0MkJFH
OcP8X37jB/tkcUuIb7ppzDt9Ayy+scL4akPaFHSYB70S3cDCgff+4blDIOnA0TNLU4LRnzQLXdQf
dfZrZjmtQ2VejyuNNMrV6QF98OtMahdjz8qSbJUVoVhg6VQaVJSmIu3fLx4bG0nI151AxJ9Q+H9U
MP6itZahUhYBRUsGinclM7NALA5bdS2M7J2qm9BB/jdw5qpmlJR82YNxWy5k9wrliTy7MIEywcAN
pGu4MjLkjObpe240IDggehXDFypWPe/K8xEUMiIMr4N4QEPgF8hLfUEB+6xTnKXY4v15qM5IBc5w
becjzpg0Ci+1O/ExVx2+rM1ZGlpfSuVFGMk3jR9i0QrkXGdWU7RCZJxv1QxblsIljAfLPW/l89SL
FEVtjOk/24xgOx3MYZRjFfqQjALMSuA4rBALxZvVPivL4QcyMoywsvbYq9UOkiRAR2KJbxP2WWKw
3R8eIczE8Kht4Gu66M34loSB1TA8GWgVhEctSNrTzGDVwOMMQje8cAZnTif1rWU+sDcQA1aeFPr7
e7oiOv9KkNUsRhQvO7nOKpGEvqubpYE77DaZAI/cMS6+QK0F3k/K3uqQX5YUGf9ZhYxJuPZIpBUw
0V7TWm6r64O5ZjB72ZePbiuS2S+Pa+FIHUB6iox3RmNIbIirvBRo6SzbjQ1HJWs5fjJgegDwG4XP
oXcItTzdc9GUVrlEKqW4Qm707vs7uyN5E+3CwxrCo/gUdnt7OpM/w41oJZeA+eDaj6CQ7ZqQb8No
Wrng0mSd09hb2mVasKwMLG9wi7vUdFCNoIekwSkaLcW53V7SoM87/cRB6IgxtQspgAZoDE/RaX+k
ASFBjYUJgpPL9/a2g2b/9TyU4kbn88xeDDdWsIGeE3eKPzLWU0sAqEdtxGDsDep6nwIf0S5wxTuL
y4jmA7JLCtnRjAWjXz7u6+J8DAlZmcGKTonE3R+UApFmKnMPj3GmWjk6CORrzHKtkCrWbfR7WBmv
PZNOvpr2miZf9GK4YI+KNcfNBmtw+rOdD/vgjUZvamf9k7FhF66uq7V6xJqGWilNSpoc/CqzVhN3
WnCYBZ8HQNEJhPEMNFrOPlTUINvHtB23kkBdRo61hiTzq7q4rGLiL9H57QYmOFYTZYCkE7Eu/YsX
ESl6vr3VKgd6Cg7U2TMzsg3jTy8p4NnJZ6Z3cLW5I162e/n/7hw0CKNBZq13DWyrDd+WZ/1il4OG
v2PnaupDY4els9OIw3xPpO1JX2UVIuHeZfSx+8UanRFMMabaT8GAQd8Mlvdfo8LZ58PeOAjg4Hjk
MWRLv35GKJwd/4CuTsKoUx2J9VCGI+l9Cfi3+9KIf9KdHXaAvtW0NGsGf/w1tJOkOEZSGGjYPlzn
js6WzDt3ZsIPPJbEOYcKEc5YY/DklZ5ow7QdHm1YlGE8h3yUs1MYICDRbu2myRuEYy7O43TQqY0E
3SGl8dPbD/jL9X05fKb2vsAENgRSChGuBITpnYsmOyyWgMmqD1kg4aboeqaWXMYJHJ5Dhutu80Bv
XoWfWyNSqqVb6Ee1ovusQuBrZe35Pp4MhWUxohhdA25C5c2lsFDKtDiAcP/xwzHy65hYEOIQOuTK
fNsLsLc1GoIi83NUSgG+3S9AJ9rTZ0xNuvzke1Cv80S2Xo9anP3mjwYOPxN5yGR8a+6pPpsPb3Mj
Idy4O1HG0Fn2c1qJwl1taaXVqU5eK/JOQpDqNx/0PqS0rH4NvciEyleIyhRP/ab+YQPtuUKL0Fdo
HXB/FMB4FJvfcmLwFX5gRC0lqUkyadI57Gy/z/HYIMc7BgdPM38YmeGuUzplSwAKjnT/wSKhP6aP
4R83qQKBYihihvA8zHck1RDWOUk+N3J1rpZDhx7LMk2MUU9o4aSt3nEq9/u4uuPjkzgOagoiMyBs
kYDwcf1EHINqWxZNFmSrYxqZ84BeTsMDr6ASQG6dbGTD5GeOiWzd8S4UXQ0RgUiW/DtHfW6V/VeA
hQZ78xK/NslVQP75WPLudJ+slczfpd+H7GtGMQ2enxTrr+FICPkeEvAGMkFRp2EyGY9w2QvO8COq
s/fK79mH9XkGlLZ6QVCuW9aBwfpSBwaXFHDdyotyClkY1743olKFrBjYfrHFkcAiFmePg2ty6gbk
SvCyIQ8N+dzsvK4B+Wy6ihR1E7T9Z455/S121XhttZGGeU548l7tCGzKGavem5UtQhSDhi2eNAQS
SAxRU6SjIBW8eDP1FMaI5cTXY4qEbDWGFuDeEyDsvfgbvQczH/H0ZyouriqzRFKSm4bhAzs5t+F9
+RmfB87l2lbhWFqM/NYuAPzJQ9zgDZS9KVurA8Ms0ENoIfJz03iqvnsxOM5HrjoC2cGv01U/oWSU
9d5Eew3VfudN3gnHC3uSFTsGdoqh/VAqy1bcxcRFYfrkoQgpNQrMux8efsruVZa4rdhov37s7Vuy
pUQqpWMiyoatwbeSioa7c9WelDqC8P7DVIoxRzDuT8rK74xkdFCoFNMU0M9eKyeHntkDsuvvd925
goEMwHmQNnzsgyWvPqDVUulgJF41XMBeQWLc28aX8KEbkdDR4uncf1jcz881soFdW1ccl6aRhEeh
RGnJW5sUUapw7GV36SeWv9p9pSmYxTeZxMpD+IECZsXuOFI80r8elakzJ1IHRWUMCm3EprZyjS60
s9Tg2fN4fc/VgLgCtsoBLV6Y9z8psrmrY2FTObrrP4gXfhEHqwWKM6IQvdfrYtV31gx+2iSkakzo
Vx/Jm80zkpi/AMteGKErAMl2UKwKdj9ILi7Zo0cDhwn2BXTdMRbY1qhBVwP4qSPZAVXewCqOh6yj
9qVWrjDD5pnnuK6h0iJ0mmgPtpWHD51EkfReR2Dz+Uc36zFET6sqXNHDobdDY6IQ994w6bdlcT5H
uVIgkBscNQK7oUotSCsdYQG6qgP9RptvFZaywO7k57xhUrEoTq5RxJtRDKE0UQ69sLSoxnAfMr8V
XbRcgc/GFuid9bxBaoAM89plnjX2GWXNLn6LgMG1WSsbOewnTeApi5LLqIbnDgggI01bbkWQekrj
73sC1X2tjX8De+5zlZX39M7ToN3TSQgzNd3xPALWvud65uDU/Ch8j4ufruyzkZeeWkUTFhiMuPKi
3fHS5kKURQlTOGO2W+4XhkBQgiiJSlZrThZ+Zv9+ykGRj3zr2ZQmLCFk3RCizCNwLsyPJm7x17Nf
dMOgf1pobDcRlL3mgQR/kJItwcMrJu0X3zFpiOfWBYgfe8vH37t0mkGRiJWG0OusBGQ4A2W1wnnX
Y5oTojkTgzo8jbPR6ho/vj//HwIsP/1+Iu2B6QjP5YL7fzS897hSjwQCoTxY15Pat5wd9z20mog4
sI86p6hxi9A7VA0CshonqIey7/FlR5tUILO1YV7pnN9hIEGxVPGTYLkHtGgfukMvVb0v/enlgDx5
WKzdUby3BiObj6/3z9LWTd8j9fujFKoFj53iAtAuEY5XirMVxHlRrKlDnbPI5/yBbTJqyztwWKOg
xcpTbw1Ft7Lj61JnHAJlrfStslNRXLcKzkRj1mhsCtZDVXTQpJKnqhe8eTcQGHp8ZM+ILb7Lp+vv
F4ao791XgPBbklxs1/00IwJakbYBHB5JUFrGopPsGDaGGwUyMGe/7LFTYA7ZWdf0N4VoCCy+1mD4
+TmJ3CdWmGzQIy29G6XZcvEUIyPlMz8zwHGaWwqm8mj11B0YEG+RZqExqkqibj4nr5AtiJ8Ol2ca
JF5XAcYN71u8nNIfIZlCFOz6egxpUZfspYGXgs9xcPr3BTcZgn1+kw93T5uY4MEbt96mzHhg0j6A
YwzSw0n80Dt0zt6hGYatv9y2aVYissOrWyYasOU5UH3Ups7ROzm4kgXuHCJffs51oFoq6F0e017e
PnZmbHxVDjY9KElBY/pB0Ymk+fNSq/urPKxw/cbMx/ypOrYr/fSJgRbpKeV2iFfvUg4xai6HWSgI
/n5xko8VdroNNmPeQd6u0e+FrQZJIqg1uZavsRns0xaLJ7AUTg/Hqa/ic8mwGwzU7spPzKNdT0ue
uH5WH1BXn/LZYGHkNP12PdmPHth6LM5RcHwzDMVIk4qQmQRMo/LBF5K+n4A/gl54kCxKMf6SfbDE
3S2cqC8qJ75U5udmSx78EF93TLwmVWD68ROpGWKatchMrleMWNbQ3tA/OvXFo+jh99RaNSudeoTe
jYUdzJDqIraXApF+2zx85Hhjkk1PEaGJRplXHL9gcJeQ3pkHHNQD0SpWmwHr5MgtqSEsFb1k8WV0
9jgJZGvztcQSSIKg9wXvrBO5LF+cWGZWm8wceVD+N+h7h7OqXpDMVlf/clXJMTPMV3MtrR+Ech62
dXy2oL33OLV/S62U3IzXXjVMKq8PC8BgHnkhqaW4IlfDsj7IiGxJpHJqr+t2+iuVt9ue5XYLpa8Y
04veeYf1ExbG4p7s1+u0O+9ZYvgt6zKeSYWocMY/iFgg/Dvz8QxzEbciLPSiZDArPmUJsAizVeFQ
Sj0gG07B6Ho9eapr8Z48JH4NQZQyTiR3piuBQpQXkpyg1sUW0a2scW/A/D9PLLjsbFVa2IlXs3Tl
zu/2uURMNk32D9mlMwgjwQnneWdQIYGFVeufTqSjbP7a164z3H4r+266M4afMzm3mANNpPy21QRO
5j5QdbGKx8ytGrFeuVVYH7zQkvYISkjJHLJhXid94gzJPegJFIpd2W83hgrTNopi5PjkcRT512l1
2YxJE0SygANqbBi/ZaMwXZmyU+GWD3HzTU8Z6WZFz91bR8CI9aT6NHtr73qEtaEtyv+N+pROYb2w
I105EB07b9W7EAlejYcVllm3F56i+DNDPRyPtDdJVJI6ykayfaZchPKwwKyB424S5/cASLI3DTRg
+K4imYKD3cZYEMb+X4slB8mRpO1fafCOkXkf8Cx/IcbghA4jki5UpljEyHWAYAsuHpSXBJVMVbVl
BUyK+6fn2NjAgRQz65DMVB/LmnPonCUmKPdjGKNDVAX+UA55AooYstgZOo3fPw72uBf38uvqZlQC
b+jFIH51Yyzoth8gNW/Z+skNNMB08y1xf5lchSLR3+KH2qiUg/iq8gMjbgNqateJ8FNDSmwWU+2i
Gl/jJYmx8/iDogcRRJuR5yFcUYswYpzbfFeysGFmTL3FfTQ0Wc40dlkXRnC+PWuug/dINCnoRyrc
509qKm8E2LmcPSJ0F08W/W9aSuCqstatDF6/clv1eBG6kZ+ZvUjrpQMf/3ZW86kPjEk0iS+mbDCm
+iAniQHWsry9IdaLhzJnuLwEAN2//txWKgMObDN1zW7Whw4GrlRbWu5A2J+nAwxmSCfroGj64oBg
ifQT1xWceP5+OvlK955BMHssvnUks0DVe2FhsvO4AWNqDBnA7MyMzA42nngWI75HHBHX0x9qcnuC
UfXxsJwwDQbOCa2PxswBRGZO9AWptgVB4qp+aCl9kdLhN8DGtjVen0KzNTsHIwjnZYU234pX2wnk
osiDLNawvlu1TJX1oD+k1d0mWW7/iUdVloWIKU2B3rAbwJSp5K3l5BsDp4RNEYxtFfOwsK5RV75/
t4Qyr5LPQbSapneim2ohzyiRfuufh8q+bSFYmh305c8T9TLVPnP+80sM39JbE+egdFOLOiCtZhGR
EvdiFrZ1aVc6DD//n2SBb2uCbiSUg6wRXynI4szLRLhkUGhXKL7m/32L5OkNrPruYRSokkrUHddA
wOfdz1FYjmopiAb+/MZBBvHfJc1WseuKFTuxsCSG/GD68Hucng+/NcbyOsx5FRbvi10l8kVissEg
x7tBqFhGxbD3TJuVBBIZNR0d+8b0y02KiRrU9Wf5fiCE2PxHRpwROR4xXuwcmett6hDK/R3IsDzI
FpNs2TpUxrr5CV9ajFpD5zkxkGEEkrkx8DClQGNiWkkcNQs5p9+BBGQTY2XGldTnGRm0BJbfdaYl
ZtktX0eWQYI4dR3CinvgaITa6y9v+u1KCTYHnlbng9ib84iJ2vtLqrbzBSrIxBgiX1CXCTsmBNA9
6b6v9rgs7fuVqVHrG6d+U3g3t24LB1mLVlTwTyCsPndPTAk/CXoTaiU6A596w1HCj/UVgNTave1m
pTfKPVBwTcDRiRA4DvfnHOJwmnaSlCzG/6mj5ZB56u4GzsSaKlXgXw+WR3jzHVkghOYFgJtPqDp3
jlPmjGbq3MNRATOoPSSTTHNXYLZPMfcPMU89PjXUZy38j+uCePfT3g2P2vyAlQ4USVgnX1Yi7OaY
70T78LEXl+32C1z9dJOQOZI6b1hR+cTXF/+H//QBVROgMrmRlEOb44xTuMxNmqAUT676R6uczoZL
z6phpM5CllVrN8SDyrXTcfUCy6T3NQwJ0fx9FQyVPWwK8dGgcoByGe4cH41PS2IKoDOvlvmpoMsQ
dU2EZaYG+ePdCMbYOU0pvXq74fsOwGbWxRLBG91oDIVa9QDBf3KdQFpEn++HEgDnSArwOtrQ/s/M
jQhNoVvnQUIRMJcPKP8XL5A08kQJqfcC0IMZztsVHtcMIHPu8X/G6zBJV98Jc7HOGFaDUMtVg6ko
RgL5nSVdr1VE+KfsOh8nR5pB4+wmFDKtjVd0ywRXWkKD57G4PrTqLn35ONgJAqFse6ederRtqk3u
LBjiwfuYS/xK8I1exXrcEkUTmnjgzIo9KK98xWSDQnnWxXt2YlUufEMoC7U19UpTn5ZWi/Rttg9r
+GqaBKSrR5+Rrjz987At/dl2gmmfqXICa/ukAigRS3vK1qkO2NkS0vqX33C1z2YzS1qP0WaPr4Tv
1fNh+9QUcZ1Z8v00criyq1RLjXIQKzI0yEdlb1Yij1cXV1feA16McpJRtTvbVsG7fhiaArH6Jq6H
YiJWJFe/rOC0rR4LZHIQZ0Afuj3zFda0O/qQZtLsOFMuyqG98CD8gtbINRYOixZJ/LeZxZuaLxdR
JbuL/SgI8oxt7DOQIlGl4NIax7gYxBq/vhisSWqr2PIcj+QOy8hDBUBFEbkPTfJ3XqU7E+DuEQ+J
L+U//dDlf+NxfnbtKyl5P44U0yvH0PRxFAfRCkWq7Av5FlpJ86YidpUFt3U0+BnCnu4cu7Fddcd+
xEqG8xHk1nJtbqf6ptuh2Sum1djRL36G3lLbQGLPF6UZBVc+hP6BKXMQ4gITRbJaleKudhCqYnsp
FO/R6KrrqthBYSHxbWH2+i0ZrTN0uYXp/+TfTZR8uN1E3C/RV5uQDuSpmpC6LNl3cJKlA9NNAAEZ
LvUq5ko+NbHDTj19Cc56H1CW8oldk6NX3F9WBa7wotKKLS1dSgQH/Ywv8SyXL0pIbOSjwjmeU/KU
flbZJzH8qwGv7kS3tXEz+ukoYropB+SWHZvswbH84YWTKJP7Zy8d7jhl/6fFO4Dgh55xrRgS+txG
Qw1b8Pr0u7fsT0UeOmsAFnlIyBd2+Uq+CJodDVr15HQSJAAWUwhy9gLyKOpGytBUJCTDKsjUqawB
3FzF5ZcLPdg/JsnwxjRDsCzA40FOf2bHomvpKRoXxnN03DG4DjUtFWShV+AeWLoi6BnnpKKZ3cz6
UDOlw7gV/9YQDQdyuLg7tjoiKJrZNlkbJNbUOnPOLtFhZoAxbmwFwl3pcjx407uL3ILh1u74iwMp
6mcCabscuh+DAD2dC9ueRsbDaktoD0o8OZVG0ECVLIB3O2Ri3hk5r9arwL+REprsVqj2jeDLJBD0
MeBHsh9gO6w0/87Zz4/tiExGBpj+jjwu5WlJhU90zpr3V8mx3ZOksClZTmlwf5m5huqOwVdcTc7N
dDgMRO6lN8uulNF8r6EVq5/YHggUTf953NsW1dVwyhzsA2v+BqYmwwh4p/2DmNOniNrZJJ4wC9M2
W+Lk2iLKFthNUzXaWiSh4yU0ZTHJ2OuNshE5uc8HGcYyhL/yreE5a1YbgeeIfTHj3d+MpJrcFWbV
IbK81EXO8PQOS+LTNdvfO4UvVsV/2ga6sSWNaQFWiWzGA5TumsA00p9zNGhS38cWyRFU1tV2WOue
MjrWPz4seRaIX74EKeQpNSZzvsLqT3udSuMHmQxH9P4RotWIzhqibgIcK7/N0O92ukmSRP8cmsXb
KlgyzHh0f55ZcLl4gr/nmEAWfQgYat9gtnh2pMvzWGiTXv7KSj4FkngmSxwqN8/b16/cvR7gAGfG
kEdUTh8WWnCjhu9xQb5iHUC21C4QcLMtT6FmDPQtmPh1u6xg1kAelOvWN9c8MRLHxTwnsgiL2wTS
FxC3HbhRJUp/oSIjIQ1tCU7Rq3A4l61kgDxtArEHYhlS1Ow8k67y8sgdkt1MIU8Nha4lpTIQjvEh
4AOUZ2U+iUfWszJM0W3WCsGUvr6O2VKVWti11y+/rOduBSIKQTpIBVQ5KkDf6tYfvwnBzmbjWMYA
SkS0jqBzz9d5tof5ZhK/c/oeJh+6jTCBefarIVtheXlwEaIyqbGq6W96E4aVB7OOivqk43N4KLej
rbX9KfR1Hxce+33TlUiWhvC2qH4zVOoYH6Iw+Wp5Hpcm87J5pcYoCmJo4jrxzhldZX5l147bZRzC
cNfx6l9dEYO6sMpq0z+6rk9dTIMVRJT1NF5ygd8UDL6/IWImN708DKZ/8Sch9LOATW+2zYc4/fz8
n/XacvCP5xd/hfb6ivq9CqGra4nQUFKPU+lEvadPxolukb0Wx3GPFiaZHuLUSk/Hv6GHBAno7Hbs
PRLxcSDauNirxvPUNfVq6mmHlSaNH1SzToO854oasFSVnmYbwzDIxZ99EPvXbn26V1EqvnUkyyVB
5hzlksUS0EmpxJj9povFa5G6fadyMAKfBkP1GrG5YXU+q9L16Z1VxFSNTPDtAalgY4HtkVsxu4GE
dwN98u7GIO1SZf2gJhhCrSnoccUOQDLIOu1i7Zn7FGrCbktHvw5qs6LX0nhLmYDvM/HgCVIW+zhc
448cF1z+3OXAXARJPZfgg6CmFSnxJc63T0MYiXqLtpb2z4IJP6QLn1E46Vexp9HICP/MFWnbdk9G
0HgQwjQinAHsga2AB4RIwTMm9/nkZv/olCauz/k7rBnI2swcLd0cSmMonKW/AT6c8VRZdUL4Z4uq
eKbV4x7mT0R7JYHQczMhN+M5FEYq7eTYNTuCLVgMKDJahFoEpvPfQPPXEWvdnpFH1gX+fQHiht3E
qrRHUx4mNvWZ00lTMu/WiX+mE+UeRUtHllXsAVCxN7jDTa4Sc65VQY57AXnLNHlAI6050m/3p0EG
/SvM83KclFQS1kb34vjJOkG62vGRX0rM6tUTXc35M6IX750McEdmDmtVugIW1rqndDp1DpgjqDKl
iut0Zod1K7IazVJIRbiOESfQ63blo0FTAelGnth4zOIiZ4U3a0NV+wJvFLRdXyoylJp8q/VWltsr
qUYFWSHCkAlteaYC+FekabEGbbvVgbWia/wEprG+UB1JtngHgSvEzDORy1d9JDsMwLfHMTU5wpLG
YEoAWZMZhDk+a62593CJy1ZsKcFHXhc1uzRrhkVCkP07opoSgWgn3Mdi6uqaAknmSheKd0+tlbNE
lKfV9Sz6C5ZHnOCwmcHZ8WapxKfj8MT/slnrinNyPDBMNt7S9BqrIt8X3y1UkNnHYuf3vXa6JGIN
E9eeHIA6n+adi7dGUiEnb75eGtkYxfApanuYKLNU0cQBH485gkrtXb30Rvx8dkYosmxWM6VRZR3C
NUVz/25QAMGYu3PoKxjM2UwkhCupQWziq2FlveOfMuaroWNwSfoEmeo0O5Bnkz4C26W/g/dtznlR
E4p2HMsFIeToEZg+u3mHWa8i4LpItbciB3Q4RtFKU6EGn4sy8Xz2dKerz80UM+29wF9TDUzVGMsY
fm+cKSz+JwkV/KADenxxM5iIsZ5AHq7PoPhEEmFq1MoLvBEYjslbfBZlOolYt2BaGl8OPoPbjJOD
V4X2/NsQkJJapXEZD6oyK9+ONWPcD5YYnoOlsLF/Frzg02lqt6rNgOxbs0swI31Cc2MxRlBkebbQ
t5qZlceTKknVJkZy6h3MNg1JLezW+zYfLuhYaATmGgxyNwXlgQTjeEcDf4B7XEN0sHrHuXO/w8l0
tM6Atfs8aGpNEEqzRr06SzZqC9D3S6v65/cy+IWlJc4P/lUWmzNv2uRrvzrTp3+et4GJMrqONo7B
Em5dTcC8s8Fk9aqxPDYGExbYjd+I1KEgTcIK3ug1ctAs8sbnBrf5mrXzBB25eJBCpfAJFI3Ho7PH
lFxmwLqpod1xQhu4ExOyC02m/ORYOLNnzVsLbO6KAn+cre56iZoF6sMsX55IVhFb7oI/SsVBAfTd
0/XOelhRW/3ErxUv6ooqgOrJnqoTfMAzUSSSmzw8p2JMM9D7soYLn2sAJievqKk/8E3DEXOLov4E
tNrOBH58AJG+M7lMXHkS2hcr4kNuvqlxRLA9Srbx857x5IOOZ7KIdkhkPizRR9PFHmi0p4MI7Njz
2/yqxM+501lo+jWxA0r+pUxSjcB0JpsITb08nzg23i3sGKpYKRYI14GWePuHoUKQMjIMHrns3VJH
oxGpMCpUbcyP2LdrHrIgafrgLGQcCOPiQTPIHamUDmzSkg6zFnxaChNVxJxtqzXv5Kbj89crCsV4
MImlKa0dE3nsm6z7klsgqqfX69fGcP/80KIgLZAV2QDDok4fb0+ITqdAtlgY7+hrhkdts0O9SUnR
9TvHzGcmqKvAKNUD6x2GjproKRYdZJUWPxziwszUVkOKLGLRuIHDntKgXe47hvJZr2wYnWNbABcm
aPOY+FoAVCXfgiUMeSIDlPke0n8Z29fzXh5JmJ7C4WTLGSQzGPNvZruGFvWQf4KhbdQCsYNYXgep
IpowNCE2WDcDUAdllgOCqVSY0BwCKAxcgaeJRBDI20x9b2nt1eyfb9fG5JWc3KSjNuYkJ5B9/iOS
6Auwb7fF9ogKqUGhM32P+8CzpneuUe4hiP4RC/6l82p8h2DXPV/EIP9D5CL0wkU/fbDNMgvaGLrI
JVU313IHYdMwmHPwn9DIqDNQF7YTOi02woU+i37NUoanoRysZln2BEup7rssCXKWb5Egh5NmgeGD
NgF1T5p+wQiJpizCcrASrL35rmmq5eFxN+puuQJ5szi8GeNB/whrqsv8kWRvMcPdLEwrJZNuayii
e/tN4MH1MLrFdxxfY8aXltVg3sQf2cNZo8ZRImoxXVK1pR75A0JZt/dh3CGfLHux8fCBZDLpVkyj
SjiiY9b6fsBShIQCfUtLf+r8ExGhVi9hBAvuX6+4Tj0PL6HbcOPIDzO+UVO1C55Ug+M3d88RK2xF
+0Z1CZSg7RYD3jqfiuWBeGMZ4rezz1E6+bPvlxgYJS97kTjeouuR+agfvWPbCAPj9iWNYJCtSobS
cMzXeLTKFWHMKKQxONOgwQSVxif9Kdpva3Oy+IWRvyIZ47D6IyDo2s0+qnIFroa2KD0Fh9m5umSk
gHUsfkjxDk9pLXqmrlyTbp/9cljX0S4W9BLmodGNtMGXg98WgPgJv01dASl9Cj2SgbR3ze5zNnsN
PjbMxcOVdWfjGbMc1cigzWxdXl/nsUIwAUEfDiTT4ATONRsaxPZT2gEwke8jz88BfcSqNyVoLJpn
HQJMMpx7P3SM6XuoIu1Eqj+vDV/3HQ3hbTMv8HstTYDO985hUkEJuiqs2dPQLq/Ij4HwbNWCurq6
bcRM6JPm0ZwLR7/BxDCiX31cz7QWMQnbj7C05m317tSelAcBzJQufOWRf8441m163mOblFhK9VYJ
QX6bxwdLvr/v+IrorjpbwZ2CwYPZMArEKF3TmOGkKM6nELfIvZzk/4qSU1Ckmk1JFv1uuBbSHRLi
EkbObJCFSdPlb+9jVupCfw8o4feTw+UvvVYTaNZJYWAKsq0aepF6lhgMWg6ppmB/xY8jfLY9FL5F
YfUjgQnpbpJHp2/94LtLKAqjPs4N1uQC48RgIjJPUmI+e29BVYvLW7jgoNuMXjCeqlocGtk8hxCN
U+V11vk5NU1mU5ScvicBzkvqP6zNc9P3OWNTBhySG05j5/iYH7Xm0kzj1dzDV3fpQYAQ1A+NiHqw
ZSz0RkodBmSPsJJzhO6WEKxqH5Ett/uqqaldyGpVrNXXif6q2K9D4KA11x87B3neD0EpBCGYexsL
0SH6MEU40kugVWIYvYgAZrCNAy60rTiAGBHMUHFfIbZhG5IOA6+2iGhEnLIR5pFhyrxdLRc0ua9o
Q/75JsXVksN8BKoC4PIhS6IVYw6Rejyb3ZoGlfy6qywogVBNK776dZAEsjzdqsgkkyGW9O2pXD3I
vFQ2VNG+/lMG5YOCdFG8D8asgOkPHFkMGaIS2LLBfMfnl8nh35E/zdOChUObuvzV/tgsj5E8+8ir
fib0h4uw8Wg9TYGhNc1PlHDp/N1kDSu6CktensAuHBm0y75p+gJqzmMwq96OytjFs2iBoLE1WfGN
AmxRtjimdzNRnW8s8JPGYc6+NWQxwhQw4GaYMdplZ1G+OdHimxPR5igjomUa1MZUAgrb4LpD/pmj
be5Wt0JuErITMrSIvauXeOoLV/M4q2BTkiQ72g9F4E27M79pbiont7nSFUUVhkDdATT+C4jWwzvh
LUf/QyP6aG3xlD9kmfWz3oryrMXsG3RYVi7ocBegWcCRyxkfQKlMfF6W1uRibkiMoa51T6AADJK3
y5EIBTHlFflIdDjjpHVITVfg8BtJQFYrz3Io+Ve4/wEb0X0Voqp0UhS0o0ubw5fei5kt2zYyPtu7
aXvVuy0Vd+fJ0r/5MZOSIE5rcspbWLfzM6ImuJoQvzidL1UO3Nc2Hk1x3EPCmC2UOZhTlQPIp6Dd
NcLID5rp+YRHoA9wSN54Bgo22u/8YmPx0JTlC801nVbbKG1+nEbH/0olqOCkxa1ThALllFOXctGf
GAPjHJfBpW3YUI39rCfbsuLth4RRjdhTl3nOI681UqdQPitCXs2IV7riX+PpCyxUtl68jOKwrlTO
TAnGj8mF41HmkjuOpSEwxHo11bDQqSui2UfPunqq9TIxx5iEVII4v0SB4gB1NjJMUVCaAYyzdWSu
w1imGriEkqqFdj6lDKHDEqzwcdvNVRoBQnIoiPKuyWCnjH+ayoyPFKrue22zgI+PQJ8Jiw50XH6l
nUDgHWHf6nkz3mOwZloTQJ6k+a1WZaarezuQ0I2slkrMjB+T8XV2VMRxxaiyjWn8PjXLwHurXzjl
cy7F0d1BCjphSaBl7TzOfzgQN8AhLxxP5vAaCL32p60na21skdsn81NWW+Qr2I8nbqQYNGj40YtE
0NYSQbrMle0QIBwSehusRCRvSD3+DkcmXza0Bi8rkyyRjqnBuqW0RFBdB0lLdvfxIJ7gq3O7jQaE
O85lQsTLvmlsoRLD7cbLOEHJ/E65Av4hD/qCvyx6rbc5XZK8vK6ZwEZZ3GPFJfNhLBX9UDIlIu2Z
YEXtOdGdIo8ohzKj3S0NifA3THt6WucYlZbzqcYSpj6lFbwRo6aImp4eAgPisNScUxeak2+K8lJh
86sYZTM+xzfFDYOO6TPECbqe20cLXPr0Kp9Tjj4qemvaoP0Slo1xwd1d6VpI2iAgD/DTPAd3yrpc
DkU08OsfRfeIZVPGHvj6hmVoloEIhGYCjSv5oH9ikXVS914hGTzeG1N9MyI2GqKLMIiYNFqG/zsY
5feAY6depQMADZPytwYkQbWGwEPoE6E9W8w8ScZc0a0uph7hN2XRHiZaG+LCzpTei0UGim0qfr+8
KxlJ3h4LLROmVco8t0P9MID9PejxacnIajAbvBkXUPjJzApkZKpPUOwra2MSFfQD66aDh7ISocV+
oaIku806bEfqwcpkdETbZnTc+ueoz3Uc2xoZXX0KsGk4J1MwXMkbp8QpixS2r4xYLlZLlwpjl1ox
2o+e6g8SMwDOTD6nOGEIMSbfjsjJIRA4Hz7Ou2FRnJ416+1FLO5ykyfBbD0J+B1xK1oE01rXQEuu
K8Jt1ansjKJ4eyZRXmp75CI54JUIF6bYf22l4whDB8qVTVCdl0W12L/0GYbRau7iPwV3Zz53b6Sn
89pbcogW1b5/LJW3V3gF5X3MqVHEDAsMKXCUiQ+IcnIJeV0nezMjMT2rR6w8tm61hSlPb33OZmof
flJ+c10D3UCFqqfXJdzpsSPM5EkWaLLkdJoLzZm165HZI6Byv6wiyDrOO2LvHExWsFBj3/Ryv45h
nhMymUINvl660yLQmWwri37lRRkP2cFEjUhXMiUSLChzyB+Vx3SBO8FiJMHPhGMOx6HkQPRaKp/O
+ibaa1SIbGuypLJTwmkjM2NsjB90mXXzq+yNXEXMDbRPgFq42cqfLE+82pYxhXWOdVaV7+Dd6Dt7
xlX8KQxchL09IjIeMVagVy9byQWJJYg7UIS3J9HRwba4P9xk+ZPVzNdf5slOj7KR+hEJQkPeqBUe
EJLtlyd9A7oqv/mmg5naeazWlFNt8NKBh3F3FzzPOl5WB2gcbJqGxYWrj/o+sROjIkktiYgZ4T7V
z4k1w4cnZw2vVmalKmOKRoHcUDIzAumJtoNMINvyubi3vESuQUWAqhfh/a4o6wxOZK70JhKtJZP7
7+T/1Cg/PtIQixcGZ6wUHxh+/1hmj9fuX3AIbVvKMhxNn0N2hj+hkiZ4ldFjVfVGXH9da80GnF8f
h9e8agMUlEUcwZWw912ALERlPQXoqLjIHKd3xYHVFtUd/XZ3ULdDFhBlnvuNH/NR8mCX8/bfvHJT
GmuuH+/qMv1qLVRIP7/Jx0IdHnrlEOvC6/eKY0eZbpmmX1McXWQguBIQrMyJ00+4XU5LCdGL0Fdx
T6xmXHddglL4DYOjBgHhXigqo7zX+vJcJJo/3LmlGaiMQBHJu1iqbSsxwRx97HV2KQjkYl0kH+o2
Y86NcDXi5TvotG7o08ArcFVZmRekvgSL+PQIxd7jbcf7VEVy7K3imW7AhuFDVBBylJx1oE69M+4y
dI+vQqaSuwEbKigAGhNJHNrwVTeQHLdC8ZxuauZW7WlWkpkzR1wtI4zpp5i9G6l5ke+s0fKKNKkL
N9b0ewPj9SzCEifm96y9EBpt4dYUwsE7xQ4j5Q9d9TIOOnXHJ1S5YaTjd8lrr5vepnhdZZQ5Zveo
DyxntBa3R9tXXb/u/r2/sdQF3tVI/LRm+whhMWJe2AcUfJgAMg4XvrYnyvLyCj0ipzv8xh3fZjhh
TVNVGuJ9lJ0x6w0Bj+6BJeWLUmui5z9Wf2U5y3PBI3+vrlKGiaZc53vclfX7zpbnmWx+Z01brdSH
dE/wyKsLIpXae99jSfoOkkTngj+hmu6024imSXkncsUuioVOqSnaNXEYbox7cYAQT6hsNtLYAvtL
0WfxvqhNpNZEHVzEYLgfqh5Hc6hp5lICeNFyqpUC5XNmi/MsgtlUk6vWaog1JDvG8czrjatv4iLs
RRN0oxmDxg7Aq9meqZWpp6NUD564hqEbMC3cur3I4tgx+5gv9O9QH85mknHKkJNyQ0PeVGukW71B
/diN2PXtT5cRN32tDCEmG/3oVnsUuf0Djwqeu3erz3kko+2vuT48rd6SiIpzZwS/u5hbnHH2MwnI
J3jk412zLbzvb1T8hRBPup4oh8MbUPxu3hzSvPb4TCWgUeeVe5xBA4D4TS4hdxONLKrSlikIWUxD
Tkl0ZQaef5guntKlhVxDGhpNx3kORBaGFhSp4AOcbulEAvNrOXCUaqXdqI82hpvpImhw9pXGcUce
EPN/MK+lOMhp732qsYHbTfepIKizb9A1s5Vc8y0dMPiI3359cwAfqcmgvF7DaAAZa6JogVynhMJn
T7T3O3/kYGjaWaOjDWe+A8WsDm7SzYqKMuV3pGvaPl/hF6/BDNAQRMwFX4FMFVk7x0A51nhcuMxk
6MJeT4UHLV3bWU/30XH+EGZ4c4bItBx7riq8QutMbeSDdDGpneTVezoEtIXGa5aSPAxNjJLNQVzV
+5JWHOINzAk4wlT3OW072eYSgWipnKYaJcuRFplCioAX4NgXP5Rt4hdVBL+oQrY3psYYvHybMGkY
Ji0+YjuSFgzfz0Zql7DwZ+q20QcbNzMaeYil1SN3kTXOsVNljTcw3AZwScAfMKM/B80jCRRKGb4C
tjSiCnaU2IC9JLEKyAOnZ1VruX/zGemvR201UNwkSHQezOGHljEiLD0XBpx5UIcTU/4Gr4ndhulj
TdVnDKBEtAngXqk0h1sNGwF9gwV6IAKgnnPEijvX/uKJ0o9N8US+ifx6rRTAF+JKGb2XIh8hG+N5
CJbpdFth/7FQCaGxIT2OL9+h9ZIG7oTWyVdsYh6a6v3qvbOKHoVewLkZo2UWozBmvsDYd0d/zcLr
F+Wm4lkfvd+dvzoYVp+k2rR+sglW1Z467nUNwr35gsFhltDRawKgNIfQ491elMSmp5flq+3dIL/3
pMLF05neD2MszabPSnJOJXKGEYngxq3jRFhw4auf2bBGkqMwBiK1bhoT8Qw1AoIZp+BaOnDd8Dpv
sx87mT7sBdnwv5P8Wu32XzR0Msi8Pa6mxrn1ptLn8qdqxaAQNick6+wBSYHuIs1YlXv82xTVo4Em
czm04xDdbUelhVGD6q8MzdY0wEUwwZIiCxLD5abpXjyESeBzIYFIf0E5sf+b34NFlBnUfIk3eNhK
C8/cgKKe6J2VINTuW78Vc3xB4vXnQ6CMu1lwI9lkaMtUWqsdHIxijwGvhgfWulZ6kV4CfFmqWyfZ
gvq3QMbSKym5S1kiQiSXv3fCgksJacJiMvX5kByok4Xv2fcrTkhfL2z90ej5kJtklH9F/ljLF9dj
e612NZpRiqbc2MPt2W3xygNRJUQSsiRAoLTBUTyblTOe10LCfnn02kxOcjR3TOvKJRGddGoxfz5a
d+UjCZfigl9BndkJW/lu/kf1rmMVMa1oh9MY0nphEwV0wEdDcLanGXEL7sL+aQkvtjyYAKx3hvck
djWLo4eHHUt0NEhMWBMCtQjhfjGIS4J9aivfidbvlekBqeENCJjwS94AKjQpMnZQkT+98rPVmNTg
rgXjf/3Y6twO34ILpDgxDbWbNKhE/9Vl+JZ+jhXpZGWQY22fzfU/fRNSQJqy7Rqxl9wIVXp3HyRf
IvVvNyi0qWrHdSj2n0YF9iiJSDvzLtz3tDKvMBgie/49ViNhAkZ19p2LA+GjSApuGEmcstFOmZ1V
cYt5kJzV3MPgfLAs+FDshyd3oQq2CYxRhCep1FWQog/voFnG/K8pli3fjF8sZiMoSZyEaIelPSIv
DiSTSGnY+Dwia54MgAfWjP7aG9NJRN96UTAw4vdB+mk/TJlRT3fJlG+bT4O4cd/qHgshcjjoDLY5
oEj8MTd5LHbGgKzhLS4alMowg9VSGuvfE94Mf0CojOZgXKMgaz9DMeFYyZ8vBnfPDsloeEoE2YGx
jSefwMv/YwyotK8erV2A0230ieykifE0SmcDBDu0RpRCIoPIaGf0GWHZLO5EaMQpYVZDIETOCO+C
8RiNgv6xKhPZXIsujJpfpF9BkL+4j2nTwOxZ8nC+rpOB/OvY7eLyJBn+yv8KmdZEiuSfhlyv2hQt
aa0JDQ426eVkCKcgJCc9QOsgyFavWrj++4xM3yiIjiD82mNFEz0Yv84v77E4DcJA4eeS+fz5vcfM
5G79Bz/G+d/TUBilfr3pubbNTpoumHukJSGrhQWqLSGAbzk4cYCPcu6WTnCVv8Xj8lbMcjCwRMB+
9H+JV98tTcF1RZjDb3AOQ3rFzLXTpYMCLoyRRDbiVxHIb/nzGG/pmNk0gUpry1DM+uraNHmolY76
CyndxVffzbgSvdOmQuXut0wNH0C5M30nnw2nI81m7aLr+QdeyNoUkTSVe+u/Nt3S8LkUPQSXys4J
SUs3cqtGkfM5PY+cp5/0TlZWsHmmIs2Pxyl5+8HIIkSzQf0R5dEslBJGFq1eBCMKogpVZIVLLLua
x8tLkSyWA3Taejzx1kcCTcjqv4tJkUME+2RZfhaLAm7uqyBP+HQMYc0EonX/q/dqMfOaU31Uh3ie
E6KbQdIVRnqHkqzP/zl0H505dgI6uwIfkhx4ms+bsQiOtjx2Lzrku36ewY2rQGlzxDf1WU7h/tvJ
R1MUsdgZiA8qkwWnH2vOoO+LH5xuxJXIDeaodeNExJNMwYLDW87htSyLrrTzIGiXjhXigEgNPbap
BW/Y/F8BwQ9ZGjmLD7Dk/5hPf48MF7pJ8PVtQAIEWQYPeC8W+ubX0qxXtkCjAOxbWEKwsB5wISGR
n3+0uSrzQInTcrjmp8YFxZtkhgizW7DU4qQN5U9LSUADp9T8raRuCW26sadZHrH526hRH1UxsFrd
dBrasLIQOa5JNmJ9AqW0t9nq+4sYi5X3Rq0U+FXShEpWL2hPJA7F+1r7Tc0BOi6O3S/+RYUFvkYg
DQMXlNu2Cdv5/TgvJC6CyTXmTKHVstoylC7U55Jmw7Nsjmtn3z9+masxQAV/zqF2/+Fb/szXen9Y
iS35X9b23gwc3pNt31QdNPUn8GqMqF1sTyhr7oMra8xxs6SV7J/6XJPqQ3JvXYbL6PLMZjIJtjfV
iqo99eIEa8P9Yu/BP+WPjgUiqjeDYLNJlxLsYXJVWljfxty1vt68KtpsBYAGTTiogG3oLbS7ECHC
/luxJNOSzpWyUas3YeJgMcZXkBKo3tSADLNX3NpKVcPfZhMbyAu1sdx+Xl3BJJD+C090eOhLEvi9
AoKvXXl8sheK2SL8iOdjP2x95v9mYNdM16VmOLUS9rvQ3ivxH7Kx1Aq+DjKZZ87gpUDmbZ3uWJXS
H9ZsoPvtsw/IXCRjkbZfZ/z9PvRm4UBDM5jdNFCJIjtTisHOOCRA0OB8xr8Uxs1CYJF1hBFB43w+
rB7xC9aK1E+pR7Ig2IRgh4qfU61XlH1dUY/klSTHNn2KYI7SKZINEOElWMkLgNM6ejUJ6FGAQbzE
o0x51hkYtQAC2SOufGlIx+soHpK86BJd2+Gl7QSSPIMY4AK3Ubf6qqByDShqdO/S6gdl+W3io0SN
dxH6ooXiOvC4lrcnSQ7YbRCds7mMNWPHmIag97Mx+iMYl/jPMtmscRjhWUXIyE0S4YTUIt/jSO8O
cf+yazRfRuSzP8spDB149JcSvCj4ayJSBasvN1yFu1HgfxdH6zNL7TLG7E1MLlt3r2bLRLaPENNQ
BXAVJjrkrQzyFxKnOx7Qy68L2QdHyY4nLBXt++ZsZ7P+PZMVMzHM9vl/URHgRGXSxjIaiii2NmH8
ne9bfohuHJ8tBfI0KAXjISgFS4lqsiIhixXndUBQ9jncYCMyMvU6MmsHqSKqLM2tZw7hBjvCmDTg
QwBTf/gjvud11oq0OnTK6/BvVeP5Wz2u25SSBsuW6b83K8vT4mPpefVT96Q/r4MnzPYiq/sdToNo
rNtYJBoIxUJkj62TIwplJO/TNA8+2qmRPeQeeYZyLXJCpgj3Pv8EFE/EHz27xObikHAXm3+4zXCS
Hgf4coskgIehPqJpZF1HixDavC66n9gOlNVdUusF6Yn+9XT4Ll4joZRj4034AZG8mNQSDw6mGXFh
eoRJlV0zWA2c1TfAyHrXfSaNa/Rtp6QQKU42O5sUWfUptU+mhzlhyl1CQxyU/l5cTK4MWX3GTlb0
DWQ49dOFrWJUppxaf+8YNtzZqY8DeL1zMDz27qm6Q3H2eULyKzI6Tzog68EScXdeK+f+f29vK5Fz
cnDeO4I/mb5cW+exSyuDrviSlWcAIlnBxk46b5HWCiYdBNOP3IK7uuu8TLYJxX0cTXS1IRgm7veI
e4OttW093YnFbZY0T0da5SH8KWZFP0EP5QZh2gf3k6IMlyAf/R0Sf1IT/1E2iPPL4JYkh3Kh+JP+
BGVQOe41CKxM1LitDR3jAwDofUwWAN9ehScs3BY01K4TDIhwcfhh+SvohJ/52D9szOwOXwK8OPMJ
bLOLXktkcSKfMOC7a7ck17uYpdHbeDxvrk3hfoMmN0IJKx7GEZqNnhKQ/i/rv7cZ3LjQ6L0RW1Hw
/MdQb53k3H3k+xXYNvsiZQ3Xucx+vaTRjFEcDoqYB3kKIQRg+xxYMKZs/D0tBskGOQrWICtQSCGA
0V/Ct1AiUpVk//4aZlHWk4Vaf18ISuoKWBWpZR+Q8SVxkkjdgMSbovxGa7rEL57/lkB5ORpTSAnJ
GQXWiI43m7lkulsZQaOF3QjDr0bNweBGHiOh+gD4SadGDQ0KHgG5/m6hgctlMpFLkOQuc74Few1t
yyjYMtqJZR4VTGfEC16dKCyN/Sf6V65yUSaGM/RWjV1n92aJiSNPhgIDyfkynOvFNpKS8zbdYI7r
DfYBU0/skGAO6vk02SI89XFcqWgUQDyn0UT2kONvKPLcYPGsWyirAD5VqAKMjBvcrDRDa5YSst1C
ar8ZWpJlptbBwAuvszxqzXOMgdaHO6vNZRwouEuws9u2hAvY7IByQFk371NB7aLbsAkcZttNPYdX
l0+hYhLsX905Q/qysMVvcA0gMdkxPfmXMdKgW3a+EdSJgUZaukBdEguYjYInVdBB7jUP0wTdkbZv
Rm/Y+PlkFqT1KlHrxFthHsvdeuk8PTtUTe2QyEMavEOT1uMnZmHai7PzVyBauw+mnBXbdnybauOg
GR1VHfXi805i+WoVhOc3z79B8kAVk2mBz0zpxNx2YSPeGnhl3xehWJkipE0TPb0v+1vTvjlaLw6x
AfYxg3oiKULh64sviE5ebRMrtRvqjJPomySuipXW0l9XEhxo09tiDHXr+rSDyHIUGtUuXVhAIGgj
poYGGai2/xpSF8q8Js5vw5GlFOUnaoAIV4UoyNq+dpIYXE2uomudzsRi7gAZfuCMwUj9DJM0stEG
usFrxJr/cLp26q3dMSbYmf4b3rf8EciCiDsvhif/W94PSN/EWFol9XdvTbHBQCaNXwU2XDyyUvAY
zFFTz5p3gkzMdSMslfcmpWV1k78J8K0Y3/p5buYrlSt6pTqKfu+17Ojo5+YH+nYrKXGmPHMBAfKn
SgM1kuezH31BWAS3Lfl52szyTKcpDOhntk9ZyEFYjfkGONse58+8I4z1jF3RH/35lGA12ypWxfMM
eULE4ggQ6xtlaWGD2i5y3ybuGxMjhVGB5O4oHry7xy/trafvTPQi4trvFP2hhOIPEjVs9sTNEZhp
US0v/VF/UOYwfjJyFkH2DPWPviRfTM/NLgL5mTAetEeIF3LeeagRah1xik0fioAUMwwgvJPhDHaH
C38apbcsbKGlVd9BobFW78jlCvnJ6R0Q+6RQJRPHBEzWmOSrIzJgpXP8qg7P6E0szWMWAMTO8r89
XoZToJRf/a0v63qY2cY6Xh0piBo86NPGwwS0RLeGVD3EqBzdmzcpapeilVNlXDz2V+CiMdtnebtZ
pUlxV0W1DO4EchyDLjRuJt7BXsNaE9rNTzULHPaG3NWegZcn3eZviEWeAQvQRNPkgmqNIJP6hyCn
r2p7lwBSJuDQ4XHjJmPAnrDeO+LiqredNjdKUscA3wqbfSbi8slNgeWd40RDQsrDOuOit0yLCKZ/
0LIwsSYw1oqmlHdHN7yF8YAs3HpxLUBwOTX7/zvQF7M1Atdi/15RA0CSBPvnVZCnRiJow6i9KW4N
np8SSaJmvwrcuAxrLrC+N9/apKo+661SUuOf8rFrYb7TeFxcBR6GFtGrhRx08mxSz0pfLXKFINqd
IrQ//lXYimblZtOYJX03pHlSiHiP87FOpWL7DTy7KEIybfj8yvo0R4045p6MqrkUlPgL4S1LuUNg
DDeDoSyOA+2VOurJSg1AcH9IR1zzDyOBVkARNp2kDtLdZp7cQ95I3qgKcyosKBHU/tdyazX4uoKq
ryuK8M9Nx6AVAZM5v/8cCrYoAgKJoEx+aIaTS1q9o15x552tTYZd4xAaj9NFGv63ZuDspJ28fKty
HuFtUp3hw2G9ctFHTOK4SSW/JMjal/E52M1jI1m5jQjssW+3BtZt6FI9NwkjCOVb6GtZhTEbQjMi
GoYgLvSAOanXbmvzwao83iBxtbvnLeGnMQV3uYy9xJB9ycYnYceF8cgVd9MWNj8Q5nJKsDXFkrMB
+VGuYIXHGYovKxEau8oF8DzSy0hFU4MvJBM/ndbTng4RuFnBGm6SZDVQmxxuad9N6RojwhbIHm2x
TU9X+ZgSzQckYUL9h4L1u4AuWNg9g6SwSiN5jTCFqt3gcvha748fjOxPQpE3u6vsIrPjV4CThL51
x2BiFx7FpnfrsGakiF72TeAaT1RQnEvva+pW0rMGwb0xYAQJeDuc1526eWJ5Z3RavlwQcXtSMlI0
2KcQxQY3vCnwiH9yj7Rk1TASjhn8Yain5Xmdd3E/5L1zUhh0IE3mKSfCKMGZXLg/RQVPuFgo++gJ
MmpS5eCgTNdLISaonz+fMvueq+ehPvZEnh4wpFSvviPMzy0n3izM+y4B+UMc5EtED976iycZC3Fm
UjUQXRdRzsUeGLR4THm4kOYZHnlA7OhZBOqkrF+dpvRWBOtMTdx2juoYbLFi481JV1tHxzfLC3gK
MGwlLb/061Tfpdy9ncLwAd3CkxlzvNZ7b3GhyvJFyIudPXwMEhgDWu0O0igE1ja7CFZXsHf2eP8w
NekdKLtGBuSgr4yiCo9M95r2NPphvTZ5VJeE/s/yYselLGBNdtxcX/R8uKtFCWMhpDDNsmQ0fvp2
LCt3sci6VhLwFh0zNJYopof4O5ryEiOjqsHxuJSpD/oOHmDdSOmsvKv5dEREaa+fsh5neGOQZp6X
P1dFW4JbTK8aQCU5eiV+i+EW9E/BIROtd58AprCCe9iv7YYKHQUT/FwP0gxGH4e8R0Zn4OkNOOIC
pr91RFKs/FnR6KPcmSEZUBveJTA3CbjNElQxQIgg4lMMVQTxHqXxpPN7pVcDt8xuPPAWnx2MWrlI
jiSSc+wiP/fCS0JQ2jIPID6tBNeWK0/im7spI6kiqjI8MBQ4TGNsv2Fjc1/BA+2QXlpzPKiBKZjE
KQgN5NmKwxkKHLtaXNMmiCzT9DDiaFA4zp/2vUoMkn6H9BO8BK9sjW05h1MwqF32W5wKXRJrCYTa
ZpNfuqiII7oFZeo+6t1593KjANXN8lqHPR0PgOOonUJUgjzSaq6Y5HZYuIRBqSmsyBIoWR+/nzEq
v/BK59N2v2SKAamizb+7coQxAmChy9zo6Z6pLgjEVx9ABIw4KA649mM3SMOyNzV8uDI5I3VwO1q+
j5+DGSud+8zSEcfSujKz/+q1jA4D6TQkjVTVmBTzThb69/UljwCn8LIc1YoCtmyGVQ1V3tPxBaIH
+w8M/KeXiCfq0+5YxB9zSJP/7lB72hVPPEG+/TDUGbm+DHSyjnBj43BhMUlfVcTLNvlCEVbTWmt2
nJNt904sjjprNvQfrvlcvpITNXR23k8kkVk74Bon3sel7J8oSBgR5igjGFfN74Td2LH171TPUsB6
V7RyIkvzjLi2ucx6svduhXGd9yPnqMkSiPLJ5TdPRmFoCr1isUdJIFq0514Tw5lyhF29u0DVvxea
GcRu8IVbp10M29Ued3nvU9QvVQxbDOAF8BOUDCPGBgqHj5AJ6XT46ILsvDixfx/0T8jyaBy729rp
/NO4kt239Zu4Bab3uDDeZooktioKEmJpQSK7ytR6Cq7I4gLyn7Yl985wL/r2E5QBiiudVD1L0sRy
MZdiNav43pSxmV+z8hElM39Jo2cVMarxSckVktRzNkFaRq2Azo0nRTrxGD0H/UHYGynw2VLIGPas
EL/ESX6ul42X/bSsNHo03Ygi+MPNlSTlSMZPhEgTE+IGEWeXFJ7qQ3kEcFXot40OZcHxJSbAynTN
qZIAVntLedT5ysRgNC5W5JQBF6TVCHAlqdwaMG/zoj+GkX+nzczMlxaqLcwI4iidr5XsGDM8FEs1
LrhE+yS9yWd622fzeRHlHkPE5n/N8noK3ms6R1yAbHF5lC3TI1GabENMY+sUa7oufOAeyTx/xO02
sPxE1qlUIFH3jb5JoZcPpb8Ifc9cK6VZ2W9Uof60WNHMTkADpHL0X/6+DZySTZbLtT6M9wwfBUjq
Vg963YT4K24puopO/10f10PGqNsQuSR932JmPcnAQ+SGo3JcL+dgIAmzbxohdE1F9vNNp2VPdTvb
El1iCi6muqIkoLq4tF0yUTPcCFvslkumMAQIVoTEl0Ge17EoaBsPMF92EZBtusII6m6N7YPaN1n2
B6UrDcHF83X6i5htERzSMI2x/yqELOycn0WjHxAtVUDC+YSXKmckhTRe1OKjJfCqp9ITGtMtqJJ5
fiLAg7nEQMHQY8gEe2y4JkLMR2s9N6TyJzU3xctrP4pz7PNjJqYcRc57UZ0MTGrqqGhWRwwAyIIy
2RkGbpqmAGYI1oExIbfl0uDwKS1SNQ/J5j6gXydTJUafQLwuZ2/qaZqWdi0xG391dm4cDKuu1EzA
vOGamszyIo9p5+vYkP3N9R7powWYmQQ1bNoo1MC/V/ZwgcrVbh5xwNpEWA7CeFhzT/cgdbdzdEQn
o/OuVUErEZd5WorhQW0wx2zL0Qkd+q+5kRppLWoI8zNy/zmqnRoeA5VVuGITO0OcJcfNzTLWj5EL
jV0TLQ0Xn7Rq8wcO5lrxSqQE3gsod531OTe07qS+RPXHrcyKeH63UlgBMr6l/aLNV2ocTsNKND5W
wyVkSNlF3SJIP8LPlV90BxhLacMH42JGa3hEKhU2ZW1rKpb0CDysiWuKna7G0YJMS33XPNziRIo6
E5IJeax2SbP2j3oyYeg9QoxwAhkGi0QrxxUJajtBUE8EWU/e8C3nyGUTqBXAyIp+AX5oTHsidFK2
dzp6nz2s43Gke0KHmUqPxvBxZAUpn7gVh6x+thXczwW/0f2DoJdqeFnXYVYV0tgE9rvpN5pkrRf/
ayU0BgDT2WzzG3ffpJAlHIj/GbMFz3OdIkn5xR30W85XQ5oodElsqbH+LFdTMI6PwUDJGl02octY
vCj6ihWDYQZF6HD6JK/VUyo5O7ZFqjmCJnHG8Hw5Ul01vnEcKi4Ak4Iq9NGqjKSAzudytk4QMaUL
RJVVNzuhXgOaymAFlg1hrDNplnQzYPw0ythw1Gosl6Pu3KlfIddjzzVoMx+mA2wDqdXd5OIPHAoV
Hq1nqhcUFrt60WvKV+Kba/uj4e4KKImECUEDrgeQ4NhAUWU/2GCRf7y5g37pSpb4Kc08NvR2E9bX
M75L2ExBSqyW2HZ8kh4JXp5e90f4LCwNDSLenGmn44ko2whhUf2HINcLZJfoOsRpISxz9fDknM0J
uS+2W8GuSwlzHwDhHZCh7LRMUe/WXsxOs1i0Gc/UMsTjIrYHu4a3JFLvTNHdJP+wWvUQ6z8eH7eQ
Ey7gacSqjWtw7KsceRzx5mYfmYzmi0ie7V7hla4Gh4zcETpdrhGbKLe3uC96SGXJgK23gUU2TE22
VrDXO6aUiYFulxb8YTOdxgoaegYE1WwD9fubStHdnmjFA2a6PRso+/mpW2AEmLDyjuFrJA6zhBpF
a0sLjWH62h9vzYGtk9qwWfqa8vVwXPDgg2EWJDqroDIcvqfS4hn3jiR9w2KC+SP0zoxc9DzMF1Ah
IAKRgEXqUm3LwaDg0kUMfSnZUAItz2FqimNOcurSB2wT9cqGgReTaaIIRD+1OFR6d5F+/AX+vS7i
xCwkKSAiReGy81VcTz8fazDoIJyuzjSTwJBBsmTAe5hyUY1wIjVIMFdZeHwR7bw9StuNFmk8PMqU
XdpJAx3R0n0aAlJqq0ZuGSATmiGQl+6jLSNVlxAMpwnZyQiB301CJVEsnHkvgCFwpdYOHhoImTox
WCEPnSedOQnZC22WkvUAB6aGKQvhLYmjpd/j7rRH1OTTLryoc0Ibxrray9Iz/KxGLIk27CTtVyOk
FTw5IMqgvYY/tOESGJj3UO9XRUg0N93EkGgKTpSAaLCazaZBPtL9t3361EPqw4Tv1hq3sJEkzogL
m0N4HaCwh4oDKK/UhYF1k8Wigo+Zj8jLhB9e/N77ihPqe4YE+f8gMyK7dXZgp2jWgyWS3Z75uzdw
Uht9nsV3azSxNsEKwSBAO7tW4qqXoFO5qbKeiRYJKdwdy8uBBD4UpGWRMgNguZxobpsHhnMELmII
nTGlDRyiEpMJpfzAXSaIamEn3BVxj3boOKhyKGIzAglG/dFUS0rrtJ9IEKGANy5w584D0wp/B3TJ
4O7+VIE+4Pg7s7jkirFEgoVDbPnqbbTJMlR44UQuCFD1UDv4yTfTQuBaw4qzt6bZTxp1XcdlqNDx
IDLZFuhubG3ZhI1OMt+LF6tvyM2y9+0zSvzqTjUBcx3h6vmxAIkhDI5hDt6xjNxPZOpiUNKiC4Cl
Uo+Vw66cpzec0vCyaqQpCtcpEp3qjlwHAvqjnKU1+2Y8+qeR3mnHyp5BZZEvn+O6U4v2U8hdikA+
RF+/NKGAEPdyH5YEBMHmioNKg1pKto67pW8M/dwFomSTotgnad7tWAf0ru9QNBLAPdAirZ31wsgm
vanp9BGckN8etcJNvlbC5j3BdjjbaXG2e876ymM+U+cSDnaTbz134rCOAQaketJtXnMYSwS9rJhU
zRzaT2kdKlPu5WCukzMgA1H2lCuIAfX36jAbp4gLv6zZFxk7eKoRh5c2BHh7BGnon6HMGuVCl6Va
Yiar1alJtIZqM16ZH07pCFBrbg9vus/WYLEDT+X1B6onjUAf+6vqnoZ3LAt+y71Ea9DVh46gCInt
sDhK2FrpP7pAXDISiFv8SL4qJp/EoF0+x2s5TxKr3hLP2D7Z1DgJIZDk5iDy7GdIbLpk5FdfS76r
oWkxiZxSPpQkMxIs8W8kjU8aH2C4y1R8gMDhmSUvP9ZF9aOcB/9WPSSzW9MZoLHgDH8Ae2AxLA+B
Zee8gP/S+DOMxj9XRUo6BR4r/d8PqctFv/rlv05bDcM07GTUscXiHbtAaNjjwmrubSig3cXaL+ed
a0l0RPQDsxiHYmTwASIJkrON/XosLlE8M131m87qpHGvnx2YhpFsAybl2XwIKFFdsgLrermt6On3
kIGa9bsKG1GpMhH1B2AMAn/1b0gdecWNpdFOvv85DUzuJ7mlx45ArQCWyu78VSbOSiKb1OXj7Aga
wCFMoa2+0rNTbHthxXH5egRoepnsVF0zdYgCIvGzqclMtEBve9un+vfOt00eukCMYJrpjIyJC1aA
RWKpOjD6u59vwuOWFhRX0BSDVi9fRnRDKc/I/mZncv9dRhGPHMLHk9QtSKNXCgExUKUt2HP4IFlD
mA46a4pbZzPjlZ+Zj7iun2pHeOiJQHu0W6LCLftWVSqdI1MFcmBWXD+qLYPUQbPdZqs+QhgibOFA
4378z1SMAQv8LfUTuOfKJrzZQXNHR6Zv2QD+SqiA/9yeX9yVA01O9Mzx80reOgiLGJH9sei/EXlW
GHvAgi5MdLUDRaUnpPofxyBnDgsMjN7VbzPVBmDzgX0pdXgxmfgQ/NahJAJ59pE+wAGiQu/Kxdg3
Q85sHl1E3SrfFmv7p9r6LvYtZ2X5BMF/OEBM9Y415ST0RdSGl4H0JugsFpxnLZsvPoMiI8FUghdg
qBPUd1VV1IpiBguXe0aNeZB/0M8GnJR/BF0ey3gwAXnR876HaF7Dcp3iKBWbTS5zAxss0mXhMjci
+cvDfFGYnOWlD0hWE8aQRjSyDtXxucdD/qnHwr1UuGRAtrPX4L3IZRr/r9mn0YXgqxv6xCn0svG+
LjWaFH13rEhJzzkk8sA1JV+PwUo3ZVJGWfkcWtyqfYx8HLfI79yoLRjX/kvPf2QG0iQbqyWm8jnl
2+cWJlONjW90kUzc7OS8dmsRRKslRHFxng4Ov8XZg3dA2mbsYc4C5fgh9EnSbcWDZokhj7KT6ovk
sBaLuausyqlqDKpAGW5+lInFpb2wAIamrHqyhRUDk8aD87zUTvtdLtb4y0rZSfvj4/UrfTe5HXSV
UYZEy9wLuD40wQ8137Sx8/3Q/HXtxKNH1QysztBmHdbTSBysMEjjaXApBBtmPtwZWheZWqRlyOpC
2Clm71FbzYkFB3zySV832/hMt2pe2KkCcTsYIW8+mKdMOqO2bCcAi621qCbeP9WmKIZQLYnEAoy+
2uE3rHoKBXRVvlyLjNtzS3m7VxYDvw7YVJffCB5T/+nAPbdyKMrNf2zc72n+JLXb36nSZU++mb02
KV4l9Ij0JomlePS9xqvUPxDK5UWE02C1NmuPN5HErxJtyCKk6JAShUeeMkx2UYXcmPuxBAlZcSf0
YHIKshsEByAIPGq/bkLofWWQKdIzD0wumLrJilCLuYa6WvKH0EADaucIqpOjgCrq44e9Fl7+zMD6
6oWRCkWllR6AnDoRHleq/Le5NljKllccZVGfeTpRcNOTJ/ghyyQnb60GqWVrtVMvKEserWywF8v8
CYrNqeAU4orcYqJQ5G2R/0ZV3aBQpG7k/z50m3VsRcZeBZHS7Nwr1J7v2uMOm5z97/4Th4n6TNY4
ePs82Zh5EZLeY48ch/L4HdKJ1aNM/QutZO6eBLQ7UGGm1uJOo7w7PSV66YgwupAbD456VzMOU8+d
fJDqLDjLD1MSUMdsw4itsTu7OZT9Ay7HbTCiGDzVLtJjbCUHs7GoY4b5FonyGWq7Jz6pegSHOSlF
i6vWpJI9L/Wr0PyZJjU1r7gAgA3XGp2ZNd8EANX6dWcfvpRMAqcxVRZiQfAZ6jXSIkwGpkgqf++E
CVM0Hfj75JNERmslj4KuvWRxwgbDalWPBrjRKlGoyjTe/BmbScKX76fvSFo2Zsdcy3cWSmUV5Xr2
nYkTdrfo1gKqhZRULqU7k1SpQkPUwqc20i4ofXblWBgMKaP3cgkb5NDMepNFE/uggs77TBlIbng+
yEUFRZQEGSFEpkTm0Ro2lggXbnF3Q1s5tZxqTSPAIHUabrBWhv75lM0cA6lRbjC7xogGpgyD0hr1
JEX0N0hDosuewKs6AMzEEbDk5z5hpLiKgFGlakZp9G4oU8esKdVUK740JD0V1fZrtK1hUO0eGfIv
nuibn051ho9ihuEf0HwLe1Yyq9z/XDDINsCyq8d31o5vZl7Eg60RedhSTRdP2zgHJlmGglAo+O+Y
Rn4x14oiB04d6sLx/beC1NRZWpzUAE2Sqh5zXaPsjXgmKnlVg6jSF3o07BmY4HjgrfhkvmvOXTcq
SmT+z+209C4KHNnNVj/4zHpM3E1wMFQnx3napmwsRoy2iaLVvd2j7pv0vhnfamMLjQ23J2CO0PNu
2UpVJmlffoyj7nvJx938q4uYtae25tGcG7WhbAT/9EYR2iP0Llz1iSoPksdbZT4Mkgg3QN8qDgUa
VzGhIOVuAEyrkriiZ4eFdCOy3OZwBMn3aXGkwx/UAi1J/LRAvvVHFUaWRl4JgY/ilsmqSeKImb+K
pj/hP3fPnFz/C4Ls1DP7qEEJ43DwqMU5sIsWtAbcmmit2tofudSukYKSXhhChK4UvwwQN5eCv8mw
sM8cVgW+wwjLSLvhMGVs2MyF+zi15NoALMN+ReiIkfKva6HQqn8JNhBfxQncafvhma43rcntARxF
waJufxw74zg/ovJ7htPbkJcrm7ErL3uH/K7+bAa1TA91JFtkt2aryxFe9zGEPXucLVGh9ylS6slC
iMJqbTgKltO4vpdsG1Qu68gd2vJii9/jI6qHv0tXDoqjKMKexByiKDyQZICWLP0Rob0Z3ydfl0Tk
JA4pt3RxkGl2hr4jiCKkEDuQu6UKbOgdRfyQmr6zgyPQ7OwDLjsOT2n8hpqOAlX51eC9DXnxMDnn
M3eWyHETVJ//HVwMJYYB5ZvMsgPC7o1PZz9mxILEvPiOaEFAL/g25ak3JPkdIJILMi1zs2FJAW7c
A+0funVPjTtpjwNK7MfgkHhsu+sGIxm1hwkZgsD+txvbu5rFsSeSA24Z839VqCG/o94p13wbA8ke
F5pSrAgG+/DVQRdvdFz4WQNAHaA8SDux3UX+Y7s/RajlyHNip6lB/JuQgn6UGsrgHjhcqxZJrMpc
jJJ06SuFbkvPtJwbvkGbVsgLdhgl0jTY4UN8OoF6kG2yH8WJscMihHN1TOsvR9mQvpSZIi55D08U
obwQfIagm4XWWnKoaBXxoixqK8jjpilD7Sk90PtqqXKAH8ZJySuZ5pLeGn0vUSP2rdKZvYsRruUN
DzbGnKPH/ULRJTb2A6e7xUM9gcMFEKC3P4V4+jUnSBtnUSlW7iUz7kJ2q8xfAiajaP3tGMP4NCE/
if+hKLphG1Afqt1Scrw0ST/FbBtyilwNSWMMbAHSQnPjlUNr72YjkdkPVfCnXgaiQVO5Y/MR650u
HSJuJwGo/Hbg29Pe6bd0Nfb8cU+kIl9P4cKjEHqVsQ84xXbYXSK9P7+v3ulUldj64JQW6kuC8z8e
3w73NjLQNR9MsemCqd/Xck196AFnMjxUgzfRCfqbJ3O70gwFY8QpUZ0ZKASKQDkWvxpfuN9tqWUg
YbJiH5fZRP7SzB9VCxKiRHeJyORbOAT7Mi9RidmrlvOdoXEk7jYGJMF/UQ467P5WubE1q+0wJQUY
WJ56XwATyQVRrhfHmLQc0Q9BjS/huT50kE1y6jAZs2Sn3sbjaEGfMyjrOCr5afxA/Y4/quCIrvLV
MNnmHZsp7lnFKA6Z9KVgkKcsCMSw/j0tamEC73wnid512kf3mz98T78Jk7aEZWIUvBjCai373KMq
5UHGy/N0mti2Oym7XDyRs8zlD3BVLi+ZxbAjjgPbHCoHJcxEI7/1kYGUhs2MC4kwUyRTDjYHSw/M
jsEuuy5s7b+K+/HMlMdEEKvPgUDP4k+jPm/mNhuDxU6Hugj1v/UlHp2754rlm5lnM76pLVQ8HJr1
scXF9T2WkhtI1duPAMNm7rLYrw9m/lDLFF7CS6ORGEVLFrlaxxErzOSDLaMIMxMlfuu87uytAXOF
kQqrZgLhA2lpRO3HBeJ0KFXzB83EIBMo5/ZCT6ZVSKXWbd9o8qN4m1ZVUCXm2mswmkxxwa9VSd2P
UEYVcfZ13uqkevxC4M3f9MEJy7fMIlF6vT3z830ZKRAlDi+F+9FDV7nDbXRvwoHEOQ7WybQmCqiV
u+uHgH0F4pdQDT7LvZn4Gc4YWYUlXtVdaL7Fp5pS54DVF1cf7SxNim5txMGzGgDxV/yfdmnDj8RS
fLdKeGvZmfcKF6OCi1W2aH98+4Pqagn350gCwz2buYkm5rx/cLxlIjTALPWF2YLTKiNAF3RNczG/
lR8bwASpHEKBt76u4UND567BYfY37/sxJypy0XZYzZfVJnSZ0bwrglKY9eIAq7/yOogrrpSpBs07
UNVicZ6Rhy/HUVjezgFV8sZGTSTVOfesElsMO/GnQClRFo5lnZI7C2dwcN+kJqcLcXIWqnEzbFHw
+s9JCSZ78TU3oUIOllr1IHORM4/Tg7tNmnayAsanfnUMHxxFowkdh4lH+TTNEe8K8/Fhqp5qCTW6
JxO5rCkTCshzGQoJYma963CQePrVwgfPsjG5EM6VbnZn63NWhSh68j6sbVccN34CDq6XLuNkVOqH
dqn7xdpcBe4MFBzAlD7V+kGRVJZ1qZru+xEBd43qe+6akPZ+JvxZYgIxC/zkZGTe/cB6aKSrdXRk
nKc2wj90pHoIHwa30LWe+Bs/qdjQLwGH8wNeKt7U9j5eBGcBE2Id6vc2recMWvdWu8FnYyVkQhpy
dpYg6bfMs4xB9rJbuio7Uu3sobJKcYlTZf1uV/+oHemNpIZym9aaQa1YOIH7tFscPOFUJ7GiRyWH
MeR9EzBdkm4Bt42txWPqRSeb9PfWrN4yP2A4rxQL6KDF8E5Us/LubHB9KuqevfcXJY6XBGazRk4G
1h42iUDzznvP4E4tkb2iP1WfO9C9H0CagoZjhZYgthPpq93lP8C6s/yNlmX0tjpOJk9wKcgrT6FW
svk+DuHiRGK+iaiyMPYA3BOBnH54Yo3af2HPty8MLLBqpXnIA06JZ1ARuer+y3J3G3eKcNdhjHuF
LD0jJDNRJ7YRxCCaPXqdW9mybw+1HMBZtxOzBaN98eU056/2BCTSiUY2RnZBV+sDN99LRd2614bt
CEC2khCIa8hZVff7qryG7Hlv8hzwg2G08YHtABSgoAi89lZTqNJUzAdERgHonx+Y2s9vPXy5BMfo
nYbDGPN22t2SBv3LF/HH7LIQkTQVvX9c/vdwUjFfpfD8AVZzknEeWplCr4Cjv/qpgomSbyI0qs+l
O4DQC+zu9Xrr497sOnIE0nZ8E961csxMjEL3+MkDjTFtiEPajUBMWfQLFsxN5WLhyoE2BXuN25UZ
w/5jeQoBGiR4rWuL1hIUlkZ6TD+IBI7oJqzRhHdSSucDmRZkSZyTqKKFrchHqEln3le7coKmgtlu
H8AXAO5f5sKaj9Ar2rFwt9hO0/XxovjKYdiG9Rzk+nJLfmQlUwRKVCZ57yLKGW7bPtoHM7lNNFg2
+JGHtbWjcEon0W6T27q9m0D56bm1FmKcMdlKBfiPVGcQ0KlEoN0kctm4FQbjnagN/OroYmMuce4e
dygsgl6pd8xaF6hEN6U1ynE8CLBUV2W0W17DvO0Vr+5E6u/K3NXlKb/hZBSzfS1qgaIxGSBwg3NG
syQ20ZCYr3+adXHm40zzAhy0QTO2YKvMMLX452uESubC/YxMaYH46KyX+RPuJUhn3oVkzJFEvsOj
t2aGr6lr+hMg7Z97yQAFZkNgcesT21xXBcK4hruro0npudm1XMRqSYJ64j6VW5hFq85LTZLJ8Be0
OFOx/VSqZ5OlcjHYDYlqr6UK2eRSKUbv6Go9bkZdFOcn9o07/JVEvNuBZk9nRJlWzweafqwAXFHa
wVebdMsFQXz3QFaKkOyRdKcCZlHETh9TZf5X7bJqKiBTqGVa0RypAyQPlDsA5id7b6s/HkU3IVob
ILafW5i5olNq6iBnzti2Xv/cxO0ngzLs7vYVGc43IFc73uL91I4dv5fhc5pbrnQY+u8p+b0NG7F2
cQBDdRuXE+MxGaGw098ujCXGjnvUTm1j0x/f/1tVL50CPoUEXksamr98zJlQYww80Cer+upRrENh
g5xE5NJIgn5G3ywlASdH0CuunLw5dSj3EGc0i0gfUP/HFr8Nb88z8ZD408Y/cevL6rGhKXJWIVZG
h7xMj4IdU5T5c1JoD06JqQHAgXTbvg0md6rCb8TYkX2ig/hw/j0bT6xyCMPm4aLzdUH68Ec09NoF
s9u1L0ifrolf9z1rpYkLsaD8Q4S/pebHjwNa/0LzXeUWGyTPbEp4xW+HFoyxXbCIhAkrBRd0OvLi
/z8uKtQdmPQB0+ziCYGyh8Ntqz5jxEdb2P4kdeNo35HGpnZlUj7m01Wfso5954+m4Qtvc7x8hUc0
Enju4Q/ukGl0Nb/wp3c2CJw2KP9fDZzQYxJP7PIxAFvJ6M/NkaiNgZOlzmoekm/NfwJj14vH5QY0
DvdqAIPbecgQiBU6qwI0BuVGBwM0O+43+mR/Luxxmj0a0iNWCOoWOeUAWBcc1y0jltoQUOvlTcRS
0h1AFJPqNOTg9eJT6e+TpN1wajCQ2rYKRIb5qdCld1sdChJEceAeU0lzo7NoTrIUZqKyU9r80Ne6
rF27+CPr1FfDLdZsykf/3yOqgYwtsXjVBhQpKd+9/Z/cYdJ11gy8T4vIxoZTCnb+6nlRL2DwjfX2
9CkCGV9aH4wQPYSiN1ZqYkwwxOiXX6zbQ1BYhKdV/S9pWiR6LRKAgpZ52dZ49iQ06nwBCPryot5i
6bTAnWCxxMdrQOBH3wm1fWF9DudE+YrDAz7FI05S7Xs0qs3nLYRJs+cXzerikS+79n+nmUcZo7Mf
IASdwpvw63+XJBLJM3AjFt+/bYQ44VAvdXg5/7vD3KThsHKFprMR0SARF1fSiWmVg2aaRYaovMGQ
mevZEIKs7DtHfgJDOhrxL55GiUuNLidGVS2Qcc61u+9ymvKUm3xcQbu2riMqJhRWUzl2wuEiQp11
O+Wjr+mT10zVgjCXVOJWeXxxBSy2NZ7Px7mqd3xjCJK9KE2OKNSDwhYx/n4IBttm9yF/z8E/1Rgq
Fbxj/8KgjFfW5iCN6S97UD4EX6PGBfGm/sZ3Qj4G6VUH8Qo/cah9DLF7P04wvadJkcfHyINx98DG
X8WjUCoJAMi/Z9fD0OUoyuq23s8ionZN5yBF24krH7umOx8S0DIBCaawPR/KaHKQdFTUDbI2Qqus
Dbs73IieZH+ZbTKtfAwRFzBpEUYLeCC4hYLIxolIOByRsmKtVuYPcoyUJAsIIjjxO1ws0Mq8muJs
COu00Ioj0xFfATCxki60S3ryE5gbKFHEwANzTNtiF8ldt0rRux7EQ3C+42UQfvo140xlOOKUH5wv
MeUOv5zbGQw9uwwa0WLHesOSkeYRpiKZ03bPGphyjw1c7kSQMc/++OMsEovErPNB/1oXkxDeBjrZ
wLVW8b4hmJOvLlqevGNI8n91HYHn5fC6/iZRQyyTYc0gfK7ql/0DJeHhLefVYzxGCG8H7dDC9c/9
HWxLbj+9DOsBJJwfkuNJg9fCyvzGwm5KYzxD4RpGdR8UPhFH3k18XnH2Vvi/IG/vatGAZPe9c4HS
/H4QfIEMIvbeQ2TVD6RqFyWbwKjaXKUjq6cG6KTQNtPlvJjYs1nyIm2aqFiltFy6jJhc7XVkeuYM
5kUMFBCzNR6GCEkknHVmP7Gkn6MZoC6hI8euhXL/BChqRcKUyxyBS4VziRcHL+UXa4WUFZjCqaTa
tjhM9kp8AOzH5f3m2qGFjoL9JyZYlp6EQaU7yedVPIWPgrspbIYuTETWg+BsdEJyuiJYmrgEyPFk
/LB836Vx5ErI314GRI982NW34piVKp2jHe0vgdgf8Dbo+FvNpXL6KSo+HltZ8zOQ2TdmKz+ZEsAX
PU7leOLSrx5ECedOZQFTODaEOmUB5pzMu2m7XBh6P+xLZhLBSUygjaIxzgiHibTJkPdspH8j+Fe8
oSC9oDHh5XmxcUmnZM7sNf8MsL3HLTl3erOclrPRhgGti/v8aJCnqsuT/k5oINoqjmlPuUvsK6XH
LBrG50LosJBBbRWu1wsSGI6ess7KbPknVWJV9Mn0WIq9pUUGw1MeWGYWPcEqZYqeiibA1ZOYUviU
CwJ0pcTgUn7sajHMZzVn+6r7CbHsEIXP/YqVJeRwfDPs2pcSDvrudpVO8VaG7FP9yZ6+LFdkGfjh
AXJh5idAQFpd6w+GYAH/F01w2000MHV6V/2lmsEDUym04tppV4jp6VBbCaotPADVCwlOTGPVpfVc
J1uu3MJZ0kIqtzfIxUb4Dfam8vd1pnMQlm9Ip8XRM6tV2YewGuLiXSv/b+1EGw6G9F0exTLU9rT6
zkq+shvflY1x2yqkOp5NNCKX4QRtDouEzk/bEkGrkWxXlRN+OBKXOMhqNKRw1eMzD+Dssta/SEwM
NbtFZ/USCK5KVD6kiXx275CNX5akG4lVS7IcjabIDHYc6pgLrzO9vBY1AIeyiRrjH9qZaUeyGxSz
Xqj4Sw+BD/V5f/snSsaXrfRek94hCGLV0AMJCy79mbgkRKfI9VpjVWmaMY0blOorC6NFTeOx1jNE
tvFRBJE4SUWBE/joe8pt0M3d0JrFjMOXqkKYypOgbzGeio5JrztoskVJQB0saAECtYJxWAvtkj+O
XxlMciAuxWFpjrH9Te8ViUdfRjNzAXg7Ne2FwVJi2R0DpUr/qKEC1osgFg/MUdmZYJ/PnCeMdgJh
bf5Fu2dRGPWWKf4hHSHpfNfVQgqdGNwH/eA77hW/6LLg5TaAUgeQa4qg32GASaHj/KCzfefG+bAA
+BKLqODX3llw+qpXAw2kKoGAEcIOfdbACjtb++MgI/Crut8y0+PpFo9T/nL5+lPg6+2HeziPrzLS
GtrNeHmbx9IPo3/zDAbKxRwOhE/Wfjxig7yBaiBS+t3Yx3Pa/F3S1I9FAVkKyTEMZ2BCPo5T5EU7
ReoBC6ORH3HG1PY4j/bk7MbgkX6nPQ1Yj2408eNKWqvb1L28E18I4OzW0eOw+Hsnm1GLtnSG97xa
wJrvamxDSKJkxQ+hBSgEUnQCTa1SPrbNDA4x+xd/hCAKLkNPTVKK8hRwCGV5Vw7ly0JNBd6RHDb1
CnAwHOX4Wst105SSM7aYsmNjIdQfVvz+yXJSjZmlR5mvKbLwzzbWJO0JvfZVAMcG2zcEqgqqtqQc
se1LAx4clnp+NAL1KWxKJJ5fJaNDj9+YR6pWeBJdC5ijPiXBW69UUqueTHQSdax2iJnY3SDv3FzY
zwJ+f7cG3OyHZnf4luS8U8ru9P9vlmwDKZPeFVGBMOYLP/wl10V3swSw0EJUfO3E92/I4gdSgDqj
IHRcukksXpWBRTAaOQswyW4kCcscUR2a/7h+LrxIiAsla8WaKKMNsM2V1xNA2M5+ChXecb8Ljmrh
jWvmrFinWczi4JLy7mxprph9cEX94hCU5/iDa8v087Nuvgw4LFsIx0iq/Jcmv+uoHLkO0VBFOAd/
Um2G8310XVbPzJkaUv39LFsWt0WFO7/QjHy+PPpbgvVNxyhDKGjtwI4tsE4Cc9UyJJRSXlToHLZB
RUWV+bVUOLb/7j6HjvoUnzlB48ClMfc/xquYs3qxkk7bXAOsQG1Lf/i7meah6WMCeYL+JpojF8C8
nvGuiCLhwMIHmufSkjbOL6rHYta0SJHozDLazud5dWfmcD38DlugaGQSSuuNZVOlLIXCq36wmq/I
twtCMfCHFKAWSMN5pQB4UN1KGuRAl67Qntjymz95C+F+v6vCz+NhASHv/WMzG0Ryq81mPjKFxiKK
1Ug9EZZVhISdUVVXaNFhZjAKVf7Xx3M5JVgKtYRrb2vWfe3rMPxScHkttt/zlo2pj72svc0lzAqc
HgncJ2cVvR8n3e7vxcCKd24blUZYsKJq1Ihv5YAS6ViNI1lrLZ76cy1m0GR4mOw5gGnN6n/ZipyK
2yqm+8dTTRk4qoQYH1JSzMGtMeBrGRYuMPqRh5FzcO7lvbdiEgc+Vl+eb82y0QocBS2KQSjRnDnA
t3YsiYWfazgrHcMZIenbKYTvWQtl+GWkj/i5Ea9dcQbkTTwtW5+GjgnE3Xk4+7oil1aVc5HS0fQU
OIuuWiUuv8/kCU2O+NAkDY9iT2+zVTnaC9VKqMNlVUShfjA01ml2KWFDclI+KSxGkhepqEL7S04/
Fx85eMBpdoynIGG0jWe3ITS+/59IN8FJAF8xjCxkVMXiMVXH4jVYDatiH0RU+6AEjScu7ogimj9O
kKGaos08pxn4L6xWE8Z41RrMzVGWuiOBuWpfJw3uY7XaLXkg89WUThUupg5xvpvqZEfThUoFHZ97
/mDBJ3vL9G4qHIU5RRqrJf9BcjYb7OpxFGYRjMAxJ3flPe+V6EPd6Qw/A/FPd02WTkL/4J1ctWXw
Zarl0gG/UJu246hNmcnJ+H26odzvo5IDW0HLpw5AdqI0e728T1fanY4+JTuAYBLBApc0EHMyP6FA
BikLZx6BoynSuH4WqX82yfxmzUA6VrbXLymPz4wZR6YY+gWQuuH5erXbDIAlRa81V8umY4sMnkiE
VQAI9qLPanAtUycDH36+JKK2PdrnRZ7Otud2oVxT7fXSIhb0vIEnpNuSUwf8z3LrfDIF/G5Ojkg8
5UAnGV8E9724bExxvYr8W2yqW/B1DgYI8r/J2S9HdGliY1U/xbMFEz6fPfcdPWgr7NCFifBcQFm0
c9CVL9uPSjUUAHiqBxdPddU+jALDWhWBimb2dhGwACfyS84iyKJF/jkd+Aik/hMYHMqO8lK9ohRs
L6+LUK8zQHxzBZlWPH33pRK5mtts322elHnYQInGpKsUDrT9c9FMcXXvA0s3H9JMX2z+cmNwgRfc
V9oJS7Hxn45sIfMgzX84eeCvh3aqQvogzYmS6/k0dZKxa821QZSxLg54TgPDV2rGsCVbRsLh694v
bC059zAyaQyb/sJV2yZz0nppJaqSFs/RvI4HbyjuRoTsDvqdXSFWMDMgSTuJkqGq+SoCKfDDgXuo
Eca44X6xBUvIBDPjBGapLKP6iCZASiTdnRCWFgIrTh5C9DiV4/QAvXRk5wmomRj6ofU7H0oJonlP
sStoMkgkGyVeXUmbCB4vTOnDBczR/a1MYHaRbevoCOEzXmDkUolI/5aWWpoZBOtDqB8P3JmQKlt7
h7LFDQkOdV3wTZ1OJuy7aW9yUw+4TM1o7nhgsu3UUSg5QS+lpZb94wYOpOU6W8kE3OEBHyBGOrV+
dk7fR9kd5Mup6l9Rs8pjdnnHuHmnNuumD4Ae5f2spbLPtZOaOUkE2lagfna7c3qBEgr9jRqN1gjZ
Y22nliHqcD6k0ApBiIpu9L00HsRNf8atYI13MI8dX1c5eM3CVApTXWuLhAiceaDTTbrCQyQ4pIlB
tRbE/+C+UPeEaYHBf96ra7yfK0GB3zCtlGkNbu07brzeU3Sm1HXFz65wXsLrTaAM6/4Nn0Rszai3
ZHrP3w3L1WALY3x5B2YAm+z9nRvS+rULX8msMSRSZ3wjFOm8MLvhAhkRvk1G/ru7ivukkBInCRTI
GZ5lNi3ZJCXPc3H1JoZ+eCMeRTAR6lArfFWofvGnmDYDJYnIm6octXXDxjWEn+pB/Jst6pOyCNwF
gComaERn2eScKZYUYi7HNSdrKJwFu8FS3mBeMcrTTssOw/7yrtlw9xXIS1pq/635bG1MyE1LGZBs
qbi6LTionPwVQ07RU7ZQRw5AyHjqJmoMLogFGkonR+3Xgiaip97fJKZLNPeCxXbvpgjF7bisibXb
xIhzCaCRt07HTS0HgFa91dW7k82lFcW7izuBTIS2FuYyLyIUvtriBs0VRDr57XOW0op1VtArhAT9
E4e5hYM5T6vJ8xFEFGJ63VM+0qhZ7e1b+69mHlN/vkQL4HWYpGnJaVw/gpA+rvgAVV5s738VlW4Y
Yd0WwktcR73/8mP+0OWYEQurmBHD9Fw6YJu/fy5EW+4ACBXVa2vvgeaUsFcqNOo0QbJLlGf7dCm7
+K7+K3yLNENxCg+fj1Z5ifUvHxgfLpGtH79xfozFUMcYtPU+J7C3Mz+tRBPpMm33CTDbV/gKgimB
5XabDdLcUnaq0oAtNNdb6dDG9Cg6R1XyLNmmRQMfvSfVTOw7eUfiNXFp4m3WJnaTJEtq/i/Jqlm8
b8X1r0fQgTQBSa33kUfsPmtNGVaNziC5dOgHEZME+SKahKaONB12GPNIBz1etfiviJ4Gtw9xky7z
PlAL8cV3lXWCtT0Jv5y9+0d2N89Z6BEG4rD1Phf7NDNiXSUKTrbymgkkyUvc/Eq31Iye4v0v9jyy
5fuL6xvvBlA2oAmTCrouewkn3ZuGu2026H9IcxPYw6YW9ErFywpCcOhVV+w/i3+hbQlKliTVk29R
oLBtrukmo87jtGlCXOKdAfJTgkneCP/18MQYUqcnIvOPFtcvJ7f0RNjFRlC2MHUu0yzB22NWd+4A
ajKeT4A0lETsWg2XsjOUsRbWxQ7LsFOIXrODgBQMHMamZz7WqFCMCAgYFx5cVlPK0m/WX6+BBbFt
Kma+zV16v2Pze1tt3XtIPpNfaruBdjFBSY1upA25XSzIY52uhZ6SwTRGMcialA7MnUvh61p2v7Fq
we0dqjEYXb5WA3/IIxhBB4VPAjJcW0UNU9LtIiZNCG9FcfFh/R0+hkWvbNYH9JjHTBr9mg0ufz0Z
Ro4MZ8JlbkP7PNzpki1lsXuTst+M+ycXOsdVBhpxlD5QYd1Zu/tWTxuBRbwn/Uu39n0W+DjgXX6J
FzxphGrtn6PKJ1cRTuhQWHm9o9Ro+NKyAbJgW+fSoC6V06GHiZo3lYtj1xyTNBCorGueQZQEuG6U
bzWemDMCgBuGrluexVo/6pzdXNXf/QQR1Mmfio5gFEyfAXddoejuCPqJhi+YB9QdpuioNrTmBCPh
d5LHOS85b/WvbnPqV1mn/U94GjPDWu0FaXpJst0VndlScz0jO/WH2/4+PwP3CL0/86CGz2GXTJzm
CLS9hKdmC6FTAJcmnrV8zPGllrmK12xsTciHZJ5kXzm1+jp57ndtW8bipX1T1vGVxylFXp5GaMn9
0y5RBCbdtmJJBrDBM1ppzmi9WBExRB8Qw+BNKKmRQo9wE1q5yI/RXCdcPsWWJEi/x5itMtGuMWDH
9k0S6DTISlRCObjPTG7c3gvUUk4oxO+IJCNXIJGLjkM+cEIBUJ+QiAo0tBRv+Thto/FcWtBfeAOA
D4LZTonaPbQuI1+AsKC7o27uH8Xhhmc1FPelzSuq32C+rNclGF2U3DxaIrWlsuzzTlf0+ESXTgHF
xyR6kAYcWzz7HRs8/nztvdMDdWTPlEwiGitKl1aWelwqYvmC0XRI2AiIs0gVKsNxrQbvKgMRmQvX
fNjuBuAKR25Ve1weDfkaJlbx/BWrOUVv8BpFq8GHaI4DX4fp3gJZ140uLXua+9POeBMIHccWgpq3
W3VB0+J9c+W9bA+3Uyh/UC9UA6JkM4Ng9NeOTZEhwpFsM5+ilrsYUHQyTTP4bwXSz99cFh3qB6kC
o3+o84mddsJpRjVQ02U6jav01jIU00qfjwVp85LXIUgRQ+CABOFMxC2MKmtnoIyfoqMBHp0p0Cnf
FOL6340EGT2Gd1vsN5AK1oGnyE6cK9lA7HX9xUMZPptYOEtCwPxXsoh6Ey18bfw7MlAZ/S5tlLiv
tVrpdZILvvSrKJzGVb7LRrxGp/iWAsqhJBr9oxHgkRVcuH+9r0gbbIgfLfNodEtSKswx2yeyyoIi
vc2QCN9b30Aa3h9qLWyrd5rFsuuiKwuiQpwm0URl5ClVknkrm+pAQoaWiqpjfdZW1z2j1BVaYcwv
SfbrQB/w1UaBDxeyP8wBFz/oCPv29U4YmxcJEdDIOYIaRvX9bTGRMvi7vB4HlVxN33eQmeHPyCcV
2NvTBId9NuWCYsswUpWR4SYkNLDszJevtagbh2mxC1ASYNaSn12N/bTud08PQopfxU+XHKsJ1ZFE
2BpyBykgHsnOmKX+gwPbj+BudxirKPOaqvZL4p2WQ+Y81YxT9pqM+VCij/f90bHaVKBR7ES0Dbo+
KqZF8Zhyq14HoPd8W1PPTFwo2IPJGrZXhc5PrdWqUBDFJb3I2192JiiTPQWGNxW2MDOU/3ekcfO3
rtS8BXmzwUGIS7PkzWEY+NpbhasXN2/UG74Tu5T0ppHGz8mFb1/zJLFKzpQlyvE1IYj6TLu5amL7
sQWGhzMv/6gATz9saaG6rxb8Wfwbnz4COChH0Z9cahUnNaqKNXoxn2idJnhuUhwfpNP8Rbw8Y8AR
y695p5dWWAEfaNxprW312xpCyv03c8rlvM19KUyGt1z/DFAD7q54burN/X8PQ2XzmhHwE5IfD45X
Q+kQzuwJ/2Ug/X5yKTxDcy2lzyFZwhINJyoaOfsDK2kJjjEKnoVdOK+vqGDOYDge5JgXnF8S7I8V
Bj11TmYfCoY6wHFjLND7qdQXjHsSGE12kqjY94pY+b7qwyTVsD8MlW1UU/iQVbnTdPGl8WmTI8V7
NWjXdgrKKhtbXj/ZrsUx+7kOJiDKJlc3B0cqO2w+29z046OwcsJlVooXSuxN60odaRcMqsWD75ka
LuB2cT5pbc1uZYx6Cg46K4RSfjYvnDNTGLo4UheKWoqYm75YheN1KWHefuguuGU6nMoc0B6yP5n+
zqDAnJh0P/B8/V8ayXepFJEF8luIbezGeuKpSst944qu25EWasPuTIHT9zUXw0TA62MKE6EsjFuF
KWSD470FuYv1D0JE37aCpZirrK8Dr4eFKtPCGyT77h+mVLu6dvNRaocksneOoBiwddPgttVth0gL
o92dAM6XKVLTIZmo5SzGueCkLtrooEn8S5VAo0r9WmUV33ZDYn9jN0moeF43e/dD0AdPV3d1q1v0
6qfki474rmiJWjayyaWlsCRABxZbonXzbMyJjKw8gVCcOKvrd/2UL/gpaLNP8TQbG2FoteYqXfjh
0JgzKi21dyp8qWHRZNbRhLDF2b6GaAtJAD9NQS6d/wTXk1O+auGqF5ITeyT3QWG8Kcxuyj5irrGs
7cruexmsHkgVgukm7Dll4QBu5SzV5rmXw+pykzGxsJJU0pz9cfTQf0URHkEhwDmAP3KIVqnX/7/n
LXbF/yuGQK2ATqCzQvyka5XExqmN6G55o7h1vYoEow3adlE9qgIxUGcCP7RFbRNm+NOihTEG02lr
6GZOarlAC52nAU4DnbJOVPwshzNaBa6HL51w93EyyYx29+HznBUwDLb3FPCtM6pnQS0VFYsXfCOn
ua96k2mYzVH6GHjdw44FFmaCBeSRFWqac2sf7ZOMvmusMyguFfciW6Uq6ri7nPeyXRIOOIw1qcIh
F9FQvXbuYLuvWgl4pfjuzIQ/ebIrCzOSM7YSSSbfAocqtbKkxgT1Gd7dCX17Ve/SgcOdrwz8OMka
g6frhY0DYnaigzS2CdaCbsk1CeUpujtbQKA+Nrqb8T8qxcLLPnZBNqIWn9dwGWGKiwkUUNVF3vgz
/+PquG28jGfsOVOdet9FPdg8VLezcLjTd7+gp+abWPheJ9W1Mh4ZtIUvsBGvpBXFIl7Jf+NmlPna
zAtZ8U8gGCPsz7D3k4PmICnVQVnsZOWG9aH7+QrnjJnDJbNI1jiHxYeCf9UCEwziL+aP3CC3eyAN
0VxaX2igilaZlOAeSDTg/Hbch1tbYGoZwDooEIjz5MkIPv8U9Rqlg198ywS1A2t2Y4TSD4ZTZ7Fj
HFavRY2NJMMBdQ+c8i8yJQsJfV5WvLoeYqyK73eC1TGfsSAsn6TOuox9BD4uHI5EGB3TRL5eVPKc
c0ng1k1vAjT5AYgdptUGj18bMvGEtIjsuPVEc+gDOG4EJJX9CUyse3pV2GWdelqbBAjYt611vupa
PnopyJIvCnzBK8Edzil48ikWwyCEg5LAnm7EONc397me6XuWSy76FXC8njzHvTu2PBkvNHPhLlo8
rMF0rCsdNYzp6mJaaBAZ194x1CaBISrgZnqWUd8dCuCGMbnWF/i2rILFZm07wxzC4L3ybKItevuI
Z+68NRNMjasUbNgWgugmC7ZUdN1/Yk6gsJlfVlPQxO8Ck0g+ONYLBcrboWqyY6eBbo/yPZhv2zld
mZTvWiEKowaIssWxVBBL1YGVD8BCDAF2Gf304Y78deS63Wyz/+oXyhtoBOueye4jM+cFHHAb4tWq
cYC1+d8weYz0aOuZMW1+VnIs6QSSnjbJ2xj/un1p8dMQ+gPZhnKDkFXyaHWvv+BzjQgVkhPMuJY7
MZZj+qqcQFPnQxwCVYO3oW5u+5aESwnDDZnpbC6qHbnc24Hi2/I1FsAhJBpEurZj4GkG4t7OXJqy
Legn9kMc106nIeXnfj8XiJvrkR0LPpc4ueWPLnsFmDOqC+1MgC40oOChnMP+dPkD9Ui1+jGwtvkt
+iOfr3U2Qq4wwyERMfx8bJzNknvv80oj72O34zUqKVtEx6rjNVlVH+q5n9czVUZllD5okUs5osFf
Ha5c9Vzzxc9DU/V5dNbhBmF/X83WOCGbOICUOS99TxwZ5xTKenZZMp8/7KtdMBdferIj6xa8cIBM
5BEq8K3ozEIjsBg3QUEXBd/zxof2jeHKpfgr2UY7rvddFRURK9i2L84HTXHSyf7c8lMwFwQnUa8b
7ChDZ/RhuOVD3DbofK7gc6mESPDSthLStvKzE1vFxWREbwH2PUiLq9pO7T4gKs+WwUMoO493iwrr
r5gUtIzz/NOTTBDs7711yVUQKO082ZELbz+x2ToDMCwcdBGiPAml8vL3HiLQx6k9QUMbl1jUxhU6
YLqhGQsJlUaKlvz6aj/rcixw7fwYlottUV0n0DzWHJAO3+Cvtc9yXQq8wJp9CmOsArBiELLwNN2i
z2oHXAltFK5dLHfybB+jDsZ4CtlzMNzsBLmqqUQzoem+QAcUJdBimpFA3vXH2zquUf7FKOkLD4ou
terVJO5bsmYGNFmRzF1Swu9CM+FQCaDBt/yqMs6B1YlshMrhVkXoOvuryk9Wfmh2RwKJ9HklJ9DR
JdR8QOlsXGCBSaT9Rv/wGJHZvP6OqQ4wTWZIgXbp9n28DHK2r14xRIrph98+cFOr/UC/Dto5FyI8
mhjHEjPILSG3BXU30NtJQ6WscrfzDUhJXfsPZmqfu+XzbBFT78tPnuXCZoD/kOExhjLQL1gyOugR
x/MLgD6cXCtyEMMBS/gt49/z5dBw6fhuPvYiwhVd8sIQGiP+TnXOS1f5nxmpKTfSsWM7nE5esvB4
OXufRaKBG7kPEmgwmwTiEZfQhcYRb9q1g6NkJX7oXcRHE+u4uFqa27WYRex7bsbQ+368kdOAMbFk
xqSOLvvT+1vOyWt2/Kd05WpFiCgwhH8rG4yg8BzMJ65eJ9VEbICaKbX6AXtAyzOkG1J7sqGpNmqx
HGzKWvjM0vQEarsFQ5XigPbq3B4dOmQ0INI2t65LNigk7+B5YxbEDliKKmOzwxvAmrZJgYAKfbu3
0lJjH4qninRJuwaUE1+MKBajWnKAvItA5gX9+NMHdAse9D0hsljvm08j0yIexQmKrWgbA7QbcQ36
oKOGeWL5MiTy7unVBDGdAnrQfeIcQrYwkycPitSQ+jlI/7DQNwdnf+JvJ7Ar6roBpnNYsjRO+KeX
J5K66CSPgsyloqnUJWn8c5uHoKeUXl6fO81/GtLRqg49HBcHPVd1PazxvPUJ6b7IrJjmZ7Ifc562
XkEW86h+ije4of/bbKUc87jUuSC7yUgQQPLvBfHDh1Y0g3cwMbt1lkh6mTBhKVt4U9yi6od0W4l1
/jOz3iMf2vYYkjhoOuQIhvjtykarxNj/PNE4A/5kE3Gbw/0F1Y0Q26HtEOIp+IWrX+JF7x2RIrYg
3zpYG1Y0UrCpyiwWQXjZjjEVhqMcJZp4NQnfA/J8B4RpwkkInLyHKHWWVmv9p8tYi5EQ8FOYA9w6
Mw7zAexCOGtmkKbK67RNx35e7g+83EGgtOn4n3v0D8AmQlgfwggsA1iCZq/hJJ+4ZAZbKS86EoMK
NNB4STkIAAWXAQwxMmTLbadpf6rFi48CNLGS84BNN2kyBF1dVQFTziJzopaBfnHmv+YSD8zQdeNx
NNzeQsJqJPUexVIUtoBpPxZdw8N4r1u7M5WfA8QFPyCrdQq3S+7l0TS88a01mqj1+fZCxxLIBSE+
qrZIcL84FRFT9dkygSOF9W/gpZyfCXTYYjb03ZWDWcJzqrBhMF0OuqCwEnuwtmMtF1iWluuhwPCZ
t1bL/woKhOZdV55R0vNDsKISTyfg/S6FrvX0w86IYQWF/qYMqKpmqkNMvaPvF0g+1IXL2DXu1eQ9
RfkRMLMPUn8GjEyhW4pT5c5O2aogNgrIcs6eWTUQ1z7lhI+y+pygWQlH9c+eMLRVBBop9edLHdo8
mGYdvkVlMvw4H2zihrzXWBF+p02MsA/EX6HKd3cKQ2d3K6qmHCgA6tDvApzWiUiVuFYNs5dxCIX2
JHEslLuRGy5iauW5YVoBU+6aMRKnK4q1kt6QjEMKBR0t+jo9NvBL5tfuOqm94t/35x6XJQu1dR6H
b8Q6DbVH2FdxZxHc772rF0dnIr13m8mlb920xXET+C1x/eH+KD5X2wIx5vzRtEX7Z9m/ZrfrHS4O
6Sreuoa5zjyAiCU24fGR7JltgUhEy+KTJjwiofLiwKo9g+V4b+1I0hiYLNxoGDAHXdVX4F/bbbo7
jgvWXFoVwoLubFBekI4CUbW+yXKdSm3Y7evqH6rhXbxkT6N7iER0sX3SJUT74xpo9BTpCWgDrysX
ijfV1ov/qCD1yO6oAIVPcHf8LWl2iMq1Be9GM387j6aKU1lW64VoiAkPWNsWWSdw5T2GbOF0m350
nZ2ZpDscDQ+CH1iFZInhXigC7CZ+YFh/kLgfk4vsHkmQrIFeoa1o6EK29Lar7FkFev3WhRjjRA6S
bXa/zRAMFRwKYRGhiwbbACXVSqUtrnv5HMWXC6WcGYtOUXV/Vv5oDnheQ879DL2oSMoUayEstw3j
sJdoYGt5/RqfdoMVdaCR6eePRSvWVZYEmXPVc8gDTFS6o3Fd1Y0gJDbBKFUZe55wsr5KTgAh6osv
M7oMwzXulXd/JorIOEZPiWTre6+g+SCrXgP5IgdUATPYtHzK//hwwtpLIH5zn39yphUAl1vfO2AI
2iZ6aKhV6TfB38aKDiob1KLIpHwPJXBhF5qbRLly+rMDyy1y/gCL94HBVz1206NghkyUfosKjF9k
e2s6c+g+N6Rkx0FFxbYcnGcTEep3PApCttrZb1pkWQQUQGD8DB39qzpe542xvPPkqksn1KWPSR7u
vPDHrc90v3gxZPmN0uHhTL8uih2ysgS7VbwY3/JSusktnUgMpsRMFG45gUMyeWvWHpxIeI56esFm
Kyejz5ijVjKBvWdiP3fJSv8wTSg3zP6n7pcHu2jpOAixPo7yO/hSaHaJQ06ZvxZ94VcvgAy8dc+k
vMtA3g/LgpHfUz+1aRSWYvejiFq6CcBi9lFzivNTb7xzg4i0BpWsaxxVoM7FYZozwj2zaYw5imXT
UmJ8J1Db4VMMcI6O3z8K+yYBm7qYvlEfrImlAwSYbuQ4uNs693msiiacTj72Y9N0i/APmMxcutid
+N9AGFzZDS9cXqv8Vb3o2aGTpS2sCzGNDoczHNetL5Ct8+fXtnRjlqKniuj45M8E8ACl+pFFNeMQ
wXCHT1fT7V54s9GHVm18OEgnvP0B3oQQ7r82JehOahbYzIqyay0JOm6xYNip7qqzjgvWM43teXb1
WL+Loz9pe8+9D6Jcp6WLu+EnVgA8ygoMgPPZA0sG3QOrwomtxLAGghyu0Yngvl6UMWCDoF+4ekSL
C25VZhrojzcvYcoiJdj161H2VpnZjWZ6p+IlyGeTedmr1tR0LGTnsEtv+CG9x3ZtV8BK2qEUgAQ6
QzmtIqTPyw9OtMhILEXtJPjOty7kBvs8ws8vmAp0hXNOrPsNINvPU9xbjA+mPVinHdw2ayV1tyk/
1rKnSIEJfqMRwVz6iThh2pXavI5bpxazpEDw0M9HzEc5lE1VyyFTqtVVLA72EzvqFmNHsjT2iAR5
81A6xHa3hQ9mrFx1rg/CeSR3aK8qYPaAyJPE/t3Z7XicYweXXcgLtmerYab3fx8nRv29x0ubd8we
RNTLnCJPpWrf1zthrNggtgbfqs4Rp4yPx6Do7yyxilJ4zbdMnCjCsJ3QvkS84e/joGd0HJ8pstfh
u0yb/WgGLlVTRiLLqK6n2D5Tpdd9G2nA+NWwiqDPTirs7apqbQHdcNXe3iDzfoTZkKw0aVyGnU0f
OnjFo2c1FSY/dmxbH1UEdRTOvUWqlLqxy3ecE+gj71K3DLiI+Ny7EEvfNK8TUt2xtEnnRGRXg0p/
hm43M8JTTO9CYkpzBVpQr7bq+QbEnSgqF3LgGSX3A3+zquBioMSugx74I5P2cYNsa0hdmPTXMfOm
qkEBTF97N4QI0MVV6KRhvm912/Mnl1S+qfLaBrkw3yWwa++kqMneC0XH/fodo64DXLh6UQyYZH+c
ZpfGavRgFViB5HuqZ0FK6d+yuG3DMWJzq2hgpEU49BI0PiAdI61jdpsb9lA5hDINjGXmGPG8M8Bv
sy06+LEEb6PjDyEbknXlGPJQkMIvIHeDKzI9bB7rmWd2sRGftM9ORytxSVXFDXPSyZxyOwCbTMsK
fAFgy5dSp9YrnZncFpvngfGumxsw9EYvRKEIBIER78uDM47a0ck9OKE8j2d6xUCr5tjxwstBbMLr
CSsASNxxPLSKT9RbutrpFEzIy9bXcKooX0djRL4gR6Azb13XIa7CnHncdIYUgcGp6N/ls3hgS/Kh
1edIBKNI5thRfLy5V/e88VXsuFUu6C0EeuCrcJf7lZzis9aiPf5d/fisusgB3hWE8ra9ftfI0PMj
01/ZAw4q+JjXJAVGOeplPceC5R0L0xBgOmkeIdecCa95Z82kQvzbujKpQdy+twsglzYO6dj3IZ9i
b27nf0KoER096uqvI4knUGR3Q6ihOJ5dXCjTFfvAlVIHILR3ThVKQnM6x+s/gb2jjL1EPI5h2F+U
ujsYDK3Ptlgts/CpR1aoPB5s8jCg6p47tTC7IR2S29Gw3OBzzjSwjp+t7YeXX1C7cMsjLuh54JxE
o2zjQQqvGsu/Ro4fJdrFKqwFMm4vcWXK8AExfD2qBpBlNFW8WRIHh4cOmC7+ZkIyXgMtPwoUuEdI
ycCCCCfquQ2i8qcdQtLjV/aUtIzsFQO8gQUOMe+CasGgKDDgGon///V87LCszkLEX6kfl3zBqyyh
std2xRfieR/no64iW/Z8OzKj3B6yYDkvGTYLB1Fy7Y0hNYj+9Qt3ot1D8TtVWYLVKi7SdO34VecT
yYyaPnFUvp7roxQeMDQbh9t/FwoE74lDrnr6OVMlxWMwwuROAQdrSzSosLsEiqggunXkxcQqQnT3
39EXUmZ5AgXL/ViRzTnbPO2Q8IFOw9ne/EURYHBCBTjH8VEvKWkq/Cx6MKpOrTiLfz+5Syo/90Mt
1l9sWpwBFKY21kAYBvN+7HN/PxWCbF7yz4J3jYTGfXgBgMkpJ7s1bvZfnrYA72Bxdgh6rwXBLIOM
9evau66T5b8aK/h0zL3+5NUHs6ywkFGAeASsXyidtAzznHxsWYC64EUXAVbW7GtyJ65FUQ5O3CDG
kQZOvNa1NU98Q01W/PSt5kcq04B3kKGT2QRmdamYefwlyXpmVoZvmTJyD2ErsfFNZ9Q9aXztiUzQ
g8L2Kas607OomhuQorl2z0kVhW9yB6ER4GfwZNweJ6rEWlZiTuT6ulzbkFw6C/lfdk37audzYckW
hFAlRp5kQ4D0fevA6xzUEfyJKLYiGeM1wSH8p6H4EUZ3z969aUjBwST3pWTKG6Cm7JnBpEuvnkMM
/+5Q7rlJHYxHSxVIorlzitrocemitthP1dlmvO4YlmpkKz0dxiteBZCobsePU16xKLQm9ItDtjnq
yCdrA7aqlbKkwhfqAtC8e9/dn5AIoSg60v7Oe+N8UWwEJjxVYf6S37nGiYveAkHVpmAtXvbROCpf
hRCuGSZaq8IC50KJ3e2O5NwAP+78YYqh3B/yKvQ57dOYRHfiLnqHU25fMluEAA9rDbN+7QTCEtMu
esrqklAC5+SuER+5K1XLtQwp/qnRwJDL9rmHUCecQsltkmn9EsxpiOO7poFYjso/jduUwsbR4SnR
cnFMAFkDuEIcGYyky6ar5nZJEiIokAxPbqNFQVdaAOtTpVyNBBz3mPqpYCJcGev+bEqg7w1UgCpa
i+h+oXQmYxDiQzfzTUj+nMy3l7Rxtgu1HrsE9Hl4Cx40KEujxbZiM3zPAxyQh9oDswtXX8KV6p1H
X0Ym+gd/MUkltbaJvaxfSBbKG6JQSao9so5pd9bw8LWkDHBFngK/DK86lAKR0ocMMtDkuZQNjXCq
IGP2Qa8ln5emfypt0x3M3HcvvhNEYuwft8IIFyJ7xQ9bVh9AQA1cOykPHfl5UvxM+227lru9H753
G+hvzD7BHvRW7LeqkqvVJJhsu/JJsaKHiz/8i6+zJM8yuvYQiOA3j92dz0pUdyvp4K8FMAcGkTv4
RqE8WyEqBx86Lqzz4np3RYWz+Mj8KrUazbMh0MjgK5bYMeo4lihSlQ7xToYxvZs+NwniZT+/f5/a
Y0AIlxyM1/tGmYIFv0zb1ZY+Dhmc4LbxRWWdZaVVqJBnXAX7iTootROGjdvf11bAYCErgoAODNXw
NAjgV47hcWLul11jF/AkqzdUCtCGQvG7EHaRSPidpLkFgMdKQSld9Sv6HrF2ZmVGjLw2pJhVgW0o
h/QaCnwskzAcMPSAxZ0xvIx4E9WxDm8s+KPgsZqFtAwidtHWqEeHIIXp5esGbUvoxZqH59PbgNlC
Quq0diC8Sl2WmhyukpvVi/JR7MBY0QhrmjUKDpje1Bw0R2WVx8q1tpKtrj9B2eUs0oJMJ7winJAS
akc6cd4ppBC1F5TQNYL0XuS4fmgrV4wyUwHvbZriP5lFxeYjQCFiCoqr5/hf13W/twYant8FtVEU
IXU8b6s2xKJ87fjp6RHt6KDORxpjDwNIla4eqyrR4NbkBRqkfpbR9YUi/AtaOI1tyEVuCyYUDgV8
R86500u1vleehz0VtE504fSMf2TrrJ20QNe9iVUA4dxT8AoTOoi5yONl+55SxVNcKDR12Eo5qBps
qG8m2Gfx8Fvr4ketv/7+Rg0gytt6i36FBo1pzvxdFZ7aJQuP/YCHW+VPfPckJWUiLxXymI4gTN3V
U7O1LNoT7lWSxhtnoP+6iE5350r7hcpuGe+DTD3PaLDLqS/jMIs13ddZr2QOjqXyg+uG17vRkeEK
bvImp2kFafb3CradereP5trow/dLVOOhokUo8xotbCjLiwkLrjDMQSXXBxLiENMNJ+24UyD55Xdb
tdfJ5pUqwThLgTsAXnjndefAW7vVe5u1gjkMaFcb9Pz6ZiDQAcjJLtkeE1JAo3F40TaRWIXaO/RX
1lAG5g5X4aICADaUmVQ1VV+jyLJ/OLJZUIn5qd1lq4sSTaQu7XRlqGhONHYqeXy6vBp7b8In9bNt
oQyJjJzXtYYablzYa4HtQfLAYFLUyc0qpPkEULmZo8JFtVv/H+3NfYzRoq9aOI5BWXP32fbaSFsI
BY5CroickVHV9pZUJTyUZlpOQevpMH3TT/SaCK8NpZNGgvNr7oF0aObBCQuE4RdfcGnKNKT+/oOE
AV6KShdLaGnvJG7nOjMI8VNvfZYpX5qtJ8IGg6jgZubCQlF8a7ufG5vFxtD1ailPyYX7ycELNKas
jqarSRCk1QA0Yjd0R1YJZI5gHmcYfKW/xU1OgBUBCHMJ0pZo7prhMvY5o921YSHQyXw9LPUvVGhn
aRPgBh825hQzwV1l15D/TyeI7ek/cOFBPnJEWHwGGH4JBzYI23BTnX+TWFuYNLRQAqCZVoY3+3Wr
Vf4sd97sOMM0H8YEzyUFbnIybP58NI2RVmlu6dzdfeJLlqoOZBlexjPZlymkEKA++E+IbecMBkcA
mTPEE9eXh1q4mN7x9WVP8ZROZUaR/iJfLerDS4Yx1GORHiLSpXoJKkz3bbIsz65WR7GYM3q0sZy1
6kujQymF4o48SB8Nm0ixMwH8RzSjyKU6TWsbA+5bKuYGObIYs2/YN7qxxOFAPncXvaLmlkzoir2c
VKWXB7dSTgJhVUJUB1Ubn4uPAG0jQbH37rE7ZGSOedJ92L+0bQKC0AI6Zu9l6bU17163cJUIOS7u
F9NyOp26IJo/PVfUnhy0Fvu1bicifJ1TxGgtB9iyXM9gVH+qp0k9+NRHZsWw0KVrMsPJO7Sldlh2
DVUJOaoO4gKdXBzvyVHwp/sVUi48eNwO9awDcXXbp6ry5pVn46EBKKIRCnSzL/ymfO718/XZN8FR
HIHh+9Er1BT6RZfurCrplEy1+xDExnrv6rNZEYiuv9YdiChOTbchxTaYEWZNnQ8qP7vI+6semvm3
jJUf3bHHb9tZ59E8XISxEWfNfUIDeJhEH4zd31gBGh97Elv93UgnvN++6oI8VleBfiCx04mvUUqY
zGG8X2ONAzrRkyPLrstSV5HZKwsFLahk+7h0GUcjX8UmjOREZQURN3+yM8x+lvQOFDdDFuIJOILu
eAV3BAkoAbJ6PqjT4wWKRiKw3WGxWWHo2CtUO8avhNGCOU5dnHk5nC1W8ge/1wNed9QVNZMDeb+u
DdnnaYL7xGqIYh3MkFSQJu1CTLjFf9w0QSdmr/DhA9iMlnSuDYasa2iFRkQ7ZniqQYmm4MY8NWoi
YNSD4oFB8YOAcAErcDe+OOsrqoMp9ZNjNeapueFpHfgfe3x9FQOG0jKZ1Ti2Pqg8qIfOChVmso4G
WFCPnNIl8V1WFdmyHxoowQScJN94lAt8eEUo10FjKZ6eiEDJAt9DWaSzetLWm/Gyk+aCvLQdYIzA
YmxQ6c87oUzMtrdGkWw2iq67MWbF8h20svGi3ZKTKW+D5rtvRiff58dG/NsSAkzlGj9p3wCJh6VR
MiM65rsxjaWRlQjoZYaMzCzo0kcq7iDuSOZ1qUY+iWQMpsPFtPmPEhlnf32MWLrfxuJ6GRYhSeTK
2YbW7E5CeCeV21dN44RBQR5ZDtJquAej8/3e1fF182Nys8VhXu59nNWPc523CjI5Q+Dz4EGN39qc
vRafJI5htzWhQYGI/hr3ejmA6nHXpTkhJ5UY1ASUvSCovITAb25BBuZVOPA5+lRUp397EiXWx8FZ
npl/5MPvhxM9315tx68gZy8isjxejv2PnBDfPCDOV2y3IAn924L2Ye1J8RJlryhiOoTaPIfha+r6
JjLpaHq4aT2OoxQvjo4Efof+heLp0q1yv+xGKiad9tXAQtx73qz/8hb090t/QpoBZRydtMqKT/6m
VHSp6NgqvFKbm2rLsX35hbK7/AyaUTUfMNFangjroZPrSNmC5NM5tn6o+jcI+RtYOahz/afiGZF1
1VpX6PC+8jE2gPS1cPtZ4om6b26Z6p6D3JClt9NAKu8OZrJ91HyntPNg5FivCQU5betvGH+EQF8M
+q/mNvsAz/s2wnT6act+AU0g9F0PcMc6Oy1sX1o7MWNp+jEwNEcQBEp6eb9r5iMD9CzIAX0PkxAL
jkays++BjOeqWQ8V00G6PiC222s7VexOi0vMvi3PN42lVWBV8IxzY7vPu4C6MPb1LSITI3sRj0/w
LrQ5Fywk9orvVCKqnLnFUjtpr4dLmiBYi9ESoc0tJENSFIAvBJ9+MsV9qDSU3Bu8IGn3e5czGt5j
/0MRlahx67A9Jos0h8t5ZwwklcRvjs+7k9msDPKYpKhwnG7UpKC1NiLC2pTon9UUoDR2Ic8mFdvU
3jdURC0IshzDdgUy4JUwXqdXr8jkyZJvujWEl0trt9Ikfv0dFLqqqfPZhIO74FAvcYyMR8J+CCBr
Trjbd/g/7wGfEWkC279uD5ECQiwz5wBzNMevWXs2rSHK2868q2DPzmrQaDN3hPZF+VXL5172NfCR
j2Wftg7Xvo+VpBp+LFkVz0h9L7yiIU7z5ny9R3+8tft+j8hIulJxaY+3dhnLyRcaPwkKs0M9wPPu
Pk3r+77ngnE17N6LJJ4oRwU99r6gQJLiCtwiucrrFvmbZRpsj0e0AHFpm4UfyoZ3z0xFDIkOuPrn
2gKXkDdas6P1rp52NMEfy9cxEB+6ztd4HzOuYByosZhykM3Ss1lEgcd7Cxn2WbNDy/h0lwC1NIV9
pzvr17zXlDPVikQH8h2O0AA+3Ql4Km4gWXA8DfC2yrQoCcHkQOOkVyNsV3IfXQS6BarOPFgjMggO
McVs/FT1HhZy/syzLfk3P+P2YGolxsDs9rJ79HNkAj4bnJ0vT8bQzanwv/v1nWSjcyWKEpudIBmQ
5cgPKRtff7PFzjZm0vTfKhnNSZMrTp1BdHMHtwWUYUISdktHeVvVvxLDaEa/+WZJfsTctPyyTzaG
v3JtPpV6dgDYRXfQavtQk9CHqoSyxPSibHfNyz5N0XVn07rsNXpCoFk1UzkEsotu04FE39lFBK6l
QiLUPmNEd6UrjgF38Ix6qC+oZ9FQDPG2+idTkzpTqEV3czCiIqG3MfEN6/bxMIPo2ecveSkRt+Ho
YyySj5yjumQHH3o3WwKvCV+xeNgaMCQxQ04qglSM+03y9GXM1LqPF5nILF3gyjFXtPCgjHgspHOt
5zcGfwlluxwtec4JBo78958Ns5G/0KXzXm9PB1HIpYM/waQXL53/4Sm7Z08oT6OBPQCOKspqm7sR
SA7DoBQBwEjIR1OjDvyQ26L9UExtJwfMQV190McTJyP0ZzPDp0vR7OfiBSc9xsqkAvyqgoYjuQw+
vDlufAWJ8JUuLqsCSrv7hnuKQhyawX71l6YRiH1Jgq9sBfAzSoPkN2zaLCQzJqThhyC4WIi9iQ9v
vkY6+fvDC/37JFZDnb3Fn4YQzDaUo0NVRjdUaY/fuT8pdSNsTUS+iC61Jg+PEOIzhY/1RukTj9b2
magYDN3/R8adCA9BO7X9kfwdbAVB7GQJ2KrWrceR39DhJnGuDwgmowbl0xP5QeyoGQN+lQXQZ7KR
kBjRBTInScZHVtX/6l2ZFPMZKfstcLqTZu7wqkkBFX4wq/1l2++lL1VhCiTNyvZg0562YmWEBWbb
cc4FM1FMN9WXUVyWFElk5Sb9q/35bnCi7qHL1trHHdQYKnojndPRxbAksGI0RSJ573INlAhjKbpJ
qAt0n6r453vK+tTWTyowpvTEqmWRlLjY8muWjXopfIkEYvHV8mN5WItt7HmN39m9syAv2glgAlbE
iWV5y+zIsB68HS5ol6wCSjPcz0EVYHsiawmdv5h7OJr6vfMHc/IRa81WoRyAgjZvHYIcfVqw0Wwt
TZTTDtwFemviCgfNDXDD17zZCGgIm+5znsWR0eNivOzBzoCgQwW4Sl6CfZb9P69uxJag0qpe26tD
mR0SWSaClBM9o/exfkChzM9O1lxgyYVC0fdPWYaSqm4X7UPOwIE4pyuG1Z+CXMkv+0Gil8dbtADk
RAehZWs1pYn/WfLaol4D2QdKhsNTAMU0B9ZEz8J+lh94G2vHiKzVCpjBrB3sUcn9E/+tuAwOimfj
qjHPX31AN3jEkJuJugChWFxDCvUBdChPwmnvEr2mvhOPWu8WTGkvzSvVvqyesO9i1YgdFPUIh6ts
Fuv+uz4MidOe2kxmgj9NpyAaycfLVsabgNYCYx1jckKvguDyq+zz8tY2/ZNW3mcDJXFPkjPjWb4W
CKxQQgtVSzD9CB0iRK1JyASlMZFC+F0wn3c/ejCnJVYGDrMtHn10EJxmsIohDCQtPsy8au7+CsuY
pao6sPjGLRGCct5SM78NB+x843W5lp2zyfNZ5C+KjGtn7TX6ELB1mWAVVaTqZWffOlwfilFztTeB
OYo+Vt4MBNZ1u5qZidkbGdvbRFGQZ9tlp/bxiRxplPK3nzyy7cG4vyB1BoqrwMTnPr32sHRbv2jm
VBLz2h5pssCwR4U3t+wRJ5B+Gl0tZ7ZPHTFksq3z6qOuD36LTN9RcNjBLhCDgZ49vd4jS87sb/nI
wX0e3IwJOFVWB0Xw0+x8xErtsWuDuerZeWkGLFDnP6bHrwAXvyH0k9dvZEYbCGqyLfEuRpUKSG9C
uQoxQ6XVQPo/vgSEljDw3wTUmdvXxJkUQuW6vndFMbW2+fWhsAxZfEgu+lQMT3BkTl4tNJ+aDZiq
scBILpkQAkJPu9ZEdDqRgX0Uhkc0Sh3G6ZgT5EjcPXplJYBI3C6/qNvYVEDFrc5H5ZucTLgzFxQU
+n4sNWdilLsI1UIF+tkpbIwb4z2zhjNNXhtipDcU/r97+z84rf6ymmPe8h4QQp9Rvb2qlMjcN+Ly
EW2rt5K7hG5Gc0JPvkjsxJyIrY1lxyDYKUq7y+RkKx/VxeOWyhGCoHRqpsRswa3TT0gBAymQt+TO
mfGmp+69NKWBQvA4zlhZiQeUjtGo0h0NE4upd8++TBlDRxz5M4esyh/m9Cow7Dxo7tg7DtGcV4ye
y+KMN4vdMsg0/KZmGjQ9b+B02Ray7fVJjZ9EUFAFM0SbMcffHfTslKqU4I8LbOD0379vdtbgJf3s
qhTH7/hxoJKWiRLEaeTdBGbdOjTtFa8W9HEpbd8XWTust+uibUaxhmen3h+dkRoZwgY+86wOYf6K
mB4OwPar/wCd2LoLNPkw02IXtv7/7gU5TBLw448NSkt8PZh91IWJZMP87eGkPOzngINvNeO56w6S
C6Xcgh4DrK4X3TjhP8AxwDj+si32B5F/K1HpfaKQL3xMgY/txht7Wfs/4rrv44WPZRwtS0FE3BF1
E9U9IlYoNdYrWZrAuRMCn8OuEhl9LBALMFvZ3NEwpmnxQzHk1Wt7SUBXS49f4eKwy1PVc7AJewDb
bV4ABuVqkdESbCcLQWFPoT4vM7bpc5oj9Zt8PXu7FvAGtC1+cVIykA5uVJ+HzUbftHaQMuYrCWw5
6/9vmx+sRLPA75rYQriE3k1U5mjF2InJps2n6H+zQ/n0QvaujM7BZaNwOXFEUGm6HcoHTKav/n4M
K5MiXrVGylCB6Yh7L+uG8Gx8YASQ3/z/fi+Mwus8kOppKOaISbdEnd5ehuzQ7x7iFo4Eh4Oeqr5B
aazgLRdwPeGh3zTA39X/qoopcdnsy5cNOTimouOhdhwiQzyNcGFnNEDJJTHGGJZCPx50YmclVX9p
p4zwzlW+i6HmljCKLFb3RZwf63Y4+d+/ijH/LFBLR2rbgKqyZaEKAzwdzeHWPCTQOVyesOi9oOin
lbtZs6G9oOQZupBqQb0kxpDrnFDT+w/YudTMBUEdb8PYOVfnrGIuXE60oVAHLf6iJ7L57fxb/UJR
OumNsBmh534Fj4zYYF8g8d0jWaOWt3QHuhTdCEpERTzEEkCYXEM6vIomc0mSWCBcR6I534VW0SEI
Xzs0ZW+R+XnZaF6+a1qT7Lylgb9wETyu4kCNmekfJaTwJXc82i+Li5dzcAh0TH9ikClBpnSDYtTH
2OwDmmvBpyfM7ihVnqHFii/hNLgxNBBfO0l8h1F6l4rhhpI21NWnRMK/VRdYR+w00NVoqoSlGPhP
kTh3pQ286afllYH/tP04F1VGTatnHzRBHoYgx8bdf2A2WVJLYHXK4nhcAM+/vv45mO8QZQsrhl/J
gb+UiJt6+TMV+AmACrBY5/1MFQNmwajl7YVHxk6Bk3g68cYqDS6ZeSkVUhtqwv24sTwzxVNJPrN4
+yjiynUtEWX3DJk0ftsUYY+BnWEkbrrLWhRuEH17yYHMDNH2qBhq4L6kDBTL2tTJAFFS1NLXbKy0
GfWDgsGllgR7TaSHnyxmziOKiPwSaJR5SCZdJ9CicCqTl4tizmy5cNh7HUPgxy3aeNQEhagi+qrZ
IBUWWuzY6INSAZgbTdPLopfDl1MGmFRHPrWFxMTDzrNlPuwQukejQVZ6fbYKipo9DsxkxNroyurg
ZGtqCXyLcH1koQ1Aqaf1jyypHjge3hxZa75CCroMl76d5LOnh3nfeTelUlbeAKoBPoALYTd1Jghm
20mBQ2vqW4nzpBb0/QtDC9htiCt2p0pN7rbUUiimdsedalm2YT0GbrhRwA75y11DIb7bv8km8ScB
YnojtUzYEJrziGbEodsxVfikaE1dx8cwXU5Ux56s1vPTpJEcRLigRkNxLPetX8rdiYxeNVZI1fjn
np7K80s5PSZAH07eAKs4ygwPu3KR8V2EB/nH7upVMvEkf156lUaxUqw1/V0dz+OylY2FBjJy25/5
ziDc3SdhOuNLB2Mlm4V45pOKiNZA/AnrEE6NhKmcv3GqXMK3MOoSNUxibMvMrNWQFRqYQ24wmnGc
08ZSQoKrGS6HksBeDo5MW69WUcjVD6A7ytt8A4+4WC7WgA+aF9wAQIRr4uCVQuS0jrMAa235Knh9
EdwaLf8WUxiSGf8+GR2VZOT4k25TDTyakXdUOhgHXJIZMM0R03SQvpIigs7D+hqywuTz652apC7K
rB4dl5RjkmWQXlnIP9pPQ4WzAG3jAS0wH6vkXiWr4Wu4dl/DXP7fpVzlQz6QbPJygxtmOWFtHoJj
41XIBuag5oZIrkPlhMSwqX3Zu6j+qrMXwpOCOb87ht2KOrMe3T59zxr2wxgtgDWlulLPZ8zov7qS
QrYp8rVLFsOqVk9C73SQgl5xbTKh/z2s3O4sqlNmlx62XA2dISJ9XEnTr/n54Ayxkv/b5e9Rpau2
6cfySuSjMxBlDtJ+AT733zwuTTTbWKE2XDoetqCa8sG0F2pmrY0Sgy5mgfFYIg5boqIOlF0gnlGi
ABfjeyWwAQmXvsc1MA8KEBT0xFsiaphIHKIiDlSaKUuUGCkLRDQ3D4nC5ivzGRMQ2MVdgmi9SMsR
mhsyxugRXLp9hwYG4ptvaASBtXYvS3EC+g6JbrxqrT9oYCKFbBlY9M8Lfd7UAsW7mOUJx13IzAIQ
MFKwWcgAR1AhEXeQA/Ydp6OCPuMCCL4hUnipkEg9nJ3EwjaHmUmMWb9UJ+YwFQpnyhwsl5yjDBa+
u5GOfqgqYYU+xu0sfKbp1J+ns9wrdUtnn7CTDqjnsTjSib5CcvArXWo2CrZUvyUaKZvqTPSLhn87
mIFB2OFhVxsOv9lzi7+l9Um+FBWWD84byAp2XdzgGhFWorJVrclPOywdNutZch/ylFkC6hY3DbUj
oW3SQgc5q8BKo1+EKhcYQGdYs7+2OuYoZYKgM+53wIm0WxueSYZMEyZVwHKVmLNtlFvaKRST0DdP
YqGxY0CBU15etv8HCkZlVV7xTeYHIx6tgN+LqLnhP8MFt4eDm80NE1sFukgAr7sPDQndP68NQRwP
Q88Js/vLUnTqPXS/2hz8Lr6R6qpYeNq37YmGhuQ6JtLp++2clsPOyiJU+mawAM1BxHz2PFktU0vZ
s9nrpW/vsNrLwjjueAJ8WSA+aOBCnQRBcPIi7pkSGJu/5ENRhV0dkrQ/rGymEivQCox2hijkk2FC
RLbTB6AfdzcV5jyWKV5k8R/zZ2S3yAmSAxDsL4Ma+rkM1cWDgvrvSTcYDqmvc0MSaeFKxpw31lCe
bX3r9bOt2k+8pewpT5Z0y7uWWE7QW5a/ogUewggxL9vnwlrU6gjvDwslJ1qClktdDi0O36hrde/f
GVQYO4wwbH7a+aQtvfwAwOVPday+cLhoZCWysyspNJi79+90rqeaEg/9/9onfQiJmN9z21MnSSvr
r7eJLd+T56ZyUOaPRf7K5tr7hfeDnQsklXad8gvhkw9MZLK338P80OTCUL4y+HlhEKgSc0SBwCDC
lWRyYVQbbl5bREtE9OcCxRdL9HWf68l7PKQQeOwctheB3/RFXYpu8/mh3HUBVajUWSwxzLXOzRqr
nKObeEZRIEWKdvSxNCl1SfznLA8mcH+IccrM94G3K0jvRepZTIY2tcilt3LHghrOXwrUSZyf3y4D
KspZ01e/pcZotyelPRAU1l6luS23NbCu+N8Vv93Hr2ko+6r2FvXhprbI9ctnUdygcL2cVxKYs7Xh
Xm1MZqOKtBH28YmqyqTqpi7kgHO5sf39IWZPXoKbLu7zriojsMOW9FRWacjXGp5wfCqIPcxYpKYP
+H4rJubRVy79HZYthQ8+8Uj+8keb2dchSQq7Qpss2yeplXJoA4wSTy3+oDjwBubZLpgaS425Ss65
aygwSLKPfuvk32ViuLvJ9E9LYdBtDMp3JehbB9idwsCJsy/hCtpkHCPGNClHZF8v2t7bDr+1b6/U
UTJpqFmRESpr2+wW6xwfIej1UNR7P0fozObtGrf5t3KXNsa1nCw6Yqy3wnZdrRUoTJq3xZWonkCP
XSQ8TeT1ePyHGpjPJd6/oZoSFuG7nXkoCQttD6xTI+aZESIIbc6HtYGwpxkpjDAE3vsZQsVmXeVJ
8BmqRZVmUYuoyctOM2MLHNZD3jle1o1nVHxTGcM6jOkfjzSWJ05f0FeJCrZmf7xRFNwJoWEKBvxY
F8ju6ZwWfTV3FJOjayFrfy33NY5vWNMvnzRgohTOPzXwbm9biGi2OO8EnKI/0D3XqyB2ycPGhyZC
+K9fT3nhTVyX3A/RVVv1h2HAeh4eFFev60aDQXnqiQyn8kja0GS7iO6Vi8NpiSj/769CHjl+sYgc
r8tsUwmh96K1LARrh2+cPAc7DIN8zlaVmV1968IRHTCihlKGxr8r563MxqNFK/N4jNVi3Muxbnyh
81xXStANx2YpVfRexZGWe1L8v79TCMzbSzZvXtneiiYPTKERZITWnPOisePQSg/WZ0ykgPXoiUAR
zLO26kW63MaP3UJlyHaVG9wRzumkyt3Zq5R3bQ62599AAHvebIVrRBzNh8MLm1PDDXGwjuQdinmd
hMbf7xpijNtQcsnJhVMkl80wW5zicWJdJM1+432eyJOq0CJAsjaFM2TT69uCFSLdp8ZB7JXzTBk3
0kvnlbMtwtUJ/36MrVtab0PCNlZ3CsFGBmsBYgO5d1lz5gk+gP6C5wagqBkwkHZMEFQ557iI8iNZ
BxGGp1yFaiOCSHY8s5Aqkuuj3jMlTtkIWtNcdidvDBqKyM3O8A8Qi9jfcDYOT5zIXoFNZCJ3WKCT
fnkXjHLQTlCUPF2LOe2+XP7jSPSn1qT35P0I3/0XSDnArnbFf12E6JtL14IGckJv5MLkfNdZJO9D
r7worcUOrrcGpJ2EIjRlYea4kmj6bxdvGGFx8XAWH+gG62o/cp4bUD/MP2nMzvskonAn0f4pA0XZ
1LLqFMWajcwQS95Et1KdPySAkE2eGyHFvVcBqO5JoL5Y1yb+PxJCTB5MUe+JqZssFViNKTrb5vmM
yYsAWjZTVqb6grXwhHqwjYvLjfMa82dN1a5U+d+XsY4nRFRsdObFg2cEzfzeuc6o2M6CARY3cR25
mViOhUDYl/I3N2atmaryAYutZG4j0S/Qh2CQT9xZcykbkJK02JbUVfkoJuhrN9hTCQp/+mSUhQQT
0tW31o6JYL7fLPuO856VeaD+cX1oMO/N4CKXd8moyN/7+JCD368ybLEmxxo3UzHuWgyMeHtp82Pn
kzEUxbgvGQ18L2mNHOjua8ogrYCic+1rNMERNivs1L+EID3UrBfevAK6M6UWGisz98nhKtdp4rRu
dFl9eVV0rtluTEtSGZoD1/L4oqDRSSuZzIU3dM3u/BTl073MkQWHWj76SsEg3uq+NPaJm6Y3FJHu
M9FpYqwrSd6xTvMwQd4nHro/uQLJRJw8+t8Q+DGekRg/6QQ1QzluLVQsEDMwPRclOtf9r6OGf1Vi
6TdX7FVbLbt1O/jXV8XWscJ3zIFQSX+ak4LW6ex+3uoBNvEOlFmqqoH791IGGHp05wjvaDMEPX4Q
LbPXqHeDRUmkFL4kwctIFKmMMIc+Hjme6j65QMNo0Sad9Ur8Dr9nSlAG8asW0vTLwe0hD1QOVcgG
g/ly+W50jdKFuDIplBY46Qa/qTUA1Mc7wizn+wfE/empumSvSXpFA45ctz8ponWc7hLhBy+UcUhm
CcRW9QH52XuDd7AKMaGoNj6LTkbOV6lXiHa4MITFgPh9jTAjDIh4MNd8BYyRnWtIA7I1Sji6JsSr
swWZJZTUt9LbYF4jc/y/Ko2idYpvj2yVvUqZAujmwN61JBJiDvBQMLPcokUC+r5IRCJjwbF7gSEB
BQtujGpoHNYtk7lUi37584t0wJFYI1TyvhI/Y/mmte++6b5Och3P6TKwBCVcmtXyTdv0EvFsCjbv
ueNwT8Ag4zXKj0DbM65OBFMzIsk7pq0revNmBEFRGDCbOAXMq7hn9DeTCrG5Azs7aIXg6o8kHu0o
Qp23QPsX8VjcN7a42kgm1AfwTdI0jamZW2CmzDhh3YbVxz+KhiIzH/lInAjIOM8Dz5syvryZVeFC
sP/ngl2PNspxX3JASd8EPOe/dyPDdu2qvB8SYVAtwQ04/5vSRejHnyd92rS03nTULvYLiw5StStt
DTXk69G6R59KpptzMsp63JCHkl840th7kgA2FxCpK65Nkal1KysA4ShOk948qF7jCel21Uq5uXGd
hOQgQzqjx5NM7VuExIWMHAYAobP7cVoEItDuR2HPHAp56CRnfnX3OjJduU8BcbNIuJEtm13KDZrf
OO2TqJ/JFwLyEvCtf2zvTshVhyxvAysnVHwG0OUU2DzX9xaf7YvTuFUMlqc8sYvYEQJmBRJI6Qkf
rc+d9EkHnpHcB02FAGciwIVg4yztqiwWA5tDHzk9S9lxXqGHc4LrsGKY+Dw+pEwW2Bxjk6Np3adR
ZrdTTFTsH0LcW7p2JxkSMbq/s4jkeT8n0z6o/XaxnUJkgoL/mwyPLr57YqASGnBjt7OuUiIg3Mps
bzWBAHtegNuCgKVR2McrTCNDF058fhJ51hMK2a0OtJdDfL4HXTjDM4BxiUjSF0e/2HgTWb3KZOgG
icxZsYuTzx1RWprA/bbjEd9xU8hWZQCdVfXVltQzXaZ+ra8MuBSS2iY3pLa565+Oa42s+BQYZ9tO
bUWvFv5ZoX0dwH3cccE0HADCJ/Isw65Y+9OJ4Hum4sAJ3lncbZEffK2lieCvhJzhChgIWf5UwbRB
HBc1Zag2eRUyF4QWkOhdDt2LzqATMA9m1KIzLAcdpqNBiC1O1epeM+ubpwh5O8rhkofp2nRdvhes
qbJl2PLtxOVKqjE5yWf2YA2zkJUMn9/UlpTYIt/mLXzUgt6V4zEWngQjfslApvRcVpj8KURejHoi
tqxLonHZP4I+xi8aph9V6ox0k7HPPav3J95mq7ggSiGfZUu+ERiqXwpJo+UFKJgUH1i6gPnicJTQ
AYBhe856FnnMmA7UzJyuo57Yv99/4AHgAmP3TlT/5vGrZOR9e78N60ft7n0kZ2C83Ql27PbzMb0O
F1IWJr+hJAt9MwNzkj6qf0zQO22Wtl9m/C5hzmaaL38rHtK3sBibpuHoPV2/KT3vOd3pM48kqtmy
Lq6NHWGz4pM/BMj1ZxdEFBBA/tl2598rhXFHoRYqvxjD4Md7hHcWYUWTlASbC3RAJVBSj13dqLuL
dALPEZe5C75RNQqcW2hriQdlviSR4HidRfFRCRO/l8yJC0alFuo6ZkDYXi+M/yZui9kJ1vwO+3rC
kc/7b9wTwQfs3IRvahYRH2P/yhEcN8viw0l+lUvFAiwjr0gD+kOV+fdbmqsP+L7eQ+aNnwLo5NG2
4wIxQqFwst49nz7zxGbbNIhnRFzdbUOHVxuLB8FAOlYYm0P0KntWg+1kw/w7GaBlMCtlg5GWLz1R
9tABInZ5r9On1xB21t1GH7HSu0qf7v0Q0bMtomtOTXdRvyVR01kJhh0tq9Qv0CQJ8hSRVNq44yvf
HIqsCl49l+BVxmuo/1iEUTt7r26/qM6cQTbebtIumGMWKpeDAlZKEiFtf2gK0OGDsvPfZy2Zbfzc
FZcRHtMVSXUnhQUT/HopqQuucTUwHWFfYc2ng+PA77HXhS4DTeGfIegWuEvqa/01shdxzqmk+9EU
7wTKkM2YW3r5GbEqTkzR7U0/pvGQ745pWcuwgehz1TBo5FlC6J9b5mA27MeCdgzG7/D2Eck4Xh4I
rEVD6NMkEof/4MGT2Uea73CSVJalSpnfLdWm2JjqLVkkinm0f6ZeWDcysdJGOISpjbATK+3tcR2G
K76zj8o/zLgxm/5KhzIQ/vM/6wMfgU6cHIGBdKsHTGwnkUL/RWQBA46vm2ehYTOq9SPb+MVTw+Qx
dJjXWEiXYoofnzLZ1FhMxHXrzu8zd3nswH6ftwLaUp6kkQm4/ILbJy8pVM2Y+Pl/IDSm0u3/79Ii
secMAe7kEUEYoCoX/15GePbnasgLONEYNiI2WE49nI+oK3G6T7JdSOmf5DIhXhQHTMwgSV3QfxzG
IDZTiEaYu+dygXUh6EVvcliRC4BFkIR9XIymrvCAKLbvSvm9YamjaEKSjYMy/pDQszLSyYt9DHIW
R42Cs0fzlE+aG9C7FjwlmgmOo/Z4zWOaQRV5XH0DE64d/oAOpcLbiX31gOzkqBbO3XJS8ag85FDp
fiosYJGq1NX8D+jqta9VZTkBmeA6WJIirFViDW2kmGJKjo2UgsTUHvpijP1Z45vloKvXGJhXwY5w
BrVtzLsTfiLOqWpCSyBN4D9MkDHvNeOmpX5I2kwIhfZQgsiwFqE+UX0/qOh5A1B5CrwCfIg9YJFO
/8dBG+I9OHd0bmvLvDiPCZQHUdvJCyfKTdZU5sQrlyyUI8nQOGYf9Pg+jnsd1aBv+WtkIaJCpC5Q
QgNCWznrExoWA1ADCji490TggRgiTm+SkAoyil/mHbY1n5uug3QQrQ+g2KENflaQaZF8FRiXYefm
1v4wgxxF4u5jr8EcscBfvSslZBQfDNCwI6FpLU3Z6dPcTFhaQO9d0Gw/r7PjVG8hpM3RmiCORN8D
YO3wCFO4j7VtOQmCntAMmmSXBZ4fFzlysEZajBVvbHzBLAgc8/CzBqmuYJdznhPNF1CQN07fGsn+
D4vIHr/JKl4iMiJTn7oc5+vzn6WTmqpECv09w/UTvu/4zO8cyjeoTgrn3s+du2W0/nBDratPaz93
gQgQSrCxdZDTcELevEgorbXFSxvzD4NqOKCz98laJfM/SnNXtdRn0TvH69UcXuyWJokAaeNxlHpP
i2iTUOS+2GxcxKy2NEeQ8dLhbq2D9K7rvChbfMcOZ58mQqhS+G17pYc67Uo8f4wlJsrG5jGhgAhs
j4nkoH7nf5hEd35iTONxGtrLPHVQeoBsBZw1QU9gpXSMPBR7bFI+DppPjs3uA9cXNuKBMDWNL+Ml
FWF1nESddnBH4JC7KUF485+z4JYSubyoFm71etI6mpiFgH7gNgLLleog5oVYhuAbQv9KebbMv5e8
BkybRfwTjuXb/ZulKhzZVpRvaXqtNIQU/JxNRuOeUZNyjerX7TPHA51Ijdl4tguaLBpI/sT4Wzxp
QxyQcWnxAMsNlkmVHTaB0g87fB3YI2OohABQJOiAHWUCjZIe5iVdNdI7QAI/fIlMckpfhVyM+1JA
pY+r/BJG1/cen1MJLMasqNxpWxIzJTCHVCqAPtrpEO8/TE7XO8dBtvDAUiMchxacoN7kYGPbUQt5
vKSlwxvavQSlcl3wLXfvFU2kU3LCXV7DrfGj04m5dN0muHZNkKwPTcR0d+eP+DZa80EzSvBsvGCP
BIsZEuJEDSI73X6bbbO2E//S8ul3Cpnqmmc5Y1rutEzVqU5zQfSnNyFBEmrSxL74tJ2PTI3U3tJR
mTvM58pz2cmwr1hz2vm9v8d2V001B/SZ2OYzALZA54W0K/+sL/70IG+ZBC07Qcu7IJK1ocmnUzY5
rH1aUlDqVORw5fs+BX0k5ODZvRKt+8X8TplWktiwQ2vqzcAkCHRMyyD7KrvZoagLulIqCcYif6uE
BJYxG7Iy4fl7bOS1Z2ip33ku8H7Fd8RwYDivq2snh5dspgHkh80sg5Wsy2GPUH1ZhohEc+u1wU2e
BP26jSTPV7Sh9RskUst/GAN3v0ejzrHviSkfiE9zEpQw3ZbLmsSFuugjN4dZcwjXZh7pcGBC4ZVc
rm8P7ASdEYzaLW4n/wlATTLxW7wwm/YkNmQCaRgHdJ+1TZ4A1iibZ/WmuqKvQt/x7PqfsUaaLzag
+4X3c0ONxmSAffq3E1/wkwN3B2ryi7dZMZkzwuUdpZJYbOSdyujYiPc1ZzZrfuXRZoFQA2DR4YNE
4ELFrBWfvsEJ2r5AU2R7RRfin1tHENEkKNqqSpEbrLB470lefKi5tedKw/JIMydae0s5bAtkLQq5
VV6uxUgERkxde+Cu0SWcRC2pSwzS/Snxbw4q/vQgzmTTAO8PpeNNtwKZr20q37fktvtFya2TNdGW
qVtcqDIWO5LuJeZ33GbKwRiCL3CzasiKKpaDrlu8NTtOyYUmlSaCJPfbDu74BUQ/2BqpSPuSHdX0
QG1TAtUMTQEhMbl1M0xXzt1s9w8W3QAFFKvCuhV9bWRQ29czKxWmPmpuhnReSG7CBOV3+LXi6pFB
U4VtrUNuOhCaFQEP41FGuSIPThQmfEy+BPS1Z5pVUv40AsyN94DwKh5mxaqQqIYr1ndDf9zeFk2D
r5dYgTBZsdDGZEKUS7/i7aywNRzEOZnOeT92B+k0Qs/GAnoraiCUK72LXitDczcBmV75Nc8V2xDh
mQdxtB/corInCDd+aNq0jvcbMOuyGNZn0kUhuioSKubAVShSS35P/SpF5Jd7J3oOA3xXnj59buju
lRgMMdz2rElWAsclsfjRLGcWk3BxpYf3HCU6UMldkFeALYLDXyjDGu7a2p8A5/o+MzOetgRyZ6/b
Kgxg7PKUs/mIdAgTmMhX8+Ifx/dRsc6+3ygatBty/fxFzMIQ+b5Bgh0COgPG6j8bGXq9gk+6dwmR
b8TjM3uplR5U/iUy3oLs0mKvlcuWsuQkHJ+2E5yMSeU6uxPHn7UD4uk2xkcDnQGi479o/Z8Fdtg9
1EHmod1I+NAh6fPwVszhRkdyJ1fG61HAcyLZ5h9s0y+ooF8jNMjzfRZ8r1z9WTKhuEalFzSIHO+u
EuwrWJk0Tl1SYNb7MOKy/gqKI+oSn5cnq3TXjz0Eea4UyhTXfGO1nCaRQxlclp/6MGwu/1bDTs2C
yCdzk6Ibc08/aaxMZgxqiILe0ZLCmMd29+1/s1v0XbNhrg+pQE+BWKlKgMmkVppABzW4I7j5/9Jt
/uOIVjAuLZY4MBnDK/48sL2qkmbhPxwSO3hIWfW0wWJ/FInSFiOxLmNaijqlWy/Iug/AllLBlV/f
j3OL8uuJua7jT/57lvQUCDfCWXKi41y6BGjgEp+j7pDPDZW9h6L2Ll1f0cSg9jdhEhS0uOW+LpbR
KXep2ufTO0ioyBZiEOZfxwqM+rUc2QOjOd5yyL3acPmTe5C1ppAy4ZH8rNJhoQnAlgYC6Awp/hBZ
1HtdnhjhvmGuj7KQSAJwcdI/TDSTUQ/AU6g3dDBWQ1Xp7yscqvbwvlyTLNogbFCXO31mi+2SgoPg
D1TFbnhY0MFEOMvPO7BQWvhWqyftVbuISkFqVgxefOs/EfbrwVmfjzllicutIGemL3c3cjxGxHwo
WLU4PZ/djDh624j2z2ky9denloIblhIEdGb+qtk1hZXC608+17ZQonKGvu+ZeuHK3He8j/QP4tod
GlxeGYN5Yn7qpRqfxQ8H+kPlupeliCm28KOH2u7ug9ErJU2z0tZ4VPohgMpsdLwpXcnyl8CpzICc
44g2uwJIgJPLuSgw7UIoqzrBhTN/+1QybzrStbXj7L0XmLF3kUfSXVfFGQ83Gmmr0ba/xVGOM3pa
CKf/1Ozx4cXObsWONO9Ur20KEr35EAV9P/QYh25Yor1K2YLEE31x4xSgtp+REYdlLTMr4p5gds6E
bfiAHeF8HcSohiXo2yaiCAfigeBCjLC1hFJTf7O/BfimZBCJhvuY4bhbTpxIorPJ5gSidV8UXSkT
AMFgs41IZbOIsYTSBnEAMEV7rZFNGN5sN2n4sgP9EJCv4kpIo2lNVK56MvWCaKF7d8amcjz9Dg67
zB96CF/HFKVW/k/7VC/yyqi1gtRx/0Wy8JkG0vMpiPX6H02ejqszm4Sb2FS4MoKtByS9lTCb7G3l
k9HBPZhdK9Dkj3UW9UkDdah57tlP+IdxoRllnzfNkAmVPeKWHCB+j+N1HqZ0NWW+AGAtr7cRX0mA
Sc1DrmydBoSmoo3ZE+Ms7z9wMwJrazBIC6TwG/gfpzsJS9g1A+IbhCrqVq9l5i0aeLEAYSBWuTiF
70jC7QYtPrQ9Wf6uViLPw7Vy5pEuXJEuLjjTRcHjjMXCSrZrDj604MEixaW+cX7SE4OqsBVmURYO
Zv9bQaRuWcV6MgOmxVP/h0kBs4Rakcmv3Ar6tUzq8URE/i3G+0hVmxj4hvkOQ4jXAc4AmAc4kZBj
637t7AaAn3tNbXQkQTU1fdvKEkeGTtWzWCz8YyWTw+2gvkPHZ8wi//XsRBsEfaZM0QGvW1+TY0eU
zIBVmpoZKRtdLAkS30m7kGhTndLJ/7RFG+n4yCZwEuqfHw5pD94cvXD3aat5Pjh6GA+amoICqAUo
1S42HlMoYAafA9oXyzseHg0fD5kO/nyRKCWZI0NiPzJ2GJCBPAVN5IdpiNlIK/J1hHtX7W6gfo6H
9CRN6FLVkKFNsqx+d9ZR7n027bukFxMJln6qP/jfXFa8eDLVqU7vleiwyu61O7hCP/fg1sk+7k2c
XTu38AT78DYSWeTZNCVZJI2R/LTpOrDRa3WNPFbdfW4Nxuiub1xRECPkLaSGAb5KNcnEecYe+Ic1
nUSv9Zwpi87M6+krrieqo54qI436ONbZ4S784ZJPecz4YQfJj6SvC9NkgX/xC46MsocifEnjhN8Y
fBhBVqAMlTMK3i+6VuL2VlzkQbELuIv0/R8KWst6vRhsACVkwdSlHqrQBFw3t6hP2mCt9Ut7W8Gw
2YEYi1W6H0IHLIKyjf3/C5INl2SFa/4PrdLXC1ju22+e5WGKFkGXx7cs6h2DX9McXv0NC3AYOi65
ZWSn1+qP+dwMog+CuWg67i3ZTn94FGNRFggrlEOVFkTwcApVmy08RnF4bWlSkCYZtuBZlWCqCPWs
8u2AWMdwfDmMdgqxADXy4rzG4ZO3h5MKrMgoyJRmEANe5ReG9RIZTc+LszxrBGayBJGx1vhAadDe
XznXh+aRmCeuK5VGpwAgfbP3d73AL5PGrVAYhTe8Lb9nV4RKRBXTm6nXwmyLz7dpt0LU9k/Jdz/2
sswKwPGzcI9ynILZ3oHAfe60PPY0HNALYr+U/1LTaYzV5e3JJzuW7LAE0ZIME8yyIBX2QxG/3jLd
SE8ByKueV2bOIvtKgR45PR5UEdN6HA59fpQZeeolZiuq0voXwquxVkhgW2KYROs/UbIOyTmiOgij
PSLKtPjUnKakltflK/q7Cpgl59D9LxI+Inf52Fsw/RmU8rYON+8npUD3dXQJh1pQqxtaC6w3Rpq3
gd9B4+wHPq9ojRz3669EX3svBbEKkMNHCSUWepHRrw3xbQpyHmqbp8fIkiTRetxjp4KBB3vDAbbB
GANWAHLT628kmxCs4kzOnOKGCFVdtDsEIgVIpTut57LoHhrRdgSES2v6UbiC0lQPSGx9M5KBXBUr
Luz7FPPBmSKBCMbh5exJuGfwd5e17Ndfk5HGQNrTOCIddsIUDNcPlC0/EKXN9eH7ZNDZvSS4coC+
suh/bKpA5wOLtRw1lBlbEsTsetKCLS5RxhQ5XdK3uzWFvkdIXr4nrhIepcIoudJ45kUYUKLoxgdQ
Mx2q+3SP0bH2BRKEzSR+TyU3YNSYZgdNsukQJALp7nT4p+ktkZw1PVRhV5mwf3MDUGy/21NM+41D
A1R39CjIvGzpN1uo/ztqcHceB6vlvFt02YpIvvt/LXFi8Bb51GiWJl4FjJAHYgvlIGffxveDFkku
Nl5nd8sAWizMpL283A7kf3IO4fxLYiDUadLQMvIlwjkTqDZUlkp+HfsaSCYEd8pN0W0FRecWxl30
Dzbzu7XVKyHOQjFdHgLYmOhNAr6Pc8uaEDhQk2q2P6zEPl3WGZaqW4TMlF05HP8dbpY5Iz336Nd7
lpXxu3IsZUVLH7HiIVHlGnL25vUAT8imUe43zjjh2xwIi7KpWh+Pb0CjHJRnFNdkdd0fVq0OimIa
4Y5F87M80C/hnNHASPrryAzQRzXVg49XlXBnKM98Lqa9vu2TdqsHUuf75r+1E+Bo9CfAVrW1h/Qa
cJmvL+TKe6SbXMU3fcQGULUzDjpOm+AG0Xi9Q6PfTtTauxqD9QNQ5U8oV0l8yvF5zZlCV+kks2gZ
+JT75HWVOvIm1ILnNRsSLQ2mX2eWnokmPSJWnQBwW5hpzFftdbMBeBH16pYcOFbczRtgAii95RVb
pOLvC6RlnpWSnxyLvp71DM3IVKuBlrwWMLNaMShKm2dtIHZ+s6pTzZ1qx6ThQNe3cBd1EKASMI6c
IX0Ta74MwNWQCKJB7WexczrT/QCDrg+rVFM/d4SbbieXzTz+5+TuvLd721XMfQT8MfgZb41Ik05p
jfba8QADT3XIusFiT7cnCPVWuynmtOXxgt03SFahcjSyy6NARsgjEZXOxHvXw4SOqrh3RFnSJuAt
l+GZ+vwpyDJaWwkLoSM+mQBiVet9Xzl/tR7M18tkLkylsOvo6e/2o1f6GeSLjYKzBunca+fXA0qS
EwyaAfiGBHTL9gF7bRD9QxRzDSPXDdnZFZGAIj5OoajQjDjoOzgZInqVHg/2txyO9m7g5hESGco9
H/nJjgkEHkwR7GIUG++lL3d6X5HRlx+s/AG8iKeNt2JWMvoAVOuzA00wEExdV1nD98Y54UUOTOfl
nPgrSAeoy2g4F7+nmz+zj0lbh0aWKZ50q3clixBFOklmRLt9vKejbo/11Qk7gRSqfTfEH864BS8S
WMQD59h71oCCebV5Q4EIZ8CzbjHphcxsXrXcXuK0mYqeFecCkBjaJw/h8v5JT2WEEU9yT+MAusfv
FfhUyeEBnJLPC2STipBNnxVViG+6GuxrJNZhFsJrMyjf3O35SnvR9VnRt6l8D8lm9MbkHjzdfsrh
P/VvUdY+N2/Xq1CiNKCVXh/ZwEvg5TFMpSswrbkIkTiPKHoE38CjX7cLsDPzczkmN/EmIuuL+mwB
OBd8OI8qqcRjVCm+/slptmq5m7xE9h/2a03ee/b1db6ReoCXvVTZ5FHyvFASYG4zNpwrgho1PewP
SxiuIRvdBpwS50MMewbo7eaWYMrpgmfBAJThJd2KWkwhLQNhDtRBQBG/00P3ge4tIlAxiWtGqZI0
+sgBlNxPz9GbEHXywYeY0UkErK7sZEut8dgEYoH07v5zdGxZHaIAN8nRZ03+dtCTfsK0apaSjlTQ
oGf59JTDLcnaOJyyfL1cM24CIFTi73dXC/T7GztJJnZh7IlFNAz8hVOGOv64UKjodfjpDn539e+/
jgjUnFvlFvMZO5M8GhoqFNgiDgJhJ02EgYKjgQdAaVDwR1mzN/RdXpxF09ofsk3WJ3FMnNoNGtap
IzkWzBLDcsQsNxBRcPitEBYek4OtCmOj6nZWutq8eu0It/ZiL8sukZ3DFW6nfjJeozgwLVRL4eUs
TnoL8uUIaC5wsSXN/7ozRLHgv9IldkfpqTuNgb25wkQE9JuXsSVToMeb1IZFmId0RE7vMTzdQOwK
AKjFbSFgIVz+xx2ixxVj01BFR2emAMwwJ0TFFEIUw7bNe/xXa0hg5FuScbPEPVp0KKh5lffkihld
BToU+jI5bTxoffc3oLZ9xEP+tHYmk/GF4v39RHUH9rcvKyppVbdmSuG4BzAROZfjZ+/H/uAA4YBP
XQr0uPcT1xqQodiAA8vPKsdVk19SOJ22wTksAaLhnx/126QCyzn/Gn130fe5lJxIVrb0agt9YwB9
e4w5Unu2VtQxObadlQtSLngi0p/JG5sSvC5OS0s+Y7tHCx/GSnWAeystEvueDKxQC57u6a2ein0K
cxDwyqxCp1Il/XxmJ2TLlyLx7rJwZYAJwYpHzxtQ0VUsO+A7Bsrn9r/k0oLZfms5JaKMRfHtz8tH
qa9WQksqBdgb5SAV4AsEdyoQrc9pIxPyTvHmCiBE/YpiYdm/qDPdVTPfOLwhF9SqCjp8wEDX6NpQ
p596WzRV/epL4d8V5MqtoD/D4sMk7BNJqCrahRIlD2qknI036QNasboGfYn4lat/9Q9E3v6aybsM
DlQlx4s2YWdMoaJTzhubRO//HH8hWAO9G+zxQasmQ5RqwSDs6tVA0Rbbx/8Oap57xdu4AQh0/h4w
7AtLyaa75U1KCbfVvzCOAL4gXIN9iuJiEOAt0OTPEXsdaqIjN6KxcXi/KnOVQDhxW6JcWH1Ho38U
BuqIMurLzbmDkk5lXJOiRIroTEJOiyTrtH5FVBaFGuhpvX309W539/heTxYaAt//XqETw3tZtxLO
EV4kul6L1MIrwuoNdPfdDP5zSfJtAkfx+xupCUtQNPkZwnoRs/Vs2Wnt6lHyd1vpuB6R2LqZZAFv
p4k50dsGBXb7XtRHRdsH6GKn6g7S0IfLEena7swoKdvftAkzCfjwckhcZrwXlkSQeqDBiSRkxems
p/6RR7vyg0YQZyrPY5hC96hFnz2k2flrfW0X/iC3xmx8iT2mScvNRqtf86hlhzse3bvdknXxP/st
mxLH9E8nv6/XnoMFrXVSamermgB/j3G42FXHK+qMvMUQ2h52eMtwgCmVuqc+Q+0nqvbTuCVP78ge
NB4Fu/nk2287T7TVdPO5Qd1fQfHca6aDTrCIUpR3ar8RO1Upp68bPZFoIs6AGfsbudoJfxYM8mqh
dD0i+izNltHlga/UDtTb6I2st+rYC1iydHa+99EEsnuEkGUxTSeB+V4t02JTBMvycV75sZb9ikm1
hatFyeh+Pu/3yXXl4epid4hZEabiqDTVzV5xZ60L0hgz3JmD2wCqzcnOz6s/7MLTpYR1HyxWq64Z
oTbKz9h5XUMk/gNBazjRIS7TmgsBQVkvfkIAWy8v+4H/cRd/hLyI1QVdt0iWFYW/8ZLwovHVd3Qa
IEVU+EXXvn8VcZO/DEpHwmo/pGoiMJOJCU4bR2r8vnMrwSjB1pNC5DZGVhmcDhOlVmcGnvqr7zBA
27Pi2NXxT3IYJp/VxeoaMUZt0R6BOtb4Gpo1WJN/Bi07B7H+y8i3zIwt4cxKew4y2OV/HyCxz8A3
RevqeCbmHwIYByVqRw1R5LSuM7H72rTdap/zdpNAi/AEpE79xP2kjBBcTk7R/t2NxEh1YkwXPChC
3q5s3AJCL4WwMn2Q4n52kfuOckna0q2eUOJ+msNyKvqwV8iInUrc7tXdVmxHWj9yic/4hKL6wdgr
4DiZpEBciqAAGNXkgskbx5UiRoXKxCUiJ/llsIqxo28NK5QWJg+KA/n37m4vPSNoLlVjLlgRTiMI
IIDv787JNMhgpXrXt+r7JGUwvjIG0+CzELD43oMK8Z7tmG+nPpGrzcWp+hOwBwxj+jy6ks5FGjke
OkYteZwPMDV9sygrl992USz2FBpg83rG1MDyL1uzhpOp0O5DAcac8uV0HfszsN0BC7O6daSMuh9S
Y+MWucm9DUKvVCSqQ8QgT/USsVba3v/JFKPAO/7ozkV7qYwq8U2HScHzg54pwMn5muqPu8/MHCRQ
3uQEkBF7qxDtz2Q++ZAdvsidHW5M9/J8dYI/SZv9SMa9VjiglLtnetggwMQ6WwSxEgaHQW+I658Z
TctEH/9ghYJ7SPmwgksilD41ZJmWtbJOuFnLrq1qlNIbhDhYICM4eBAabd/nBqa5dvFpU2Xo52j8
0bdbdaIA3FLZMCctNLP2mXQnLuJkk3aZwRJzXvOaybTX1mc8ziOBbN5IpdrzUAdirvPOIGE7sv4b
Q01B6omV1MpZMh9Ll140uZUX6+Ii0dBcqWS14PfPkNpGFXZAijNJSQBf5bu7pEaShYlDrwVGbJs6
7fgVpq2TARgw8r7+z5AGq1RRrsu4s7yRfgEbsUvMH3B+nvLD+YlhNR/yDDdi9GUh4bshe653iKWV
aqLgq3Wk94aaaocKVmV7UnNd9koOOlWCoJjrkEJLWgXtjrLCelenYrMF1e+91cTB7qvNfIhIYM9F
5hXk7AJrergS/V10MtRV5Q0YUt39FNBJqnoxd1jYJLP453I/xEJCyZf4I+bMv/5KpUT8DoKANX33
rJFe/JCByXcGq647O3T3QbMhx5Z7/lYYDWW4ih2SrN+2BEreGkY3QqHONQFKkZzC2IL+I3m4h8/t
T8Tou+J9FOoQCh6jik/Yp9PL7eTdGL1s87jfZrnpm02+zoxZilIG6MUGfPhDNZp/d5fxUPMVujxn
Spr/UFqFTJ9mxKfUHy6gykiowJt0ANXtqPdWFu3dHrcoGsWpw4YcjAh9aJQMt1kFjVthzE3kfmQp
yTlVdBgAgeQoE62ODYLAAH0IBfVlYK7CIUsj4n58oTx9Yymp0OIkYYpOgJD1C0BUXv+laMQZFQLw
mzOi8O7tYg79s+vLSMUNJ11OCMNi8rXWONPbwgexTJEl/SMj4OmRZZkaLVpFmfz9qN6dfEPVOOyL
X5a/NCWNeVTYRWfVRJhpb79Ulz/SXvautPvWKnwD1oz3kCsSBesPkNZfwB1VUy4FQKgn2my6CFl5
KEmZxlYjOjL7SDsF4/cyjRh0iBHNLWQL01arbWSTHPGtq72+W8du0mYeamH2RrwgpWVpdZgrJvTq
fomvEE4bXIcJ2ZojA+lvZXyK4+vNlatf1jd9UymDbSfw31t2oNm+/1vZAFbSPdWRolaR1xS9xL4m
FAKppRcyN35hWD1TNcT4no+X4Lenwrii+jCTUJuFIG1c51OxCpOqDwyFHBt6Mi5JyQMczRP2Xnif
Df1FSzEkXhqL2x3vlWjhgNzXal8avQsPfqRD4CGVTQSG+18CQKPXfMJkUSAZ1C5tfdTahVMS5qHp
eZuFegz2Qfi8M2MCq08F6R7MAFEmaZkNZpVlAGyzFdGzc55j2wZjC66Bdo1J1n3v9w2gdK4Kv1o0
Z1wCZNndPQnUm1ea89KNfQJwVGtE2BrT8zIYuUjrYRBjP7kPQU5wbx3EPA4AP5G9Dyj77JrMN3ui
ozq0pBpa7zbJRl6csWKG3iRqdI1rn0cFmNbNoXMpFUOyb6JFlbgvcQoD3BsqQESdaa2xAQ12foCK
xeOEbcJrg3Yb+6TOjFoCQSuaKJQKHqYlO8oxBQnrmS0yOIjNHctEkQSiLofIoBGwhlKZxhoMb/yw
oYFYWSfrH3mBqEUuYFeIZfHxQpLE2COquQgpPZQ8b2oxweWj3Rn6e+dFbM0N6rna5j246+4Fuoef
DvdQ2FHfJSNJqZH5Lf74uPNbl+WvMqKUf3E9qthn+liKKmQvKtY3Xex9hRQz1/gt0EhnQQjCKj9b
Xugm9Qf5ba2ajRoAGq7VbiBr0JfKdXjrd6FSTOOy5JMKzJdFMCeInmQgl1fKGHRXvGw4UqLELHc0
TYhvaWV+70BNpULIjL/McbKxnmDNiYceDgnHV70PfoJ4vfrw6CrEMxGPlVDbqMPPFQ8+shSpv++p
2JlcD+lIA0dSoqbFnPGsPimOptEd4Dk0qCdqGNCXrD4h2ujYWWHOs3c4AduFyRAhREQ1+pcfXdVY
Pcm1kMs3OMpjs3mtx5gfkPbZvupv+di7Ifan9bmDhPnIO56XrQ22tD590qFEhRgQ/u9jW/oJqYwJ
PgImVmLwIS9qjrXkUqW8odAGizefqq59qeRTiW1qdftTGv8abtiH42mubLA5zvRSMx7o3mZypkJG
0IaYN6lmd0UKWGmmWdMK9aAn2vATn3Y6gWP0874aDaTofL3+InLhtfRdG6vnrNZ+Eng8cR+/4lzO
U/hTuuhHRL4kwlkR98B5OlTmoW+e47saNus/ZcMZBS5NX76qs3HZIy+y+z4c9+1Pq0CJYOwmYisy
H0zRygzPZk3/XfhvWnmDeIQFNJE/TVPCPxN738G4JMzv1bHhWWav/HQ5mOlm5wjOGkjJGUumirFf
90FHKjiZ8gpHfLWNorD4IjQ5+Y6iVAtWHYP3ii9bYpKWMshw6ulWJIyFp+xvEQsXoO9a8xUdLCxR
w6pKmG7ocFdF8yv//wU4dT2COth4vPu6/1Iu+nFV9lIxTLtw++fFzq9qt93dfiiNpF1e1zpQ1eDI
YhY0powgGn3rKHi8rI9sjGeTbxGty57EGZ9LzKw3GLSGqoKhOHDrviGh/3uR3oUo2nfg7jFJ1fe7
O0YA4TrakdJfZaO6xuSFz7GYIpaifOhLKT6EeNuM+GHwJpreBTgBuZZsqEYG7IvAWcO3BzlHWe90
NqIwMUD1VOPJgo7kzBZoWoifTeBqLAZHZcpI58WmJFb57vFps3FhGDAsbNyGIIX0yNt0iTUjUxVd
S51gUUrGiail8wNsbF8GE/LQvzOWsPGxZXqCcK6YjMi+MUW/cyuVnniHMxQfburxqe6D1h4vDVeC
zyVHem1NWYGB6zdBmE9LoyXTN0JdbbDpx/L4oBEJFwanxy7+xL80kyl+1xnSXKMQx0R/VhJsIoCK
pxDFHmmeY6Gaz3VICAM1DhRVwyotEMXN9j1B4ZyPQLzmre6efKSY0mMayIQLj106fnXJrfCUGO4n
0+1Vh5yWMNUfGLCeepjrYCCQSIWQfpXQ/WdeV9LHm9XS6o0oavaOWY6+jhhw3fOk/qLKa2vHqlZZ
8SMNd/Yn35n8pFn1wfA/Ulgwmnd7jXqvXljIOMETQMzj4vgZ9JDOSFLaYtJTfVI/A996nW2G5VBa
zQZH7PRIOqjtA//G5PraCqcN9s3KKHrcQvoJ/E2480GNtoSOjRUX+IfXUHiXh5XOKlQM/aSmO6NV
fkD5kwrygORcWFAgJVf0aC5SSwLLWhGdN44VuMqM5C2zTwIGCU4XJ9EJIUZR9vE0uOAKAyiOEP0q
yNByPQzKY57i9ST8xiGnYbL8av9ENCcpPFAOkKUIX0vPhfrSx/HPTsEOhcA3RS6C5CcOtJTeE24Q
847Nch8iSBxJ17n+LoveRxOHLX9jaoJuwaDEu7G/FLQbzPSKYMVvyoK6RVNoCgcSAUcD158NBUYp
Kj1TjwarETLuZCUCjd303UXRVHbHYZxGCYil/dAAzcSWDvadxdgicXMwQOb9dZtMVen2+KkHEHml
x0fFg15uk//IjzNqzmfnNB1NXbkWhbK4vyz9ChM+2kqalcwPmkEWJG1oKPiHlF9DpLdLe+mO3KvX
MlUkeP8AbcIJNJOJVk6LxYX5ypVz1/NpvUgcV9WCV++je4Bkzv6sGpb3YUvh/g9WvM5FFzmvBInp
FWXMPfxOZCe37IHJBrLKri/kre9pegKI/BIh2FCLL5b2yQKSAmRXPHnxdCPKvORvqlJ6Mi3Inuc6
qrW1kJ+H5bvhRLd12PYvXsOIfshm3etR9Tj8KOQzVHxgxW/72iKwO09rD66jHJ81y74l4q4NmokU
D3DFU20uXbG+S97D1gqxD75rP81w+Z7L4JycuZIha2ZtQw7veVo7epl+bDr2IBXdrNfktjJgbBUg
GlAcWsjl3FxIbeKjtHKpe/S5LN5P4B9YNpNyMdBuzUyBqlZmOTV7RQ2uWrpFPLqZJprrCyNxZXVc
hjWKYgFwHGTnZdcKNmm7rFL9iUjkJAAGcZFgFqsD8qcM9T/VkoOv5Rn4CSLAakvzdkGiCi+qPTKl
ZadwZqF7WipnZW2OqxjwpiOTXzveJ0d0ss+GvOtGTCuuaBlYyBIekdsCo3FAcjZtDKWLQIYpigpG
xHSF7QqfW4AYCtk4o6ModhItCgtpR3qzaTdI0/xJ8wm0jg66Vl8PXOp8MNbeH0wE8edd7G9tI3uS
j6wAQ0UmL5p2G9cx4fkgn790G1+rQYi864pOW8ggqVj0i90RgPmZXV1bE9RwpBpT6T2RlTAj1dCD
gLmdgGBBu4CkvvDhGqYPQ4bIHUI9DbmdQRDnAjvzkKu5RfbDr7p5+0MbskFqX3yZxyst8M4IHd1K
m4C5id8X7k03Kj6M9PBh9+ztkDQcNqeTh7MMDMWKc7It50VMoLytoGVwWSYywCOhxpARWP7kkiyF
mCRijE5iRUdwdx/0s3I0gNcsScqMawMxQA0o4Ecl9YwAgabd0OecIFq/buDLagZQvUw6Ynm57NEG
00P2CmwKghZsHXjqnktr+o3BSx3WaCt6UVzg8dLaO9ql0XsJQ0JOeaHUNaKMK3nTBr+deT2L++dY
BApQyx9+ECb5IWvz6bNmFAdmlXwDsFHUUjeRkBy0Ak97fKCWgX71ELxoTXeMWBY8U5LxBEgEYKuX
/+y2KvSq0fLnmjYFPu/nteddGUkCbz+BIjrkF/cm/+DSmzaW0XkP3L4If7xxnUK/AWkQo3WiLu0c
4xpSyGLxy4/o90ajwseufhuGoNKOhAR1lqp8BFfOF3QXMDsUXeozm/vKfy0rgDP0RrmeAnKFE/Y6
lVY5IaKHHeuzR8iq4xopbaYEc6IXQ5NFYVdk+ql4n68yVkcbOqQDQbknRoG2cPUc6huGgoNvNqY4
/3yh0Wmf48tGSAU9vAzhE0A2njpOsydiOwWkmTdae9eCijxPfY56oq3/Yv7CWpTtxwDN2RvJt4Sd
NH+eKhfM2yBCSp0QWvQn/QSURpqIsKCJMgakfJ/A3kIRX+04kRBTg/1D6n340UPILMvGdp+IT3vd
XAeyQIGTE3O+JEZgbZvkbNANEvOJ/N62e4W+IAxgDRPJLvWQGBGmgQfiefiTsMAePXWSJwgUIkFd
VNcywill4Tc+x/Y0WKGBS90UN6uxE6SkEowxE16sw6Bl6Jugid1Ofluy3E/TRVxpxrl1lwaaij3L
uNmpJgMy72Op1t9Ou/IaUvpmNrNU6+RzCyh1FUaM980LVyEZeQvqVRC3U7r0hyb5hu3x0doCJgRl
ZdG9w9MRWmbc9/MwATn/oPYtLu3qDjQe4xCF24NpxmV6xuK+HIRxJ+eHXEeRy6yl8cngveEad3f7
MY6PsCn0CkicNJ24q5/ahKKV7XJ8Hd4lOC3vRQ+EUIm4QX9qkI39AYJoz2BsX5ye1QeBtpPu4h9T
qGaKBfijaQ4dpSeRks3goCSeIpA0dwTr3LRqYSR+r5eDZRTOl091Yz+poaHRsvu8ljc/G7+BxAxf
WUIXlG/oFSrp/kpnF1PiJ6kw2+m9aEpgR3GYhnb0HuZNx80SwjhXaCKvYyclEVYiAjkUy0wPrXjK
H0CY31WaJL5csoxYl52cJFNWPLMpP+Y6VYFgw7hJ7oas7LuFsv+aUT9wlAe0ONtv65exQkdC+ztr
hftdLjrHd27DGj9tpAxbPPo+jLnGQYy21RGPqiWXOIZ+A3pX+lQRBGcQWZbhPcbHQSVDcFhkZC+0
SDOW/SEz35aSRjksuDsWz+XfDblV8dioJplMqMCY6djCyrzy0I/Bzi+Dp/CIVU0GYRaCGqS4EWo8
KeyNi9BLCqs4W5YhLh7TzoE1czaZsr5DxnmJx6dbJld8HcYTZpVzZx0DbAtT4Ku9W0XU+VbdIL3Q
Xesz+m53e+lFdfafV53uwOz0xvANMcV+oQF+De7lJn7HWBGKt80zkaZU9hxFFFLpZeb4xlDIqpR+
bnUILoi//dGDiENgaFtf3s+KWqpU1SZToIjIBQZ6m755VLWy0Sdm0lMSEO2KTMbwul2ssepS8YkK
VPrKJ1yJKr+fH6xj/koM4/eb1hR75x77c3F2ceCbBLripU27/jZyNmOgadzIgwHcxGE7Fgt4d6fl
bQDS7sLmLQXot4WI974daFod7I7mZ3Ko/zWQBjvO+oO0sA3I48YPnpZdz8xo5jixkI3UybeVTbpr
0Q7D24Z1/CNSHh3LGO4dZtRqu3KI1vrL4Uc6dUVN/YfW4BI3uXpJa3jfElNLeyAmgZk+kHVevX7i
yd71QifZr40dmgkEkf9jQV/G2XD19ydgkidYtTSC16gsgDbapcKl5eiy5U6oLxPpajiy1Sjzi5MX
vufDsPEk+crlZE1brgXBxNJsI+93XkcvlNBFiy2TRW8kEW9jAllvGUYHVl+IM8vHHdve3VbBPaob
GHsLpZoviKM7CTqilUT1Ej8ZlEf8ok5PoU6Wcm/UNoSEqJW3Grp1C9ZTxjH/Vkbhq7WNJVOGyp9h
OCO/tk2uj3PpfkGI7iay2JVdX6XoYOnbOuyp/6aDuzLiUbErV9M9XAJuutUOULeRPZ+Ti3xRDIMl
iugSpVXayh+w0pLOnCyLsAcGBCvJ2wLsQjIB96Y8kS27w7O7ad3Mcnb04q3C5beOfp1ttlsdeWsn
xlnhbaXyJ0bJASlzgK0ymaim3xssGKRatjXFs5F0gHEgOMyMrVPJhr4BnkIDc79cZV3FmV5B9jIG
fQak3ZoUFASPTiSM4+YZhtqNBnaCMwzc1K8gYCk3NQwUDMzbDvSH/hG3K50Uj5dy+FWnTvFxgV6B
aQ0uNkD78qffW1cnDnSgBtUaaU/DEDq4gqetOa2XFcZ4+0D/CaKWExDvisxc9N91baRCe6c8KaPs
8mq/csOgYALjT24O0/n1nO8x3YDJATnA2UVFSlhNqX9CKh/qWF9kZRJxsmVZCrWPsEhyuJyZqesg
1m0lvuYrrOMnxSr4Ciicz3MdwAz/epB+kkvWp7Q/lkO7jNFK/33Hd+3a8VDXedLuud5fIer44FyG
xD5mckqdFEpvoLL4N0oY8CmXW+OsKfcC4Pczq7YZlwgGC4BC4+UzvFPaLnGsWMO3cXL7Y1jOEdfY
HrN2Byk7jwtLs3LgQeIQTX7hD/ZENGRZumOVp83PnxWSFOgv5b7VBiSfDEWGwy4e5rg26mmrTgxE
Vo9oFU35IdDK9LbBux20NyHbzrAte8UVl6sbeVnEA8PUIuypy9xLmdOr0YkrfNn5EZN2HgZDOond
rH8cnOm4rwzEt2JTRbiql40YMEp9ihL0JoadKZJzz0k84TDC/mzpagwyx5PULruBdV2sA4Wl0UA/
nndeT+nAUJvlYgZTv+Fi3YBIpvn6qmAhQ2RNaIMk7lftt149YZEQ+3cspv4Q++xvlayxRvfI53ZQ
B7h+6lMhNm4bYXvWIqs6AyyEkzQJ+4o8B3dtdwp4FUkOvm9RuT9SyJvoLTnJSQXTCFub4pu3Igp7
cmxp6jp3XoX/zYwUwOgOSCf2NhRN6KJWVx6Bk46A5RAukaJlg9UGxMuetv3VxUX4D3cK2+tvoUvb
HRBs0l+3GaEE662ZOEOe+A+CXaKyZXh5c9LE/NCeKQxGMgLLA4Xs5wj5vdz05NtQdoD6FP2uyQ/G
yUdGmyRW6Ha2LRF9mLNoAQDq5Nwj/kSTaHjcGPJOpaAkfKAqJ7+Y8yDxpT6vJYL1HSLvZSs5dTxY
KOmZflKkjOa+/owttH41KsE+M1GMjyEUmE+8BzT/X77mXvF+/qW+GcD9Wqo/7gA6Fwiyw6LZv45S
QnqhJtriYaPHvGUVJsN0kABdsk6TWhkM/iLDqzjhL1l96OJiOvgaeDQoDb4WA3OWjItnyBFpxAw2
ATVM7npNty3AlfD+1P4eJYSA+hRPbQZOps3vZsbs/TNe8vGGBncycoXSoQG8pJmnwMitDXxmQAHP
mdo7L+KrHVCeDEuAePJm/7QtGPKQC2+9qDZzvOums2RBD1eQNI5S6KZx+tpoLEpmPNdzkkCKMfiS
xtWcixpBzHl65URSDHd/s6GGdkGyDBvDbM2KW4AG4SS13rnBCXXsnBDQnd3kdxpFa6LRrhs7CQfl
9KaEBXoNc2pBOqYg3Z6Gf2B9RdJiflHdgY2g8wFER9r9VVP3Mx9FDM5apjzTRfa1gyCB14r/8T2j
S/5sv58whBZtZaxh0QEcfyfZyZbEzU9xeTtQGvMt8dwB8NbivjRmGBf+nZy0LX37dB23KaXxSLeA
H7PnmqVgSmZLWb38FHgXXtVyMtTJWUasBr0ySzDLPArTu3ypZ7je2LAxfll4L9EWOFf/enKNSiyo
Xh0x1yWi5fjBvnJNtWcnQRWtaG5Eeh96/FhEVoXyDHLj7P4uvVhF+eeLBYP+gZcGRfzCdlKto/gd
ygjPVTc4DFxbW8x1YnZZzoEQLMkQ3TJ7s2iGoa/5JXHilwBNg/5uTIZiw+SuQzrs/EOjqarzjfVh
9XjWVsm+BvnA09iI/dCUHYxUJjqzFQzdBeWzO5mKPTADRRoZtA0EJdKx3oMJS+KuoEK6GR+4J4AM
/jG9YiURItHUBKD8+kbIZNPigdS87TjK++2bG+XSywPPof9Kstn3nuvp1GsfgO73uzHbvyJLNi0u
4GRS/6CnpsLQbDZNhTOiaXVW8TbFC+rwCF6ze5UbEkynq2biQp7+vVidXCubcpBiKK0Z/VO/IZJg
sG4+NU12yf6geCFPAGg+5RHHANslE3T9wXB9U/9A9z84bR1U3zuYFAPyPeMB8yGFMLq34mhbEzku
7tqkhD45wEwByvS/4j6bJRxo2e1xVPKlndyvqgZ9dvmpEKhklEPfhgCvo5zJKXFNSgh3k6riNg5e
FgEMsUxKQWU0hu1aMtHB7OFlJ+ftu8fCDEqM/BIr+UVgwgxZEHmjDBKFhCzwOHQYz8qnSbxSYUk9
JGoAyVxFktkrhIjLV2sKHyyFJ413nK8gRDBSNZiv2m15s/xBN9Fn60pp2aqTDoPX2wIUUFZwvI86
39rT6hZqCEgtcT0sYoFX7aABJT8koenOrT28fLLC2O+105YAOf0Mk6Dk5wBf0tGkX2KabJFqR4k3
QwFXcHbshKHKN020SxIdlOAbxVj4Rj1dCpPwLko/B13gRGvuDSJwGHyrgb7w8hM02rO34fOfq6lc
EKjDh07+wPX0+B0uaBoJggWxXOuyl9SoUfhyTGytjP/NZFy1tLUUZaXOFwjVabcuglzmJZYfPtf5
wKw9N4qnj48T5tOdvBImLZEm7zzuThBk36yFiGaY5InjoAtVwNQhA3Bf40iEww7FIV90RdYNE6QT
kW8ARSGx68JgzNBP04C8aEM6tVYx+ZfQzuDqo7QrF/6SKeivniGLSKitWdB8K0ReZ9ltq7oLxpu5
UhTFJ3xBLgTFRMNXXpzR3L+eSpDr2/5blelQ4Wf75aCf33xp0WWjlmpmBORI3t+6icR36nmwEXVh
XbWhO1KIGxrV7QfqfjvFrPbwdqNougNJAl7DkaInPNaY2ce77my6J01y2ZD4kP4gjbqrIRnbQcwU
fVxTJ2bKG3bOtQwmsQlWQ7Z+PEMjW8vhz4tfWaSHMr+RQExzoD+wcb2DaeCWJyN5abMYYAksJlcj
So5vCwF/q2g+y1adp74pgkWyu4/UEXaDmnQIYC64HG+8zw7tNa+QUCcRoycrIIqFY3MseAqD7G2m
WeY6xl4ur5+pq2aiSzy4DGWPG//Ylq44+8vJitK/BqITzXGFOWs2x8XuYU1XWPin0iefRjL3LGLq
sP19gpVFreqQzF/xlW12Hz40sTH3Gr6L6h0VFFSn/4A10Qm7X8t5udp/x7f2yPjrw4yzOoywIYts
V5W4RAG2qmMllL5yf4JFzptn0Q2BDgNsCMfs0mHMB/NwNpHh/e69QCfqwUIqfEgXF4kwRiKddwL2
9e1U/s80TizWb7dAd9HTymxILz+81DcVLJwNY1NYif09Iu0ckkP8Dv+EPzuxGY+ImILX+mFP4iZk
2ZcL3V6Ysj4YfuIbJjyU9dd5HnsdNlvcx+Dg8/7kvImFeORvkChNfFfWhLzRQGvAj8WMxwMGK7BO
Oj0O/FmJXMEfGCWUe+4hHZPZGZoQDy5JyMFTm5MK2OQi5ZBiF4hLxakqFWyXGgVsr+iOgzFcaip1
jXgDnjk6ts0TVOSuCYQGdYkMwafecR4BFb4SRiJck4XQi0gRDvUWOAi7I6PR82Rl+NWAL2HwgP1B
uMNXwsmGaWKLls9LhiU3KCO805USFjy8c/PzW02a/vY3I43H9aAwVcLwaQLTEQaG50pNFuO/MgD0
tqSGoGYvx/1mk7TEE1aQsMr1cm/esWkkhq03VQQETzdOuKWMKqmZFEFLDbOCxn8V1EF4nNkSTXhn
TPgDOMXwPf2lpkuHpJ2ZfiW9nQdCdkyX/Vug8p1s8YcACD2QBmsMu9tnpfW0Nmu6FPycmDKBi5+c
bBhZjgk2SJgMRlURTKPpXYLfY7OpNQ5Qps9XXTwoA+eq4flkKGrMpM1rLr1mUrA24VoGSLaEbX2f
rGm15WF78E4anTREr4CxZHuc3PzS2YeNA12LFDB/GdrbSrLSBqxzpwNXvN40W7TrcCAPfg6vwjLU
yT7R46GSY64dJ9PBEctRTO+N0OdxOjxa8/1yni0mFrcK1nKk16env+KXsQ1dxB5xW512rNVKJXRx
4hDLQ5ub/UEzuGuBD3mQ3H1ITN+xdhQ9RONMgdmVbwjug+P8MRpToP0vff/LUMzN1duEhoQazA+5
uUfl1etE6LFV9rCQoPb9Sl3FLhHvnOcglzAQDqbR4XZ6ZJpYSMD0EirXK5T6SQ7azbOBv0N2JgHS
E2x+InAoFBwJgATPzrf1BNPsP4bptMouZM+tRHekLGtf8gb31wjtSych19gWxtHsuYny6U5NCin6
XKS+8PskEMCfkoW8PuHjYzriAZbzUtkJd8bRqmO9GSkHOZ5n/3xYB/UX4YG7Ijgbr82yDbpftRFv
ZrPS0WDdYQHRbUTVYpuPj97YGiSATUNeEfEM7I6/54ItxBSB1WWZJnPB6nHkNjvCmBnMgkZio4C4
SZxq94d5VPy63Z+usPiH93o3SPLcS2J0uHGH3eKpLKbBl5f7CLPZz+BXwtMi0hAFsmlBU0vocG9O
+h1J8UVBu891Lhd/iqbJQCag7nMs0uUtZ+mO93uOJRRfWOMdYYbD9VKumTS63mBDsBkKpyeCZF6s
1dVtVifDnxoxd4n3N14m1HkFRdKVue2Cy2s4WCgdwrAzcHrhuD8NtrPRDj7kNODkvZ8Lo5gavH/X
wpgFMUX1IOOSpe72BJ1cpmdwsMRM0KgvCHlh1P2K3d7dMtZ1wRfu0PcpC2DaLpu17XE3NbDlSqIw
nrnF0B0J4peE/SnH9P0AyEY5LGOFmt3GUiBA06ajv+09w1fOnpEsqb+n+c8iyvGMOl/fRmtpedmp
6xDk608wq7kTG/rLWvMf7wFWoRaHOqEEl/EsnyrsoGTzZUAgfkfUYe+i91Q/7QSG9QFXan79+iA4
9xON0ZFI0gF3pnp7gz1LKSdhrGiy5Ddmk3rceOB6UubUrEuf6wUWGUiwNisRWxLDrgO6/oC7OLBc
w+umnbnG0VqHFNKCkrOLBDbYQEEcKJ8ljuFmcIx2+URD5w92va88lZGyx89x+Mr9FMj8AMUFGhBw
KtQJOainTF/CONFbaMQg3irdeSyms7L5/D0UB9en+JDuYA+4AgRznuoENWveeUWbMsl0DPEc7cbB
iV2rRxHm7HpA0/1oApdpDF99r2Alstv4m7h7doUXP6IosG9iOHkkSsXLNAzMbo8KFS9imRrlIb2j
f900AGnvlJFul4n+danImhseD8DmwgxupTUweSbQqWtGvqEZ5U0xPmHxhoKI55BL1XmZrTLOP7gD
ubyHpEjfrEJy5Vf20iVZlnX2bVgIPNQlc7Cu/NRliZAndpbwpj6sDmJ3yeVQFoj4ewfuB6lwI0/K
BqTBaxnTKveeN25RhZVwvhfO9lsSDFPxCc9h/RCFf9kR0qQ4xVkIgiZRPYfE1qm3SL7t/pRJTa0x
+7Dyu66OzujxPp0MCjlVXfuJNjnYF/wx/kbqs9EYdOHFy7BRO3TL9QuQgyvukkX/Io/kl31NOQHh
K35Fr4UUxRrxT2Xwm1OQZ5IbNj6wa+XPpjqfif4svybRZ57QiW6S/RQS2bvVvLlciB9S23pXgOly
w/XF4wcOxiWY0pFNIztI9AqS0VhbkJ5VR98P9CRci3vUIBMdSlL6diNhECbjRhOiLrfKpKSd/vns
mhOr1/znE210bqenpey9eEljY4b1n6rZAMs9E050aLyTbRDCvofloNX7FcornK0DZO+D41sdp1RG
Lqo1Lhc3I9iXCPVKR1QKWArqReuTcA1WwPIfU3/40FYqlYzaBY2LUpv38GUrTg+dkDSCJItaEOau
/PuZ72ML+skxQFwH2+cT4eWcmePg/MCkdX4SEmwZeL91S+hnvGvEC0ck4rWNJX0YuK723y6Cb/dO
vNzHKe3wIhGwf/x44UT+lDvVIZlBKcJsCbH8NvPGuRZXX2qWc2pnX99VmXm/iCVcOjewDPL5d+wZ
ezXmLBPOB+tK59xXjdMdgJVDAJ8c2N4MuTnZOi7wMYtWc3hWEuZzoIusWBvQTrZB8qRxUh5C+fcU
k1twGrIC3cIOg32Innyk8AD22hXuuhTFxVjCtj+10GHkc1VOLiaGhGIOM22KuCbWBku+tePKy1f2
5NMkDK8D/xP9nkLCJXmWkx78JcUhFqcVpLRuHR834hY9zoxTYCESx4HZOAnHxGjstV4ayt6/eSsf
UXzsLUTRhOeMuqbzuQtTBz5zY7PnCr8V1MKIyAvRvbjD6tMYc4bWWTLJwmJsibSWIANuzh1VI8xp
vIsemDDFsLNgpDp37C+g9JBd0xvbI40IU4pxNoFDXE4TmLQ9WnmI7GZb7peylQg6f2Y6R9b8rzTS
/Zo5x1pKrS4PdnQ8bD9z2C2jO25Vl+Anv3/TdMGlTYnHVXoEi5fRZS0kdymPz3FVkYkzHEYHBY04
ic4g/ttK01FRlJlL3R+UsFcdQiKMpfj1hH1Nr3JTDEX6cGb4piELugdmXew67qd0u6VtjrLw7nJa
wLL81hD9VuhZP8D3s8V8tk5ZbVCkmSXXZOjeWahgKy/YYCjyZ/eMfjJQ83Xl7kAhGrHs0ZaLvus/
GD5ppDtvAtV28YVIgCNti3x7/DDrlo+k30gGX0uCvbQ61jOrq7mkUXxk9Ex9DaoOe74JQW+AOQKg
P+ajp3aqmisRBD6GlzhonLQtW1l3CT65MbNXGBGuKaJyjs8GmrzxBfvVV5AlZp7qJtLcYRTfXE7I
t9cqT+7RGIKQLrwDfZLvFkHXQKsWuzABatL0mFvX1MKpdZFCwF/i+RSVV6u6m5ciyhAZP44W7CYx
BtsvnGx0UfShoF52MMwjg3bVGPadhzz9YIowEbLf6CxroTkxtxKWaTqQf/WUBDSMNzqgHbjiF/kp
rCu6vzAMd/mVxlBWKvfJXPmpi9gUUomlzDcrJ00o2vwO/c90yzniNU1QZ8GfI9ulice4QiEF+dgZ
xaBIcQIz17RYWLx5OLpFAlr6AFFe80U5w+EED4G4f5AS0VnyqP6S1bvoi7P6la0dmz9ECXav01ft
M9ncSuYOmYnxS5cAMGuu2IZLkqu5nAnPj4ttioPvNCYui9D6gclfG0URCty8fr8JvDJ/HH8WRYSj
cgGM3F6USRl7aQkhsR47PXHek0n5yzDhbZY4X6xYv360Fev9tg8s4B76/nPoy+k6SfoYTYK7LSx8
xkCJ9jnhJ4cmDNNHBCiZnGU3+yVwkTu/YBeRrlGOhCxsx/FDNC2dbm6sourbs+1G4pMTXdzm/G3z
LRKqyniNBNejLY9NttZaB7mNul65fM6ESXvPaDKVKu4Sd4/QM1wHZxCPlQwFgnusTjnG3ti0TsCu
SUAfQ//OfJpR/uOzxQhe9Oh3w4/CjBMaZ2Dhhm9VxjXN5SgqBNojyPTE4e2yAOkZjGVwNd0TUrPZ
rYWPKQrzH2XAHiAcxNVQFIO8bCFRdze7PzIKgx2tVjHArR8bud3SwdsRFGJ7rccd/F0ZNUKfj49Y
mA0PFgB/vy2InGiKYaBY2hN46m3BNaFPLecC8DkL1txaHDR64kJnr3ESKtBAbPNt01B5ve10OwEk
P5Kb50OLu4fG+rUKfmeQ+FN+nQTpgQGBSCAuE1ZRPUd/DtFTNSaJU9NJb3AiZR1iYVYhtVxP6rrK
F76k4acFrFVfsZ9x8B4LevVrayEGIli6Xh9MlLTPW/BAIEVIanOG8FdM5xgvFWv3W/RhaI5iahXc
7+GilA4U5V9kSSQa6Le6cDrgWExoPeDxWnOjlHBXsD8cR9kojj/SWMzarn4NVofPGyLv3Fn8/6pl
rEgj9tDtuq7VI5XWmZveV+ci4GqxqXYj3Wl5f8zA11A3MID9E/EVSt5bJF7oNmx5G3edLf3sIfcn
aAxBzpOOvIN/W+0Rf5OpyUYDCliHx/76+x/85usDE3jh5Dq8n4n0szxUY4ULNacXUAtPYg45lN8n
hB+BAaDaSkLZl6UVbGSMPAIjoYX3WtXZRdlSpXtSbwRdCVsl5uw7f439vvrwqNd+A2AMzxarW/Tl
EJZkTfYMdtV4SedE0TAvbse4QhJRv/ONlqWHWaCij/14oa5czdK8vdh6N2U1w1slr6qvU0qXzJp0
0QDgmuYvbvpE8eQgJEakA/81aRsXTcUB/42XWyi+CzBSGUuRVQ8PWXOGRNcfrqgidM5VSyGB/DYY
m8LNpeqXJ+CznHATYfaE/tO7lJ3fBHe/j+ZmhMHUtZT3y5qEY3NSPymqJGtNeijxCs1P3o3oyFIq
zjC6zyEsvTVZgHjgRGAMQ9fwl/q1EfZI4/PZwwyo65BcUsMltSth3Arcxkfs2WVsK0sGqPbdxEHd
BLkxfFZIUDm9K7JC2FasZiOlrEzGMTkhw2v3F1LApjrQA0eCfqM2qEj70TPjY3dZKNe+3ZRY+3E7
ljUMjzbtwLavgpNis6S4dDhsrO4T0UarLrkXgD3Vt1LGqnsWutZAY45WJRCzs3Us8yoOVkI2uRTk
T3QrmNmHvV7SeSfY3JFI/iQOqYp7/FVhCUwtqY/qKHESzsDQ6YtFffp+vpcfC+ct9jZkEJP/N3S/
riycyy7jgLo73DFsp194qBYTJ6GRNRUcMw5vLvQvw/iQ/+hQC9MCr9W+nCpmuTmEH9D9M0t4CQa/
iN/AmyrUOfBNKzhNIDbNvGpAXSH0oSEgP++WYj0s9eX2EH8xX0YmZ7cpzdOQjK391kG47aH32W3W
9rvzQ2t7EWxGRMJBzj/p8YN+ZtdMQgsRtiFiKJwIrjjLHQDleXpfL5wojsb/iD1MctR2QXYkbn2E
0EHW0oSBAMoKJnJyFlS78JbFiaBuO6k73DYa0DaOY/DWs+Hj7XDcEvFLIm0ZIGGSZofZ6delRzuJ
8B7SzDmRaI+F55cCC5wpQo0cuQAIbDb0UP6D83dFojCdlIYJflQwOW1Dw72voYTD3ulhyBx6rGPQ
YaB7OumsWEJNxkt5XgHmy+krA8cyxUmGqUoLxqipLwmhPylyu7yeKR+j7R7feLgwBCx8ogt3hrS2
pyVki6KIwdv4pkx+5ItYd+waBO4vVUnzmaiBX2Ie8BLKwupXZMqdqnYsfozvKz0N4QwL7QLypqhj
aSf5nJREulZ1pMB1l3r10rtGF8qvjLHMco7MytndtFjdtf++l2vg3JzvKYGCvArTFGeFgLAmnwsG
nOlWLmEJ2td181Vy6ST9RuGYLaxa8OYmu2eu56IbQaBsFgjqGr6oG14R2PZ9zLaiJiH98nQ/QTSs
TbT473iy+JpXnVzHVQliKbAgqvoIIKRphGkwcgjcU4Cj/+JbWhtxm/BxEXTZpqJlVQqoHjE+Q6fD
/VcsfV7JPCukIXU8gxZt8AYh1//z2JGfHLFM6fghYedZFXarwpjIa/4lxKSsYCWKr5FrUEGYuhm3
s2dGT/1CyJBVEaAeGrOdce4j26Kbk47RWdBw5jVA8oqyooLNOISGIzzo+hGkEmZT6vU9Y1/Ec/sH
XY5UzQk5sbPQ56dKSDdyUSVLnchIILGtKV1sk64Xib/n1ZAr+bKt3tQr3AYG+yy/qZ3zB+hxLbnc
SUVA/h9RaNm9quxUzv9CxN3DFyz248wrBhcvLT+/VPV4lznAcQe0NciPs6AS1E6P5TQOn6Zq3ZBv
rYeNE+aBN0cEkV4IETGLh0kxoyMaZhLU67THK8MABbexx8nSyjBWryOM9+gPuFQMwn4UMBqBQa5h
iem05GAlXDQBQexGDv1NGTaZpfvYGyu/JA6105Uelb230xvWVpsd/vNtRj4PBm7Tdqhaq6yLHWMe
SSvMlvhMOGzWWn1JALP8oKxQl9sIeQcixIg98idl3iKDkfYFEDbLo7ekrSMeuLLe/CON+hI5AW7g
5hUbS0F/7Be7DlnDgKdWpAFG1IoYBUhu9GnrnRZJmOwCULPi+fHfgN9Fqz0SOOmQJnorr45/eIR6
euJaovbyCrJRuEuNdLZQidU9UIpWMdN+r6krJhgxgz9pWlCu7aowa0F0RfXMAcEacbEEo9kq2+Ak
+9wXp7aX3rF7P2RcYdwShmP+PfUYX7oZ09+Gg+S/WnQU7sl+0X46oELoq9Y0lsq1OiDh7el3mXbn
ErYpyKJN32cLkfLu8f++5+BAUAM/aNaBrrEKf56WkSw7B6ICEaSySmNww1FcM42tYUThbQJnkc1B
izL92q4JWUtmpbZynYBMLlEM4TmZeJAgVJtqSdbJ9sCtQpHNnRqOviWRS9rTDmo1MS/7Dh8A4TWP
3NaCpoOjzPoxrAbwnn7CpDMSYbnJvRJ5C0IvgV2Uuwsrger5IxqtxpOQfZFSzxh7cDl1vP5i1JLs
QpolNrhC7wQdWUTAgCSYRhgPjpgcT6nHtx3VAc3UE/oY8wmT+Ng1zvAHoURV0nTMy455J2ZR7rJ/
0el4Fz7JJKIs+WVi3Gbvj3I+/nTop/tFU1hRp+aK5CAb/GtDU3lprdw7li4K5wRW1mOW9rKn64F7
SW/jnUjw/Eydz89EMZDAj79KFCqIJsvLTpPCh/lzkzdST5cWeoBe6K8ffgu+Ct76iSMZAMUILn2X
58OWzIbPHNnfjSCKyhv2vAF+VVoaWgULmDgoyLfgl9BiGuRoR1DyxKOYWaBbunipBCDOQ7FvTr8S
43/LStmFLrdvRU2PtW1HC+/DaucGD4MVN6Nu1OJSJD4BkA0rE4TrFBfdxsdDUgD+9XM0FN7rxpeS
jnEW2BlP0ltZZnEphtZra07rI4P+/f9JUD7wCOLn/IbjmHyPvskt4J1W5TWs8mSoVST19AkXLngA
/keRLHs2fVt51ByzDloV6JqRtum9y6GS8Uky/qCRRYLoj8rsyWSupW9ZxRvS8A2hhgyjCWURx96S
Bv4yhY+WfsNE5hJK1RW03Kl4GoEI6L+Eaemu0fQOqWs4IVzkIH3zYQ/yGpEIrL31b8tz1Twp0jvB
cXsLP1294h9jlF362IdZ8xk/8mPwExcxK6e0lWf8lWnlJHEV0bVTJ35AT7KU271FwK1z659Vxud7
PDHJN0rtUljNNHC2b0lVVpp96F9NszEKC6zTjwhpDMUPlwd/JbgLlqw6nJazWsVyFD1zhLjj6sFr
oHcw9EI4vrQZ8+ID/jyhP2cGurily9sDjdA4L/JPwPumUxalxK3703PBRPt4K85Zr696CX42bvik
B+W5cY3Pkd2iuy9WjueWc5n26b21CUMFyHjOkw0sFUh9SXkAjmeY5Uhz60D8CLHP7AH3qTf6zJ+/
KKhoKwbfR/KrmOYmAhk/Jcv7BgG5ellO54KEMMC5mi0ljTuHtlmELxa6lzkQ8blMHqAlKdUi7nSs
lRuF4x0gv50lU2zdWzQuTGuvUiN+twlPveMU21uKhutwwMGf/YGlDN+Qo1rGPpUctXeVBUb1NqG1
hjgMFiUy4VtwyVfDwXRUvEf9z4koolp9nYLrSh51jZVPqVgLdkA7qQJ/AemODFw30J187rZSN//i
poj5CvooqmJBFYNHX2+9ARNlShV3D2tvA2Yjqw4ifvu/18hmTJ7JBejAS25m06Q+uv+15H+2AQva
1kRLEQ38fUAQ7DkNyR0hT/W6XNzJfuYjFgiB97C/DH1ejQRs/YCHgIFMLOPSDwKMxd/A1HTKTNLH
lfAoImkrhGYZ/Pi5I011Fdp6kAM7PZ5vmKm7bb1FsrE5YG241GNMFaxHCnBo/XRPqTmFEuLadBP6
kMZZWf6e6zDJucslRWJd9mvg0bC/kQqdaqsMl6iWntdMGAHoKfJQ4DAvL7DqeL3MuU8Tnc8SVdCU
I4W100IH6zkVv6RKrunp8RI7NNhPFhGYBEMgX4/IscrIC7iU4CTV9b5KGw/PF2TjxyUfhpnKWkgo
oDIK8VZPNGOXiUGo+GQjecARC/kIyYw0QrShqIC5PFGbaQu3W95dI6io52HUrKAEh4dVlk6JrhLr
PzdPwTyY9wDHeyJsiBPT8zfTPOgagv4a2b+lMYmPthhqhX4VAzXlA9C3obaRHdYEMnSQSfjlu8YN
ecb7hzXz+GTjObhNQtJpwF6MTNtBxDLzROXCSQHmKbbiOrgmhzJegbR6UgTNeCCJYBXZV6LnaXx+
0hQGTIMbEE8La/OasFHwNa39+S80SEAlY67WMrLO2jyrL2K9UIqLt3W81uNBxFGVCqV4gZ1N+Bdb
svjrOSIEPeg3/hdpDZQ32/ZlyTz5yURGaCMZ8B7wjCRv2m8FUBqLWH2sOgR7BkH4rhzPHkngyQ/i
gQehrsqogu2NrmxAVVvjc3HPGfoz6SHcEaLs+XIFep03ysit0hMhIulxmY8qF3mNXGgOgvR+aZUH
ycIscuBa7/02i4XMI0JXWv2x1ePSsyl+fdJiJDepjm4L17ASjnpbd70iJOEX2vQErGaarKY1D8Lp
14McoEQDICxHEg2x1Be8MW6MG8DVAJgLvzaU4ICyS97pU49Hyqy/ZUQKw0+Afx0ik1vtcJQQ1NQA
6frSmL+K4EwdxvRNI1+uWm7fQg0GSDmbn5tNWSp8uoQWXtrcBFeZNG7HIIxMmxAMzNicpo6fK4Te
We+kZNIsXMdIJ1sPFxRHs5+V6LudUudZ5Hm+XblBb3nc6dbGYnNx5O9rNqfkuM2/5z3P+F3z4Oqd
9yntfdVMcvvO62YKZpBz4SLcajr96ydckP9QSJm6wOmy5ehHomKnEn5KtfXwcKRulO+2eKlEWqRU
b4+216U+A8BJyL0dvN48SzHFg/l0iqvHbx30Fi+9uk4L5aTtfoLBZT+d9MsM8Cy0MQ7NxavFOYjR
CRiV+7lNn0tVrytfe+k1IXUyDgAQsNX/uIe3IXpGFNOKIvIFDUrsT3CtMoslsEpV1Ek3G4wm/uJN
Q8GWPSV13/paRZu4KcfsZZGhjFamYNqiEPnWOnsDuQQJfOxRcoXA6C0JwfEE2YUb1TM9ltwoimgS
ncjSaLWmFoGpXFOPEhdAmiR/1uKEdYezB6jlJyYumhJoW+wBqyY7I/HYaa4waFCNucBjfy0fD08l
5BPAGH8CkndeZFeUxY8wtJo1py1IXRrOO6JZ+jMamuHgtooKzB7WaqEFVWL2rgkezjU40FRJtQLK
PdQyNcSyQYq5Nf1LAuev4rw7gMJcLbu6hKMFmivjXPOuN5yRz6OsbE5yFMG2wO5LebLGd/g5QeiR
sJ9AZ8OeKj0+F+KrAaZaqdcQgQLpfwrk72uBnA5tgUaxbK1yZhwifc9zP+rOQVebyUvYMrf7BmQ3
NGG4XHK/gNEgA9gXlhKmEM7O4kwtvnMtPNOSvRiO/9ekIGCcdjvWyn/qXbE7xbFckg67sJho48vW
t6hI1C1E9QQuxn7dJzd0qoaweuvvZw7ydgrDZz0wBKRppYMg89JPCEwPJuoZl8xAZeKgsuQJVagS
HAL6ifeUQ5kirTJEZa3bxq6Xen09rPZRgMRQMTVFahpiWiBCKFjLsBUFu+V09H+biHrM9hZy5bE5
QrEIvTwu/+7eWj3/yW6z+LfQ1ZNghitvFICpRs/u1iglVyF9neZGz63yTdCLBnVgKiQ72GRCEi45
2GcF1sAB9ipzGsoEb4u89lSjrm9p5AePmWolXYLnzVItUPKqoib1mo66vwPCwtfUnK+m8aGCDehg
iqGMk15XLrRrTjoh0vHVfyQMVv5We33MpGjBPB8TxVkG4znbUg6QtSRyJR/1DfC65KW6yVRlvA0/
UATtbVwAGMeQU8YzHSP86hcU2j63f5JLDJ4IGwOfw1jWSqHVGPqnviPS1ulxt6OiTio7LWGvIa/K
NC1g2PiaB0KzshWMLD5n3GIR6QPKD6h9Jrz282PVBQTzZUjXWOmcm6UxccWytWai2zDqGS4UQ5bk
8+uc5ZLGLTG6dTsnAHRXfbE/kk5bCy81cc4bn+Yx8oMJKK19TaIl7ozX+BZ73z9jME+iZOYhK7yz
qMCgRdAWx653BQEtNR5H/3WwmDJYi2paVIcv6+gHB0ByJYD+iW3va2XaJbs3AOBWfq5BchXbFaaw
ItjmCNIPuHZC/taOtLUS0/VNdEOV0gtPBW2LgCZZ98a17rTv9htNVZM0rK7VJQgn9DsxDrgSJ8pJ
kA4porxKz6izfxRaMDEGArM57daLu2pm45Xe3tSER3PIaFruVsn8sQTLY2cYa2iezS9J5md3ReE3
1b9FcaPZm6+pV7ux8lKirIE7GzD7C8L89z94a7Ar86p9AxyJ0wG15qCwj+w0UQ9R+jlbKPYd995V
RqkD7VyXnFmftxt1QEVX4U6uT4V7WHq33hgAn7OHeOMsxregQ6yb/Cmpi3BFtLxM7iZLhGfFfPUp
px9DZx3rWdkGhyw6QWpcN/xt/8KQ5RtABjOnuNmS0uw+16vcFNEkQeA3wlUXLFdm78E9nRghzwcR
xW/ScIEfBJdW0fywT5Ltx/wJbwLevpe0PsL3oyyHeInKYkyC2j+XnYkEQ5CAQwOycD49N5LTJAM1
Zqhu82pux1KuxGo3ovKFl+4qRHfshJ609zmCMARA6+YWD4EZxew20o9w3jpC+OghfzWGulhZGZ3c
0Bj+tBFxmH/eq2MK7E2Zr3mP8tX4Afny3Lq/SpzQ/cHsV3vKNHiEOFqhLGuG6M8KJ/1hkT++PLI5
YsqQAGRlDRmm9T9XhOuJmUIuM13dk8TtLTVUGi11orH3lfYaONXn2Q8YpsiMGkWq3YDaSrtlLwY2
zSZcYUVYxCwlOie6O0eOSlsR9gpybUv/SXGjBdULCbhLO8xBwqu9DUbnKIQJkZ1vAShasrFi7jbJ
hZnKGuA0PLORnmO9gtHsTkJ7xoeHiTGHr1X18tiDtu1KMbrgqZkXcPUeg95h0Ww5SDhJLpUq+PQn
tEOMn1aaGsLzeN/fKwCQkbHMDJNdZ1REdFmdpUIesZNdPcNVLNx2h8iGRA5QuS048WjX4yktNisp
lPNd3Y+/hDKJwIv8GG81+1wEOLQyqBsAAGeim/3Ax9GYbgkQNLczaeQnQeMPwWSbut2HreYwxSL3
qWRyzj3mOtaoiDjLNvQ72KL/EBgHhRrOk0UUJd0Xe2bM9C5/7u+82LhScj5zL3mD3R2XQdCN6Uf9
EtMhwXBrj6ZvABiHKqwUj5z0nShuKATULJ7Y9Z2Q3IL6MqFZQv7W5mi+fyYuwJs17/zKJkBguRdX
8MBjTr/5n509vq0wHyR5vheYtikIk+yn+EhFy+YZHM/XtqM6jGcMmid35fxitRKk7ahJ7LrdVgEC
dFLxIDq3WW+ewwNHxe9iULA4ZAY6s76JUvsMfiCWK9x+czrZC3/KAFD5KQT9geooLPJJixmc7359
wsK0dgmvQLGB3lBbmUR/t0sSZC1rw5wtak49jJP7BqhJLlQU5Yj1ZANBWc5k3nu9BFHpr3OiyLyT
G2U0yo2+3z7mmgPpU5UeoFRAJTXg/vzrvUhiPEyYxS6xhSxCfyVSE36N+7Vb4gyfkwpZzkME+M1r
4RFXz//KH5S3iwt+Ip4dIlAZxm+piWIIcU3c0xwr0Pu6Jgat4s2Kh4ROOPV2SsVLr7Fo91Cs3jr2
0uSqne0NYPKvQY/UWZwB84T8IRLWnIhxIDAInpMrrcFKuQ62SDPWh93eFvmj+rKYQ25+Sfck0zig
OAm697BeeBuKHlwUY0CZ31GEtLXw8zjtwuIKR+B3gc1SSfZMLDpF1l8bmMty5G9kphfbZBNAyksy
GSlchof7x/DREPuj636jubZv3KT8toSoJtFFMEeBOylCiQzH5OTZDjmGAuSv+EaOO2R8+ivHcxMf
HkMiNthmcmIugQPQqFNzocfF1asf17zS5OSyNPAYWh4fvyDAwTk58cLo5SPaQbfGXAAAlebc2z9e
ZwgwJ7rh2asMbNgFA+4BxsSiLW2x1jR0rYRKHfV0v9rHizb3wq7I/BFzDwOyeKr1resUDZN55a0E
intjp1a4RLyCXeXwKCFUjfONyrwrZgNkWgWnxpiNsHAnG4gEYS2If2q7NqB2bS7sSgLeW3q0eu2V
hK6m7CbRY6/F0CdfWU2x2kfye1bTH6f1cU5HUuB+MczoJb4yVNLRTt6ot8JAwy3XsrVjWWbHuj9b
17d078RPk13y1XG0yGMsHpzXyicviYdzc+WWWslqOWjPah8JkQZ+qP+d8pGU2E86P2rwr/WNbRbV
6pj6auwSLoJr+UqhtpgbY4KzeMaXcF2JzbGBYwvwXCDvbvlQyXpdAqhF8Yjg0UZpnKdl4i+3SUYx
VzKZaqGTi+fcfYO9xTcDsTQfmcUWGg2me+voYwcBIqFeTl74qJYqDkdIt+ZbzfzAiLlEc5phg0IT
H2Noa9LW8AGBno0+0KIPakCj18Ki1nbV00B0pcQiQRg2hZMEer0pjjFFD0RJvGfqZ1u35h30oO4Q
ePue8xwRs03rul/TO02FiYvgjCjJR90swENGLkVE7YSS2eCLNYK9Qf8p18GTSceScdjOLAGRVvmV
YuEBJ17ImObPhL2FjJCsbq/l2u6ksh+oDwoFxnKd5ekldD8saw/MA7rII2gOHR3JtNWg0j1rcCV4
+z1nP1CmnzGd0odihV0ldr9xJS8d3OM62FBz0V6USExUmft8HdhJ7ky4EQx/eToSuL2M1Y67XSlx
bVju0U/WxQlpxH3qPZcgddlf3p+xtq5JhiEzjSGhdrnWV5unIfhpQENWIRz1hmzBNPHnbkV8qnzj
+qH2C/X3wjigRCb75J/S9pVGPlfc+fddQHFVDcjrndHOkyO/OZ5K74GeVLrWlW2HCKyW3vEL25HJ
8HgaTrzuruqnSRm75M+YpwW2nNICR+RSgAxooBnfYPz3htoxAkNswx/7+aU8iJGAXv1Zp1er0FJB
CCt7FaHCzu3QuyCBX42Mk18DJrdRGUZ/AJlqlfsKaY7NSBWFZzNpWXJOO43fPZ/j8QjBOpeD+wUU
nE+ivYxf7ytREj1NBEMGSZjXW1S/A6/NhivHIWSxWXZh6G9kr8rwTLjQ8koTKW8ctI2NuIPhlW1O
zT63oRu5sCU+0Q8HtiE8YNUgYRgHtDTJLzPWpZC/SZNmXKqiAoVnBMhxJSD/DZ2n3SWbdBnIyAVk
GfOKMFsZr4kUIgzjdoWCPH08hMXDMwnVs/SctYfvOJBcgs0qzbyxXAYs6u3M49nVzUIbQKf90diE
/rT4wco97/r2lA7YBM6RsAxoy2pzHZJKqhhLr2ufZV/2eAJrWIMhmyY3KG87ZPVJtB5lA0IAvZap
T00PtdQkjQFKZY2RYiaYE9mqWt1LT3tENnarRqrqbL+LYenxqGEglhpGQlKb6WLvbt5PAvYHr6AX
4HhyuHuGqJ8PIKM9lV+mgd1vpwXC1UkHM88V//lF0sgqsFjf6Fi5KgwY+g6/N87Bwpwo/g/1hVjk
N+1g4U8IgZjtuuoWEUb0o7yJLYzYMsWvfl2hK+wdhoGEUfqruNBWrXO0F7kZJwbyC14hLXDJZENg
6nVaH7tOw5Fd7tG8/s9KOg8fdTE8YXxAQZXNY71UahZU4jp+NCaHjCgEvqYp4+XSYeLyyY9b+Jzv
/inLdFD8U3ES4Eaf96WiEKOxRF52tvfxTm1GDmX8xHSgH3Omu7sNlYry6xt7g26/UwpFEpx14DAo
OK88N2wpftnjpOEtnH8lIUaoiP4N1tYyhVeudpffHavs1wo0R8+cs+gyt+zvjFOeYACnLastSgeQ
nt/ZqndX7n/miKn76g4X/k8Z9BOFXsPIQEO2SGmwKqiXqdulqjI6nw5Ne52Pwyj3wkmIX7bS36Bq
c2AjLD8KHbpGaqj12u6bvTVAPQJafn8gEaOD8KfE3sGwz4o8xtyFWqIAKpfp/oUVuktyTzAPKQHX
XNu+ZZm2FCy0mce7Ts2/WvENHKjEFCQ0V41pMGqYYDLFptoF9XjEnPnZnSCHBFpZFGiE6FU3sK0J
m7OrDZp8nHCLH3C1YkkIhU3wU9/9E01CWZPynsfty93O23HnMM3sKU60+0MX15t5dqopY6e5q9t5
T+gyMaN6JG13RquWI4KDv8ZA31Odcc+ONXE81vy/GJ1tk5EkEeWJi8IEYGx6Ss7x9qErS880hv09
U0LvSNcol1Go2GTXA1PAfdKqXR+Zm4w7KF7nbpK9BtoFUhZh7Ihv3LgZa1LJgnFpgfgww8AbC7A3
1YEvVg3dAKv1YWLC7ghS+krDnlI0cLjNHXfrYvcElXG1k7JZmPZadcUIqHn1/e7u4HnPY2kAWojH
i2rut5QgK7WXqcq0/ev3FQ6HCZo4goiAYIX/UUOpRdnDUKUyusNOYIoWG8aMu/C3mfCLzuna5JBd
jHglZMUZg8pHTbhI34m9n4BiuMryVVHn/02bk73zW8g+svG9ifuqH/44P5giD/tkSAab3zUDjyuC
cXAjsdbhqgukS8ReVlhzYKDHrPo6EKnbZYf0f/5H3roT57pzEs9eulnTKd+ajmiAEfJU+1s2V2v1
+ViFspy91WLrASkPLciqf8fQhrWHs7VjhKqaIAKvFaCiHCwGYXUXUORUjZp7tRechNT8mdxt56vs
cHpY9ULyjmI7bpuwfaTjBEmG0WDFfImSV01hL9Rdf09VyTBiPbYu+JMVhQ7K0y3U9Uwh+zXyEM7U
XbIWbw1q2Gvx3wdBt674W4crunWqNsnd2YwHL95sya094ckaA8auDi0XYjvBcbfWdEVfEzKfuSqM
N+6+S5T/TbCmlwkp6s6ir/vcQSz4sEGkwXAPDDUHwRjQZ+sbRX0ltqpMDAGPLTwKMF5oQ5eH+TpZ
0RPkHkSuAhEW13gIOmS0HEGDp2ACSEXpPU4YyIErsqoUhZnfIDAszFyGIwVaGTSe2pZYVHVvIJwL
ZEHjsbH60/b0CjHG+wavaEoPc3ggJNJpLViZQlcYYzRcgc3qHr8TlUiO4PsFBUt2wySBxs0pCiSa
s/jEIIrYcXK0I6zXrU6ZEZzlZjpI02AFSeHxNbYIU+Bpf6B9rEILMsJCTQR5YIajnuP0qs1v8r1t
IkxnKVBjyMN5s5d6hzHERBtBQ/ZPhFqUTBEdy/zlz9oTXdWcbsnyu4/0XCRQRc9mcxnLrOdGO4NE
WEOe0IKjIdUujmD4HZjFtqV+5CL067Mp8MEHDA3NYRGE5Y8g/FuzjF0MgwtS5DJPkjHXQpxpNvAo
58is4q6lNFYt4SNOKio+p/l4CqWFE/foLKqLRVhsJsBf3cyIz6um4PhhdGhT+hWENiIViChsPdKM
uZK2ZE1WfMEryzX5T4CMbpmG6AMeLYWPaVdK/vMqpQK5xXXqO+VtiDI47l8Y+GGiQ9/0OKvfq+yC
G0vNq8WwpGgvPSMEdRGcxE0nsr5w6FPBr7wDBaLwi8jdOF45kZYfSk1KJ4TUnN9lAWLru0WaWMgr
v1/xeWj+e8JgyRkbBnW6se32UdRrrUOoGj4SO8Zx2JDJaSm5g78pBzndqOdywDEHLH3BJ5w+V5b8
QkSVN9yNvdod594lHVceNMjcMUMXYid64DvhtLoqUfEosd3OnrIjynLMFqC2L1ANKAjzwG2+8d5g
SQvS5ZKlxtF6IOghjdeWdebZsxciaeKq/2DyOBDZA01VijULO+GhhWsokfgYlmzJcaPujwrldfKJ
Ki7ASI1PatokoDqPBvgVWLvSZZArl+crAkkUf5cQP2W5pjHZE0QX4LcTFK5ftcymx/ZeKK7azh+/
4vMFVseXzg1miz64nOLqwTi5H1sGNASjlLgQS9yvIBAEEhvi3wdt9lISBQMuje6u4igDtUDQ+JTs
gCgbGQV0pmMA9xVqKnHQ2aU4M8mtkHs+c5rqPPYecFJla3ivmx0tAtDa0wQ4sfz0XbTKbhgqr5Ks
4y36IBBmeNMwCqeMjl7fBUGU11K9TiWZ7I3yTM6bZK8944n1iC54QbARjm+s74/B61oOiD9AJDZW
v9Imd/d2gfVxs9vabD2B76fQjcPQ/1Mt6baip92Qlk8BjX1vroytTRuUGU4f4nH2FbveBtgw2MuE
npdC416QZq0pjDO3nIyRXOzXOQ1dNruH7OMMGbcv44TVYjVtIFwcDkOhzY10+ghbIXBUism5QI0u
fseySz3ZQdxaEWNKJ+AKatg+aanSgeaf74zDjXRrLNo0HwxVGr74L5yHh7FWi7XmyrRIWW9g1fVb
72gQ8yOb9TuiXuXK96gLNbX9vC4fuNAlbbT+aFrz5iZEWPcvIULUir0V7YxKO0ydrAMlA9pS9xwJ
0fpxbyDVwnXiWjTRuTegpNl+RLFIGKvFSMLD5uCpP3jk4+fI868VNGG0Q6ls+EZKT+rWoxv5bgVm
HqZEhysCe9H/j6fcSFJHNuLNSpXvyLFZyk17swKnzZD5oaRzd+POAAKKGggEzSrg6szVNSE2MPZD
luk8xlc4PKOlqkqnxOZg6vys/NXIvoiEzXZdI3fpzG4v5YbNMaiMedD9/K6VYuQ+wVpVwVwC+HR5
uVahyVnBeyWsWbNdsBbrjpbdjsCR62u3bvriagM4ZUXlSDFoT+Mqikv4lkbhVHX5uRqwLlLmbhSB
T/EztD2qf975BaJ9xOcBnpJVvx/gFVJSThRIcewW+6rlMgf3MLWD9Uy+XdMKrW0ev1e3pBnSDk+W
xo32wC3V4S5ksr8DsA7ievn7d07U+cJAnnru6/OF7HA/xTmFNrRlr3NeR44RZ+G9YmNJJ7/DH8uU
vXs5triFW/J723eh5n2ZshFau7C4BR8nHzI8va/2XH353DgXO0FyY99WevALHBRn+wZS3cuCbAXd
3k27B5wBI/BwEQm5YY2Tod3Yr/Of6jntETJjDkF/AK2yJh626ZommT4CmxZCyEKVYn6zvNHU7YEg
LPrNpu1xERfXxxxR9ZnaXb6Q/TqAE62f+O1iGENSJJZfrBq8zrJsFxQq9TIWai1sOhWe6DbYDtp/
yTozsec1jV2x3CjL2ioouSBuQJB/J/R3TKcG8fivqDjPj2uv11yfdpwtSBgREpgWWWtBHdi7CwUP
JLlgp/YCwCyH+75V6VPC6y+c1cWM1osf7H3qYOEl7rJVVP5DcOyIXFFI25ieyXEx3z7Zi3nezflX
FxD+IU74n7vtciz1HPacJCCLTZ7kHyKJB7lZKJyJLRSIEM4rjhbpaBYF1jnsd+bpYBb9nyczrSJX
tlY/pLXgYd+AkOo3tPhy8tO37cLfJr6hkPDXHlPNZesX500nrxQy+CmXDonHpGYHNqrytBgIrHCO
aE1KKJXe0sYs/pCLJs324MKiQor+7n+UAIiEKNkk5Bb3dnqnm/NlSXEh1rcHm3me3FVSRYLbKcH4
Ks4DEhVRXaBRKeE5jgKSJBLtBSmDVkEcoMCJ8cGyGmTyG22RaxdT8oUG2GFGiHLNAc73rhLOhqKw
G3Lc6mw6aICwclDO7E7Ome2gLnOCwxAFgQdstyBRyyss2ulwtioeHpXeX0yrf8SsWJ9O9XtM2T1t
EW5l5uWeFs5TLd1VBiJNKcNJLD0iV8tHWBrwC9IcJqiGgP/NFlmzEjZmNSdGEXntxHwsukPl8d7U
o4oTiohJrFdU21CW+hZZiCZR7fYrCrl57firu+yf7964I27LAunL+lkugojv+0N0hrNdlIjjLhO7
Ue6dAMbG8i3C3RbaNeCyb1yK15ec9FDAs45Xt5uYdCiWMflPiaOoLlBxRpkbJV3IqB3ojUVOM3dc
Yl6v1e9Z6UpTDV+VhvkpJPBgEiJYGbk14LXR2gYAtP7LzjcGK5A82cknxJaHjlWYZBc2L47WJQuC
2golVikTNneil8E/LqanadIEeMMsW+rwJcaL0f/3u2k9FHl1A+6ijO6Ng/S32+Z+rzbIJxyMSTsF
WYYu+nAEtvbVGmw4IkRONL1C6N58KGslWMgWBL1fxl5hAhlthoIwZ29jkjcUAiw+ysdEcvpvf68X
tJUHnwNUm+RmR4P3Ahtn7Oqb5RWaZ6fMB27PUHOLH+q0p1TpGueFH5pktbJ67vwm7sWZXJ167XIq
/t53G8sSDPGQWNiMYfOEm5ACxvGBw0OXzu1x0TOCfYC9DvInWa+Zf0caaryobvA5JIKF9kcBEFzj
Bxq3NpMMq9ucUvDfDo/wkFSVoOB87ZBJwZ9kIG7hSBJYMIAtUR6uYIXeJJR4ilgB70WKKllGlQhc
0o8xGy5Pj2c/mYecUQ9Ja5PsSuIKtfvL91u7Bnk5LnxETXYFSwmLYE8eIZT4ktIZpUsWsWvBK22D
Bt0dBbanLNbavoAjGAVsutLUrsjyxULfECoXcn3r4+bcoLQNZp4ARiOR5TDeBrsy+RYc14Zjle1U
S1TMJxwyQPgBo3wYvfYy5/VgmYWyjVtqARSJv7FE1A3VzRBav95k76nFEcuFDp7fwCM3lDPnrk76
72+A6zpxlNmthRRqqo/osSmPbgl7YAdJzA+4okhK+se7Z+5RsamIXRlxSVWjM16mQUYWPCPhl3VX
En1BD3mq9Fa3CsKgI+WgBERymC68Q3h3MDdvjl8OTX5f8ygi8MCakAhlf38vYj78at0UYFKfMlfm
7qbcjLo7yH8MSRN6uLCslCdhJjL5/9oeVFkosnXRh5cJKPP8R59/ZwZozkb4/VmbhDNEXtwC7Fvp
R+8nnz4WTb4SraIWg5J2Hai71MGNRfsnL8fdpGT94ftkASnssdRPSsoJkTrKw6xFDgGr8XeRftt6
+e/R38nKzJRZOH+sRftQ6HxqOWyHL4UjZYXWWsJYLgacJ54GMRmUrn8kfR89QkXhYOvhxOLJ4+QL
oeljlCtD77J560GRTnSzVWygtqBQu6znZSHmBVzAo7lrIYSxTQ/ldPKzu8E+c9QTdmY66GwuD1IC
xDRh42wYJ4UHa4TvBGwLOh1sPLO2QZTATYU/g7HyWRkiX87aL2OInQg73Bgs9++zNnhDO3DknGth
PSiERjlyqAClwWp897yYtx3wZZgsyAOHLlX78blHdPzOAz/uSVk28JzN74+F553WlBwDnNKAkrot
z2DBtb3jjRsgC6li4KJ51+HoF/6t9lDqATYS/vfbpgiU080SSSy8bCXKU97hdPA1MTSzBIpfI3+8
vhcY1ye7B6+4Ubka3Gz47M/qbXLa/nm+PJ6TokFWV6hU+4Ul4TkcUgfvJ1+xStJiAk4q5ycxdKNL
vPJPqP2cdgGeN6BhXtEu5i1hWlY0UWcF6z64l7ZKzPp+fctxtT2HvPcGkYxO9gBdoL9fmr0SYyhd
olVKuxUDkwRjXODYBYqu+P1QFNB4cJxF/pV9s4I28PwX7kxAu7lK9e8D9rnlsxmu0bp7GPTDS8or
Nwih7qyo8B3jKNmDj+sqcjX9MAa6uIYcOUMzxDPRbEAwswk2VNeE/qG+1XjN63maGw6cMwSiFkl/
PniWOi+GcJsKj3jq2Q4m3jWSX0ilcXvAcvkCdYDIFqOXsvW6HPh/dcK0xbKyxS67HqdjOaV3BOU6
l4dqT9lQYjHFMRPWOdCa4yTqeapSEBv2HGbY9Aa27nkW5d0/Z5peGOi2fQ5d8gUmsM3pG4qnjGXH
RMkMZlJ4iMlHBkYZhVSjqUtmPw8S4bqSCeN95b/5IETd51Gk+PXx3n5ENGRbKSJnw0rtAYvl1EDn
3riQn3MAQlaSV7N8cy0k/rax4ALyuNrm/dIDB6yRGzRO2Qmeht8aF2LFiLx0ApBIaTTpcwB9mF4C
dKPVtcokkZIIcpqRZtJZ+LKHmHtNEETlaXItbOUpLBMCJb6+oo4u+mW/u0KSZx9hRfccFvwWScEp
i0qa3Ce2tZW6yRqdsTgeGfU/9CZu3ZB9mdIN9so2QtwIxJT8VV0aDuQ4CDAY1wWzIBv/YTD6Bx0s
hBEoR5auwNhkbBrz//crzRlV+k3hWx2JA2R8mkGmQNgsy+BrYOKQlwidRCGxPHjBDmUj0+gbyItF
57nM+1SeG7oDSW9/PBgfdchu6J38mnEJUKUU3Tfu05JlbmAGaFSY1TTdn8jd01ddRufXIUdpNAIV
xfC96P1MLzq+skxSt1rKvFr9+L6UuowhuRO0q23Ie863lMzZzqv9eZxVtDXGnRYEftEmZsKNnL3P
L2b90NtsSuNDPp0QP6el1Rp6CXz3WZel0fpCWTkomr9B0qsQ0IuAaNl62+0JOFuiXK6tIgMMsAgy
iiNHRY2PykA9QoJnycTbmY5F5hF4o1AuabptMAP8kjDas0sK3Ir92o2NW2D/+gvsI56iiP69mPN9
iIJh5P9le0k5JGPEATpzXf2YdD2M9hTjWw7e3eCT24TF0Y/zmjovdI//Qt/Rzr9Pp2dXZjzX8zyX
mcWgwHx6XA+honyBoiUBUP+PlRXEyrvjsNerCv76sGj3gJMl6ZLudlCQ6aiwhcZjw6APlWVZFuTS
zNm3Y4tBB7nbZiSIYx653ax7sU3p1bxsoxDu7WRTvgOrDiefj9s2VajKiWLFV9ntQxxc1rU4ZwEz
xgtl6lqrbpA8YQPlTrjvrDwrLfAfnJnbGMpi8/RYTb/ni/LqhkSpjFnU6BHhhwqDnWP9T6r3BnCz
7VZ45P79ullO6zEcKCa6Yt0noi44Z6gGhHUKu7fwtm0Pk1MakCrgk1zDFLHTvta63f0GaKMDEOAh
BycrV/7KSpv9wgrMTDv0V3bde3JrxPMyoY2jB8PozDoISYt6XPyW8Pcb3WqV7Vld9zqMyM3LJDGs
lCIn5KnPvEvAoWsXo1Uw/JZI6MizRRi3TIrXU8N/WsXpEJ3tN8FgfWig4XF4eF+Uu90GSuHkwElM
w2oCbpwVE+reWYjxSL0mnAn64L0juSfVRRBeOJHNPual5wk+YIihvdv4365xkUtfHOo+lj1lOm1D
sXMt7tXq5HbtsMfwjQvvleMflAYvJ2zNTQQkei/+DrM/n5p39+GWzv+sokyJEm0dGZ/tN7G2RhRH
sefhbbqwwFrKyTI+WwQ2BeoMNz8LhVecP1nJeap1aPgmehC5MO2mEecMwWejo20vHK2lSxmz7RZF
8nuNL5EkeXL6/TDZf689lpzwCE2PfM+MtqegfI7u4GAXSZJ0M1dZCccaSLR7SI67DTLd2nnR1dNE
+J9vUV5mFF8Nm/GYHvZPZ2t/m52UH3cG2qovpEECKL0lv9nZK/UsyuvjeiHdDSMJE7Bb0LLUer8u
N3t7wd0sWE1/b+vYFDHmQFwL8ayb3XOH7z/9+rOe2orlPbjsDItcj2OVP3KlHdVvtKhOrNOiLvJB
JEuHUG0vj/M0nKEV/om6t4TD5F2W9sd1caf9wnmkgB0w/oBi05w+CAJJOeDh4Px+3YUCMWBDhxzw
T4RB9CMadID8FcW2/TIQEZkRUrS1pQIrefHuT5t5UTIj+68xo70t3pEHydotgPGjeiUT8vk56bE4
c2BgrtKtUyOBx4V2mPMSgnRISys7mhIo75SJgU/Ioh+rMjVnKHHd9BhMEZkQ7K5Hh3Xrr3vlxc09
IOdqTpeF7soyVnHTHlmExRVG15rySlQ/Oye6ulO1dlq5x51VliridCrzYumY1WDVmGl2dUCxs1LK
M12eqTQ1BlAibjRlLrYCTqh7cEplfhK0x/D3ItpQ7z2rYM6NpZ2Da9QPdbj75ScURV/ZbT01Z+bw
xO8+Vt9AGKNbcN69JwJqJ9UUREHzHJyEU32+M5FClOCordqCrKKwYjGZGUWHgW07vnWycxcebYLv
VzSHD98CEVSnuGngN48DqmQOWN7PJKa7NfmXYGErLc8euVuFEIX7fS5gFxMxnWriHBp77Q6mu1SA
gdc7AN5SAoHbuDE+K/e4AxFPsFL9Mpw6bIGjRCStkoXgYABNksJi46nRtXVGOGQmMgGBCkGmUC5H
tX2OZpwyqiJYfbquUSoObArUNg9UOFvByGp3VeDNf3wynjeX88aih2o6IqCvTpkT3iqplLEKpwvG
2/cYnObQ6dxtCJ7QEAhQBIjOLPQtKiTwjspqi76aGk5i/N+523zLEvnuYT/GhymwHC3Uszq56bZc
WYZapPft6HM2n0LlhmejPFNkVnUFFd2VwvjWFDAy1O1T7mI2FlTd5GAX9Xc1cN2L+tKggdEoaESt
Mn/OiHrjHk9O8FauCs31+Vzi6wbTKKx0/EOHk0niCpo3xKZr5i3uV5TR65M/6soIC5ODdGnH6hPA
YYczXBxGby7OscqCVoSZarLW0yYKZh4rcVhNK2vnxxI8kwPVWszQfKyvcBmeDFOcAQUvHazMoHBx
HcUgbxkqSVNzAFPRzxaU1zVkKtsSrk59Ts6TU2v3hsw25DSz5ttAVJMjZ/617Z9j+y3+BgWzQ4G4
DVgi5+fA/iMWCjfC7x3DoCIcMBe4PHLrfx6AY+6/8ztJU99ORO3Wggr1OK6c1ci2vjQju6qiea5+
oVVKZFXVBTUnuxUOd5EPvMkOLP3uIvEUlf/5HW/QGjapUJCkwREpH8DKeVccxC0OliKjB0jhehxQ
AVMxkjWxPrW5V7XCVjXh3nJg79cVgfQiMG73xQDLRzjycJ1Ux3n1TuBCiWoK0O247cfOVzb4j1fQ
m1MBN+lpjpNPNbZOciueEXWmIHnCiParZvmgCmFD5il8plcBPxsF/FXzOOR+6zd48tv+TXyH5KeF
hg7jTMMMCGEOKL0EVwKA6kl+W2s/700p1PpFVfpAuRtrzTRUPseXVIrOE3anv5qkCZbhEjLMc20V
5pblOq6kNS9ib7lGntGkG47UCL+1xMurj7GcIjjU0siumGMYZFbJHXZcwCsoSW70sKmKHQVL92Q6
eem0QYv05U03r2jUBERCowxmnTLgcyk4f3G1Rj8+f2cJRJqEByULiU1spVOnWobfN9ijzLy2B4t+
IZbm9TAWMJFTSe8xMGw7oIcTTZp/SaLI4h/4I8MQ7SH3ogGzq4ly60NdgHA2YD8A1FpjMdAL3P2z
Mct0o862RW16XV4QNXcSqShzertNDWOmO+2WqiuSDWsCj1VE/NR9rd04im6CNN8AD6RiwExMxUir
wBobmz4VNg1cUa2fOjgQJlIi+fCtszRvKkjHENAtqWvXtFP5M9dL3xpY1LdptO4DILTlMav+mfO0
OtQNMos8PKwlu89N1bea6Dn3LnBEi3OxVBxaX11MJzwdwG4tDfCrAG6CSPBujo9JbxMDAfIvdXWw
lL8Sh3qsT069YYySnfPHiDB61TJSYzMAROukB6N4fqzhRcNVs27eXOHsoR+ZpEguXrF21CDfnQl4
7rMneLPWEsUbRGX4/unFqMabhhy65CjMUEystZxij95fVltq8unr3Jsylqap9auZJpvXI0GyZArX
oCiUJ7Sq2b9Zf7WWkg1E1pL4QJyvLg21RO8irMrAYOo38J/ycTuayHbfLKjopRX/IKiXR2Zwi8lb
2mL3yq9TeKzU7MfAyO3SRkgMSEm+Tan5m+4Z2K4khQpADJLL9p3FEcwIhYxNsaDGuLOoNEZ6aDTF
mqt1JNqFX9pR3sykqxu2TtUdOFgMcNuyq7Ild9SPXOFu7I4AOQKMF8SU1Xet0FqyD+lJTLU1GFOc
b5pYTPQcS9KgNBuqQTHq/5v0tNIEAfW+ufDGHY9PZ9gPdtt5Mrnyde6808G9NCMnZD53cFOCcLSn
obnvl8eYRm/VNYeDq5+8EAgPaqRwagbvnp2LVFr9CNt4vkwhFiv25tEDz1aXbIB4k8Wtqu/UaaQW
CNWxbARdPhU9SUcKpAsEX8cb1H2GXeAMGu9+AEkUz9NCYNTsPozpFcf+vGh4Aq/s76EHa2iob49a
J+IqxmDx3AUIlhDhCKQtbQjraP4O4N8KofVbXNB51+CCehigwS6IwbRa/TYuUsnnR9XTguWQ1NQ2
G7JRq6phAn2w323aPUfxybmZd3buVKYbts7sux5FudmjjuT6gshVMmGlMJ3tBgoA8dOlgCqgCzT+
oAcu1FFF3tAIOvoGSTbtFdWPjIIbQLOTN+NCxWMqLgtsTCLPsJxaZrlEcb5RLnpC7IFLHrPMUxNn
PJawgXdEsUOEBQuOFe8kHz0oUMWByZF6xE2On7sBMsdp3bZltHb7m3Y+pipd+hjTOqwpOW8BwcYi
PP/TnwR6rnCsLfxFBtbx5M6eMNK7ACNjn/ST78tUyWo+Jrf+QN6H/QNSgPpCScYdKubAABAJAA2l
erTX5j/Bb1jTuakDlFJkMKEiWsdJd4Xh026eRiPC3REluDhHvxl7i7rRXK0Mn7Ha75dh6WUNgIAc
aV4Z9inxMqKbsWaX5nr1P2+aWGeEYRMpPyChgA4Ypfjfjq086P9rW8ej0Y3BUDC1zv1xLSmPTy+V
Z8MDKH1Kwb+81LpnZ3WuMwxU8H80yqsK7WkV13But1+H8BcZDovcrHFTEt/HL5acrEpK1tymAILO
EIC0dwHWjxdoPJtKA6/m7MAXXNKAayBDiGqfoljknHtm5a/MRuS5sbErbpi6F1OewRkP2oqjARhk
bXqQIEr85zD3Dc96LTUheJk6Q2nTx9nKoJxHWzGlcjiChmcKCPioIfq2MV93aWFKyV3eng3c7G/W
N4aDeOyqd0X6iwH8wZ11b5b4z6AmAZHY+i3XGcm65MrlKiKvBf8mWQId6LNWtgXkoxpjXyGxcI5z
JUpcyNaT/H3T/+igWQ+VVETQkq6ZLO/5Ci7JF3U9Ts4j1mAWjmehLH/Nn3UCKXmYJIDxogSPuW02
SE8GzD/3BzUSf6rq1CUpzr31tV1v4xpz7gv521AnKWzVFRzOb31QK9ZRVTvCd3/qMO9zxbCSJT3M
vPUMIZoLxeBSGHVesu3rrvBcGvLO/fOl0T1z7r1FHGruYomJg+OEBP8CK4OWPN8qCBzshtapW/Ce
zXWWEB83ZmSjpcquIGlFTUnfDDd1NFyOR6hhY206PwCAEWLP9XGdJmTBMfm+onkp8DxGus6pRKVj
4m/aWK6tYxCr6g0GCa1/ph5q62zMKYbrc3Fj0VfvDdbV5n/yihU6t+TIkpIBw13VhJ1bqd2jUzdk
mTVuZVTLjfOZo1M00FLbLIfBQYw9YUOeTcbKPwDfCE8LNpPNILsrtNrPL4n1rFcyNVP0b9Yar9EY
oMBKH3Z39qqnd6MVFBHf/m3Dnfa6NWYWy/AwspSMKYAbp/TGydlx1Srtzeemew9rtoAvRK61vnFl
l0BJNjcfC9WwG+SjCe+rRti6YpkKJx+WGi2MaPeKf15/yxEm5Pxoyz4R3nBLnidFB+Yh6erBXXH1
RzLh+Se0O5EqBNmR6Y4IEjOOVBrm5qr2fEoxyR+eq3kwS7wVKZ4C7VUTH/X6XGB+mKyZBXhg9Yf/
UXM1CW/+Iy+Y7r7IGhxSIg4v1e/Rpupvk9pqOQFg1YRjPaulz6y47m4BpyatoIjlrxVB1kkbryNE
6JhgvDqZujvMc3bDUlUiWPuaix6fSIf5lzSfuA7DUo0hJdACx4Sk4K5MlnJwQphhd0JcEiFWe9t9
PHkdM6Am62AFGk9LXxqLBIMAuVRWQ5Gkv0cTX12OhH6Zf9Qthsf4T/dxfJrkQvNRit+oSI1+YOTJ
v8Yvtnuj+cLqEhDNowg1ZtceABtJeJlXTM0VVT0qMj2zkkhf60+0PHLZKCMUUwQoRMAsW+yvSh6y
7DuovMX+JglpwFsb74qG1iBjC6o6355vC2np0JrmednVplTr48l+Xo4BJLo0ZidABKNIeHozXHYV
Ne/8u/hShhdB1gjkzQjKNiDJyLJYi0ABS+6c1HU/pg9Q8eo4d+eY1Iu+jzanQ6+qY9iTgQiOzIPx
iMEd6zPgmn4+DKn3EZXly5uElRetPRfzwpLmCKuy4HrqhZsBi0bEpUy7YmoLI4cn6/UQbLtSNRrh
nb73Hlyw/RStN/GYA09bvFvPNATWvWslwmD4TDAMIMk2CfU4xqpHNxDmWOAv15F91I+iMHWA89hK
QzRKiZNNUDCl2bZPLcv7KhafLXqI5E16OK5oqDocL/w+GQ919NtFeDgPTQpVwwfoBkP7VUjPIiuD
K6JA4AmOeFy0uT1TYfx/wbD5xmAUU9LeZTGXnbczymBHx6ApkCemJ2YQTROynAVaKLFUxFDdXG1a
drcLRTMppqhW4EoV0oc//4D+hLIwXFrYQXD0Wb2ydvwa6HnXRLwiQ/JJIsfscm5AycLTJvvWNIYC
Jw2wsIJQUPihMBoklUcuhpGJAZx627BslQlQNzpAunXjcxxM5L3ovpIFmpSP9O9RRTLFzAbDANRy
Li/PwLNAsOCJmeLmDeVNZq/8JH0O2CheEjeVUBLEyE2d9K9BSKEL4NqF+Yl0DL3UtxroZSCtxOq0
P3vtRbV31k544U/ebfNKIfbsDeHyWnt8nZ1K5sMakzzsz1RPbAgx8fG0kNWSmGmtzV6wcpuOQwiA
Av6kROtHXXQf11ZIWDxsyeeUSlzCzrn5tvbYys5DCk5k4ctuMp9TCrFWSK4b7BhkNA8pkOK5cbv4
II+oTAn8g8ELLbCFTzIuk3nmikvi8m7tZ+3tFv9k84vYOl8PVo+re6M8k93tXwkU+Rp+LXa2U8+Y
Ej4IbJlz8UK4qepdE4G3bGxz6jUiToKxyJBZkQHAEaJB1Q0M+1R+vy1RRs9YkCgiV7EyXjYeypny
HY37ZbGAbJvylFba5IG3EM4jk9wTmV5W4bCDKXtHkbHbiKJgZbaZpNyfLhatGqatENUkIOhwNU3c
X2bFuVVt7FD+04OWNlnJYERpbpJzalnlSf7AYg7KoTLebfqNb4i9qwvdVctd1F6MIbY8ruxFFxhr
AnVkFHZMPXLc3UCCMS4QXToJIt0OehlCxtTJrfJvvitPSyvlISfohPdrZ2kBN9xPFEA8TC4eeJ0E
LNnmwT2ZkW20eCNCECUQxYjRWcpg897huFHue2AM4qbN3CFaT6sRxj9jEUUucj2YFKJ06TGVANEU
8UHKz8V9FMzp6lRfyJz8/PCQ40ZNfGyzaaGHswsNQDkJd8SNdmlyAr1YEGLDYz4phLgSMd07XExP
DleMglwjU+UAINRB9jJ4A9wXjk3ua8u2ZU1yQVFbqnJBtcv/zqGMRW9HDCV0F+VOCwThnHqWGK+u
ivQzNcGgubPnBaHt2v7RdWMupsBwYdwpmg2+68fZBkUKEJyPo8WY70w3/Q9hgeOBR41sMqe4YUVJ
+ZDwQF6wZPz2aAJ9YtHEjbPfWquExtsb+ipMzaqYAQ+7KEZJKYzmpgJwI8RkHggR7DExZACVUd2Y
+0YHOwlzelQvkkYGEvkc5iSPXWRAMZ5Y+J00NqOfRl3Z2pllg8uGhFbjnyOxjdCjsuHhVL6qovDC
E8Oxbyc+IjT55vnCSgBydMXUXwGDabEdLgyCc9ACH1lBmpnqnft9X0AG2vXZs+m3YKz9Wk3bIfBX
s1zJhMcFE6XNRnGNbwdi+U7JrW8mHMjE/CcvDA/mezMZVtSJ/q4tHR2zDBtYdl/IscMSit/S7l5p
/ne0kWGF2gPKA6+Fp43vtNkOmfjC8KdT4JzZg8rgeyrm2aokwsNOb2S+Dpvjj667hE/uY7IFAT5W
//CvBsQIvIYsCmFYsiyIqNnkSkTqA/CROOkuTj/FNkWb70Wz+1e3K78ddhXEixX4t1ag9tyOph6I
B33oyVq2KWU0Z86UtciHzUZX+RCICcvMsPj0i+H6hH73y9lYhVssWjoUGoysu0VXhkMVSMvgBb8c
4xUBxBqYWC/+X7b6NaB9DOtNAjiK/npd7vqn9YeSQlBUoMOynkTpWmcwnIruLb8fKF3fZI7+17XJ
fhuKAPUmWdqEr18FBkAs31gLobLAOXN0wUmM1FpPkahxARjOLzLxN0zbu2mIAZA2+lsrE6ZKJYLa
cf6npJA1dbQ+C/cr9T5+QqBs5vkFoh4IpRcHoB61StAK0fsCWFYpT0qtQHA7SaKiPOpsjBrda3KQ
804jx8KHEY+qPqAu08v2SrOXooUbWs7AUSar65Oj1AnFjNDuvoELY/C32Yn62WxuZYk4PPJpEHkj
u6FQMu+5FmPxdr95VrdBECjtbnNv3WfzLWPb1bNPQ39RGNAVI4oKe2PhdO2zjPkqDLtbByAr9AQr
Hzqva/0TOuVD1OL5blApwTQ5Cemf7CEbVByh0enFvmGWsS5HxB9Y+PwhNje0Uqa4IEA56AhwuJLB
YhMVZLod86tbA2EThJj1haqFZm18GsYxNonRruMth450TFsrBiHZcIBsbwaj0wRVkwZVsc3ecHR+
EPTIXzfcn/S/MxVN2nsjait6M0W9TPIiZ5stdWAwebLGLg01yqctmD2Qq/9H2x3wcFg9WgtZ8lXE
a83TUyJEKnQbCEjnssN53kAk1Ov2eqeLEa4gWWpapKQlU0ARXdG/Q5JFm7294t8c+DEoiqz0222O
P/oDc2tRAwQMDTvB9F3r8Cngc8Lp5ga2Bx0KJUAFyMU1GN3ktwPUcH/e8/Iy3IfV8ftWWhgVjJv5
MrITqJk1Z1Wss+TuAxNq8Q9Y2fFqe/aaisHEazFNZx4TQVXAL0RUhdaeTx8mXzz2Pgf0H84FdVuA
QZgkC4NB7hxHcKlSdiLaxTuqY0YNXsAxu8KMx8gZUJcBfKN56eziGUKXKmSycBpBINWPPMV9xAqz
m7wG21h8IwJxN7zhSE4L72C9nr9PJHkAurVf5jB5+vj3VNEfevtroI5O53j0yfAhMI2YB4yFkH1R
21iTw/8/LSF4Qi5gERNf3tvYx9Zvs9fAsTJLy9d9PqRXr0dmPgHwxhLkvNRzwQbzT0mjTXusCe/v
BPHSuCgqeCjzgqNCn5k/NwZT5X/GgRHnpic8YjF7lWGnyzRo9JNzWacKenI+IDakaa5S28/Adk7X
CwhqoFefFkCb8sFHiui2W7xj32l6huaVQj9Opr1WepFbqmsyTIhFhJbqhTmlisYbOePpGnymyyI9
gjDLNk5AwJyreUWJ88s0H9EjoPBRNkotGHOqipME5wcOwSr7KHbNn6/s1OZEs1SasjrcCoGHU0s1
KsRcbTN4/4osOOqEcb8X5jms5+vkMABVWPNzvczJc6dJhSbvJJypT6/8d1NTlfgS2FvsJmIcF1aN
K0cFPXscuPdzjocfQUqa2AO6M7I9UutWgFzV3dGniwu/GfCuSMWIjzp0AuILpJCCOtsiv7TDnB49
qVyaMGvFdmCTwqVkldCO+R+i6oYTcORoRh/s3NH9jJD44FUKlym521Z/vIjxzn7jrXGxhqOtlruB
QoxNiS8+rXlR9ovTqallQ7GEiZdy42PC5qYowARmaqWdlWaGzdcBUTefIxmTSLhsD2A/g6CSXh4Q
s+StcBgcWVV51ckowG70sVGPawnCN17s4WQXuaU0gb2YqGVUC33+BFpOrHNfhRVUjPvPPmrpiDt/
KSXYA/DcIYIvmmYC9q+9zzgJebhtVw1PhXXIZwJfDMjy3MfaVmo2yyU0iLm4MsoVD5g5DVd/NH1H
Ickrjwzj4X1RiKKzpUlycJ50omps/7WtCHwqle/c72HX/1t9ciljFkRWg2FYSDr93BHNCARJORmS
FYf+R6u7JZQhEU3EShspNKBCxfIHr5zdLWJXcW2uiFRy15QYNtE9EUJeTqJ1/fn7li1hwMn5KiI5
XpGvyJRY8pK0YbqPdMRpUxgTghH3C5839VNquK3WuG0NhSmo+Voriwt10QWU1sQMFRAWl4gm5ocw
S5UvFRHYNjRqRVfrJGLIU0K1gpiSJgV6miZz4XUAUW1KvWHkS2347bwl8jfX6+RGkZdfFzg6l8b1
rVP90OLiNWryOl8y8HJVhWSzeEkIzG9OAus7aSElGoogywbrBEr7MW3+C322FTpucQht4UO4MsSe
xMiEKAT5wHMAUIopaZfIfQJz7n5qTQ5Fh6f3sRoQFMLB6U2oAbqwVcnEH75sGUURHgniIWi4rkzM
w3HkMLy5mt6YAthC7KXkfKaxZdWA9fORSKf+3rG5fOXNFYSblFOEGGOdYyffwqNIlqMCGwYa7UAg
lQgSLdJ5NWMDcnrFdHfeGj4URWO3GKdPJgfcxTUasMT6ar/375gBqT4Dpt1ig6sL4FJSGUXr5P6q
YhxzdKYAvYL93wivbMHW8uUzIR0L1j8O3DBLZKn5dnBxtkelWcTZ00ZxH6ArezbVqQI0RmXv/qe1
2Syosclf/PzKIg/Xhrr4cEWoUUyDRWgh1pEeTTECsSoJO6dgpsSfy4Qq2qCJ12D/lBzF7YJ+EtMR
IYgfyHhcg8C67qBuPtDp63uUykbCyEbJ1okkLV8GUHdXBfZv9lhIohDlnSYhEwdvxLyMHczb4TJa
Zj6XKY69w6hWFFWdCBNhjm8zayFtkKf7/CYXyv3PUy4YAfdlIwslWwq50aYBvABmdDkhbsj0tDZc
7TcO1O/KW3phDu2wqc0ucepvB/7DDs7+SGxzX8gDTYBluqiPA9yp25KYgNR3ABIsU8NY03j5FqJF
zvaGptVATBWMEV3LFEqJW7Y4JcyRT5e4qdHmtNu9Ua1/7x028nmEwhzCGiiI5x/4m56gfwBNvJ0Z
KRCYCLhyg9Lu3YreJIW5xbjFzbisf1eZIfpToxQgEmrXHzgcfMq3iRc0Fc1gRW7ytiq6C4eT3IFl
ddMTJoLnE/k06TZTLxuHmFNutrZQh3BJmwaysnfwGv3G+YMudS+BMf2OdPyaiAjqv5V7P0qn/dSJ
MnedU7TEpizSKdHetBZXzfoPK662i8vhriDyqLzQGkj4UoiKqanV5k3GiiCQWdOfjzzcUk+BoMTk
ZTIzS9OANO9hfesAN+RqOeOyaKXDCv5XGVfErJa6BolEgQ3bh2FrS+U7IcDGvtcAD9Zt+4hqbZEf
EH3z8rOEOTXzSmM93a63vq3j6j0VcqgNSOUq4uwAcB1/y8B6e2wHQzbHHn/ce0EqzI0HoPxzSRAe
YHD0N5RpdyEgZOoUbtFxSPkC9ucykxGkj581Q7vNYGU6jAz47vgeZ9Qto2Y1VujuUpySoSvtByE0
UoFIeajRbkqWpr+IHSVpIKUUeS1VOkrYPmDVHQBI5g3arCiVP5IjPi4e0tq8PqteUirTWJIMfBF4
MslJg71KpiEpvarmezdFtrYHUdCAg7Hd4AqTv0kEo5Y2YHMRU6FiOvtMjeHoYP0WFNdmWVuwlXgX
HeFQQyhatc1DA+GxDk7mBBTh7+vo/VT271iwjxWYmS+DpEMItKnyDHNn78xFKINFK46CiZb6iUz1
Pn4iqBPlyizfvATY3x7jTItNXrUIvjMMGPXifiU1y/CqD8ShX4o9m2lCpCXWO2BQ5zkjwPBi4NHp
ig8CqrO1EC4rDGjBsI0Q54dHEOm4T0dDHw+DD/Qv7KmUhj1y90xKo+yMxVzVNoGgAvDOpaCj5sHz
ioFQ9FvnEyqslmBhrV75TcKVxzTbALBTJJxVr+XdVOFPBHVwG2Ka9H31rqA0OYwd7GJGwcIDbVlO
E1sNqNXdIHGM9+VmNkEtB/Bw7WNQvrC9ynRk8u9tS56V9ZW+jHiJbIPrx2OZcYB5LKaBbfoGJrqv
Y5kCRPhAorpZgHqCzYCRLOgGm8fmkfFBvptxsUG3wqhf5OpkbTe2rm/VQoJjsgJ64LQUHrHDnl71
OQhMMYlKRuhNDUNddx7KmkInQPBfvbSpc/NViwn9DwXx+2UyyUl2jn03iujllIahEpwlyNwGz0Lt
PpZPFdW31i2vAy92K7eJerkPV7FBsAHXmV3a0eDb3PnREeJW8PGULN7vOmErGM8Cea01uIlT2zyS
c0K1rDGTMSxbEMyD7aG4ZX+CLlxM5+bVNqpCm9YYm+gwVSMytOlyWxaRcZgbpDYos4peJkCOXW4B
HKXh1TmndiscNRfu5dEdCXjCrftKodbzkdGcwo6zSHyRIosUjUdhe6lmVor8y1KUlnvXozW/Jcv9
1tXsv2mftqNPzZ4CIxsvNvMN6IFCrqhyaei5o/Rg2BDbkfRbDpCZ5hfh6oXeKx0lRMjuu8Bf4W/D
olLyH8MkZxo8/zjenblWT+iRrQodaTxk8NAWDwbIQOtgvXykEAxRZ7SdQFrtdc6nfRnowyfEjd+o
EtHlhp2lo3Rq07tbnU5Km5TBB+jG0mNDB/8qHF9znIA4ld0QXZHFMSZTF2LQZX/lH0T8OuxEJ9h0
HSba46qoqbuJieUCdPXqlXdl99Yh1R3Afm/PrlJ+4cv/tCMba0zftJ8juOU5ML69qUHGrc7B4i6t
l0qkNZPUyaBOcmQKdatgBMbjI4TtGRvLy4Eql3XKcDfectafzQ3HjBTiZyoO8MEkibNxtNN8gQND
TZEopHPivJuQzZXbjv2itYIVDduh3MXnHakphv7YhxFYtULUH1tcZEvvVYJpJkDIBj+Iz8Z2dBVP
8fceoMyRMeU4enolsP3uXaF0lIA73fMwemOmXsxroIgG5kOICSvgKbZ2723c9aEgM3bZ1bcqiYQg
yWgj0RXykuSwdVCNJONjHproPQOchF2r/R9x1b3HjT/rRfATbNdGmlxcNWRctlGYQPzxDfVbN/82
PMkLxobGHJGfE6N8/n0TV6ovdX3BAWeN8X7HxIv6IHhc2kHEjAl2JB0oX6wINHN6+4R+VY1EFGuA
8tTLQQAnKGqHyUj4Or3kS3jM3DPCPW3DfGoaEchB2hHOcnugaeg51Dkfla9ABdB8OUSofPkoeJI7
RMNQttlEeb78Y23OxMesusHAMF2F/nbFKRtZNUj0fRPOFVyuuTB5Jmo5qeb3SG2YQ5kPlRS8vxLl
HOwBCA2sGy2nmjQukjHUaQTdBeZ9Ju/MPxl2F95KcGSMcb20zXDCRSuVTJByJ/0Url6Gf8WRsqjE
90UACgLKt8Hg3osm19FwJWjICQDB0rDacY6yyCG6/X7OzMv9IHML1K0HXpLv2P3S4zpdLisz6etE
Bg48+mz7/S8z9w9T9LK5GeVrQh+68mdloy6FRTbjvsYpXQFGovw+/bbsbYE63lN5fh6yqDW/1l+0
FL1HpobhfwKqy0dg7rGoWHQkvLI9sY2Q+yitGWCV7km6AEVtMeN2Gb8qEm5ux0fRKoihz8Iqi+QR
vlbWmE2PNCkjtaSWkTUyA85KEBL+ZUCg6QAizIMYLHAnpFu5PDA983UFxKQdh/nTLCbhw12DKeAh
ky/LhmW+PLjNJU9U1RnzL5vb7Iy/XtKohmnbqae+Is7ojEuyzkfuxpjJE5P+9cf5MKRFVQs6R7uM
XZjE43j/CO8iheMOGGVaHzboDYIsCn3aCN9N6v7txGSeT27fL98y4biVWO9utRFDr9KWEde3cdeu
oZbbJlTTl+AZbgmKSCFoy90retZUJnDaFcd7zdaX24YBCFdjCgg7F3XucJmeDqk8dAKLMRNGDakc
MdswNOyD6amqcsdpgt9Wd2e3Qq/JjQK4g6slqeQzZ4st9NuZaevVhHOiMYNuLLMt3jzzVVpeBqgE
Yg4nsKSZNAXlINdbE2gns4FUxtadPAWoBpHTXFAztjAb8FDMlDcOY7jcSpo6zNlyeejdXbI6hRj9
Lviwy17cQ2mFCxrz7OkyV/0MxGuwysp6XCAl8gyiv8g4Jmcm9mEvL754ckaXOpDfpGTxjBdrEWYY
mBslUtc+nJIxWMishBGxYeGjxtYtFhJJIGZTCzYgXXqc1LVcW1gUmFKTezPt8nU8hti88g7/KLQf
IHIPqKrGDetPEOxvXiLjh14T94EM8PCY0wENzdAOTDVSuSwGnpGemWp2lJ6CmZDDfaIC8t+huZY/
ppdB1wpsDiqtYmaSiv09LgDaIvkvu4xLKUNARa1r94uzRagScc9Cyot6vGFOm04mMlpAwI1pG96o
V2VHa5fIasuuYYf/UsiAkzbQ1F4WV9bt1Ybywf70VY3MNI25y842v1xyHjwkzOBvL99dkh99rX+2
nl2EWaf1meTjowO7w5dOcu+/1OquMdBe//cH/jUwEJU0QN1QsEgW6KkZwaj/dxhoD9GV1GjeeyPs
XDIeY2FUVJqXoGTo66qm8MdA/ZfxOm/O8277YjyEln8PEHsenoxnGQRLkLVVUfsONfKctdQXVsEu
1ojUpm7pWB57m/Cnv+8rgW9QzX6UXWXyZEll3JuztUqjXlqOS0+WKc9U+eUFvMN+bcQbSWz6BShN
efWzg1UFwiLAHTW+j4oB8uh1/eRT7dBsM7h35r1g3frin+2KgwGI2nipTKnGJMV3mfH/vZsH4Y0A
ild8S9IRvyqwRhrB0NQWoZcA2rcXkMb2bhb8HHkIWAwYGND5x+vD0m4WO1p/4F02dOgIBERza1eI
a6NK1r2Jxbg1P9MZlG9hjh28d2Vi0DiYSSiqkoEmlB3K/46lJLDPytFYUC2+BKvg4ZVzKVSNk/W7
4Tuyhf/L5sgqpmzdMLJt72ua81820IXB4UBPdjR1LSxSoCtMV3M5iWb+AU7PFNDcODXdYq3bGrJ7
AxbY5GOJsYaIIOoQor6pfz8RSEAIxnmTMwqriYpo1BtQrvqtcqq86+ByvdH7UNIFX8hIxrXS9zVN
8Th1jWncwoNpWnw8X61HRb8/BMFLDco9ZkxAfxICaV61+GOkmlyf4+s4rY5pQmaPON12o252wT/W
A8mFvz8LQIItcTuWiYXOUNGw0APq68iEnD516VmPtt1jU69R6f846saYk4N2BJYrnezDjKEPG+yP
5txmXG6nR2xvnUZYDAyV4JgOCxEFTdCrQrmDtN9NG/9zEMqZVSV6V8tAFiBocx0wDX1QRg4kauKQ
g21c9qKefQT+nl50OBP5VDww+M6xNpEezsvXeVN6d/NSDNn2bs+4nYzKEx5u70ghoepmlCSjwb3f
PLiYjxYPxfYlasR6eTYkkUKDUh1H+6SILSdKlUrcQNBcx9f0mDHbkgAFQhzfcW44wVLfo+T7K/Br
LY2S/YWve7TyyJ2hBFJ9LRNNYd/KyCMV/VqysewnihYvjiM8SzNvhAL0l4FP7+aD1/TuXMM0gO5m
lu2wM/Y7piT8gqntNXtBbJEcrbdbexHl1I+haDcrmzXgxMfiJRai9xgIyK+u1YhQ8y7omTdSI8vW
M8WxsSOYcv0/RmUm/Na+6W+T71Ih/fhOB6/ZkTJMos1ofdZs8tLvUwYkt+w39V073+eoflNjBZst
trohAVtvkgBKiDAMO8wlUnVQlYoyr3EYGLPejQwUu+orebvapz49DLryY0v/JLUSHSzUzD1HM2Vq
aBQetDAA9EWPAipevDiqMHYkwWiUxgX/wSwxjpro+4omiyVig1whsNTatmKAiOr+mbyELIb9WuDa
1gYCXZQHpy3n60O2OdSGBjEdHKw7sFbDqBBxxPzDtevQwCQOKUcWQfe1XuvS7h20xB10E1HxtO7b
fJUOBRUYgTG1vMe60Bf1AqUKf4OAqKLOSFxnHIjm08ASZMX89LnaO98rup2DrNUX+/uTHI89Bdp5
UYKcnjdgE/pzovPFuqbg+BMXiTZ8br2UY17TOLPET6oX0jCPme3qzTTX8uYNKrUsiVxJSfCXzNGx
D3axfg7gPQfrSql22HZGnshlvJP6KvyMabWRam9Gs3j1JHdFs2owW3Q6VxEWTVxIuaSw3BzinOP1
BRZaoTPoyM5iuGCESb/XnRrq0rYDo/7D+ZHdfQhLm1aUmJNWJ1AQ/x6ZLd8ZF5GJKEz8OgcG5ZDs
PpRuuuUWOiO8hpXrGM2xOskjicWrqnPGrDuAS+138zYCwR+drHiysmZNVe/N1Wom3dWL4CaIAE7H
1eK+zyLsueL1pEKcuxFT4ppEecteIGlXAWG8pkeEftkmHgjMWad/tBZP9iaeIqoPY1zdzA8DeMLu
jYITXiKCukQMjscBbzO/9yGJ3Kadb85j6YwzzcJuLaqQVWjSIotEX4hsIHeX2pA+MqlHYzQ6ykmh
yt7lX/FXjNqCOMF8vLXk3Q7xlbxUz/tV64TcdAz9Xa8GoVhFtN2/15/M0QivBsha7ozKHYw2OOMf
DwjGQuJHPJo7MXVizcZI7moYCT9kaZVkcuwRHe227WuwlGI85bmhnjBrKS3VqEXBgdx3bGMAhxJQ
0Xi5k1cyOAcUq2G+aS7n7PxyWxcOo0QWhgY4I1B1m26J+x0pjBKC32RWW/sWEjtw4JtxBO+ANm+K
EZxJDC2wf124w3yvX4vBPCd6EVuniqWLSCq1V5CjMWStOXbGjf9NGXSsl46C9UXzH/qd7mnf5m9L
dGi5Gf3bj7Oqf412YOgELYIqZD+ayQZ0GIBDQSj3sTyJ+aFBI4VE8M1DmD/vWwhsMN2e/UZnvWjg
HYwVxQuvvgVd4rFqBjclDOZD8Y1riQB1yZBClMA+s2tVTx9w4TRybSLVZ5DOjki+VZRF/hrfsxAU
6uvERL13jyu48C5DMskYzlrtllLXcNjld4GIakJc5OpTVJiMc0alHwvLbyNxY3oV9vPoYNlDfeaK
D14dqZ0ZpMZxz7FA23J7hnng2Y/GqRGQoRx2HL/F4LC6rxCoVbuyWBhY1/Hos8BzfX6xsbCWQBqr
EG6Tfun53rfcpfPkRRo3ev3lsIWOJYnsszn4FYOA6X/tqYz13aCOtZ1r0lLSPFKGeqoKf7N8zBgF
gNRonynsvYIn7Ys4+dKjdubQ44EhtRAjKpjy/FOMfcVga3PVF3nu0Ol63PCtTYcLOJMj7v2rz2Lz
eE+33QAxIzVS+j4tfo3LNsfaUgSop2YH2qz3LW5wsd0IfhpTGul0NWVoc8jWpyDGtxZ62jvGhaDL
4mkasx9PctUG0TBWyb90NjHUPlztp0FUwiZzT7sllxv3N2KzIuLwOIH6AsDEgaOaxXdOqOXilSDe
LLOzr8pRaa4gCmrmatUtjXphgC5hhY7tn/MRsElzgCTXg8gWF71EfgvVYR28cv5qlMwKjrTRMdzL
Scrju2vAyl/hTyHWn0PECBTE+viMvRuGR/TPsQAcEst//wrA97L7E5LfOzo1PRpsawPAfaIEevtb
pZxqQXzwsgCfvdRF36O3DdN2YFKfs6hfx7IwYt+OYsU8pzAsgxekjQfmtMssVHd8JqjDm/n+rQGZ
6CQvgV1nXEwdPXFv4KowM7S9FZdNH3VLgAzs5GkrMmdGVhJOItZlYSy3yUHeDipobJJjByr3tHn2
r7QyaXyMO6LyXLa3yQ36iCOYnfWolRGEjermUNKkJUBr59wl1nZSmD8k5EEFE0iEvehtlrQ+Kzxa
ficVJoDkYfCvYiJuM3lsPzNGAV2p0QmA/SkASOrJIMkcmBdhJWPRERhkOAsfliana5FZoQPDKmFG
ne+X4VwRJnjD/Iclwhf9MQFjcqEAp8dEBZL3vByEhyM/IqwVNWBndJlxRNY19eP6wXAhuwYmX8Hv
LW9UG+c9s9JDJZU4yjCTkwmvpbQMH9ZZbSwrHh/OgTkIadc9qZEIERhTJYVKU6+ItYh8hYNmBQAe
Sp/FdkQsDor0gKA6CwuOWhtr4oqb4zoedfosX/W3QqtH7gcN3nhJxC/MxdR2ymuK1qayx2xCdejh
dMEj5YCZCmgnToyXJW23iyXP9d/FiurowSIiDgqF0/5zBn2D5+nGb07mMPJwvVT5drHg0TOEPHUK
OXA7MywUJIBP89sCC8aJfDIypnvzWi/mpD+/M8Y3+8Bwe/AQzOaigy4KF7NrFePMj0M9B6ajU7Xm
z5ioDAk3FcaNZY+3G0Qdg5Y/nqfxsCvXrI6Jc2ipm60STDm5SQYleHyN/34Vf1lb5kS/0gFRbKRm
Z6E0diHmya16BVRg2EY0NPIFNHQqv4V0LejPTPi7o/FAPysyYVGgq5UdNiUMqxuSg/WBmULRnDyK
L4fdf2YQ6YYWdkQpY39ob28/R5van8FMYZmDl1gpIsFjhhjUNriVOxtY/c/tpwreQZh61Ef2nJj0
ofpModuk4ZWRChggSrgu6rzAROHMb/M2QAXNSdh1R4q/qeHAjpAiC149jlFFzX4i72x4hjdEhj93
UJ7nkA+Zk2dDr17MZ5tDzu2ZJJsx/JPNJeA5W26mcX0rlVdGk1YjPWbRAaZU4Ivj/UJeh1MBHlQ2
bPH6i+wpEDe5bow5vs90a+I3kdQCvF4+HsA/9SC3HcozQ7SMMN6j/PyhjtNufxaDwltrgdx+QvdB
mtvepv9OFFUzyHUy3PPiS0a971DvK36UMEQSxUu49IEFzIXxzVHtkZ+SfIRZuzyOZ4CUh4EMOi0S
7QDvWDScYrHHC27UswhDMxBFBWyL/FpgOtq9PdHtRqNL1J3G5qjG8dYUO9AtrdOtXg9TX31hRMgf
QV3UcMt1xpsd5AxOLm2YaXJLCnHgT4v44bvP3KXOaxz2An3EymjayXDMeiztXy4Ue+VirEwd8yBM
X2usLSdQA2rM/FxIeqy5duDJnyKIu7nxy2tDEvp5qHWG2fCEy9xXdbnPmhWOcudhI+19HHr118dY
Nu2EPKQfpnpv5DV4EXeMoEDbPRUqpz3ZoA3wdjx4KEGdAo9/20jqPc57A7LG74Av7LyMHYsrCcSw
UuX9rTZlZMQ+pPPNG0Bb+ugJ5SXeIvS6pcoiTtjtWXY59xzZY6+QUze+4e/mM24Ywu6VJPkKPjxX
TQ8r3dkMdeyjvcrsXiOrf2BAoNWaDSnaDHDOCC0s643ceLvs7Gkcp/iaFLu6cP1mzPr133R7FvJ0
Z41ABghx4hiyJzAHH6KDsH5IowCWh5LsZkjZc4xcOowp5ahQIjiTDROSIMP5rBuA+iO4YeFwaJri
uPLRHW3iSWN5e4XN24vrck0Ep91ZRod/YVQ2hs4Daf5CdzPRcENN18nvn2r/7RZFBMJLg+REMFhK
fU/6O6nXEnljRxnUNSndwr3rE+wGcoBDAccDlCcKaFwQtLJo6RJ6BSdlaoSdRgl9EuQGa6YueST2
IBFHxaLWLfPKYD3hoqe/DAVX9pFQbxWCTsD+DU9PplY3dJvYBne0dScVe0IE9KGkbs1rFj1udSGk
LUV1Sa9zaxcHWkNY6w8AxStyxFoAW52SSIoXWg0ZlmM87GLpQJAjVZYjFetVHzXmenPEk2P9vnmF
VoKiiZPsq7RFYaG5Y4uH0NwwtBreO70Fq6XMbQTjmMlPh68Zk0vqrL5oE02A9HXyhgek+9/1cY3B
4FxMkpC0oMKNUFsoMdiyrgh5FWzCW4qP7Qp99S18D4FCQVVtwQDJTR2IpAOxAUSBirZCF3/EIThE
unhuj3D5PwBf9+C7ugAtfaePu32hK5dW6+xQkEcXTCQX2Vr2FRU2f2Vn8AzeboGxl5weIwT+birD
HvfdnAaF2V8ARXEMOHxOpPK9j1+HEI12duOQs6eQnE/3we5QbilWs5JDgPsCNfbxUuGdywIV0spD
cHO7GO1AZzhAc887HbcfMJCH4Tf//JBbMDRBhyIYiZlE92GFh++xvqQOkxe+fG+nQ4P8hwIxdw99
6J+N23F7wFzBvOfe9ZV8QqtBh0M0RjJekeZVyS/HYKNppbeZxLA2SEFz9dl/vXGQGamrdh44smFh
tw85M72X8X9sX7VizzCUfLJJ7SG4iCWZiq4h4u7VNGJfAoCsATj2F8VqVp0auxfZsrEJfsg3IXAL
1W7OLilRzk76roFl1s0UaFpGNVz6i6yaXAXhqBqfWwEX+iCZhx9ceaVmBcc9LITflxFqD5b40JLh
pwiKJnfQpZY/kgown7/mQ3FUJL6fu36aNxj/JxDKQuQ7R0a46ra/q7jymyMak/P8MVDIxVMb/43q
JHsDyUHESi+NtE5RyBGKuBUqMY0U+E2OOCrRSCBmhNq2p/A4Ucj+589n/wrfDhlCeHpk7ZQMBa0u
I/aqUR7NrRRL/dN569RRcLs38HSTY01Vqsg/pnarZwzeKofCQNc+v/w5/cmLh9QK0Jugeld6Obyi
ranAUm4qvRAz7m5h/yYdlMvyNBAANJLasLIyTv69FfjviPNAAlNw/aExoIvRH7hkf7jBYOi1EkrB
DRFy/8T7Q58+/8zoGdZRJQ6zOIvqdrzToUtdo482m/IR++ct7jsKhIV7SqcTt+5NasGUHH7lpy9Q
x5vcNe6yK2BymaEqG9No6HiPCp+Lwn2wnIv7krHRDiD8ZEZeLOSaRYeL6ud8KW4y/xp/ogogn0wo
o8fqqzBQBOK6HiSK7CLQgFsQ0/7uGFYu1MFWH7U2NC34jMFvTaOi5jrMDL+4n23SHkDPHJkB3P+7
K2HVP4QAgvesW2YZL7ps1ScVlliFPchLusyE6gfE1i9gyHePkqGtHJGIGflB6S2XaY0CLmKXpMhC
+VfJBwmswgrQNpGaBQj+OI+vDPxXE5by5MoeBwl21nX5qSnNYuIua3n0PomQbRtCiKk/NdUAapYK
bbsAwSto1OvmjhFzEPtHm4vtZTKLjzqUJOHq4wdtV+gYeUjATd/OhyB/mf0SWu8PeCSrnRkQmgif
Xurwv94F9YMf/u8DCb8FKhyaRjlNB5eR0com8972zzVorP2UH44b7EDYek7FH63ynzTMi92z2sXl
cAhG4HV+hZC1I4PPOpbEe1FYRNQSqqvtRdzUeEBE2csfJW4ybiNl6ZyCsRzu7VFKGzG/8loXLMUq
hqWWMEKYd0gAjfnoUg3sbV+8uwXpoum4KpfoZGJ8YPdhvACylHW1HSR2bB253EmNNYcBl9mJZAMj
QkmiOEVL1SsBguOYI1qRwHQDbyVVEWk2oGGXE9djNUDcFPiICP7mDhcyOc64kYRV/ZINxawWmPGt
U4D+CPxmxf0IxDagvXIUDI9uGrSoGFMQFY62/NrTCSScZRsHBhX/uM7hQgZnQs2SkTM/5aRgFYoi
Sr5c5ps5ufKjkiPgaiLfC8LxPUcizyXj2nly9tHBMHk9ivySlt8wthr7o+Ag9uv+bxo4vE9HNPsH
mvTIvfai35DWbFh7IHtypEkZHuaM4CJJ9Vs2jrWwrt406J9axMcl5gozaRvH1Og3NTbM21iAeoEF
PWflXjtF0v3MEkIWKie4e6ZXeog5QCuPFK8BJqOSCqgchvWzPZ/UriNuZCVkXh5+mbAjIW8sY7M3
g+Ctv4ecHbUPfhbYu8Pss1Scyr6f/9Azp0UdxNGQftIlgDDpEGshH8speU5JKybztvP+M3qqJV6Z
DDmxzri2zxg5K4Talw3andqz0b/e7sAL7wOHqjfX9PVxLqxlDHX04im5tjYjylDuVMPG3hE/oVBa
9JkxLUBF11IsMeBFXWw6eCmmNxjRhsdshU2yU3lrgRBNumXbRKYsLARK7Fn63V17LO4GKAyYSsfk
QTGUfzgrnACiL3sNkcY6M7n1cBs1qLQbHIiq58NegdOljK3VoXGILqEK80TumNiMBk45L6C02Ong
srCCxso5lDwsCl4DaCZY0xwWqdCYta1h5nKRMkd5dVwRPK1WrJiY2JHxswjzMZQoYN2hqs4kJSIi
0bkGHVFlBrIKwwOp+gameXyPFHckFDPA7SJwXfGkqV2Go0fykqBitmqab7okYQAU3cbRFYaz57yf
aOiWFK41PECmc4tYNx8y8p9BNVZRBoZLHsXX/o/k2Keck5YKWOBqZ3XYZkBBBzzsgU6TyYwDqU2x
T/0/S0Kz9FGlZEQIBxBkkTXswunUqKT85TAkEzCeLa8+ZJiEIHoQNPm4AXagUZLts+zKaUoMW6NZ
0ATdXsB1/KK4tOQn3gWyx2ge+wLwz+v1t7ZVDJPsQrENKy0w5tab/pcEsjaaEkGP7VxS2ASUSiSM
AH9i8K3+EmLWKzeDoNHbjDiNVlCHHmvH//cAgr0sEg+efvZlHUEREyF9D+7Ur9bGnTbn2LRD5yX0
UyO9w2cLq9bIvQE2IKtYY6OvWo3TY8Jo5CMaAXDqa7hNqBM7DFAQ/bVXbFJ1NIlQr9aDqPBr1oBz
Cl6tvP5YO3xgnnfa8Q8z+5F4+u8bOjvmleSYa6Wm9nVOwRtU49HCqCj7J6cgeOMnaCPdR1ODW+Q0
pKab5niRrjVTT83j2Eoo32/ifjzXtWSxYlS1F/Lc8FBmEcyNuMN3ad/8mAVbgMMbFC4zaEfun1sd
quY1qxYVL8rS+7OJP/D0nnaK4/9699RPDzqcA+t7/VmO1gGLOKStBCtoC/GovFyRzZSXxtBrRh8K
4hFttzebbw0vY0Qr42eJu7PvEWfLnJkkCFPqD63Z5y2x6DGVo7W0Ga/KNJq0Fh6kGS4IaV5Js5KQ
UBqmQvGie9/FUFciLDCjRB31D71DmhiOMhNdYTW3tLh+JuxzCUI5hYhUiJYbOa/ub/M9eQewS1Xs
FjIoUiuLaUeOCKVzdpP8nBGRsclqhJE4KyyT9ytbjxktiHWlLXG8SSER3o4ZmoUSaB7LMifsMdf9
S0ZA4BTGWUMVajgtI3Pu711ryOP8kb1hXzDmcCujTI94PUfF3sAbEIKnBmHzNrlW+0Fsdc09odf1
sL2U+z8Df/JYnkqaw/0+nCxj//zxvsaIXUnsayWOdT6U3NQuEQjsi7rztT3kUq9VXSIJB0AswNxE
qGx0RtdAzyfl94opG+jdaanaNQpyBSEQ9isOK2eKffi5uwTfmlgvrY+wi7AkNLBTBwnFk8OAiaOw
A2Yt58P5Wi4ShEpRRX7SSC6DxpO/Bp2yvKT34Pfm7vLsOq5TcC3kCxME2fQezL1j/LWKLlL54yl4
W2KQW7yWMIfnL2AwcGeXh6w6zUeD059uYhh1XniKNq//1Ae9p+5rNWxk5oNaPekpwtzGJ2JFrLp+
26LqMbfNoIsKEtUMt54mmfFycIKmksQ134W4VF4qSsmCTwjBfbwFvlhbpXX4hMOp882hhSHxjt0W
mGK+UCKS0ShX3o5MJVIiAluLjCiUQMY+b6c+MS+R9DSiA+b8oPtz5upBSw9UL3MtuVMkXl97yebB
76EEY1ESpHjP3IStFWlLWpYB/xT+OTqv65JfiKuh6eFLC5EE3UpEwMK3lMyMDlnoLjYxeoalN8V0
5XW542weJ6owqAaGko+xaSHUYFWthS8IQDaBFg20OxrTcXUiZ0kWYCzUabGjnzl96fkJ+vTRiwVU
qFvgdaraZcpqNBSEWFJjLhMMSwfUboQeywDKkdNxymgoSjtabZQlNK3bSSIQ3MEkkfDk736KXlqP
vc1yIt9QbvT+pewcF8V48575PFNkrDo9wh41R6XscUZ+j1xPnlFD2KQenzDiobe5AG0fZUFKMb7U
PV0j12hVbbkeayFnV4DiDxBG4+rUbc6K/5tII+Zbf/E0zuYG1oHCLFFpxq7S7TMO7vZURL5uLQnY
PGnU9F6GpkaTaVdLysEbVKSlJSJMIYfYq/Q04HMW71U6h0MTMhHBpPFqoHzaocYzgMVwtwdnv/r0
amYBE22c9FPpVsSMKJ6Snv66TCPCi/xllKDqP0mmy2MxERQuOGupurwBySyLQ2uVNuqiZ4nvOH3c
tI5Q1DssXOUnzYhEf8u4NEWQu6J75LH2Xw0TVA3UmS85sQ0kEgnvntuDkREH6ztMjjnw2Fu4SoSR
Itm4TlbF52LErv4nrVgijszn/iLLY0ShLXhfKms2gtDnZeEWgDhI/UvpJ6ra60bF/nIU4G/8b93o
YvVz5Erl4WZl4e1NYTsdNwP22+qm/Np9Hnvrd+4IGMKOuC6QphVG582JvVLcaYosKp2bDUS0ix1a
t9YNXroLZ1pte+l12tuyNU5r+2GYoF6CHEDmji0t5qlXN4Zm0zzh7NN5TgEulUxfxHbCNO/AgfK5
WhfHtUT/QaMjyZ4genm+zMBcu4DzjbGAhxi7cYgfGVc2odfYSjqJaYq3HAFjwH8AYzku8fkreCUM
5hVcVDWHbiIhEIRPEWXuoz/lwZccS2ZdJ7UVmL89Dld2dmPEWbgKImL7ENlQyP1Jb3ERrL+pFKKI
jIzjEMmdfGBDPvAeDT+Wk9zZ3lXBV3R7UOZ1cRJ1tAr39zCYmUTcp/y447lO73/L0CLaObu5MpBH
+woJG5xH7WMwjJNobut460eRwu++GdDefMzN0Xbq7zLjvRztiwv9O7QTz9yYVIR4pM0RMY7px8K+
Ek7mnM1T1MNs+xXb3208FbYJW8hXwKcPvIAXcSfZn3DjX7BfR7Xak10xpieupZtmgc401RgpKEAg
XeQMYTFSik4sK+O1W81LpAGe7o/NbiNk9hmRFGtz7c1lSNQ0kBJ8xm6CGRt0sr/vBJSBe9+GBa6y
ZKSv25Vpi32jUNspD3rrwQQKs8oSZCGrpch/O0Bme0R5hlFodQQER1r+1s50BarNvHCeLRAxRxAe
StjYY9/fkHRJ7PWs46Y46DxzGodi8w4kNdCd30RYuzlks+v5ty2297XB3uD5n7qlXlLB7Atqdqoj
iawhF0I4n99O2jQp8PpEg11fw3IEnarcpB+CME4rdxFMLu0eeiv6VS5L4BS0Eg6W/ThZXGzdugin
kg3UDVXjvCtjYtIDonOfAOhZt8EOU57522Bv02j3yTZ4lheAby1l9CThbmsHyYWjDTV6XHQ3lojV
0aywFn0+DG2hHId8jOfqhmfUFruljsd+3AwRssf70OPeJb0dbuDvcytj+OHVaM1SuyS21ZrBCl5J
d3rMr96Swz0LpEz1QmHvPNN8Xj6E4dwZpkOFwjjmZGt5lH1zJvEE/Y3KhHmyDcc6iMC2GiwEpVCH
RP/PtWs3r84dSGmf1YWG5imF8/jXn+EigdP/hhVu5rwExJnF1Q1SqjsXudPyyXGDoy/arwz46F1l
l48+qFouwVPa0DPUT1squPSYv1TdEqq8QLcNnawXOCKDQ7jhcDkn5/UvDLYyNoxovXMj6mxdGgfF
umbE+E9D7gSmUepgL+URh0SRfGfoSedmE2/q4gBdwpIM/qgyL0JVNGPMvJJ/44/leyNP3TFWbZSt
3c38YyboP/ASnEGxYOdwJWIemCW4SDZVO3aqhnE+78P9C6+YkJF+IwAbFTQUc8ZMNr27aHNsRFjw
H0mSXOY8C5OpThKQEx0tYM1iDe1YLC486DkWXxoITBAzKBxTl4C4qZ9OKQ3ogCWCkRFgXYUlB7NB
SHfOiaT+EGOUlj/EhH5d8coFStSnKJ8RQsG5K3P8PCrtVfhsmDv38GnJGuzphgl4dgLYpQAbgPMT
961JHTCeZt0OdpmozcOE6G/mH+BFNdsiIN2F6/uAe6Ypu2EmqjaKOCS12kIVqDQxo10mQ7Sy9VfF
7nwV4pbOrVylGkMHEGEmawvASxTf2Gnw1qUZIcoA63Z4wzp2eNquCXCZiftCZ09tWjY5bWDNyFHD
SMnf0+wqSGuuR03gGXXO1drDxnFGlLwvojmItfHg8jg1Dn1KPlozVlU33UhZY83owdsI3nGI0Cx3
7gw/ifr/38/8yyIV8fbCmpAdK4KO8PI+e/pbwFn6dJFe+dL8jvY+Mo5MhVWdqMHHW+eRVsTUwy3P
497UcqS8GyxNpT3xybbIgZQzyEoa+9awrvUkemLPArvT2AvNOJPf5znL47amTMD2CdhEwkTiODIp
0Y4UBier13YB3OiXLwUxlNrPyO8Mbxnff6/ct4MLb4chibja5d37q7+EpjxDPG31EQa4o+zGLBCo
iVhCwNS7cWRyJHcIHQu2voH4TDyNHoxHvp8yzGuGWouO8Ci2p9Gy4f/ADFCJOFbvCrHzOBAUD2Wh
0eP2sJA6/O0f2vuY14ha0/qCgLmzKz3TvSqLi2wPNCbl8Lm5tCpIn+RJ6jSVdtyqS2SMY2ELmkxS
GZaJ1qJ8V/ImONDMJiIC5U4scb4nRW2fB0Q3uij5zIdPtjCJUS4Nd2RnDOa6kawK1yNWVpCBDbeC
ooREqz+M+4JFkOX0nPthYxIhGYPtimQ/kdPsZBdvQqMAEUoC/t8hh2cN3b0UGh5h8xDrOcwWHmKf
lPaAL9f4/vT6OX4F1z+tTHO7NXciXmcll4ju5SQRSTiB+ScfGzk4dwqrkFI7zXPCZR3avXVC8YCC
KmL5Viay6lbE+rgmm450LP7ruys6I5BenXwW+F8PqQZ030GapMeDfQSXE7GqEH7dAs7t33cIVETK
64B2wksMFQJ8atXtKOg27a24PK+EUJlhvSbofMYn/JalueTGOSyYz2nRgtEBlzsJwrT6vAwAYKeP
RQZytUd5HnOr5dnWNhQ8WJ3A+JTAwkQMoVvzHtw9cLB9AYXdH3dhBGsypBT3E1mgRUvEuT+1TJ4d
HFc1gyk+iVrGmorTEqLS8XsAblm8kSZRM3RzirLRiQVupDT7eSpZ6p1BcXCuMa/SK4XqczVbnngN
ssWCsG3RCO9fiITNn4PdOFHqBzOjlC+3z4Us4Cr6u9I6l1giD5HwsLrPQNX5CD1rczga90P5sH9S
Esw6ksF1nBpkgN2FgYylSjiMgfEXJNXx4QCRV0A07NqXr9y1Xcbks9V4XP3bkXQHrgeEVVRy/CgE
ojnFe1Gnzjtzl7q27GtbGYg4UT7r8gdeHnyaVOwWw3B+6MQ+gct5ZXF1JVVSTDaMZEd3Dbgj3DmJ
7VZDuGNzHv1nBjORXmOCPpZ+Ya7pQB8WFVuq0ReRYLicDfb5N7fZH/px4ikO7qEfQ2A/WZxtPI7l
XkqpAXktuby6SIAkwDJFIxGLjTHB9h46XF61Xuk5Vf16rF4xtB0oEohlmOyivj8qPjKJSbtREOpi
yPGzZMcf7d+i4vnSN6aTVZG9/+kIHiI2bdVISqoeEy9r6sEievaKKRIIUdzCJT/L+H7nrTRvmafB
WTRGdPabgyA8nzO/dOOoGOx/OmOOxpIvypDaVUl1Y8gUxvMsbVblxeSL7MyGs6s4244hTqtr3xNj
07bdG3z9+UICO5DFEeru76yFDfPxvgUomTy4pjMgI5xKyukmp+qc2cTPJ6ijzEsbP08VUgYVyeCB
mS7W9omGu8e+59N4ZQX3U/0TgZXYP4mjJLtQ3fpj27ylKhcRS1Q9F9pv7t1Oe0KrM3q75O6CS5dy
v2UsegTdmWTPu0JmTzhx2BfQXHuEu8qjWn3/TphDiuTMq0obuqT2RE6D6qXRyRzQ5pWTF+HZ6nsr
LJMM+PUaYNyGvxAxlGU8FOkkDGOzEbIwEWXZRrinuOM5UMBiI6PRsScsgEkg+z9m1aGs9C2bcBJJ
6aLdNjCWZFI/1GNN7wu5SW69tuyhIl4ZTggOnxg6X7Sno97+McMQLgdrJrxI8ilE2v9+d26q4gBo
cNa8HbJYyuN7TXYAZdPNkuerB60HqnzDuAlPIg6B5WrrZdm+/yO15CobRzyOBQq6Kg2dSflbRPCo
jM3gFUo/xgbYuAYiRY6/A1ZLmYe32eI7i7Fherq73DJrFtdvF7dBg6P/G0j9A/L+QClwUYrg+hHI
8y26wfKn5FKzncmm8UBjAcK22PlJr2ch41duy6VjVaxwrYmVrt1wMv2Ad9UToYgq0JfQw8qyad+J
WgngPIi2I+OF8mMnnVnMxO9nyi+Mcp+/dA8TVbRSKMtdvcJnBiXXahjmwV6IXup3yyriwYciSdrj
0zrneStnHukz9iEKVYIwS9gzm2lCKyVWJvE17TLBo1ww1iM4KGVeBRuhcJeYTn1h6C9mrw2K1rDI
dWy/hW1QUj78f8sHvmn2Kbj5wf1u7WwG6nYlBhEzcdZEsB1Y8OVwufj03B/AJT3YZRTH+bdxEO5R
7akzut019TESILCTNeVoDeJLAq/M4XNQjAIsMnlrXQTdbeBo7eTjZFjKNF727+YWkFarCRvSfzey
OuH5ZCZQ7hQa5i9GrjUNqWGtSSt9nojomKZXmxUFBBdkdZlJeIOZiV7+lpu0hAitdkpoWQq/Czn1
Yg4XTFjGvwz6EO7VgiEeaF6a6lFUfI+SKYwbshSppZaLNLyEP9WwxNsl6KQrYlnmCA/v+ml9H0+c
PXTdsjbf672n7MSrdIaJWngCBBXm5sdnRsqcyalSwIPYUuZS7uJr7FiLSK5800PdHKtOcwDtFIF6
AfEbUUEwkpj1Rfy9Jha8zwoIUr9ciZAoF9zVsnOE3d/nrYAO1rLV0cihOd0RjWg566o54byo5SHA
xqVJKs9lJA0F7D6sEXPdLivC49eMuyp/V8w298SF04x0c04WFsqk+naJ8Cwv+h+IHPlaPRBzApXr
qwNcMtUdvRx5p1oHnTGQsdJf51LB7YE3ksXnHAcDPR04fH3tPRJhCigT2jnTXNuGb5a0NdrI1c1g
8gHaBj7r6zMOirTtoeIAFsY43aLWZAAPfmR2OJ9UMysq5R+LAt03FxVlApBj/DGkbrEJLYuS1OeH
b9KBHqh5bbB82NxEIJFzjFrx/nVDjVF7WqELf8ArEPsc0JVT3+KN/VXjycitumhgFIgyxMoOdtek
dr8+bEe4f2JD+zu9Pm5P2FqfJfF7vttzuixCIe08lFdd1FdDHA/QvtL+jF0FGeTLNP5UTZtMNwLo
FqV+i+dVcGPvNkdjkTt2PWw9lqSllYHfTEczNbzMouzwjz3SEyvlIPgmZTiy6gPJhxqUM6yzUx2d
KP1iQWBi15GGChLALJXZm00ASAkRLNIS3j0oGRFplmi75EfFk4uPB1CftsUaPT3+TWZv8INxlfuz
iddHj3OZMMLAxz2256LZMoCkfHpymwXBav89ZITwDXtMhvrfdHvCkYE4XRsoo871lqlEsv6j1st1
ApTpvN8oX1tH3FD3hzCufnfpPIgNa3Ne4os8oFHvjAdYAineayynwQISjw3edfh/XuQR2LKJwI/4
HW0/IltdndW8kexBrlpzCKTjx57BwpILNx6vf25bcpVm+vYbIL/0NSdF24cPeiNjVxkXmpYSK6+M
xjw68KZ2r7GDznQulh6qiShEewU7PEHXR1vTLmn3Dmwq9IvsYW8/D98XGBijtvOY1HNb/12b0FfO
ohjrfxWDVYSeybXgYGfcotjERzD60EPiKDSLw/4cReL9Q1/AvpFvkqhfuPNkrkxs+ptTXATNj6SY
j/aHbbN8UUPTP0U+OXLQZ7GIY4zhUAFU0naPYomdGfywRtCp4AezG9PeVR9zjhkQuFsH5Uc6dv7z
s8aFwrcziwqc5J9pa4djad/zdbmZFAiaG8OfQKvyi/R2E7/Lk+gWYK9xeNQCKvOy4wqZI1O7Emfz
7Ftv5OQgPTM3EUtiNgRZibZjCNRihS2ZawBd7VGfjAeycgAV1sljVSsdb/B9LsAo8yYpBK2+/I6w
dLFl2zxN0O/V1x5X3eA64ksA0u1RYLGXqZ5g7xx0IbFxZFF7eg+60GJ2ZOuU3muKeogtQIeL6ACr
elNXKsds6vMvo5bsuyLiZxAiUQ9UGAttEJXZ5S5kRzXDknsX5vaDl8mCzHJ2LAq7uKuuh/yFw8qu
fgyVYYh16t5xruml2YRRoPJbDm0cjMN3BSnERmi1XRqTWWtnPz0yIT1WI81/FyQWomrCglqB6u0O
E1GDTdDS6swm2KgUGB2mKi9YofbSDe8ihJyq1FFCb4GOEAWmL2dryWmXaAQ8yvHBXSgJ62rVlji5
WysbxSO6HN1Y0oIirBXwkbGg2UImX+FjuV2VrNLayo1KN0EqM3ovPwjQJc6TF2iKliuQnm8u8YMO
D7sCRqWbpRrJR5NtpF5VAs26OiEnehg59Zuchef9wu15cQf3m9XV1S2MT+s1YyYNaCRgCnNDAmPo
cBAWp7InvmOwm0UY7nIy4ZMSAal9nGFUFa9DTxQLjCq2DX9Rzu/7XftRuhx0siftB2hLNjp9uT1/
WbptNb92Irpo6PHQIBDJxTMI+s+aOQp9JQcPK9PY3hSdAFcaRCfYxYk3a6eHsvL6o/wAo8rDgzHg
d8hB/OngWQdpIZLjFW6K2EFGq4ZV7wxIXWsuKJhC/gLqdkgIQz9kDzq/sexu5Bt7ZT02H4Uvb0QP
cfUVAWINxz7Ax7S7ULFOK3QzxHkf4eUxq9/xHes/g7zWO5vwnf1+MMPzeW/GJA1CbTETDsXp63BM
TSQxuTuXtHlRPYv92HSoMKBp/yEjQV7UBx5+fWARWqLah/mHVviK3R1RPf91NnQ2fVlwq44aSyM/
yZvqkm46M/Wm4IjC4dukQkCWzW9L4MNRu+CBsdWx1OILCdvvYgnv7ocSYi8c7/RxgNdjTYvhrYG6
ZCU6keO1j8MPxY3XVMCMhAHIizS4JgA015PNTBLukufeFk2fX4wUsxgEJa6t4TJIDssLVrDHOenw
qTWTSJCX8qYCkqBVUKUcy1gEffNCzclInjjFvWTpTK2fbolyNFrtF9XtRbtNFyy6PG7dzxpHGsbY
WDpMVIhMhCilJMox4KXDHokutx7sYmn0ULpMVk5bryG5CcAuuqhP5oPU6qSIS/SuqjC6RJm0k78p
Z6Zw9H8b2W/MD3XC5sDAAV8gUo9QY4XIhAQTOTNxBTHs1i0wPXIb9SijiFwwhmBaXmLiluHhKTYP
9bKix2y1VxusXss0DCpFX5p+D1K266/CrqBa0zRH3Lpdq7GwOeJN7gOeqwBlUHZuAzk2JAy1Hs6v
K997gIcea32XUfY0hrsoMsW1xhSzAsJZTOQFELFXxp28/DD6ungh3Y6Rv/nHVh3l+TmmdedZEA6X
UkGjcYdLZ9D4CDAAoFGpMxukbS4MaE/WH4pGgwRaJzEy4DRIFfe28jxBuH5plsUIhwCyyTdOJpHR
R4SWI24Rys0T3WH+Nx/zC/SdCFaJiRU2NkieRaF7mP6Ek6gMhQSth110dXMO6+pn8fJ+A2h+yQFc
ZFo16MOl1VUqmdCzlGnkm8U7ACbXqIIabwO1K6okN75BbawpvTCdchVa9HwkHfBTW5jbO2YDoZAy
0Bgwp1DfgNghtlT62nA66I/7p3nzK3t+uk8/FuCCz9/QzDdAxap76YS2AUQ/e63WVmxw7dSj+GCS
XzPz7ctvBkNIt+K72qBuGK4FcOUhK+dtptRKoTl2LBXHSYgqi7vO3py1HXmjO3Wa0II0YbItp1+C
0+Rxc00sUce26X3m3NTK1oVWWnQZ9D8Yw96+jZfxTXiQ6XW0V5/ZEaGpYS9dEVPXc5CAPRQfdmkn
EFOK0TX7dbXYsXDDc+8irtn3LoRzGy9hpoaXmAvuN8iB7Gyo4qLAW3bcqePvCSbCcgETyy5ADUIp
JcOB+UiNwljS0Xk5HsoTV7hhD0fopoNSyf0gG6Ct+93e6q09DFLjuiU+ygdNKf/+5GGBnTVMsEse
Jbkpz+f0QTu0aWH20MgcA7FZ8uJvuGuGV8UKhqjDQB+TztcKw+fCgxpcCpmdCvNPOBu77SMFEqEs
HyPF3d/6Fg7+l2dq1vydd8VQ1IKzjnV1JsNjS8jrjMMMZceU9iBzyJkLe6Yw+AMI/fSbEk4jiK9L
sUZfD7r2Ue+jXpeG6MqOA7K11FplQpIrJKVNvIJoI/gY/xQ0THus+SImf9Tt/Bc8W1bWAtoKeaPa
i7O/1v8w4vy3yO+FFLVNW4coRDo7nB8zpbhsjiBNqSvnKj3vUA3SXxrNzxhMj0NvCiQbVUW+4kEn
tdrCjJsWe+aDCaqhcyOwHT3Bn8nI336zh6AxTm1ZgtBHEeKv8Ameks/L5/ZBHnhljX8IsvtggUII
v4p0p5AAiHtlOoMowfiTIgOJg2O9mHVWkR9c2w/HSliuQXJynzA1x1aglvjZ247vFsuyydOs5u3j
NwpAI/QX4US/OgPgYoW4ALeWZDYbvZjfPCM6HOEcCR6k5OdtUNcktMz022WpqynIy5b4SQpjh9ej
ldbLgpqJoo2ufq5tLAsJ64p/Hw+eXcmzA2DH0TNeaOKmZSOnDDkaV6QScymv12kknst13kL5Nxq0
JOIvh+d89P8ebOB8WAChIVAdyPCe4JRoROu884jBSjFC6SjTJIbXboUip9I6Nd8KihNi3ZcirkxH
+EZDFHd/6hvPr7NuCiolwyPSd7qIR69e8BBYIjb85xI0sfmdJFuR+jllYxg2vdEh/aLASXdLhDnc
vX8kk9Hy4bzTrEUY2WJXJPzG/AHLDjkHxYYULA6IY1hSlzC6LAlsfMnYxD202jedVkkzdAbIGEfQ
pzaQuPffvg/vEAersHTjF00xjHAF14N6eplLb0G4dVAS7WVRInTj+1M7GGV5h5AdoSCJ+6oaNNZn
T050exjNDwWkCjrc8FAlNdPUgDmH+NI0K8qc+IantG9IN9O47hmHk4NoHQUz2osv8ZsxviimpcWA
2/6jGHeFGJgaS90jb5b5+i4MiPlV7WX7r3jOvtPeXErE+FP7fSoWs7fyjxQ03iUqSwWBXuDu871S
4tiDO/GXrJR/Kaj8onfy7kw4+5QDb3658iOlY756fcPJWPs6avkNTneg0Iz2ABOP5s6xJcr1o/Ey
kcQRpvK69RDuorAJFdkdKCeFPToNfW6FVIfidKJfElqfq6R6GgLD3+u2vvnHYMu6c5WoFLmSLeZD
C/z4H4PMTFEbkV4s6st3fx7xS44HSrDF9WM6gU1K3Z+DA6Av1AAANf6CgAKTjswb/0zxjcOsTBcY
CIXRY4iIktgWUXcSfpX8W9C74UL1X5Bfp/1YzirbZndUu5V0K6ZNKTPK/dw05mEFAPAVagm4xOdo
S2ZdmszSWRsEbZ3vkON2qK/wPK3ts7RypdTatMQ28gbSQUCQOVd/f4pU1JbrwMXlhyDinnb8+eAX
V06xgv13c6eSCK02jJhO+F6Tl741DlpaGmp8vWMlr5HrxptoI3NlF25H1fHZY4Eqx3XBpafEx3Ov
YomwQP0Rs/LWOF8XX+WhTktXj9j5C4VaR+IYJz/ria5aFtbIjmahjqGHmtIcYlhrCl1iSNsPxTmR
/71qhSwIQ4AJR49a/0mGZTd2lESXWS9UWiuoNMywXO5MRrn0MSly1nANbxT+L7jTJdDNs3fhMUZJ
MGa1IG7ajPbu+8j9+6UZfQCpvog633l7kbaDSdmZqLkmvb1XvL/1PDPzZ/MZeh9ncYitTA+t5X9o
kPalfeluOKqzsFP+ST0ujcQm7vcMz6Zb/QoOVwkIfu4Cya4LqWcY0Y+//BzuXvM4j047M3ASnCbT
ooguwqZ9N3zb/9qlEkSfkNd/7JTGlKC1FjjPguv80BV/rczm+uZlfSnj3VBKa/1Tnp6M2MOgZ6zU
U/VyqZeRdQQF2vl8emvVw2F+kaw3nzAKMVsylcpiG0M+8Yi8YjKNdOpOh3PQ7AQYs64np5DCmsOi
h9LsXMCaVCV/KZc2NHQPb6lhQ9nON4IthA+xBQEcuUN3YcI1X/EI036MIcJchVleti8SnbH4NTXs
PgtCLQzlu6+s2h19Qwb3TVHxkZuuQusIhZnITpmevSfkoBLyyH2gF4wVxyOCj1TPfPN9FCG64fUj
WZIs/mffO07DI/NQLna8sWz0eZ6oWOtLZRnRW6rQ/utMkKG395+wHlcpgHqmjqOraB50zOhoTE9z
hkz1NGU+4aauIuScMGe3WZVfyyPpRRxJ44UG0DOifLAIA43W3u3Vufie/UcoIRlWKw0sNY6T457Y
I14t9LYeXRPAfHgMOa5cCvQpVZhT437j7r1F3Gh1gQtVU+TFejao2muAXFhT0uzTI+5sGqGCfCRL
YO7PWJyTWl9qRrdEvVqAOGQX6gQaeSADRPqojdFqc270KglRBnyBpNZXRByJwsY+aNv7NUvN9CfR
AAKkEsJRKrcODep23WcsjfoX0O7Vkk62H1gHNUe1E7ZdAx6BHNJTMKIeWeBCtxgX136LEShMPC2g
8rxVaVKVKMPbEmKqoVYo+cew6inGZi3QHY904++Gsl6R4zlnNVA+FgLkjgU0OPmHqBbntCYcZuQ/
YCsGxzMpnl9+gvkJ8TASdmKfNCcfCFOyTZK0KUQvUCVz5YB+cDC6tlp8B+SMJGZY+w2ca5LsoQuG
Vg0+zO/Ec5gY6Dqq0a/uIDvOnMRawUByShs/6SKhERuvDdMkUAHbB0gARNHuLly9oUeo2lZZ0VIE
usW1RaEeE7h4f8hmEZL0UPpcKk8+nmlxC5GIeD+dtg6A7tXX5qQ8gSegpegsSKVAQ42nNCzBhSU/
qZHIr0RXe0o5hZroxiGNHDh9u6a+QxWqqHxvkBDhQ1VLFFzWH7eUS44ocbvhSC3mEJ+Irvv76Aj7
xNg89d2+U/H0PX5DQwIkMKFGgHPrP5pLklhF6QY+MSOa19EbScMLnsgadDTMa29Nul9rlxNth4pH
Z74A89WTkbRtIRfUy0PRJ63KD0XgTtoi6J3vYV+uPuxYMe0fx87ICjiulTURwXz5trLm0sjXiXnj
FT2vQKrJ+mjcwNK3xcGvOdah2AcqStJddNFTe4bI2lhysrrEr/yU4ZoE9i3zrQTveLEL10P+/PC3
kIIobuO+0NdSLjm/KglQCWC3Cv8wY8NoVkdncH68OYtHTKxxrNJYD8mqUD0Ms88XxZQwIhNeMPJx
bb0VLcmjHl+7SOag+h6rgSNuSy6VD0BdH3x2x8/qeX6zXfjthwAJM6ds3kjr5lAnqKAlwaYribMn
yLu8f6BUUmwadLRRf5XilRSxGyfEkc8bvMjj2jryYmaVjvEFc2xDGv+qKB8RTkJ7NHSfXfjYDoVz
kleKWzLnHqye6THnLwqUjVDinoJY6ZVBpA3tFaB3eCk3ffQdTIye1mRKKiwnoY3mPtA6ycC+nLAx
dZLHpBzV9RtB8cSWgfojXGw0+yUS+ELIi0aL9A+hAa3YW/QQAc1YKqi1iC3AFHdNjinXWoY0YfoJ
ONEbPG/Bzb6O93rK4+SjaAtg3j9yXDtfMRiEhGKmydwp+JaFmLZPf6UEvi50QlDCjyLXKpQpgW5H
TFhoWe1DgrFBUfFNiXVZIphBb/Fjqc1YJEzsNmG2l6t3g5qtbH8B4uyKmLEjGKNKht2e323ykD2g
y7PAFAG4sFxO+pJ+6piX3CQlRHxQCQ2hRxsYIBlD4dzBlzNomLBj6h7YtVBpIk41DX2J6R0RH887
lC1jui9M5CqjUORUBmvxQYyKu8MNCORsNixTgdGBSE7rFvkXE+6lDwztKCOIJBphfw2VdUPU46az
4J6W86k9Jnf6zFl3hYJC0VRCFEZvWKc43DJXU61q5Dzhu35GUfXyOTx1lf9sPGSaKb61yU9R3dlB
e9ekNwW2fSrZQMyt22wvCB/CV3NfU11q4oSmxsCedGC2Z6FR3eSFDqZOn+YLrSSKsdORTYgTsosD
dSSdRUvPYI4LiimfgHljx0lsw2nB4XWI+5EHE6MfhR+7/+21SP00HXyWZppzWi6JZpfPCbppXKeX
b612QMUxctfMKoe+/ZrSK6AaFXBsXr7/4FwyvRVvkfqO+lXMJMUo5zAQx85pLBDGnKWrLCJWk5Pd
142wk9WaeM1j9zNB0XmY2fuCc8lwhIJ66S4D80PccuPxBgmyN4nJKCZtG5jKDJms1/MDpmPz92GO
AsuvRiAqsEee60wL9ilVnu01Jcs8hvqm0ALt9tsy+nWeePuhQroG29oLUbks70gojB/5UpCACgsY
EXLHYFKkCbyFgD9YiuKOG5/4u8e/Lb4xTZn3BpbKHjza1saGctzj2L1toEg7YdYovE0kDgG2EXGt
oIxKiE0aDGCvnWajs3ZRRoq6k7cGMjroEH2tn3TegF/OVVJm414ZlF/QWW8AIJGGZlYDcdCzim7T
eEdEE95EODLWwlAW7t4qacky1d809CP0DpH15enOBMIi+2vegjLMVnrv+1zW/m/Bv1R3hlng9zLS
TDGHZCPOZJf7g+doHK69fQaIH+5PwwA0r4cPDTf02JLOxlwVCOIWH4fEfq6GOQ7z6ITtCil4mH1S
860ZSvyzMcahN+3NKkvqDerSgcxgjmyuDuPZ2r0nVNPWqOoIV8KyEqBB6fwknEHK2RlpyqJRJbdN
LtMd6nDiLdhbdlkG7q224YlvtY4zSWdTR7dUBB1j33GNcUVFNSF5X1k/sGvUfDCjGCLz6EwbAYWQ
6hXYASmDhSsp7hsZKINoLqJYiXUyuXA+TZ88bg34etbaFiMAZz3xiXJ817NWtH3yM+L3K+JyiAHJ
uMWOXrgEAWnEE4euMD5kYXnWmXo8ESN/ZGUQQuv4t0TtNCWmcF8c9EmvRNxvk6fhsp1IROd9YsIh
mx68/eZYaYIgngG4MEx7gr4ZnBQCgSvb69jZ90BenvY50MO1QTOfUAHdBCzO/zyRblRabTPOCcby
sNXck1PuDmgnPyFWFJ5fDUefwUGe7VHBaawjFMQLwV+WeSBRuTZ4/PPFE89CuEHYph5Q4YGA1yfx
nou73+qFKfoo8j1Re4L9mvVR+5kD0RMnE+1Og+6eozTnQjS5eYOnzX4hdZaNBhpTsmx6fib0clf1
0onFjYDKiYo+b+Fj1Fxiwl2drek/r/+JuLJOZCkn3pyVJ9CzjBA/9quueGAKyj2mTYBW+V6n68bX
FQ8p5L5FDPFG/6VvW24WTf/yjYUsisoPRKWOUrb7EmpjUYD73EeZmZRkKeqn0KWs87q+dDFWOQvg
OSg8DWUl5Mv+aouzuDkaWp0PFLPmVxVK5MrmuWihuew2oAg/rD9i03V4VuBss/Z2ZqGHMdwW45LJ
ALuKdmyjShekmaZE3Kvuc3o70qzbFmpu41jnsgVsFXCrVmu0UFEpEqxD10UqxgGO1dsXzTWOXuDx
nzjO+Qeo3sD4FmwKSKQBWqko1Os1OURCx+0PsdLh1FZ2LXgmXutTxbqZ69rTI7CJGzxsaeIgO7F6
Nol7WeS3uTqZmhRAFZFT1T5vfGYaAyB1bn63og6j//SHBs71MvARO19zALcMvY5oT1o8miV94i5x
0FtfXLl97iZP/vcT2Wm0uryvdDvyJxru3qqFpl2f3Z7s1eh+T5V7Ytpw3RNKvenfJpNBMqwIp2na
GlNHUeZ0hgqAIW39nhj2I0sD13FV0y3NxBI1mZqH0Pdmg0jUwXWJA7zd3AOTFghtFtq49DIzOJC7
98VauAvoBJI0qx2RozDn8uNQeLghwpgIR+YXKb5frZKzL9g3yDThE66Cm+BQKnv2uXSlYYWY/z/C
WC3SN/VoQk/eH1J2aJWKuNH4Ejq6zkpqSWBXs7RX/Gm1iqKmjeXdywU2CeVEY7HirLEUtQRbyNQu
EajG0tuevWFKiBOJ9rpOzGUtOQdBjzhuGEvTTRw2dGrWKbZbuSv6MnF43uNFoakp11Bb0BYEKc3K
cIO/CY7mOnOKxbbU+4z75W/btBkGIlQvaBcth1aAfz/HimPekfPnJlKV11YdWpheYsOJ7j1cI9hF
Mqq1h23TCOZPGlSo7mLVfWhAxK3uSaVFNKYirW2lzpa+1kMdnfBbxMFdejKK0omoi4DXE/6oA3nW
jwgtnLriVr48pFsakDsWGb3vK1cKbbohKz4PWKSUiUD+qlai5YdYIYkcgzvy6WG/2er2l07FlqN3
bqVxr8glAmyi43cvfhF/jV3Zs/0aV2kpnNY4TAisNkGbOyhE+rm7kGtA6q6ZSiNhSDxmmyK4Gvdb
d4xIRCgWpdJQlxHDYSXmwuXkPkdM+ZkJXf0GhlU1MEVAzBANkE20gbGEvZG/gD4LjQUzjwAiK5N3
tXtHdNZ0hJajTlSMRqdoRJ+We1IBUhVPsoOQm5pZK2TehzCoJfwK9OfGFPBrA3VyZoM2JLxW0RW9
aTbZJRQptbJPy1tHpWiBxyQitM3G/ks9gIfTXe71J58xuXXhe1y/H6t653Ha0Hs+dA3VaiI1mjl/
wAmpbjHlZnl9Gan/UwMLFzLPwviV2GZEZms6O2nZanhaL7LlxkV/vVhJhpwLhJ5h9fpEhYCikoX5
ootd+MXFoLdhs+m5GiWlE00hlftg2UOF6wBE1TOZXjewFDVqOHxX+ovDK4UP3LV5cTzB3iIAnztM
teal+O2MWBEkxY2nKeJTlooZtvPFIVZAw7gNIbH0atCMDgpuWVZjZGdwFXEJtu2FlEeyEapulBLu
9xSOFKovj+n3Y+W1vvZCCUIwPw6c4SyzN5LTd9+DHOY2ez8MUmMk/Ts3C/DGQ8pJKNPIdKWFo8BC
v0thP2drwSJ9Y+QuHNLfYLqPM1enpDHpAHjpWFjojzJ6pb3uzAPYYxNSYZC+MgXldir83TWFsd/k
jzrJrH9UF3JUvYwBlisfXX9WvDFpZHx2JJtbzgHa70hxkSLrv6/WapaskppIIq+Cq6RIVlbBAlvQ
Fi7k913tZbJGnY6nQenUtNi/d3fgsHGQnOmjmxEjQDwO825Sidku/HGX7GLNe4REvrszPyTSNwCc
py2F3gHJ1SSzu+rLy4SiVc2ci8pclHwuhy13VB0pIa6beDe1Qu6ka8cEtQFo2mpsusuWGlKphYbJ
8pDTfxeOhH9mdVAonx4151LU0iFiJvUiRQV5JToi2k/bdOwSU0/OrcjZ1fT0xTF35gzBT3IZTyqA
ZOvryFkOWOZd8wKjxgStcILYSbyMMzVPtNq6mBAfN4DusLECXUYVxa9mNPFjG5jLSOaKpG0HbQEs
qotIbszKsxpnGeKa6fBpIsnwn55ck25BN2+hhgfyHR95Du6FHLDVs68pfZj9nhKdWriPbGGQWmuu
nGqe6/ADZrSIxbY8iI+Qfex3Kobu4P8VChmJDa/wL3zy4cqDgfcYpLN5QZ/F29a9pBr6rGBDdYiZ
TJk99NA+dqrsnVgV0Wg9tKekBZyqoBuq0kuooDqJOSPLwtkO76AV8v4XKAMHlomWzkYqlWljUnOs
Q+wAu4wgSvnce6oBhkwdV0pA0L40gI6d8ataJ67MEv7D5TwZu4oDSQkZJIDeRuNLK4sW420/DGbW
8d+6A6F1QzrI6SnUt/YQU8Km53xnQKirTXwRKlqTMxoC1to8seb0mdiASpl4Bz2YaGuWZLYGmzwU
YSDm5bPjoU3QWV0ynbIrZWp9EQe/Xvj5ngJRPNuB3wXmvtMlmyKbnze1KnRJbpN+Pb1iUjAxQEpY
x8jsikmJR65RLdexV6Xr23pfxRRzhk24t8tvGwbrI4OwUQaq/TC15B3/zs/OHL8sWfqEAyAWY3Bl
6wI+Lc+ypCQ+95cFdvp8h6+3NgD1us9ytkkL9OP2zMImOKziX6NfRuJyNzxlEotlqsQG0786jpnq
sBFsnpfSwxjZCZc5wIgWxPsqpOi8Hm0a+IZPWxlCS8ze7tfd98eV3/AqHuHuX1pRA/FFUkKTjDy0
aTfq0gKt28V9PKVLBLC2Z23EsGSwo9QspavPBtq3hbXOAjthHxA9qZmih0lL5mmJj1+SXWb2hDtU
9MFjD5lLo03GqB+z9mITXycr6ffBwbT842pPRGqtCvS1Vpo4dBWQ6glTN7Vf28xZ8bVxYSr7MBhh
HDU4gwbt2C/Bai572+QE2MvGMOxwG2wPuwqWE5diRLroPjh/JVOoRIAgBJp2rida/v4odiyeUVAk
KlQnZKCscmhopC+uU+8JVIhffinG4THQ2VWSkTivfPSh2PGMKmO0I43zXzZyu7ndGP9jKOmFm5dt
CXoTtvUmdazVEcdmL4Lv0pZfABwzuAX3IWoo5BZfK6xABaV8lJavxz3whNKcvYRVJAf/cbiG4vn9
nvOW1moAj76kq0WhTsebxYWhwZ6H+RBXigZzelGdLa81ZdoJkc0rMBmHRRUiWQ7/e9Gj4mjD633q
VTOArzfLlwJzO6smUPI0qJxu67xSgtGlCqfcytN/2uJ6B7cjcmyVaFNPwa6m5wWvm6iyB9xxbU9p
f3wmgrjOinMgrT7kBU0eVLz5bX1n32omXtBBph1nM6G3DGAk9hbsncIJ6/hc5gWnhzZeaEWQ3Znc
FKNWomFeQGS55jwQ6/ay2JKPvcfz0JulHnbBnx1t7fOeJkIVf6eaWp1BJCT53ZeVrY68izueICmZ
9h7XEy9i2uCY94GzEl+XVTQfXj/jKBWmk3AmBUQ3IuXCJkPqaOoyx3kZIVlGezC07OLTrENfbOOe
AqNUsl73NqsZ1scZobfzGom83AW3UBlImejXfVOUnvHNRQ8YKGFMsbuU6VweAArx941TKeVaIwe7
qtYfijJ9JnySbqybeZ+TVpQaXU5SDmXVaQ8tfCBkbiXB4JcIsVVNJm/yE5jeGch79J91/FVPwGc9
awJS1l5R+AWPMoaBU+cergM6U/hg5pG0CjVt6lMuXLGvZFCLdXUEP1Yk3OoIxf30+mjXav+BPa2W
NAgftjzv7w7Q32h0RayINjI1CWWFppR0er+TrusoOfYpYRzQSuKz6NwXgCDRRRDSomu55ev5J/Xd
2LP+che4CCY03R5vRnx03Pv4bDaxIbY1PQQyND/iX4mdpYa86pA2HPJAUAALsNR+kA2+GaboRf9r
keRkizgDd2ETaZi0LtrwxwR9Ru0v2/wUfujpZLjTMMMluD88/SChlFd3pBfvjnB6MWh+Zt6/+zjV
Z+sEesUSnEf5zkx68UQnGMQWtRSK6V0Tt2VddlZ5JdTaj5Yq8SsHLsSXvJRt3eERFWXT/mISUW6w
QlsUYlQEcvz/xEzfJKAk9B3opFwCYEkq5oCaOwYYCvespblJhTo+b/v5rYAgiG6poz9Ir2ZLuTNl
636MDbDkXvRMjEVMt2cdjFnN36xxxMgWi+BgxV3oGEn0iOFbG7ZjN/fZjNpJD+6+w02KpDaQ/Z0y
YapTHOLMLkfsV6Sqb6EcqSb8qHtDWu4jJ+0GBDN+c704zvAGP6H3s6e2VDwM2dyTDDzaL5gO+WMT
YSozUQFN+cpYy8Mnscz9nAJq/JchDRa+wYueQRTdaWZm5r+duxGNfvEFEw+fHhdpsEbtJHdYZxyn
rtn1h9j4Mklzk3eReMIgu/NowDVQaadb/i5wh/VX/+mYcxkD1eGtagkhM1lLGU+ECKUOCWBk4dmb
1SZhD0skSrYdkL3M7tzzEaW4T515NHawU94Y+CLbIM5W8hun3SMQC6bz1XISgvnxnFdE0RfHUGim
2zQ+49AoP3xyUIMiqMvt96r3ICi/8+k+r0jizRRWQOJD6f5iSY3agEIIWQM0Wq07IaZ/B30oWURt
jlGSWRJEABgOpv13XI7HjK2mITOheZMsEupEZNeMSE5ucJTr9UqRXv+lRtz1OQm0LOvUBKwk/5gj
BFCkNmadNjJeLiJ6/wVA6YpxNrZiDkss9cjO8YufwOfKiXxmiotutI1snLSRr/a2O0/+ahWvTPLp
QE01P3XdbTTzMwdnNlyALJZvJwbpr+ZemEA2FiYVCCkzhlQSSRp8S3MR7iB2XUVWTbrIkNVPjzmA
dgcmkAns41JC4ZaqNXikqtdQZ2YT9S6wBIZ/nRqBtfRXb9x/V/63T/IK3uLEcibDhMcX3qMei1HN
13/dB+QoGHTtr0hObpImrIQfgEEVa/n8cPXLFfcSETIXdCXIIKLAjKtQOKuuZjIvVPDCKfYb5mb/
N3gfbORZTgkS0RiYKMjTimfUIWvGkKpnvOOpVtVDz5i5r3cnBBsWvmqe48lHivxkbCOfTFTtWgec
2tTi0SBXqWgix6g6setkrPAKOtTbmvFn2CxlRUBv3S1tTBIrkP6iGt9UFvVHEOyG/j9xfNrn1l0o
V1h81uxXQIFa6TvGwnfgP7TC7GE7DTHTf9UICQGWiiZl/m2ulAki9cjXaTlrEPmzmIJ62BsGguxx
T4dUtmxpLtmZbX91dMuX+KUsVl6PimbH2CwtqFGxeiEdURsnNq07uGpz1hPsNOKwx+0UPtWv0LtO
Kvw4WQNL4dH47fvmFlUBmkfPeY57nkIv11lVm9Pfvwj0ql0LZ3LfQ67qpp0vhRRsYtiJMBsGikpZ
C4SyTj/6GpEsY+ce1xLVSj1POihLOikRpyKvM5/HI55H9RTAVT5vEz975ioABobNCWgAG74jrY9g
6CFXoix/Rrd+sSBrce9BSe/jlG/Z92IcqdLBwkjoIrOShtcJpOqZ1bvncKH2oEnaVPtsc2rLTwMj
BGoMidQAyN9VfM8FeDqHOSblmqF5UyexTtSzDTwfzrPqbyUOHUrrqaX+NU5fJ6n8KgK3sHQw8UF2
TSLZAB1mYDSi+6s2qNqMJRz3cPpKAlf+H/czwaSgRVQSDX1PhVOUC1iQ2INDmOOZX8Sj5YLf8ZS7
jOP2sfXO7SzOyXyHYFzqia9Ydzr2/XsERmD6LZOa6Ncz33bbVs7+JjBOn8f3LCCLxYEwjkCSvdP6
7qj0Q/Ru2B1/AEODW/RlNu7JGZWuQpNkZpqZoF9iNooJW+KlCF4r0y0ttF827HlkxBrw77aQeHTC
QXackD/uZ/LM1zAv356n7KSMY1BIk7S1StNx6GewYblAp33r+KJqp9hdOW1XbczHmP5BeuYqXeKi
SzeNdfdilIMluw1NJnFedFD8jNUtabw9K1XF5mOA+x9YOFLTu9XdDrahm2+XRrSS8dztdUuxXfrb
bINTgqZ9fmzmQ6KroQRmJOqdhHU6RK371cU1j93payKEvX43vaCYJgKBGxxFOGfT4E09UAQmRUq+
WufeM1RhJvGqWjX9ujUbFGH4rL2SYRw08822glFOMGqE7Rmf+GPVk3VXOZ3+5V4IRzuzFLby23Vq
hY6DH9c7bBIUaWEUapCsCGndTTGe5bgDkTeV0BLBQRBRA/qoKYeaGjuyIrVv358Oy16JVrly61ZI
c3GQXKBpFgx7LoKJ368mHlKPLkbjtfz9AFI3E6nq5jVfk1DL8XEJ89WZYkid0W486JMQnn6/hgG3
tIMjZWZABcgGEbra+jgKvAagiVjlj/MnkIZgZEpZGMIZKkbLWjAphEHTITFBYSHfo+4JqQjuVnLm
I8lrQpugDzLHEkkWXo7vQahii8cUheK/znv6/7CbXBEFiRJJ92QTicv57fc5JfKeHGnO/RnalTgI
F9mA5fBjbgG0qoEwr2PH/6y71H1XgmpKz6SWmsZJ5NCFo89tM+/YktOAnCRdpqnF1NU1885mFdlY
17O9E5KCD4ty0cTVQTva/MBETYiFbmoJ1lrQnHJ2ZZf0+3y8iOurgo3Y3Bwqk+6hqvJ26E+RccC3
ONyGAxkIU7aaiH7SHnXztcyvPPxP7QARd5+O0KHfdpAahCGg/Z3PDrWMC5pzElpDKCAHtKrYxeCH
e/jcrHdrrAGrZiDwTK63Jpo6y5eP7SDYa8jPj4RMChd170fZAPNESfKshwDXDIRnTu2yUC/0IK/5
Ep6UUKwccumaSlAGhphLVb+AtalYZWXAq53INsSFuVbMu/2PijAwY6zzaQSeu7vQBl4Q5xzplDFj
mVNY65vcbc2UuMQ5LZwY1PWTBb8nL1wPbS8IhDI7BD24Mg8gAw7NfCI5bl2Ai1LXGMOaxo+4uVZk
92nScrT5cr/baD6TB0Si5X2KAsnP2p/OXUsiiZyGyerNvRQnJl19RxGlMXQMn5Camh/jyc1m9qVK
EtG7rauBb8JIb5/oYV/uGlGajJTY1tVPlO2nMY/hzmhPETYdAJMA/gq8O6WYoT3mXpPiedwuMj/H
CB82w6+qaNpeiCRLXdBdFNj3ngEbKQ+Eu67FUc1Bdm5WRJpyw7bKGhdQM8Frk0QmLgw1fd7dyj45
rOO+mjR+M69/rBd9kgv6pxbWBHmJPnVV6S/YiFIW/ZtwIAsYlD2wBSbh7TQ/EdYowDLskSKT+kaH
DimBiyaExuhz9oyMkOsRq7YGk174WWkJR5i9UrSg8NmkQUdY+0atJ98co4QSC8HzgS1JO+sOCfn9
cOuAbvzCMgeQHUK2FdlBlwCXjoBizdoKj2HaIrL6uKIDJbi26Sw4oseYZfISvXxa3TrF6l49KMZ+
k27fGT4q0pGfpb1LwB+J35GN+QGfXl40pDzgK21Vn72eNqOJZ2xUeaoopnVgdviJ8igGVCYuwtsR
YKAR02TYcjshoXYxVFZDF5zwOXKKBKYLrF5usXsmVjCKKK5B8VNQtDXIydvWZD4UkKxxTIh68c60
VyisdkqATsikjqVEX6TmPC3AzENJMVQZ0eF208nrPmMMVE9avcLmV6QGK3cIOcd40Ses0Nb9NA87
aH+mcpVo3hQbgC7//CojqH2qUHSGk5SWZzKeot7+x1wWenWdAGeMwYpg1KpWr2ivty0XIsq7Mg0L
UCluswSaWwdXPwwSoKfcBiBMVSfzgovJfbzUJqLEFwbJWEBot3Ch37wkorRt2l43+dtICFw7Ej9q
hYtVdtEUY2ytfNGT3HfEe2Wr/ISY3N3cfoTTPKXPhkuTbZgy8K8NySBJ59uU02UeFIxaggKBtvpk
O3xa+ewWdO5WLgXX+WBKNSAgjPYxfA3VYFFst2Ys2e79fLbjEziyPct7Ws/Fo9s/ueuE1HQrZX8O
YC36Fiu27kT4Lnd3qMc+AT/WXouFRGDZwQz3/mr9omqkh6g4++UpFO8UFoTLUNcf6PSG3hLe1w+q
WrW6+XoixPimlAchbvJC7QNu0INs/lf6/xaLgkKCBIpZh5naK9xAOCcfcKG2/LPzCVWKbiZ52BFs
aFjt/pH/ryfes/EE78vWYc5eDW0WxE+2I2GpohrKboWkTxGiNRZ26j1OZ+g4qFG+HQ48ez/2duem
5XQTH5h9+i/B1RaYWjJSSoYC4ooAVqyUHe+NyYdKxv5zkzH7jz8KdoYn5m5U5juYjc+GdVilOGvx
VvzWtPzlG+2egi4XQMBYzUa/id23t1KKTAY20IfcxGGZMAWJMsaMqiuao3ofpzPrylVnck9GlrIA
1Lea8jDDeHNId1xQyQ7T2Kos80vBosg138bUMub/JOf8xRv6DOPoheWPjY77zZlATUHh223Ke/wL
5oTmAlSTthU+1iHkYOoCH/ksHdTBupdYWZQq+98kq7pJTOtnn+XlcL/MAL54U5lh/fOOHRDPdhPm
n/MSUDL7Bo7SdYaNd0NYHEVwCE67u1ka0OGp2kur4ScD4dF92pSzK9TuA74JRd3WY5bgymYxitxD
qdjVOF+Mejr3BoEyoKumf/30yLx0eHY5qRIzUupVflAqhh8249V/JeQosX7JEM2nWb2S15WWRsIM
A1MWHiEFTvDjSM+0MF/70kyDh7oQACWTybfvZ0493JdeHxZSHn10lB2v1j5q0CWSxGIzETMXjKjK
pHGkIUSPpCgiAi1C8yx2/pesKrvPGTk+wXa6dKvnRYcCA8eKnYOpeR7szqn7ULgqu0TdIwkEZvOz
QLyvupFjzGguUbqCeTG06KaMFNBZwAPBb30LyOgrfPb3aW7qxKBgaAkHhnAJayxZaJxAhIjiIUcg
CphzcjV/jwFp28UFL6NQR1mFxUmj96gEtxyjcOLNqd9+KMSaNVOvall1OGUAspwTZUXSzPRq2BB2
WczYAgoNVfzRmPwZGX/CXmwya3LBndbJkV7P4LfjhIHWPJ7pR1dktmrU0j7RWt1p1LUCQpy6zT95
UdbnQ85q3UdKF8RHoYYrZZWpcVGnYlysQS0EGI+JUrrsHkAXpcNXPRGFVyZaFpc9KdKQ3oy3KFr7
pNg5L/ZwMAox9hujNX7izHTxV+Fn0Zvk9M3gCfVlQ73mxoKnAtOco0wYt6o+gHlt8x29XPMp7y6i
ofX3ggiwo7LcRPg1NnhnQssyrmeWVr8AdG1p5R8klqDSw0gIMEgCmoWc7jxlgJmuxf2b6jWNQ97F
ERq40xJ2LMoUjLGBLkd00saVu5jz6RRWtTl84XXLRHfkCA+A4qPLYLQAbMm5x/VQOWM2X3Q2PO2Q
fzPbIZayoDw0c86wrP0QqgHrJb2FW+p0Vf6qkBJy4QkQycinxNQMlHqSj47WqglC3vyBs0xIfh78
m0UZwBj8MD/fdSsqjWeU9hkGcVCTejrtYILjAcF7YRdgSm1uqcg6dzYDm4HHhpXXmbkhtWSJVEmr
i0CX1dSlrdMCAvKOL2yjHSIMEcPP7awYn4IWR1DYugqA+x9O0yNJOrfFpeeg+pMlmox+aAxqT75/
425D9XDrZSaxmcHo4DeMHXQ7JBICSaQaPoSG0tOrtxGJupF/oBcG7zhLIRb7HUwdHc5tWyBF2MdK
90HqCU+N3h7VuXal3TQ01jM35Joel+1hs8kF6E0X2puNkB9XnEynXwRl+Ds+5Y+kZWYxz9qTh/3v
laz4W6sWQBZ5oinbsR3HtxMZa9lggXsVY2J8BEFatoTY4j9JgJfI5EvYM5sk/foK5pWFJ15I+3QY
XXESjguH15uaxBrI50eeZsHSVCn+aLq3obhw/4R9osxi6tCT8leQxfQ3Nbyx9lEFlLaSTOX+QyUn
M4VHbgUlz5LxMi7n9/kAwGhLYgoTL9LypeeqfLFjAeI6u2BIUyEaaG3ie3KBFEyYPH9oNDVyQ32M
8shDu006cuE5TsSuqA2na/HWq+C9JHv9mr4ZB7UXft7mjIjCMeyZG+74HpABm/3p3hfee0zHrz8j
WVsH3WJbAy6gWg9DqX6EoxzRBeKo1JRYtJzOncp4EWQFkhVVN6nIBjl+1zC3bwUxUKma2OKuZgSE
xKQTaupvzLXjO2iB9HlJrqE+vg15CRfh81Tg5adUIMJJZ9RAwRSlkBBfVDc518e6iBQprIWMLDyM
0KPZutBB//TxnzfPV9sFAEXFA3lG1HvJiEpVTAbi9cO7QmLnN6XrbSA1IBH2OBFA9nQZfQyXe9T1
OTHz8UxB+jfiX3S/C6OCxCv5M16Kjsmnl9XtETGprGKA2qN4IraVmUcw56fiz75XCO+xy1vymjwB
qJiLO22m0C4AuHPPBlrypGRDdTZ3cCQc4LG2qmbSFPnYj/tcKyGGTz5nhXLWOhTaawzOXSg7abDQ
XyoyX86tc25AFbM8vI3ohlrSTGQlRcTM0LMRQw2vrrh8YFGDXjKxekafX4JuCAqLIw56w46wFqdv
DtYc9ZXuyT2AH2dA+/sJUAAybrOFzNx2kVVFhlXn5Fckc3JBqPJcSnm6nkOTKEuhi0ipKErmwji/
DTAeNzKQlGWUJK7jOr41qA451JdYjGkQS+w6v8VUg6X5Cq2RmDUlWv5RHuBHLkuJtrToxPNTlS9m
rSlpx5S75CPlDwbRLcy5PcXp6kt2sxymmtfSNVrjUikqkmNEHC6CsNZM24+njs/5IueWVOArIyHc
YQsIy6LeQuoCLgVkixoC/IVAtkOouOiXoX3YqtCguKsLMcQuYAtBUAZy34UTQLkQ8WcNFNu1XTNh
nr1I2HkN66KZ0aLU+e/Yk1BKOsXbYgO0fCh+n7h7DxdvSO3APiJNInTFkPC9aXv3yUZ8uPP5LnIN
AzvysZY7fO3ioqlC78Djr6OMHr3prA66b1yCV+QBSx8npIyAEw5Ybs1FTWBSaDKEC2EcSqa1sbPO
XarV132/XAV8NJUJzH2MGjPSlCMn7m4i1KZMASZVoYevBgQCZfGJ8sEKYQQPmMXbu/BGy60e6LGq
OD0n8GJgEDI928Wspn/qxwChvRwb8oxt6qiM88aqPt3Wgm/Ju1es2wWuIj+cQ1AFDYuQuJqvEnsn
gteyGxc1XwqDFLH3Y7TI+8HQU4R/uLuV3mI0OKokFel8juMOPGRJcHeEWoKZLOk7wV6B02CoL+2M
WerJ2xFEzgko+5eorqbdfN/ZzBE1Qo6jyXEOeQsjZk6LxfB2CDj4so04v2zKPayMVjQcv3398VPj
hQ1C4WMPK2UJex6FhWLTgorjPubWAvQv5zDzXBfC5JqVMuMo2mwr1+kldeXnp0PeAX4po7B/M2vt
GTP0LE0LXrTWa2E3jeiGUHQTYZBTRBXsQEubSMyo1sp9PwsvCUTSP5DSEfXp6FywWOpi/F55WPOw
OLYG8cj2NVm+6ASxc9oshDKNFR79ptSfEtTQApI8AdDEeEbFVFIBkYOB1zis/74X1KZsJaPqy0nP
+Xz66wetRLullDlrAkoQDjFmtnnGMNQ+Kr1ArmdSX6fZpB41XuEwHlIcjt/HjwqGYp8W/fSOoN/A
lKzOJgnygnz1ersNDo3tboQ9LjyziprBglvy07my9+DJt980PuXYhve/9N+N7ba0ErUr/2jgF3tU
QgFFifC9wzg6pAkQA4AWQrAnqi1+qrSEGvq07eBwZwPIlwfClYB79eVpTavDnxkLwfU6+30kSBMJ
KHHWaCXqhpo9KLMIOgwRiRO2V6lgkGPAoMCyfsBexA9CCxwiPKP2ouiVzJHOTZIaMMwTzlJaHSI3
vHLpB1v8xLzmVHNIXWKoUCmak/DpUMvST0HS29bkdO8w01JoNg34qkhFDTUlkRKrY0iLPVLdH3+Q
+VLcEtP8strcoJuaQHcYUc73+uUJhoGnwRXik4JF3Vd4WbuVAlj0fpzsS75PFL/nriw8a7g11Wpq
1Zldprpt76dKoFHevUJ/u/1svcqKWREAk6Znxihy0KOWx7C179BUySBhWF39udHhWqT6gbDWHVFX
YyYTtmhBXL0cKy1/MnEarSHL+5u4MBYhNptmzd6LC+f8r757x5r/fSThfmBowe9IpIQNpSVQayNH
7LcMW/eKjMdV+eR7fzGE6zazJD3ed5PZnPU8d5ZZPJvf7UkS8bYyuWf7OfQ3rPzsyH2hGlHjqMYU
OHGhTXD0Y2JrXTLx4hfofBfkS2APCDj8QYmoiG+sL7O+D7d+rYhCgYm7GVQgZF6vqgch4bU4fFmt
vctyrryX7rVUYfHDRUerVjN5L6SlH2zCKejC1rlMnGQphaX3IEQn0Tli8u52hPpTlGy47nsBLc9l
B96Pckg4x2dnhJnRklbhO9PToLsbAqwiBjAy1MpniogWvblJXbnANuFQ8zgl9idUqjIBItMpUYk0
fvh0K0GE8ficvJbgn5siWqdd6xVU3acoHyAmrnz61PMpnk6Hao6VKqtp3vWqfOE49Gd4DATmYF1w
WIUprPxR+MWkHM1wP15udz1qDF2WGZ0fVbV4YtNEBCYps+sWfv0eIoaGZsvrtvA3tWDjoZfV9GyI
1i7jwwvbZw4XEc9HlP0qZPBbMp/JmFGAeCTsS7ETQQVzo69QjcZcOsqGuf2oNgc0kqARv2xSgl3p
KUaP7wQOlnuvNktHi//0FroubPFPhUJI2NJSoO9rdJ/U2bXYoslra6cIuNIfa2h3m3mTqzWfbbu2
eOAuWW5lvbuT36XRVINHaLo4QHIDdOu5dhrwZ1bMYIOBLNLpQfPkm/Tn+13noNoGBwbFxPqK+Ocf
o1uC4KAfNpBc6WuzkasuMxMp9kcDzsp2xL7hbk0vwBHoDtY6f0DgsmWZr3kToizWsDSeSuVxu1gu
h7N8narbIiezb3uKDFdfW+Pl84XC62u0mxTeYRxOcuoPZQ3o+sMjEFtCSGQlF1vJtR7myubw1TCY
wGEExU+CauMJhy4TmnQvegWXsUvj3N8EtVsIUjaNoCj4737m63zEUsUe8Oyxn17qRHu0y6xScXDf
lh91OgUvBw1KluRpIiljBiRtkolxR5n+GA8+MkbRHrz20bhs6ocAJfPUzdM0z2EjHDlrkPcftJr3
T2RmRVtKilK/0RX8yJ+TVNJvpxylr1uBQEz5udzMkhiZjnR/gNC66KD0z4gtxw6bwGfr2HBflyEI
+v5CHpYDRgFg9hwLDcTaIidCfj6SPzq1V0sfwlYqSTJhF8//l7bLO6oLgUiNbpTJZKxDsyNuzDxi
n9+TgDrLsRKb722ZODM+jjyehtyPm453kbzB9m/xGbodUVgZGCwBG9+femX92hALQzzTy3aThTRp
u6NFE3FCGS+C+ZHQ5X5kxWU/7L8pFrvNLDKVi2aBrQ+WYJDz7cwwXZUWnF0lQ/u7Ks8Ni2MJCUDg
4B4dtVLT3J6H+kwXS8PqOu37+7f+6rwmTBBozqmsce/AWEJB1PbokMC9lfsy6SUv+5A9KBXONehh
fWrarn2NZxdvl2mp5pHoVYD/hXhBV8M7+IggbxMzxiKggd0oF6sX2xFmpHZgWhyDLxzLRrqBZ7e3
54dh7lgj4wDGej9kwK/4okelIf2nTT1UdsnRkcppZzS5d+4KAXhYis7c1bKpMj+P2qjnA6d3/7X/
JCFdzQkoCcsuROyGZTLp3/EbO/tp/LvFZ6KTxqbqP6hpG5wkxhKlRq2KYHOajYrRcBCiPqAnTi0z
2yw+TiFNbHA/mDPGbeusE9vbG+ugUE771OQIYLUD/ECvrR/fFZ4TnCfxNCwZV694hqN4lotIbZCZ
Lcli5F6oDnpSVn3R1QuLWdm/6ZuwHSLtJkPCFF9VQdfzAVDnwV6y6eUIRfOuUbVwT0ndlYZlExEz
kdFSfx0s0kAvYjH7rdkmAu+BuZeAU1bGGTp0XMhz0Y2szAZJwGMze/m6GgtqIyf7shyvUH2X/8eX
u8dPbL6bCOqYbsVZ7/gAKZQmxP4O0XKyejjnjtC2wwFj9wO4bJcdiefbiMVbyDdh0PpLacIHp2D8
G7jskO/5xggxeNWbzMHhOHNs8VbQPqqH2o+x6CkyWFOc0tlZUxjAx5cfSeSV3MrpJub8FYezICT7
FXS2miGPVvRgWf58KBsaMSLhzs7XUYzMG59abr76YBbqhHOA0iB5o2F5wZf6VL1dAGdtEcpnHFsL
EbdkYINXSB06X7z19uOZLVX3aYjOw8pEuMTuAvFZvXQPnPkMParjMmqrtKspOFuveyYz8ldIwEfo
NPD7tL9x8CBQkgTgGCC6YIXsivkSb3p5BgnHaP9AXC/IW+aX6IubS4X1ivbbjatdTkNS+9d1dgqz
nQa8NS7vro0oZT6qnYLAW76hKNJP+wINoIZ9Sr4sj/ztkNgJFEKEUUpiycBPbe1JFtoMSKHxGQHv
vOFnRYI6hCQJZzGdwQXXJaQP4z28mBM1H4fRDm2pKRO8r+GPeEkNTVvjnzDixcMQuoPEgspspSyq
Qa+KBloOwvJlktL85GRtYK7eqW5jxaB582RWIyVdTv1tgvVX6G/2VyIsxJPbzysvC4+CTV3cuMrX
vTufKAAUglgThEISAtSXAIXeAjsCTy6wjH2sHIr7MhcXYkUNK5mrdFZ1IzPaQtyIO3509JYzie9B
ZAP8lueGudbfgGRCQjpftmQGajBNVO1Wnmkfh5VihqV9gB8fM/arKEB2d3v0oAvwhXJAp0q7P4Z5
wrELUsw7pjdAcY3XTqXG2uTQ5OBgBqzQCFAtKLHf0WGk7Bnxql5oh+VZoU/8suEJTMTgWQi4c1+V
FKPyjoeOyRJgs6XX6W2uMkN1/COfhvP4IIbglNKO3R6K/OxvwA+CqC8a/qLFrZcXUfGJEpxi7CHN
I+6hmIBar1/iq4QrlC6ep/okqFesFQgbqFQAJr5NxwBP5yekhPNzoGO57jrxvFXTx0bizJUoZiwB
0U7HwgGcJ1Xb5Ts46H5nKe28bfXTUIVLBocN13dOWdyPE8AQYW4bbumpc5yRNpliRzktLI1YLPk0
B/cDfAZaIJJQbfE3BQ+jbuQzJFGXzs4SiSb1Vt6v8KR+FSLcXcLhKUxvDjkYyvhrVNBNycfRNb+c
+oq7jCU8FZRUUEgSzFcDmXbz6nE6DsN0gtRurL8ybxSbhv+K1+l0oMZb23hRFPAeJ4ID48td42zc
gmsJpwAWwusW+WmPTOixFaFB4gKY8zmn/K94qk5rHEIZmuyKRf5c8cwJTasgnc9Bxq4vYCTf0wOQ
vQjvrx11KDabxrG796kaTA7FZ5tt3iXyuIgOzLbxmFggxdhxQenDd+9YDh/sKtzqF0Sp3KYFNfuZ
wO5ThPhPtQcvTPxfzKzdjW5PNUqFQgK189PcRHqvMjHECuIDwgoTA6GD9Mf6tvm7hNLEj9ngkK/c
68jUD0UJtkPJvvFFLGUf+nUweypyGp+ln9oTj/1RpGF10ZW9iTvIbbgQxy79WeVg2l3U2pPKCECQ
5nIPnXx/cTPYTFSECpj2EOboWSPlKlhEAP8usdYY9qQ8VzgwpsK2zOvaMfKs9sLuwNX00LKpAdYn
jSImfxuC9aN+JoP9s5uQ6OEwYx1nyDPrZOPvNU8AgBvNyu69FUSHsSOAkX10ZYnzPssDBlGmr1LP
nFGJJLawZC+zpHoqpHD5UqItFpO8M1lc/g5xUcBSTv+ifOJUKDRUmxVREt89Cvg3HrlC+0EyA09r
/oWGkF2tYOxTlR1tNkstTbN32pRlVtQhc57vtbiUYowH2mnv5zZl6oTNgiUUdWftVt/uRor+WGz9
EdS0rMy52QpQrlINo/yF+4dS52m4mDg+CGYwTliDXikHu+FrDvMtGx9ydE7Km5ydW0/2J0Meu6h7
Bt3rdaANxbyLGpyRDVN0nkM/o25kDuoPcOLjIgnqOgVYv4+PmSxkbpUwYsHpPIfXYsBn+uosSnmr
o3hRQEaxnvqRAL30JFbY7Jtk5q51cRTHRIR32rq683PAbjeb8eGRkhTCDebco7RFybyyjAAD4pXj
pWnazsvEF806o8XCPsQ+ClmiSkLzbWpu5zwU9dH87Zmix5A8kfBdDRLDhskM97PXvVxJ6C42kw6v
UsgLu8ErwXTmcFxwvlGsmFqLKSEtsePVa7HV0fQ4FPG19ebEEKHd3agdp4H2fRd/lyAdozCRssGp
Q3DuX0S3avTLngo0KHh+OZN58bRV6EcMFd7XOF36k4tZuhd7+q2331OSSb7dxQFODroRoE8a5xg+
eNUzB8SZ96Pz9FZ2TurZqlgQfz98Cg7bileRMByYYxCLGFzVft7JaCkkijImr3t+TDQcvbmlOzNf
asPKfqcHWovPfmIsKrLP6/lGYqFdy0tR8IWkfe3fD4cWU1DnxJC9PsqfJVunsoojVuSqxvmrAGoN
Gv2Un3rhr5UVxuFfF4zNzTenFIEUPP5J6kC1SkdIuj2W/cHPmn3DkjOn+FgnQ3YEFGqYkH8mgpE6
hZWfvI+5gpHDc4C2Ur+4r5XG8Fai2D4BKwIpz8ewQGJ8D/fd/pjr+DrXWeBZQRBfnJAkCbOJjhDh
nZ3FQvkMIFD9yLS8G7DLJng1U6hdDqZ826/ICBEWuTt6NWnNjH3kyQUhli8vfgZIFuw2B1HAuTZV
3Z/QldJ/Z9InmzkmJ3NftfQznoU9L8YXda9q2SE0nndlQsuHF9AmkvZTlLza/qiX2CZZJxPBrJ8S
D5C4sryKv9U6tOk+jqooa95OTQBYvFxk8moW7yoy3g82pthIvI0+DqHKz/xsweKhH4Okn3zvrI68
DaqrtgEb7cQ+/Kmof4C7bLwTH5cInCnU+olQxoYs0N/PEVxi74fGuvO0sDl6QDVtYgQ04CdPXgFC
jz/9oVvZ0VyQQFYxtgrsoG03VwbdH96972mn90TFNqb2jOaMSqniW75oYX9PwgxnDEQupT5HOH5M
YeOmT4/NvlFQEkS9lOoHudCKXcFGw+/wLW/VAp7ozwG0oX3+qYCnO9uCx9E4IqAUYz4QAMdWoph5
KzQ+t378dGofWSiDCMdLSR6AZjOtHpWjyouDn/tAX6qSKuuxgrZEs+LI8RD5FpBLvQZdvJn0eR7K
yuXyUS3YcxbsUt/0PydgqWGwz8iN1X5btCdYI5FUPWiEgrIPDETm6mCj/ns5GIJbrrNtusatrrZZ
+gZwbC6CYMyByYWyEH6z6EfHsEzoFlIr4vfuVuEmn6c4TYq3exZ1yNzDKcgk5spwXoH5md6o8k7R
GDze5x/DiWMgQ3PQiH787Rd1088X741jjlx8fXygtedhuW1+PaY32yJFIslpR1UpTYuYOX9fr0NJ
EAyuE6mk/ZhRc5kn9/KDAUMV5LKdvVJlNK+49Vcm7nfOu0508u7m/N4CoLQXyKWoMYvuvEqlfmta
9hwzyUko7vwaJG+VctbN4NeeTkugFSjYmAwukb7vnH7niUDGL0RkbKgX0f7G/sR6svulFHFWfNeE
Qpb/UYICu4i9iZDsogZGWq2TdgIHybzPQA0971pL2WgNx8ChgUyWZfwzKVedNBBNWLPS2sUumTGv
LrEnNTOWuyzyfschFRXIVCsKc5V3lABZlTVq81v5KiSyDY7xgTF+XsUIHJkD4dAP3k7UX9P7z42Z
xSdApNKuR63MxVUi6Hktxy9lyKzSszjcz+/e86IgabIAqBprGaRymsAqr72rdp6b0qrqVvCK3BHz
TVXOZNstxw7HPQP3AvwOT0Z2qrE2/9KhT8W3H0g+3jacj3bV2WeZaviJgTddPnfWuenS/wKoFi+D
/yWWvzn2RVjjBdZIoKRGrNqiZQgBbRNvb10XN7mWCY3/QiCyul2YxyXe3/2sSkOxQPdw2sucGDIj
hYZcvyhApLXvwHNeW5GLNef563QcJjbi8fyk+ywbL5inNKvirFrmwMk9Z5bQ4shASyue9H18K3U1
hzdK2IDGZcrUOX9vdmMG0COQEX3ZqFeAobyAxOQZdWda2VnNdYNwhH1mlvkFareQIkQXsowkmb3Y
WC++yPbeu70KCKpFXn2p0fU1lDYJG+6NDU9kEpIK2dhIYH2yoqXuo2mP4ReBgPOmIgrbdBpgsSGI
+zrAPo3ZpMV9Lx3e63Fx/ltjNa8bQYQOsZ/JQHoK839c8j36xHJ8ynJjRT35j4xHwG4PnB4vxoyX
jmBjQ7hjOFbEF0HiF2WlWz70pueFe6mEKQ0Jh3tkBbVc06yDVdxCtelcqHbK9MkpHJWADOJTLmUL
uJBJ9RV8+NPXLKsfMvc7vdKHezp+6CHscghAnY1oirK7ZZyYZ7oohBkIWUp4NCLtwJffasbrLMrb
AyTfKfo06XiFOgogOglOCEQDN2lIl9JUC8japuxah5+G4AIHSUif5y3Fk1c1Abis6A92R3imBl0M
+EZVrlNR9KoRnooduw+39+51Dd4xeQ6S5a+5kc22/ZPess8jg0dQG0my2yVlmx7Wh845bP5RLlN5
ZH0F7w9HnCfmOmRfGCI9a3ubzx3DhRMCZ5HunX7zDdDqu1YaIy2T5dA8lId5fM01uVdufnQgn40J
UEtUpOpW3zio02PwnsbUqTP0s683FHk8LAFiSdi8Ip6vTevfMKKmbc3jShqnoa9YJfWMUtMTY6cd
wfBhijjcfS4G/0HJDi2Uj1VFH6cuWCly3l+z0LlXRtmTZ8eaqUZoqh76McpME7WO2TNh368Y3eL0
0O0IXt0t/JuFnyrk+X/95mI6OQDg/CwHKXb6tH3q1RPJKfHEkrSVECaC+aZUJkd2RLqOshClaEQw
o6suq12Zf6bUB8CNHzHTyetvsOSKkP8xORoVXRm+aIZ7zMLpi3YmhiMsoEfse5yDFoq6QXzYI1ha
4dR9XWfYhUQ4cvEnIRdnoWSj2w9l2w3wHu8QirhiZ0Q4sb4zkEjhh2Vvyl0XC3Avg7kz/07b5nS3
eP3pWwuw+ROeCIKYk5mVvfeUq+5sah8zUDRYOrwfeoVX6PtQLnM4f6dkDOOLeLtDzAJzuXxvfBLF
eZccWLRV6aMgXeCBkKSQyxvWZlBsXPmJ/SXJz4R6A8tKjWAen1Hsqn3Dakt6wFeQASMb4Pw1aOb4
BLInOjU19JszHwN9Wnkgur1IPqrREGzpuOfEOsCDX/qvx7c+qJ+mh354c8N0aR20Ll5MngSEn1c9
vduSzdQJd0xnCec278+2paLnGX0YJHVJOvwG7BIzIY5xs/x99y2d58jIttFCX/vUyoP+4ywSC8Oe
oXiqpgGBSMFIc2EG2ciI4tu0e/kkkI+Dq0deeDCIjCPnDpGSk8pKbH/2dM7I4V5bCVSWfKCowCWT
lKQIOe7fnZUR0a3DR0GW8xZbGhD6RJTYO7KwvAn0wJFSduA2dJncQDzXYhJsLizPx8Gj3UnqWLYr
XV1MnZB31I5EnHEA5Nm1eOv3KemLzFGmANml8YAH2kHZ5k/JhurqwK3QDlBtjzNqqMwsn0NsEIWS
okD0JfU7cGb8LNwPxjG1RpdpREmuLi4FhPciQqv6WXs/SVQd5Pg5Bto5DZr+eDcecgatgVbISRmV
4lS//s/hcWJC9oKS73FBRiZ8PCuStVI9bMDIlNCrRfVKeN+3DfHvImpLdkNKCqXDuERVqr+2rkxW
dqttFgCb+Tz8eUeCTbMWasVpLT5eDTGUAdlM+iOQMwqkXyR7QgtgUVbO2O8gUgMrLT1R8+KTyy9u
57W+/Lc8G16QvxQ32tTdAG5tauWcX/1qUX8kQ6KTdCF+0ctpazlbCdZpRWUXKqXG9AbS83ktPdvk
KohfWSllFojlT4bxy0Ue0CB2IChlMBbuKpKy12g4as/u+h9NIzUdeIyhShUVriAzLsVrngb9MGLU
MEsTsKG81xOg582+CxlQAtEtYPOTTsKh1maQysRO80sfJcXBr6kNKhfglz6GW54p/xMcPzq80S5y
91Yun7RODQQ/77PCvTQCUyT//faTgGpjcHh8HOLmv49lVICqE9FdyJZi5idiTdtuIlzZ+O/jP+mD
IWjc9DQ+2X5u9ZVOXi6UwQXoEtV31xXs5WFUOEUvTwOc8/iH8dfH9638s/N2AhWBWLf4BwlKQkaL
0B/TB2IcTNWgbAD3YyYM5/tLjpfwIIqULpHY/xtIU02xyOt9yE1Z4TFCDrOIDU1O/gDGa/ooJTnu
sVt94s5mdC/BX4pqdJjuoYaRTc+qlcPivpdU0SWS/OLFfgcpRTuQ6x1yrTLJdPCvhcaEh3fyndH/
HpdulbvIXz3JI5RPMJ/silpYcodDVZba8sot5QKhdaof9ypuji9QJ2RGXR5RQatxK0HufBXjLEuX
WVsiq6LjirPfdpmCfLg17KHHfPJ2qKPb3Ymj4HBaJcQZS1Ai2ysoVs9SmPMeXNBYLj3a4AR6m1yc
4rXIyeZRRalQsgW+HlRhUT8knXQvL5qfgR1oxmV7TYUqU8cAGK7e/yVKyYlpJs+xJU5SDPxutwI8
GEzCAIXpdxZqI+okVPVcjhq5SP9vG1gVrE0syxW5Xl0Vqtil8sWC815t5fJnwaufdeDPNuFcUoGE
g10Xz2vGS131H92O+yC8mecLKF/NAgtSZhMclZPt0uRC6ofLHUzm2vF+JajEHuVbkWrC9FWphERc
EBnxZ8XHRbWn6gj3W0uc8U329+j6a2ec1Gdx/BaUPmjk5PG5QLvrsjQM4DbGAaMBkvguD3k6jHuS
A9QlS65l8N7hUpkkDLRqXCBKsE2V1MHhvIB1T1YBYjcG5scPyJwGb/PBUE+eVJ8HzGEW8qmZGy/m
yMdxrvbvu354L6f00CiYEcY1NxkowIOjmJRC314VCEVW+o17gIj9gTJ6vDeW8+PLNBvWLGcqJpj2
TH+DObvtbaY8poTZR5wbxSFNKasFLiPh3lhy/7Zv4Gbj9ieVMew2M3k1T92v5iAG5pOylmKxg22X
rJoq2XbThZxbW84kXe+qcPTqWP3Ld1w4M+Qb8507UC64Ro0GTFR7bZNBsZrQHcGaj8Fvnz/MFqww
1yGQyN+PQe4qR7CWhhg9fYyyWHNvi8elEGnCGKhQHrZASQ+tYyVGJF6T1/uoBFLfNmSrqq7NSbmq
EiYm5XIve0Ux24q9T3WmWZ/rNJOceUgZmoJM87dSgm+lGA3JQBVLAxYtLCsy+1IGL3ASkdpEOQHm
Gy2z49FHgLMqJWrCVU2p+/1MtZtTMat9RNL/jTQU97Bd4T9C0OpL3lWN7Jh3sVU0yE5/wvMMH80y
ZhBr1AfFunIyzRAy3u0ZNOXhrdGKj//bbq3SDZd5tkkDGCpWizyfAhqKRvll5dNua8KQ7bfXbZrT
msNRkgHi17bBEOyucrkWOasp/VqY201U3TJfHhAEo7LvF1PwbftgvUraWUqeHReKqsHED9liGXAg
OLtzUyAm2jsbJiYVgyIc/04K6Zekur1lY04ECwwPbgMC2rp1BEo6VmYtZfMsNrT4ijYofV+PlSt7
Am+CrzQoGLHrlAWOuMohlrGDNj4U5lMwPVqKKetAL/B9t2Xlepw4vzEjXRvZI7Ux7ZI5ennO4Sb8
9dwAbvTfWOGg3/bD5XtQ8mmJKEcbSgmCcOEY4dFjaW16z4pYA9fLMgeWXFnWccKEA5j+vVSU88aR
EQLKJ8it8a7Oegd/1OfjLY0ZBwvRBzcpPIOSozEUkuHXIJZrhM2OUQdRUm3AJC628Y6sUgCHzqaZ
LlfIdR1UniGY3kialqV5eRHe1RzoV45WwKy9uXlOk3DGyzdvrE4VX/rIg6T0V+MCfm25M9C/FKhx
aRh9K11ef5b0RCheZ/Xxdqpcynd/9C2IqcNe94JBtD/+zNB8SC6gbNksw9mwFs4SH4f6vGTAnL0H
8vLvVSxnlwZ/+XZvQTOdUDU6V4ga0rxT6IfXaxZE4zCOK4V9Ggi+BGrJdte7Xyi3L5Opht8nGggO
/slzmOdlX3lyb+SAPi+CzIk6R/qPVzDaWZIvWYUWVfVjTDPRh94OyxRrMMKeP/Ufr8JwoPBUUrdm
H0sLPW/orIcX6F4eWaPV8F4NqCkW+QvumkadgYKiqdSu/odbnuU+oR5qRTOYcL/2KXSvDDXFImFZ
2NbXnvokByeijpAdsRThxYWgwjaoXez1T7p0ntawmlyJpBNHNGGH70ZKZYnPYPufSGwNutMv6Dz9
krvwoElhoCeOEzI84rrZRONZN1d8AQ2MklIB103E0oxoA7GA80nGEEVCyOLkhTDVuDZPtnToiRho
dMyvKulLQ+0KXO6SvMHjAZ/OOP3SD/qq+PFww0Shtmr/chXoiG/lAhJDCUi+RazeqlzRsy6RtsZm
0J6uR2nJ3C+yTmhUzUHut5OH7wFQ8KzjAYmFbcuodKNiYFjCt2C4hA56LcJYRmT8eKOqJx8wn6IB
Xk75nZVn0Qsm2tW8gi0EmfVMc4uPVT6rnp/bE1VJf6DiQ6G38aC4whj3HVeFhTaZyNJHYh/JGXcM
/074pAimlis8lc8udnpW+dBd9kiZnWfPRDP//doFyP2LG8q7YouHY7II1N3M7pTNh5aMhUYH3jvP
2E/8F2e9P1tkgkbL13mo0BCQTBGef/WxyDEPuBFQUH5rBcYA0todb+ZsVuGoBUOS/0A5nPuQOzsf
VTVNh+2JTX4ZjpI9i0tKbIoghOACq0kFly1yJhX+zj8DEBnvPI8AtZF+2tORsacH7XHEcXZKuqCZ
w2Y5HGAuK53YVkmj5mhQOMy5DA8Iou17+kON7jY2LbHGs6XcTg7/LHynhmWUYKtgnqlgS58HROeI
3DQmJ9JFQ1Wj6WqHlNI85DUbaWpqoyBdJuQ2Jmq7n8GsrPLkKH1tQg6/AEkaqJxeyYc/4wC+Th1/
LhubUEm8v2c0TOBD9wN8OgTg6IFgTthgW2DK5JWQPlJqB9ScjaMnFyC8FPNHiR9Go0gD1fHh7fR9
EbSuS60zap/8ldQCZigwAL+Cu5MtstOwHpoMsgoeWCK20BMPMx0eCLdwspXwNzruzKd17C1woDqo
CBft4O+BhqABwdIK3KUTL7Lg2hCKbanhD+W933zVAlPS4IXc41xU5L9auRd+2WVWzWkAcuUyn9xp
PN2Dl5yEXyxKMyf7ddQPHVCxxhJptj92qivo0MCWk4OI8hoYrkI36QLZUAbvQEw0ssRkSx3l4urV
7F3S4FYPr45LUgzBOEZKKhxJ3aJN9YsFCuy75JeRjx6N0ErTOvuGQ5+Q7q54v7EZjLveyDP1xJVn
Ez8+d5OJXpZsK9d7r1WyBF6s7RuX8LLn0PCcTWB57EW9XSmssk3l7IIvz8Lz3fvLfDPzhYGKKl0E
o0LGdyPUZbjhy1GwvlGwRe6AAC+Ne89iiysacviSyCxrcaBPYpzfwBx/ALTJJuFSTl2sfWmoHN1C
Tq/s9SpAG7i5EhfJl0pHTn22nfVcEYhINKvgHEBt7T3S7T5pAlHymlCc/VaY37ZsSvaVvsFjPAEj
16ohNoDumFW6wy2XmwDMpbciI3iKyCTJPgIlm4nw+j/7dFo79ep8ZJeYdCAcXzvA8WOc3nMGc5Vp
XZVWls5sU3h3DT1swlu4va+P3OHf4jypsChIhOyJejHC7PTkE8rZXjih/prdX1Opc2QFwd27/1EG
dGRUbvK706zsiR0AoFRckXWsvDFeyJDzkG4/XbiwdjMTU2AUnq2Ujc9k9ScEgxsBUFh/cbv9fVhV
PT4a8BGp9Ad2M6ivK+BVLy9HM6Y6dRfyxy2v+EVtlWRFtUajQU/b5LzKP/ME2EJed+ux5xyMD82c
hycksTjtmsIFzDgZe9OAryorx6Wsfh1F97GJRGvmxpEnjpFqpYEQBbnIeXA0NYJE5Vz5Ks207lff
tVZ0LFJFOEWDx677uDLFyFSQUrbhWkpeyknIBfxZvKwD7RsmKMZDeshsXLjtdfvy2WE2YTyML2WV
Iy2BBDnB3C7mZWV9PZBF7yjX8mxCqe5mwVfi3866LMIHx4BikXW0km9rr4awIkqTXIV9iXWiTyap
IfNZccIRyIp2jeJtYMVEyJ6XDaxW9/9VOfKXQIWUmbgNgL38sukrzLPGeQXXrRFNmBMXy4ADrY/L
DePtSDi0cOlCr1FcKAG7YgVjCHtoNGXLKtIzIDwkteDKfiL4YBqMAlglqOG2Yy5Gv1oxKU1KXxn8
7D+KRsv6eaK5S6eMfaCnkyrh1aDVJgcMy7XDBXQauZZ2Og6rhzWOtRNgMbfUGJYsyYpcJrvcZdXz
NBEKklhiFsj9F+sd2fL8OhlAA2t9C+Zyy2jEBmvkZRIEuNmfR7Twli+dH1GI4lyuTRzlHO42w5SK
c+CtxD9mqTy4Tvp32JOz3fxQvsKkT28YmSz/4q2ZPMh3vdMB8RwYoT2373FS2RYEo/L73BQwfrT5
pAnYVsvF1KB+uj6RGmeBGBfRK2pOql6DgEg1u1PhnEJvXSvd3ceykvuNn0uQbDFrxPu6VFzQ08ah
qxnJ15k25xV8MSaStd4Nd0gm4xMZCiVuzvJSJ9tKsMvwhwQvGuyuZ8418jqoSHOv0pio6QjELmQX
4nKDGAtOuTQIbF3FyuBf4G1jflJGQxxLn3PR4uJEzJ8BBs2Ov0n6p1uFCkwn4qWctpNntu1q6CE9
A9M/VN9GlsfuII5DooOWXjAhvEWdGMMEwc2a27W7zRwroeDnzUaz10BSjG9kieV7q2Am68NBwUNc
5kd5dP0BAQbpzIGJvWUpHaLS90YzapEYcs3lrDq2gs9fbay1ZuZN+ghMpxVlONG2XGJPEQ7xB4vA
bgP0e7eHXAGvPfZ++tp5QxptAvQEkO3wArkIp9y2jwE+37j6gycxjsxh4/wj9dSQzar995Yih45R
AdsYtD/075chuQ8+v2uih7Ni5vnyDBRpqpJ4JyuY7c5IXICo5fPEfSnSMliSqEYCGNHPIhXmpqLL
F5uRL6cXVlx7sU9ddUcuwJVOGCTAAeu2Grn8oxE0AemAxLoZJZGFTr3PQDpROmiV52EoIJe95GpN
KohYAE73Fuun2CzNBU6/nEpTV9qHt6/ky5zmk6jZ7T24d4IWi7KY/sfZ+beXLbOT1+/vsReWrErS
YLlObEP+keLPlsjRI9ZXcQ9BNAiWJC2EYHcJTlortDBCzFdVYIkeipEFHjsG568rxtjvko9JmFNY
xVWn4aABjJwFBCroAjD9dH/QL5/pnQxZlR7bow1NCHufaWMbK02rKw/51nR9OtXhvYCbj0j1ZuCV
qflIKa0vNA1wg1FIqXJMhSdXehOFeF4TPK2DzcP+uOGQFkge8Bx/PqSBKufX0CBZYxIJVOQul+Wl
njX+XdMFM3l9qhe5zLYINcFtaMbKz840OF1pMPKmnb+r8tArDS1xvbpQo3S85Ba4p2TLPBI00vy9
r4/wowW19ihCTlpZnem/0Q0x+1QrdfrOvMNF43hdDOZpHKVW40PzhwlITvVlrE5qsY9umoV+Eeb5
i/CPbCBz+uTDkydYy2/BbRw+alXP/gpVKD+0n1ytHsD+mClcQFa93tYsXnT0a8K2iyRA8CQNJCU0
6dfYBj59jt5J3tQmsSkOhcBh6XwfWg3TV2gzFvmYB9wGFZJt6m7T9pqRLGY59HD4mg106CpLVV9l
5b652+I03J0KhqiS74xOvEm1Rg/tCi8a3o9/UY+mWpSd8y1SmNPNB9ADA7z/mt6ELEuYkvsWkaEI
KpNxM2/F0ZblFgSyACsUBJ2RrryEIzu3CIX+mQ0rCUekMHq0nUzEWqtxLj/sA9eBc3W3OoNZA74k
x+Czn1u1A6ThiCA5tzNhwjKD0AGafMcORa0tAAZS0u8xRuv2iM36QLnE9bgfniBVW6aG2obDQQB7
gVgXRcLS+iCI7OELQlB4oWi3dBLfFRP0LnRFQ45baKsz4kmFDdS2jJXNOvsxSwGwu07e0tawYfYh
jO3RpnoUPmZP+wiFLACfVLnCp030tYI18yYNqDfnkEbSiWL285XAM58QPFEf+96LLy9qNfONfxLO
2PuULyk496oEP3EoOW35W6p+BQ7I9h4IEqXZ1yPaR97TWbtzl355VBh/GUt4TMqL7SRv5UL2ytNe
eY3mv2XzIOcQjLWkwkE5Wv/Ol/ZJfULfMgGKhfzHrM/ATlJqatMEaWIB6GnZ2kMOzdOHcEWC6vL7
hk+Eutm4TiHl7PYkBTvn2ubEQhWhyjzK8ilJHQzlx1PIyZiuEfz8DiqL+SYOqvgO3c0c46ikthlD
AzaaQBRBwgBFrTXaGA/4nbTkHPB6okpD6nr3jPKOdPq1B7JiXseZdh0T/NGc8EXdMSo4FDLn4Qzh
Shru4RO9AjFIKYDT9IaJYPl/LUIZZ8A2CY7OntwDAip7fj/F7rZVmL7TPI0+9ZnWQEYi/ez4sbsN
P0llpUiwcZVn7XpUkveiMIj7gY2DK41NQ55p7UswxmmosRoG2vHFmxKwT12gAcsdw7ZMKQ75+rfN
OsDX95qCVRdDhkaHfhA/EXSM0D7j1UZCJEtGjzICWsSzcPV1A6Ydf5Qsw2BFY3NVed3lYl5D1a79
xtCuFqJt5HExUKldIo5ux9hNkShFfdlwMIAvGJQdLYIbUjGvbbrUIl+1sQg5ClXFYwKmbimOK53u
R+pO+m1szMF7PkMQlrzseH9GKUnKRRx5XmBvC+qq62C10b0KuAkHTQ+b9+b+Tk5b/9htp4bnskjI
5eB9DwADeajSpugjYaweisV3gD5+ZN2e7QrcfzLeEnN+Pn6YzkEwOX1HiVzk/P8aWoxTyZtGFEkM
MNscbRq3CyVyZstnS8w/e7QKbFiYE9JDt3v1ZYQ8+6lzmbJ+m9sk7C6C11DpR1RMQxqQTnhwV2oV
+VtYkFXCgcmpNMuYyBdOO5BjXDuSIn3oEYvR99x5MwLISzXcRD7WTD99dhEfEjGX9CKFJeBGILVL
0hExiI6EN3P94C/5P+axFZ66i27+d+Yw5hUMCsyYCTHYJdFhkDmDXzoogi+krYFoQ1kAN4oT+W5h
V0LMfbjHzOty0H/fud/wC+mqy6SNTRu9ZTEtezxEvJs8AzRMpivKCB/BfMjINC93FQe86xPWQTtI
nT1Zgr1OZB/bz1dNW7BpG41smE9Gw+rbMO23ouY5G5QEupQx7ydqBefhDpDfRiXfGnGDTOdvSnxX
7HJM6tUYRmlT90/mEEKzfjW6Sjnl/8Hi1cq9KAlyhNpUT92z2gKVQBwbsifqkng6QHK+P3z7TOjk
XiDt0gnYKYcvGa4fDsm1u/u8VmjKXyGVRyPEPV3kWXCoEcMKT6U2uFXuXpzuoJQ+JkUTaHhsPXER
hB1MrB7T35F1f+vKzpCCM6jHNvL7q+RavVzmbkwSSGaWXQ+KXHMpw+8s7oXSSApdzuAm5eRBM6Fg
/0g6n5dCVOhAJPSDlMLvBMV2KyvV1b8ncXLQ2UCznMMUEAiHIUwMnxW9q0cGFOyWPGk71uuwrQ+7
y/hCCnJcUZKkSv5LC1cvNWxS7h3lUoxqx5iCPd+a7kVlzEMZMjVcW6pJk5mjxGmE/Q4OhgOJXeD6
vf90xJYVjWKLSRlOPcyqWw78AgBL1NF6hVB5sjpXrCBnJCUkDS1f+HEtI8hy8RUInUKRJkmItHBG
hzTP2fzbDM3iMP4cfwF/uhnvFBJVbRuoz5zD4ulIlqCTsK6foaHVtXDlXVFgBgzrerJYQX77Du+5
owrUVt4KiUcbHijVT7uvk+2kEobYwkuw3qmqKFLJsBQUyJG10fyYUgx3bSeJicKcagyHEPErDFCZ
PqKNTmq9deBTdRopGK+h/NbnEc2tBO3PamDkuQ3pSu+gXes3YfOKV+8toSxLw4xtgZrDKs3VlNO+
45EiIo1wyemm2YRvEQYBfPYypoUdKp3fMRvWWqjG9kB9Gnx/g0PbS5IhTwCcHhhxLYYEW0Rlp8y8
DTdnaqPuw9MHDk9CnEffFXUAfuzMBgghbvHuXByXipqwfcmGhuM44pC5ZLvXrmvLH8OmFVlf1Vsa
7e3A7YZLRf3LMUCcYzHA3CET0Wl1LIThxOfcG6TrWbqIVkwkWAefTtT1QJ8B452KeIaivtH+nh6V
sFgQIIhqsWngTYcxRjuZapBHSDyfv6QfbcV2/QF3NALal+Cuje6vhwK2837yPkcL62TAOfFnnh1X
m/rrQMywv3xtIpOOnzCkvmvCDiCh07SrneK6hHf4u0y5QgueF3aNOzQLFHNHyQ6v/BBvbOIEMXzp
V7dNJE5eyieC7fUSQvSEVT6PNiNXbTQLJvB9eXFsfJ+z3tzTg5fh4gNq7SdXdl0NDYbsKdD/T135
sV9WfdF6YS7h9oyXM2PLZqvsBwmf4piW/sY3IQTP9jv3/5oiKVuCHq3ia53OYGD8faFpk6rL2klX
SVuw6h+Og+RSvs355x2qWjlbY7nzRv1tfleGnyJ7nk5mU5eA8SAirss0rVA2MDXdSbL3dO2r9J+5
dLHBkO1+2123YfoSjxB69PDSCvAaU/lBwcUo4ZKzhehu1ah46keU0pfZ66aXuaL/UGBRLA7RD4XP
RudHekcm9xDFwh6jLYW2cQxTinViDVHCSnTKq7Ec17x1tu/5ETZM72EZ14QOVPctcXq5AQeIRw2c
y11Bgkq9mWryDIkUPjgWKFhFArwsg6NYeIjETFghw51pCx82FcAHkxL7W4LDy/e40u0GAGeAVd2L
uP2bzvPdY1EaNgRGOoOCEa1RzbKdgbVrYOi/BwslGy0tCWQa113aShuJdazQB+VhmX0lqMxXScPF
qlZDq4mrgibj1NskJzeIE+W432lLCAPiT7EvAh0Sh02sWaoVcDnf2Zo0FQyXtC4fNplM4/+bp8N7
v0vvjgqDonkaUzGXNoSRnIn/eneHij9PjEG9B5yRpUbXBambQFQ1ATg2sVioQGZxMbAEdD9dLdUH
eo1SquO+zCFkpctW6VvDAaWSRWne/XyyBKmzekXKbUviLYYLHEGE9hNPPUfOW4wRkoQoDydiCObk
z9OkgV1kfXDTC/mKyY2zV4nS7i1KqPJtIZg+8I9AU/UGOcY1UE1r8d1pZdY623m2CZcWB0ZOJfh4
8dNEx4+svVEjiDmUCqQmxEKvHziRCHg75SxaaoEI0l/ITA1wZyBNNgyEiOuRgwA6m97uOZvw9etI
rjph5EjOAhkGPYAVB8HmaIp7ajXF7+deoCe6OMmxlGF6QaR2R1e1miW5cZwmoHLNrmoi0F3FhdYM
iRrd4xE3rwfESjy4cBOw+fHe/98yU9un9y749/6JrThEURvRwyyX47I61JzeNNOWcC90I/8EOQwg
XsM8XrCfx+cf+hD1xdSIYmkv2XfQkHLJ2B+RB3HqMNErbAJ350yWAUgLBtUKNvaiNC+nEpeNbkGs
ymRJvPJy4+z0n1yvY1KiMyNscp+xiQuSv/XdsHZgj4xlphjn1s4uSYERspldLAHuQJCRv/51uKWc
lXzudp2AuygzF4I0ymSqLSxswQOzuBm0EklRz5EwaKbmLWmUSF1GTyBlYBoqGjIxTQfYKoT8olb1
OzUkK7imvhXg7Y7kcFxNzrmnbNsL+OX6yOg4IvF64sgSRS0DqAOedXA83p42CsQ2ihPiLtaGRcmY
JCxCVlibGBFSHmdKzWbJXZhk+habtyGo7w1QSwj6dsgPCxwLC/kAgSMCPHfkjzaDRJM6rZMUll2c
cFsqh4tdfIcwC+II7b/aZ5M4eXrW4GzvtDDDGWLe9MirQIZOPZ5SDLfgGSWxD9wP+xBi7Uysaezi
rwaa3XeIwCVPlrTcEiCVza/gO65XVOesfu5q9mVFVV5yl7HwVjSfmp5B+MOgi1PaaqfbpunIOAQp
Fa3E2XOS2Q+EqSzPO/dWplppLXpByL5VvzXi/eO4WCVFD/j40hpXcNEC/suZP4Ubk0XZ5ozo6GqR
z9dDhuJZBoKsIA+UQpMZc1lrgBE63osMKcdwGRQ+4H/kG7jG8MKJPb43B3aiGg+G5lD11rCKyiO/
r8mlPUagcSdMaYu8on3Gbx66wbF+UmbDd8J61qbNWsUxvI+P7rOeuwOvBCLFbHsLKuh9NJ8RE7wh
YcKSP4g1/dvCOgBx9PJFmUII+bGUetL/ygKQc9oqUVge0cQJbnwTQrFOR5YBxKsh964ikyz1VWmQ
a24BwIKmHlRbmakPBeuEDlpTFMW7JcpKe9aQ0O2kYpNYWIEaxMDefsPLN9bXj4gcQdiMMWPcEU3/
fFZQmBEGYDiaClSsq7V/J1Brzp8t5T5kznVxqJhnGs9DWhacisHgTHO2atYz/tNrWFSRK1sOIqt9
SqX5qjQOlYOZ8KhqJogz/9daGizscrTYiAmE83ubie6NdqoDZ/byyPe9HZIecH8U0ubs6nM0lK24
8Hs/0Zu3Lg7QRqjjP95fUHskuICitXP+gYJM65xirpcZ4JzzH5qNvvnKh+deds5yYW2dRNNZPW8G
4lwlyze+yTrUl5Gjnrsw6RRKYz0MyTgIydoErqu6lgX+Gkf1HAYdmNhkqqMI6GqpBjiu2ROAyX6v
sTxr2FTdOsoV2q1db28zh2NkwPUPf7jkoKcn8jkZVgZjUhwlLqDpyfG0uuz/K13rtbP6er+Q4G8k
fv8pJaMPzd+llC+qyUG81/IZ7Qr0nvMPzIBAsk51b51Rwc1uQqVUUa61r3Xqz+7YEuv/R3kHm+hD
B6wCSkBknwgDstRsHlo/6oQQRPYGrDEFzx8cq7vNXa8wWpWhLnn4pXXsVBz0FHMTeeg0VBzpNiY7
H3zMe1pl9CGTGfaau/9a1Ele066p2Fx58K0l7dK2zkkmDTfV7MPTZE4PCMQ/S60wFkWoxhGu1Ybg
2jIm8aZR8uELrZ0oF38tuXox9G6cFVJQdZnxrZb/k8NKaG7Vxrjew+T1mG7muWxr/vgnEt421Awd
TGc9WKJ+wbvra9g1CA4rLHpE6LXoVJFhI1J7kHTEP8koi/d7TQAVas1y++IncjReeJVyL7d1yHJ9
CqP/rKc5vqyfB+aSLoUjND3ZrFCA66vPsYcrG7xuH3IYKzeZ0aFcqKA8l0XlMayD3LjgxuC8zovV
Ik0iZw82WAUo2Q4PIY6TwZL7b8GLq2vxJ3klN+n6+9GSLhgfkP5eN65qxeQIzUjafYx9nvDwkae2
EArOX/9uuyCLriMGbLZ554kEKbsJ+CQY5gOirOauG19ho1e9s1mD9tMyq/5rSuPFYqiN2/4JUQJo
H3+jRhdA1cFTCQPwoqbesbaN03Pnqu8joG0k06Q4ZLn13nYAaGE927f2CMSAIVnZTaG0NUW/NkwN
/2cVIL/dAlLX90HT6wXDOXjCEaztq2uK7vI2xtKvJSt1bZhogQN7be3CTkSy1XelRLBQ06jGUgnd
gUSafkc2j5YMc1tKNVGF+YrOSZMsFqXQn1Lbrug6Th+/aPrbxUa5Jy/roPLQjpQuLkPQsX+kAlTE
2RQz4l2UdvsZV8uW+9dHtr2SvIoJAh23Hwg/KNFldNCcjUyI620N2KKiqtlQimxjGnMk862xMUgH
lrOx4bdpyiThuwWBVbVrxhVuyXQMYUEkxooxrYUj35WvP2V0PMyWoh4wPnHv6gN8XC6EYGRjaEiF
ZOZLCb0WyVhw+6UuicDITnB0SfLscDe0mIZvfiwyQu2ASCbCCMy4WuFfq7jCsjcym7nl/Vgc0EJc
p5ryounv/Vzsjs95+gr/hTwJTqUkJHDsV5eFv4mEuSnjaPB7o1RbRSA1Bi3/1GeIMZtLVUZCzOV4
KwBSAwWMW1PNTX3L+2kPmGgy5qKkoo/zM4lNk+D16/csUfPYO0H/HbGtHT0LupEjnD1uVUMHcitD
egyZC3+BCPDuueQ7/TYDa3WYfqVrY6JW8If52NKVeFdJ5oRt5ICxU8GT2gPcyoXPgzY7Cxy+Hntn
dkrWsH8oFI9wnXEOQJQFVIjiZVbBYeD+QZyicy32zDJc3EP1yofqe0dj/YkHow6LbN9CqnDijqBJ
GTj8dcGfNYmhd0DxMcUg0B7bAjdwO530xoV7gOvHNZ6AMPImOuf+BR0JWG4pngXOcmjD0OxhUZFj
SmJnfjbkGqy7/9Vj4a7v4vWWlcxdUeJgQh9zS+A1p4ZoCqZCaQ9F2zxOJcTyibVs1LfaS6Z2G72J
GhwBweYZfWAc2QgbeGjYOtkXesANKKDxDSVdlCgoazTNZVFSEp+DQIhEZYiGWRKqepG5E3SPWDd5
b9gxM6W1dw8ci8yXvI04A33f3iwfVWAgZ6CPMyhExnA6jjRBHjFqTrR4DsoyRgdBMBRiH7COch9y
Qp18hMj6iyG8TsLpLGGcA8XZmMi0+/JTyWaP7J+z5baQ2GHbNfVW7AvVmpMxsfGWSvQg+gWUlQLC
4+JVlyWWw+1i72m525eBFL3M9eDwAt2ZZkHG8lneJwHW4/AYSjjSSx9Wd7ID6ZmWMv3fOYgAlWPH
IhEsYHp9WWrorq+kRPkj903UWG4YvLeBMvrmNk0TewKoveyKAU6LJ3eJJtHsujwds/Bmzd7ZrlPF
TrscnbKM0C1zQDKOenAtMnbfqqAm1QDg0AybzyUFdTNBrz9Plg836LrwwLG7fHT+KRL0D004DbXY
nP9Xgx1FqdR33OXLdpwJRd7T7hRToog/3Gmjz0gv6+ZNHI1+4vob7aR1KM4a+FAyhPG7/Ea+8hBl
eV5Rg8MkWAkwMNBq9fNoJ+em2+F7luaY9S9vlHiONXOZ7//tosobf4Rxb7eYppGDF932TM1ljCJS
rQbBOyLXAg95EnGEmWsuNgkZwJve+sfcBsJsjOLLwMXHQMHXqduI6SHOxiRnFYhIzrYEwrfNYi1I
VQWhFpEPMmwiFkV0qPXqK1uuPoPENl+ejGKB5ZcrqGi3RM8cJuDow9/v96NpK8RsKRqiYmDovgL9
WYRc44hGYCr8mocUoD/me85QbD3G4kV56SWYKK+BP9Lj1ZFZQDftJO08u2UbI/qPsRyUUBfqWXcy
7ZxOSS3BIajDrtz7pkWSy9d7T1jYWbfQI4M3Kz68lBrboY+QUmUWMigYsrFammZy3wTtcGwS6bVC
OFsjS9474n9VkB32OHj6GFcje5+HWLnisvumypYk15zwwQnIyaXcdMIn3GI1a6Ta41OFEp6kMEp/
bS/pNalezIXBfvMO1ftJOBWGeKRS6zmv/Zfq/AUtducBkk8Nj9VMPbfFWxnJwhKnAMdgdtZCLKrk
FwZs9vgof8I2KmJ0HDnfruZaLxqX3xksCJkD4uHaz5zvm5GY+cEQlz+IK1ruXoL3O5fOmIoQsICK
InfA8YxMZmnYOCSykT+WpoZWRtS6Ttb3mecmSB5EfqVnvY8V8v5wCl+Nw4TFVho4ExuQ1tzloIjW
mCixZPfhaQr8p5kl+EysF3f9vO0wthCZFSlGQ7+PslyFPrp44iolZB2drCIdr7IS2PLcmeVV0lQu
SdzJqWUrPbwqamSGDiFmIv07LlqCLo3RtpB2n8HJY65fIO8fV96sqHPGI3Yrtx1JMydyjQpvtYYC
srtHJ9lz7mI4UmuvI8XeJtrJLTB2mKJFM6qYD/Liojz2Yq1MIOUxC/k4sfTjtaBsqnnXHP8IQTz/
9wg7O5/dc/QAryzIDI9XgU2AQuqpYI7UfVO/nnIWeNtaBKnKuLGhoIzYVV2vqbZHNo3bAoW7I/Vn
g3ZxDpQelNf63+gHyMtBJhh9ISslwL/dG6KmJFcohCVcYHsOYwE2DUaOxW60ZI5JDsyYmVzZwloN
zPfEdS29I++uYoKiXKO7AvstkojVToCvNA9Q39ufdgEF5UGng/J8pcMRjeSBIPhfCh0PYN5cOZ3i
LZ7hvl4Ve1zDum8X9iPjJGyfM77N237aPTqA180mLOYRgoPfOVyt1XA9Dfg+y6NCUMP8R1inmqh/
xckypVS7x18ZxJkKphg2BiSDssvI9/RriDP8R730Vt1fvX95ObK0WcEvAVYPmtTEKVj0qcGa62zC
mzw1I2QdFM/9kWmgxoEKpy07c47qtz4xof+ul+bSUnKbzIeVvr1aZXFtkpCQAjwGrCnhPTm04L7Z
/YMfm6cHc3gTb3kSDluYAt2tv1iEozG/SK4G+xuGd7zdkAGZNzqxY5adWg+Z/a2lthWUs0vwRoxM
m9gCD/QMrX5JYvp+IKNTlZU9/fLoLcJ45wzWm6LTSa2Ke8sKXbgFX4cqN87KyKwxZITzgjgyMU4w
NEIws/TZ8dmtJFYSf+NEOhbI7bwkh/LM7bUYrF4Xn69PSPaYR0HmAsogbB6yg2Jem1nM0U/V6c/z
JJz84FooFwNIq9+HxiD9dH57VqCtQ25lORGbjqWqCN6aQKVhRhm6I57l9B2fbTEd4kBPr2oRBpfI
y53C8jwEI5O24qqSP6Yc7VX7kAOBHTtv3sdxLBbHq/91HBDQLjEXgW+G7cDFlh7cW+LYZb8hGemL
m1bnttgN/nK9GoIoTPQ53D8DhceD2VNzJdBBehJk//dIDmbr2Zt41ThWPmfUFOtZ71UYt88XHgJ+
h6s3E2b/IoXZ1rB585BNAOVUOd0w7v0U6O+zJfnDxRah+PVdlml98aXOh4OpKrU37e92FyeL2JnD
PVl4ugPbyzww+7FrS9Bur2Nz0vsCOdqZ2pqYyeESsC+uEro/fYPbmHzpGK9ZlnrXV646kbOlqkTX
lWptnKFvFYie4IkKW1HQXtTFTTW9wa6R6lQQypRjWK2MYIU2GFUOiowSnsYR2z2O01JHiUYddgtq
INQlAJZUgfn3t1fGzKFhitp/a65No7HmOPzPle2YVzQIvi15m1fklccQ/8pYsW6Y/pdwdIkRfD6p
VBAdACWbDBTrsSdmvSEYaMvUFhYGvIrZyJ7qqRgMHLCj+TOLDkX2sxyoTqZc916d+yHv25YH658T
KbOIO8LX+jQOgiw0fvMjMSAs3hJMKK9F7kqKTnjKvE8/puueyHgXlRw+J4zdqe3HSWlTxFs+XFq3
CdC83PaLepsS4AmHNgQtIEYYgHIESm6xTaj1nfIMBEfnEZ/GahLUrQ4aatJWszHsVL8tuR6coKaj
9z3rUuJx/txb+SDleS4fcDzTpabaSnMC+pJt7GGT0FmHFzSq7rEkn+VKzuIhoWdHb5DwipWtnB7A
znnPFLfWNwO76WOcbUCSDQLk2RIvM+ktQHoB30T1SMDmbsaEu/QwO/8pDBHmhC4y+nAHCIzK+Vyw
LY8ms9U2KXP/9dQZdLBepRn5y7ZYmBokfSZb23x506A3FVNu7d0NjLo70jNi2RAESyPMA0axb/Zd
HElmt8wqRtVNCvVS6tNoz6NU43uUBq+5PMPUA9lrjs0qZi7VKyLzzi5NxIdveL0Oy6rdBHjUXwg2
jhWNztNn41fvn3l4mXgeeMFr4yUmJo3PlfejJdg39Iio7bKdb5x1AiyexEtsFHDBk7k1UbusGUw8
EYstc6ChpuOJdboQX4xv8dTj5HzyFQIHail98zMZ7LCB3HDgZpdIfXLYVmuckMRbY8x98MxqbxRN
fDHBJeRfMA0fYH/kY7uofdvE+CWu7qe7LtK8/X6G0KfT5CTcCbbxDD8S5N8MjLE81S1LzvjEX2Ba
uQkw0O5d03cKPuwHuhxYnP2q7aQmGOxnZMUhw/fcK3i61KGEAJ23g2Eo7WlWWu0gnpDBTbPd4qAm
hGXyLSH/+fhwXdqqQk9+63IDVk9mBO1SJ6W7g0wnowFjxzLj0RIvqhNKqyi59BhvgIVu/XJTnrAT
y54lMsylhT6ewCPxpHlugMOZScsfaDdRskZcIu0mcIUTEjzMUIp17WM/4qJTW1+8W+RRDwmEYeVv
JZfP9G+wq45S+9fwHbnOn9+krObeI2zQ7NwtAtp1iRBJdBX2KpMZplto+Ed/HRa/uC53JFagvgqC
INd+H98m+uWixfOiHTnGS+IkrkPbQ45sMLyEe1RXoqLt1OXfEVk86iTqxVuUj9tI9dTX9TDCj0Us
yuVPJEk4TZz6brfFqRbxMvMZCKIt1Bf34DtKO9k8d3zlwZEc4wBOej/BZkT2hje0Mec28gNHNVIl
SxFk9GehWRnCicIe6Ax+Z1aNhtrI6eYKyXELAiHN829MsPE0wzPA6lrUqP8Etu3RPzK4SxNzMBF3
vivolSyxpUpxARPEDbZd1e52GYyPkpBqGkOM6bYXxz55aVWjIFcWt5dlsMcVj2XxOn9vzYBlqNrd
9pUfQhyVoeuenvdnBwsMaSxuObny87wka3J80y1YFQJdTF1PU0Jd6YXCrtw/UdiaYi8kEkK6ba+M
IzUBWzk+fDRUCPifsAZoaOcVyAGcclwke5002pedVSP+j4Mo7m9vhVtCPRV4zMa9rDHDMuVd/FHK
DArr7bhpdw6L5wrLa/jxZbK6hAFaxNrRwIs4W+bJTFWCAuBz6WcqeWxc806dQS1BjTE/01L73uZg
v4RoPwGFYy0Fg46W1xjZS3cfszIzWt9MPbbvatcIarnyFtECkEMtlKEB0sYTSVaL05OBZVZgR2lD
O2tGJLhAuqtXt6pBC6ZnSbNVrygRNSJtwTT/tZzUJf3rmnbEXnl+d9H2KSsdCxc3FfQVqH20KHPI
E5jmuIlR+AIUfvrjoA6wMjAcGCmFNffwUwtGkaGqirOpGJhmnIeYu4wZl4aDDkjFqyUc8koFV+jc
g6lcAbE1sZN1gSNmJOV7YUfGpTqifAetu/196OSoEXjdimq6IYcyq4txBtpdAcdqenLF7qp0vMUA
1IMVoBRto1y7/etr8q7aHfe4CyqUL4V3C5symtLOPukpNV2OQ0QToNl/FAwwJ5z87uMZkNbztRXA
tL4gAt+0ctd6UuEK3/8/ScpsrIU9MUkTRAfymJsxKdiTftae5m9Ho83iA4TlzJIon89UqizZxwTo
Qs8V3hs7S7WvCwDK3L/Gj0OwsL7l/45W4t4ef4Wjapvk7mO+gcKmXMyFxo/+jtaZ6vfYgmFLkVyF
1ZMr8mVvpPmfuxszGpFIsvUbNfgThzVrWn+mEOSmzXM1ON6SDPIA8moY5FfNB2Y2rn7b4LsFaZ6T
7nS6YbHzRugl4SJq9MVt8AsOLI1vfpodjV2sjlD4QxoRoRwWikBqSOLWY3Xr7OUJQY2O6y/837XY
P3Q4fR3GEAlA/Eqv217jeZcKaP6pRvJVyW+pOZSOl3BheazwQdkPjJJqNaUbrw4V9s8A7VYMEQ+d
KEh92Wrxh0xSfRIS+9mTBC/39+q2n593MxTx9SkRS91ZqgkccgJ64SmQML2hkVQybSH0PVIq+39Y
ULzOvOCQz15h9Equ+66qmdywyni1erD0zWS0ie3U4t+dwwkIrC9owtD+VF9k1e/W6vBk1HMS/oJz
K25i2pDu+WAeWPkWr0kJBmHUyjFe0DQRTFLb3TEpfZkIxxaHU+BrfYA7jEqbbyc6+txl3UbbxG7f
CF2Q3pNXrW0beOIJnoef5zE877Ozp9sf0l23/fVVlGPXTihnzSy8v9fn1kNpTC+NMTqeubT++SPH
i7MIwlkE0L1xhALx8S0DdYJFsTUYcGCMIlqGnQZhrR+NUEsOnCMnx6xFf7RuemGkTKbu49I4EdoM
LY2CqLtLZsOabHf5afhHF/3Luxwew/HlLOsfQPhR+FeXxT46Ejnmsc+TAVzfJh8sR6jhGcXYhoNu
4WwYOXBOrUMsfrDoD1UO//gtsho4U8iJhf3rxrgAVFMgZPLv/D+6Nk5gGN5RsawjyHzzPQso9ybJ
WPk3xSX8I96UVELdulgaaw6n4IptcYHHE+uFiQZlDiP7eH55AkZUZlZVnj8/Gjb1KIoq7zyp9410
S8j8aJSVkeHgW+FQUfLo3If0SRx3KF3eHx9fQfbQyH46FKE7BzZW3gO4tYszYcxVsMcI1mnXG4j/
QZMxF/g74sbG/X0/hUhE47UBcG8E19XNJvqIp0GPNwQHNZavCvpqrHM15SzopLmmdg/WeQSiZ2ls
MEMd4NmohbLSsXiSSGCrntcX6B3HtQjj6yCk3Ekd2+Vvwmu3HCQ6qrxCxSqCmdJ3PMeQm+mbiwU5
q7SfZajjRowwdame6ifcoE+BmTUNhll/IQiIbPXutfu0zu++9hj3oiesmScekKIX5gFVP15vBCtw
62mbSjeiiTlxkpMbGUabGXSz51ZeUMX49P4J4SLo5kyzzMshQA+PcSYRiDCB3QSmJtUJp8Ja9IRD
qk+8HhsoQVyrxT8mMnQZ1DpZpToX2fINp/Ds0ONPQOiUr+YNrGv+Qj8Ki0WwEzN3Gf92lnD09ek0
tE1M7q6an96sdaFlSe1IPhfhwoK1s0TWjCeTuEv9+msJzgbfYE/jBbkvKyqdo5FVqFHUZBSolRze
ayRchV6q+a+3LWpq2y15h16fjgEaEzi8McwEGGJZhTMx/CaOJzD+fW2PuEBrJoBUiz5jnHBkmnFF
0QYn3SiNAmLACAzxMmvbdhrOhyVDJX4KjVLGBHrM6dmxHp8M2naAw/gBYrTQaTLuOvcWaJoyTS2y
eZ7OKDzlRQeqJ2n7w+8AEOZmgE/NYitysqQcIt/Cr461Q7vXci93BMtGlgxwI/96VZ+C6JO6lJPm
sy2O6anTmCXn3q9kubqRMVCwO14lZOB2vuy0Lxr+xG1Yv7k57NoUrA5ZwtIjOdzO5ui/gutvBI6c
es/1iz+i1E8FbYOPOGzygbZGw5OwCNNf/mZBS0UdGkbkSYMDIvKrIRyZGVU0W+sHg8taX5ykzyvI
HoNW8xFjSjW7ifiOS0clRTyZ+RXqc4AgTQ0zZA7rovKuogVi8DqL2KJCZpB3lppM8/gdzl2lh7sN
M3Ie8NbWD/rT362+P3u7i4Uz5NVejMuIXF9uEZdf0uFlHxLU5mZgM/NdWhWKFecLz1feTxftJa93
IKU3pA2Ei8pqkXJz28SgcgE1k2wmWy7c7q1yZBvkg1dX4A1TECnJmOx2KMKaT+yfhYb43AWhK+y7
D+rdbr5exC9OFecy2iEGqKY/FkULk6hb5L6ctDfkglSpDCXq1VHTLmi+aVtv8DvJ9W+IrKhICTew
9/Cf+cpnWcskYN/pwHeXO1SYck6NNe1dKX+mzWe7H2qFVr2gZ7hF1MO6auOGby/dHps1OpdkvGTa
ExZXsiPU4zw0o8sdCBX5Jm0Ep246GOPc30+lmO80uCKOIC0/tQj2Uvh2E2SXNh8otcyfUyoWQgni
JpnEme4ux289y8pc81XzXVEa70XQzOIow981DqMCS9ItKPQoJHFXIONeaLMd2eZyhtTkQ9bh/DBM
g4ZLwXf42MtBtwjNdcPK4I7yWhr3yUP1aD6VdjlxiHMbFuTlQNG55uo8+pV7rlnuuqrZxxmt6SPG
qWkLUy8lUGmLKiYbzy2QRc3crbN9T/v0U6MR+8xXnYfUOmhq3U/LTnp0KVdJuz/2/wNP3rNIh/8c
LJ/eRvvEb5AoC9zQRMDS3oIMqVv60d057ik+rFT1tMXDbznr02pSaE6rgfMsPcPKEHqvyZ7142qk
o5k96yOmRwU++HQz4GqpBYRGirRtr0rlLa8K12uDV7OcqIJqKcHfmBf6BSQMIc7q+tNG4AEeSJId
692UsY3w12GnrZSY61RPg04tDB1WDUfqCvv+L5a1Bdwt1KqK6O7O0bITwctoQazWmCxm3ocR7bvF
ihYBoj6XyMpfMZEXEe15Ig+RqS/XtRo/5iVOC9DOFAxWN9p7M/8ZmBagQ13VGLJqJyuclAWDOmyj
167Y/1eKFzq7n8woenbV8mK78vittz0jmnVZNqNRzA0Udfb6GugGhAeEk/zslxgNkCHZVUQ2DUC+
i5MXckmLaTSxnFDifac9ieFCUJWAFrN2lTO/fig+zs2TM5Una9XemMn09wKDHUcrzyxLTJEKOhZI
Kbg8NTfWdp57MU4I5QMR/r53fHDtWTx2Sn4//63mM9cx6R4g3jmm6ufMrqcEI+IGgNHEhK3pxL0L
TjBZNxVbBMLs0mVma7C6XUuqeZ28MFJP/+jnseTKfm/O9QKzY0yFS2S86pJM1iUDkKIWm4hIly/i
tpYNChnRABUlLhrfOQpIMyq+996u2iBpNZE1gDNf5J5bSznvCGUG+XbI7z2rI8GanaTjoTCnaPrH
5xWCtSmyydOmrmkXi5omA+E2Dn4Zne+6etmojg9NZbeUJelZlIiMqPlRic9X9WcquvZBUlUKv7s3
X7CW185QObDeI91EpPGAXyjWM61apIP1pqYZ6Ffp6yVW3WJXhUKgqDdhhIGCc8E9xHz6ZUsBky30
jrPDHQ3o5+YntdqMUX5yL6v66kSQ/uWk19m/QF8namwWnV6znW6PjPe91p8eXYT+Ql3iUAn84B3r
83f1OIt6NEQ78RDvAjMggwlbxCtAdvpd0RgSr9FBzJxYSfMQ4yw6HXrOTJaz37Mc3Yi94Wy6VNcg
vYO/gAl6eKi5f1PIoIrsE5UXROlPComQd5kpaHVRXy4Mo0ycMk+nqCnMAOcbreRgGV9VkJ7twekr
Zxd6MHCy3jepHjMk/5XGkf+uD9NXwfhuUbswsltn5gQY99ftCpkdOeRPGWpKgUmMoEkL4t6FLZKX
qazULd3L4MZjvVjX7u8E/B0R6Bf70q8rjFOlA6h5Mpvl4CKEu2hu0I7ttEYBUOqiThYhGi4kruzg
bpmrvB9+WTFr6WJ1pj3oeOyvAuWRpDMcwDoAsYdAFUzB7Jc25RjewxOwR2YtK3g9ScqLs9Y/JD0u
KETesHTzaMmWJvaUG0YCsfHcd/JUaEVnPOYBipDLqD6L2Yt3Fe+vOhkY6TMIpTJ4d9L04ayBnIaJ
YGojWVEL/tD7icC+UC6z2sVg2/5TVjwPTq6I6EyRgJAsE/AhR9P/WzLvxLgSVaTBMLgknto1Gi2U
NmoFoNNKJDixpqGT1Bgm/2ghHCTQwWzP5ADmRhaEkRbnFA8DKmveCENZOZoN/ua1F2NWH3C+Z5nj
tr8F1LZOKOJBUZrHJ9W2pSuwsSNa5UUrR5PAyyETBXGUzc1Qbeo7FCkcICVswMis1rQhQIjl7kYs
/QuYIou4mVjhuNlL9wTXXT/KtbiA9eCgWxSLEme9GA1t+5a61YaNlCZb1+gxeOR7xwbxJrPY+Wls
nPq6bhh61SiuRfZRTpk1rtxkE46gmP9GpnkNNzH+CIe3OnKGTefZkP2uVrXx3AN9/SWAeQoZWLdh
1qQArsu2aWCrGxLElHxmh/xvlIDV6wblSLXgs6II5+7QxwJKN8aYO9sw0a+YdzGaeqZehLYBA3mS
DMfGkinEjs322rTjbCfdnn3HBjdiFv2/DVnW/K/uAxZB6/lhNUtISZYX10t/O50aly2PTgMyCcgt
ga2TlI6+l8EqBn+GAnzcpgbgw4hA0GbT3uYa9WovQiiWJqULsHu46vPym0mDZXkj3O4VrvDtI108
vLjjoj3JEXGB/B3Ms26P8lpsunA8aV8QcXKs4CTHJq/oxAZEFFqx8OlhjgcmyuTrHUD5IWrDV+n9
vSlzaaYwbSrJgsWqQHEJOt/1H9sqc/u3eyq7w4W2eiZLVEhOVuXNbGZyglpRENoio9mJIX8LBTIa
1d8arXFtmuX9VFg4MBI31r5MRJOAs3SkSfnAUVy8Z60PegrNjTHd6wxBA99qDilLJkk7t72DWcdi
NHfowLGNRI0szFQcpcjSFaU8NMS3SQgMz8nlWyfTD60xg3W8AYhkD85zUjoysY8PM1WVxSWYCEXD
OED205FIfED8VSu+4lbGiLEhBrRF/gNiwFjA3WUiy+EhhqP4iUiqcMKTFVk8QapyGnKeYC5cp42r
FqTSRnfBhZhiqc+XJlk/aVH2ph067koVpW2ZzLxdqAKADNw5bjverjMpD4qoGrsERhAN2O3fAoU3
/xi44S6a/eLlJUWMyUbkSO+bEuijJ0WKBJvj2IAYa5sPefW39671PqfzyV3yC1oD6oR/BqpO+wFg
vD6nRoX5YD0DztwR07Pk9QqEcflYAw1qi2FTiqX6ghSVQ5IhYHQv9KMi1RUlGvKPtWpgrztgD9lC
574gxFcwdxgCnwgF2Vrp0EPNOjBWAGyXLap0e+T8i+ME/ywV7L5FXHVzXWFahOWoXWDzwwp38bEW
0l9fthRvDhDYV02EW52/tMpZezC3gVCKAnJGp61vqjs62mTwylNzjD4oMZFbsdGSA6V26lii/52Z
XyxTVjqMojtBrxtobtsdDO4YMZvJvyQJIDj+Y6IBQp3NSTAy5+Qt125uj6Nv26hILgMyTft4U6mY
MjADJZaEKS+wBFYmf51e+a+SXxx+zLCrfSL4c+QVuF1MfZIERxDvvwdq/d7GvgQTfl5I7AYO4AYe
ucvIpHofkfw5HLmjCXCAo4bdeVMcv4M7R26VvUHidrYxEi3gU8bJrmH3yugsPguUiV/3s904e4EU
SgJWTvVcfljfg9XJyRwCvOGJu+6b8SshhxmkEbfY0NKCL1XLIliQTi4Yz0kGPyumXAtRooafQwOX
bj6o6x3RBfNAlcHjQZozHIwV2K5sKA3Ir7c43CPO7jhk4uPrmzPeIZ3gofVNtO1caT3Tvvq+JNPu
N8xYJ8br0CbzhJlvo5C9U9dKc/BHf2NZeJ0mEBNXAYm379eLutHt4J8g++7so8As8He5alRsQwbC
Oeb14KNTyZEQkMyQTVzUpIoqTqiGhDGJI5ijahe+ar34vp3xrfU6IHPpOIwN9QMjEJiwCqXeM305
F4TREioTebqp558AvG/+Ad/2Fti7LPyQ0dlEHBBnBDubNR73Bnd8Ag5yrAjPcR3gUWeFfGew4nwA
4hNWxg9NIK7eHTTml4Cqk0W+HdyFQrGbrtD9d58L34ohXsEOPQGo2SAHreM46h0s9Fhv6fWOa74/
YAbfjmVRdK2rfEo2XiEYZTH+ZXIJMvacq5ZSHBbk42AriO5CMaL2034Ip3AfWeyHJt1pwdFd8hke
GR+1n30dWt4U2MIqDlHGnVY+WWkGWjt1bymJD+HCTg5FT06rjR+z29LkYGUvP3VSudn89eom1DM9
dG/D11o9DO5vOECWbd4NvVIhVK2nD53Ty+7bpcEtfcpq3TgCvgR79hqckBrAcq0aW1FZR2wN9y2a
QQ91JPvOLuCsba2Xt9Cwxz1NsD/vCRgW+KXYprbPMR3nqe5ZusgGs60o3qTDYdwCxTBemwE/kl3j
pJhbQapzuphzR2Q2BcvXeBqGcNYnWUh1nU86rJ4J+pckdQlSwJcEe+p+o9avrVUW4lvGAEWsWzq/
GSgbdGkyL4ULEMp5BtGCyUFXSKS418TBWSZHrBbCI7xLpBkNSUjFQmQP4HbTdAZJwccp67snsXbA
e8MV5K5W2tTwFJEikYGqyeCaBz3Kj3ye5iEC/z5mlOZoRX1XZ/aXGRQjIbNxoSJ59WbnazSaS0jG
OGVcNakyzhPLnvx38U0VUHQ/WGXRbr6fNmIAsG6TyOdyMFczXg6t6lkQobUR7KO3XaBhzKk4/egK
RhZQiDIZiMAfH2ekVhZ2JVRqqB7Y/6t/Lg0uER8xFRdvnAhInFNMeZq72tlccEIUJSP9Wh9Xioz2
2jdqgry35/vu+ftgVXw88tQhshGdqfO+yNk1WXpErZ/SLuhFCKfL2mR0bcB3Tydfj4Y3pl2+23Sm
M9qyH4TpVquHEFjIQ+MVq/vq4c+E5VzWKzgVhnlqI8nMyegPRYh49Abwc22bS8NrkmP9bLZxik35
WA/flqt3fKCVNlUZJUx2/4dEMqDrWyTxKmdqAYJIS2WgJwAM5nG8QNlp5L6vS4DXsYv8MMGRbjkI
A3+Yw+OZzbzGQXZP09AOwhZyNae3i7evMeFvay3icI7RUzJj8Lupm7x8L/670W9JN5knHz+WgKsl
ZXN7Lq1vonvcQTYCPV1u214sbknp5ekHwnPDRZ+BJryQwZ9Nnj1ew8oKJ9p1dTPKrsiGe2ddNpKB
Cwy60X73DNnAkbTo2tCpUq1H/gNej9IJI/D8sForaDiM4phUIr9b7mo4TkTeu7VPNrJjDpmHHGum
0DBvsuAjRPYPEUzjgXiCKCe4kByloQxLKsJcIsq9QbADLk4P87tzZLrveg6z26ilMMtEfEcxt3OZ
io0vatPJiR5MPc4SJtFW5h8iVHwDfIyP9hvs459G7PGZVQ9lHrJRznl4uDSYg+/e/y+C0XubHX5x
lOHdK7mlmwzZrKH9+euQqMRICc9+/JtuLRlc/wbWSUA91XEWbtSfsnm44QG5xI7fHK72gRVDmS63
VZpnW+iuvdNpaGwdtxPkqramFo5kwQ0dwCVF+DBlklTTg3Y8fk5YwVajLr/dA/A/kdezUteJNzEk
uxzPqLsNyeK1DZaqA5NUSQxb4jqBVWbVx2T+DsFL1xL9tJBqs2xrj48jPrR8mV9MbOMdnTrr0SJq
Vu2yqT60Cp2W3aPu4gIXlOvH7KxwDKezAcMsGp0I7FeKE0F+Z5W7YByIhdkawBJgdUY4N3/RLGh9
+MsZ6T0ekfnTO+e2uN8DEcWBfphusHo/P1fkBrpj04V9xywauqy6+Ez6ATZEgHlwGSMm4SslUbIk
Lmc5+yR7iB2Ho/eWh43d2L7/avFf9pj5/tBB6+VBrrwWxz+zFiVYphIB+VlmyjuomkG46apRe+k5
nczFFgWhqd27MNNOvqNSVVfI4ko0dDflBrXiDdAqgjFtmhOhzoKOt8f941SkdQKfsxUMJrwLI+jR
276n10xpqUQlaBdhruYwAFgsJmmAp+mqSisIxtKpmy5FhKdCdx5GVxySD6VWfzK5cftBgQnNNZjy
O++fAbznQ5gPYatU1wgN/h0gy98tMFLadiWmqGn0nKBLxKRhgNV9eODUYHEtNV3eHoGsw6tPBTFG
L6kKaEq7CK3l2xZwpZmZynPasGhetDZYoEZDi3k9ZFxZ6OIZhmqZzy13amm9M4PLdGAoqm7/6I7K
zgx9t2Ba9dCGAD5pmjbGrnHvnQ9RhHo+QCOS/T/v3lcjiMGUOokYM4jEFdgrcgXagazlPjaGME6o
v+3gQdpampI1JPp8BPRJ/2owQCvSZ4qlfd3I+CWcP16Cb55xtVyPy2jRCl2pcWU0QLYQ36v0qb+C
VwVPDNsJAOTE0PhQX7iU5Xwnt2aY9GXskyq8kwf/exvFvqCI1ivtoD2Il76siKCtocOWAg8vyBgs
XzflS5bNPJC3X/+vMroqD/D2+/kW5LvqN+4+c9j1lQdjR+tgm7sivhHTvv7+OG5fMPmD++x6NIa+
swt+iM+mwYKIs6q2V6MjNVh1fsBcpP6WMnGLxacHQuohgmz2vTPWHqZmAC+eA7BIKC8/bnMkWlBZ
7Ig1WovI54brdsBR9BpXFHXNlULVJ86lVUv9XPuo27ACE9UKkIS8bqBEGleO36iPZ4tzGUp5wOIe
r8wb4gYWj67G5gjmLYgcVALDBZy1fkG04hdsOlM85/kWLVpHJvbqClSc/N2wk1qZSchkyBDHsF00
zcerFw0teSKxeuac4LEubhKmicFCLerMN28P+4o58IuAnU/2fUXj7GuHS5W8Hus1Ca0ov+jTLyn6
t5+GyrTBJdOQL5G0QJphMhQsHRHetS/34nykdmhQaMUj+FWxWTAMRJeDNitgbuHql5MvsluXVaCC
ltUenacxN6lRY7Z0IcMPxFTzWGiRX41ZENU5OitDxa9pKGAc3BSXpfzlpCNrrIwfQFH2rnt7YA7I
J/cfukgBEaLUdA7QgNQdgKKPg/q4dHjwpvqgbSKFHdpuytG9ipU7yU3MpjcmhdwYvLW4UCR0ke5X
Z2PppPQiJRwPrnQHeZEPshEd11rkB3lK05h3eJnDqxM/BIHKQfYVuefSWChm6GivN1vAZfOj5pRd
ewukAjLfUIW4qPewB+NryCKcVL1csnrcTrVTsA+2OxR6aSfLzanT76hMTW/ltaLkWjC4+TKVl/6h
wEibt81ErfsQ2186vQCCKn4UstzCeUgPGNcNq2M0B9o5wx8oriDfjnki0L1TatZl4/6ZbRn7cjKf
eS1LGA+fUS9gpDRphGXcYHijnxdcjCw6+J1nQm9xHbQJJjfhDNO80kVWuMfMaTHCYGI4CzopnPvN
8+dbudNrnBn/v2GeD3H/S3K63xc0Mc0UuVPpm+fQnGIqjTmZzL0zSR0oqxJOhPREBOxLSe6NEG/n
O2N78a7TqNOs/JPxbJOH92H4GM+JLHBOfp9trtX6B+jm3MT4M6BPeQ0esxJ8p0k+T/tqA1JsPb3n
qIvmAEJS2xL83Pm4R/xhBW0RuwXnwuoywqKf9/rfd76y1xopmUNSKrLIZ6IEzrYJ7EFby2QY2/V0
1YDfYLuHuEK+PxePvjnioeHrEQpvGQusTOYEgV03w11Z+5dl7nivE2kDAKUKx7bTFyceBBwJ+ITh
Xn80G3ieQeq2pOgklozCWU0MMsIvgC35BAzzq7mWxKvz7RhuBRCmYyxz4vi0OmyRqKnU65DxwGbi
L24rDf15X6FLoGseT7R+ec98GE24YJ/929H0dZKiN4qKTBQWi/I4t5aklZw3jxFfOqjxxfQgD73f
j0HlPl6pVxO9NpLpo0dV+a4Y27Ari0oTVoICOsHIFNmlvkW4QN6ygoUuLrIC71eyBfTMO4npuYe3
ZpZzp1w6kA9eZLUKZMBLR9/CjrIfdo/q117KL3HhveOgg1ySTHTvjHpHlqacXFEufyBBHDM5I5LJ
2llZ8jb5vsuT9uVt0TRcb3SXfHCyBpU7zYAwf7qzf9IrI20qkfDL4DnoqoN2nZN/7twMLK8FEevH
elKb41Jz2TZtoXFKabzV3OJ9mQxIwAstiFjJYKnyQJUoHvaVhAwsQ2MjLJXAdX+LutV23zBsG/vc
vrZso6zMYiF4r0xy3DUQ8XLe28cmUjQN7w8zjZkP1erjo5wsrc25p8E8YpQQvAB/Od4kdZVMZH47
yXPDAAewgzKNBhpt/3nIuR7iS8wmd2o1R1ZgCj9dCBwsBsQJG1ysOFQunumTXqIni7IgXP0uhbLx
3Mdf9zlbA2didNua/9InjU7xj6cere/kgbdcnHPX2RJ+lURZ1+rOOq3J4xRLiJj7bfcmM377k28Z
7lQb2kTI8KsXmkzpiyCR7XL51l5spAVbUFoPw+dqae4MxSfU21n4/MobtNGGOVwuCkuxBRdz6EBC
iRLlo351eCygHq565+YVb7vUSfc87x7ow4yUSjhFWnJnN3XEJwTw4q3E/RIaBaANgROtAaL6EX5W
2GyWnMCuF5xW+c3L02R8CKfRa5M6sN2VjWdODlKFwDqioGLp0zi1TtuFds1oHKkALVwTpya4IpaX
xEK/9UPwpd/yTrsimC6O9fFHyLwfEhVFGp/NuT2evPsJW5W7pbjSAcrJ9m74+hj8mKrf1hL6kX/T
zwgRzYW+qBkbbdu4DBTHzBaffqWd33lAEiJQdgN6bBxZoUvunfJfOV6JE5zZdlSw5eNjoF/rXidT
eUeSq9b1A6mi30cJLQ6GfM8QvZgWWYq7IdVwx91dFp5cgiEA0yabw3vZnIMrJsvRBndkTegRJ9Pk
11N0RGL0pmdaKd8KZA8DBEB6mqMFkTwRFm/wyhxQhT1wNm4DWPzBHjDjpjsoODgUefIjpr6ANbxy
9Tn1gPQtevbL333TT5wJFTTdOVoQBrZ2PB5fI1eWTWgTSq3B/HW5lcC/6YexfGsXcyz8CW/l3/IJ
dAWfbXEy+FdOcDXEwikl/t6KN3+bKmJZLdazDVvaezDIEnvCH3Ac5aJSadwE4rkB7WSsbVpRO4Yk
Rmrm1LVwoftL9rLsF6771ljR0DiWYGfoc5E37ecZBbpja5C8QDxqSy/uweMJuzUFr7B9rrUVLXhl
xuDIQSjx4iVKs7d2L0HRkQN2JUDVAlE/gp/kHF5Osq5cQAVUE7bPj2Ym8qV8qBbCAfw1dWYj0B+T
tWnVU9ftemjpVmsWfw+8LIw2U5WqJdex5me6t1Lt8jliyoiWAFmG+lEvZM2BxodaZWbwQW+mP/M2
HYV21jLtU08lU11He8o8SCs/kYfmiN76KKNRi4S6IO+N7UlTIMLAzo2qwZ2JRHNwqabWaOQNT0B/
u9ulINrmNm1XkOr5jcootdqfoOD45JyEd4otq7n4E64hNgdhR79OQHa89scZnZIaKaB1bbzvMhR/
eBXd949T5FhwaPv+t6tv8kx7QBeRAaz1pODj1ylhR2lNxbOcCXEzTEjMafMBG5a9ACJYP4TJxcay
M6uAgAZ1bEgDSrByrz/JPvsPyNVxGTf7kY4ZaMy0a7yY7KfkjJPJ1r4u00qRAxDajbYYT9eKzZJx
0rOkIPKbXGYFEKzX98LnEHMgvfUs1tCLIZWrRwX2NFkpHjfjUpjQ05XjjRk/5EyduT3zkFJTqHRk
YLNbPvaM+e/IjbD3CnJ9pBnbZSNwbaZLuZlAT2yor+QipxOLoJSY1bKf/k5aV+Phe9rD2BmRzUbz
GHypC8FFrLOtlYI2xE6G8RXKt0fGUpPAGC2/mXr2L0Krpf7dFlsHNk0dfsrNnb+Y3/6+WfidvMKf
Rc7EdtywFH39x1AmsLpICSlLIxbwe2ViCPCaTI2iq6MdU/pytB+6TpmPN8hoDbIEBuH5klmoPjAQ
ZrtDQtdj8V46SjTd7+yUa5GadcJrJZFpf/Q+5ZAuyKG72UtQt3QzGa6QLRZxBAH0OST2NK6hLsJP
vuFxFxAwmrF2x7boHTjSJ4XAiGqJDXVtorRzDLUVahjOOzaldRVD7Z+VqGrv1aS/dbeGzZk+r2zG
G1aWqqMJ6/o62oYmpcBnD6gwQ9you+TpYot+4kWey6tBy7a87VqNWd+C1gFz7yZBMc8erAOMwEoi
egkNz+ssa3RD7rj1xtTvVEi8Hltd4cfqjSWE40S52JSVuO1m0H7R8uB7ZofhRJ9WQwAnCxAO0Py2
vcIcVEy+wG2nbveUbOo13UgFeDHMvznFJeW09daNE7VFQDfhTMtjY17p3JMk0QpoSwGk0e6xstV6
R94vSaIVemez7xEeu/LXarHl+lJIshufB5HiqjKtBKMO+QUsYByGpw907kX/pbDG5BUW8fc4Gsf8
7HeV01vaCXDYyCclxlC+l+9SQ2nz+sg2rv1MYGGwEYiGZBNHA7AsxizhZgeUjNOp8hoHpGBtZe6i
NJkmSSBLEkcakmhtg8zDhgtHQAEJPOhN35HCLkGVO7sIXzo6RRKaIiksUrpA21gseurQrlrHL77L
fe9bJp8DKysCiBBUo2wAJhj1itw3Bz8YLW+jtlXoLXtOxmIRv1fKfhC5Kp/LeztgomWOCEUvsMvs
Yqq/D/HT3FvJQL5PRKRBEAWJ8gJf/CiKQKyQ8a2iOh6VV0O42GXlGpaBnjQWrWR0iX6G1Lb8Ivhc
VBCridQUrKNudRe2rIs2yhNvTujrrvDZdxhhhoXVqBGdXdJ7SUGj8NXMEIhZ9eqRntUvReM4OeOI
egt5JaTyWc1RYTa0bS8fWNhKFKTvR+jCWWvTZaTCBV8q2B30kXcgJZ0TTmXnYSv60GiZlYooyl1i
xuvhG8T3Y90yoeVCD6cW/6YzvZdwTEOT+rjmZFswOr99f1eM2JcJtHRSAxeouwDZAqjpwsYekpdZ
6vRo/p7N/m3317HDhHzgICTCPq7W0inPEnBDFJGXVQM8bNp0wfFGpZgyv9E/E6wSlnFbiFeX5Qaj
NdcsccLTPYjd5HX74RHrLtSFhmjYKxdgtdOxpnYgvYeKVLAfcf/MCFqSrP7tff6U25U0rDHDRYyZ
gMlMLYdXGaMCMc5D7IURScXV2+e375PUvooGPWI8aatgFD9lpx+0qk+j+hjR4PnMXZOZCuWjy3of
1qSZooUnA0gxEjRFbzkaa3B9OLo0ZDVhsiS7z6CXQi20HFLtyobdNWo1W3EWdm5zXNC4LKdss3+o
Y1787QoBpccIks08aL5dednOWCzP94w3i7A9DbBZQYnnt0DYNKU2bopuPmnecw8qHDzPEURvwcOd
9H1GoRg6HCer1xPgJVzlscjYiZxxeylA6pqMIm0MjLP53SBapU/QbqnPbnIcZlkdalgNdmzq7U5h
JGRmkkuM+QqWMqPE5RkDQ/9aWvjU9uiPBFgZd1vFqygdRvwUvrPMfOxd7pkzPGcOTxGMPcSxA2bN
sHIEPYfZAhVidA67FvgEiZMfBAHiXg6puLLwzc3FhkA+2qZXD/IAX8w8yS3P4/UKJjcPlnHr9xjk
YZ2bFri4WS61948F6WOkKr1Ridee7quhYP5+LOnOGlZkGbD5MUFqe148Ks1goN5jRq8CssJsh6Jv
gmYk8C8EpnLODY6H5i6dPQPcl4VhUFRUAnRT7cAnjDDX+4CoUaHp7LnXE0Dcc49Pmm4NafR5IIRR
qDSDsM0AtmU/9OTCLfTkvemTIyrMkOTUNv0WGALXy7MQ67DZ/Y7/7BwFVGKaCou7il6jsLu3mgnh
+G3xtwuEbMUM0LRnHjSBESqAc0fKoMawIAAESf5kfVQ9pzKtY3J7YGblX5GBypaUk1T27MzqKeKN
XlQe7hCIzx/YuFziCPsW76YacVL96jr76VXEATiv5CeArlA4wPXdV09IdcfTFG+xqjkUGx0WQW9T
IBCnB9+FeJ5v+Ajj4tZx/Ex45EbPZgUIb8IpuWvoNl0Rq43zUv7c3XM8jvW5HzkKNINHJL6QV6ok
5yX5z8kmPY2s78ii6tcNBVcjTwsk0MU2fx+H2cmg3G1Nd7VEV1/D+gNE+Ssp5HVuKXiBghxNXE1x
C6ofbkDi7ZASq5jbpW2ZcNT0UNrOY6s4GJrtbADrWfqB79ocFWiReIOM0qWnu+9bLidqiFbmSN4f
cZsYvBw8p2OpkM4f7SlorN+ZWwnE6h1ca9fcv6odwxevOmOoTXQmXxqbkyhT71gQDRkQ6uO56xJ/
Qm76e4+6hcNqKJiLyqHFrck7ZpwLmVxXwQJq1kYqNIvynYTbg6Vl5hBePyxlndOx7mrJoq/hSE0B
lSj5qG1T92Pj6co5mg5eD48yi5XbevQFgyQTD2lMxOg9M9qtrMuGy25Ea5FQiojTKYvSTzQf4Q/5
mlXu4BTWo4u4s0im/GeMkhZtO0s2jofWK1SrFBQYSk48FRw1vktAkZWOJ8hTaLn9LUlhGHDltNph
bTrSZyHOnqEXfHMQAXkmEjRuanaGDJoODGHtmSEV0KUnD/s7nttRs35RN6CF2qSjUeb9haQRVZeN
14Nn9BuI03JwT+9W+wIn354WGRkq+9+2CSbUhIT5QTtpTlAQeMicsRaID+SteeVAjKfgOQzJeBJp
NwaNstFroNUmzUT8eYOyU+YjGm+YLkOT7nJECf038Itxszgy/rFBBfbM44SRd/4zINywGhDJSgye
Sx+jCGxCi3a8DyF1505016jlNmSMAudp8qgn9CzEQd6cnbct7UVRullq3COk1TvRgcrYdwhQxdTw
Ze9plKLxp3VbTcoCxUll9F6T5sGjmfXHaYmmo6MNeL317lDIsYQBJB7Ry9AvX8eoy7nvajIRDNFW
nClJ4vTcloX/GgONZaYYQrHGRJpSrxAk46vxfzg09cFHUN681nIrbdgvs4ggxkUgqQ435skUurYq
ze8IAAPqDTjcExB1jthWKoFYrX8sWSdCWqDsA7Zbke62x0c76mrPg53LW+tyGrGmYz/cPmk68G8S
pNaORaqyf0Q4hK3DFuL2kZ5qLrzaXAZQJs2877poQd+HKJHcmgaCmTGXDHcrFZXABhuVDnZJLOFs
zagB4Tt944Gp5k7xdhNtldqcp/bE0iIU5eRgH62ouSOvU2xEi09nQyQFRguHtp+mUoKb1UkJGO7a
qclH0BbV7mj6ii2x4rgKoltYgbmsgryYwMYW4CijKBvgT8uZOrokg+vfdwuQVHzoWDysZGEFez0C
AU4RTChGpbItgeWVFw1VPqeN5kvisAkg6Zb88gGCLgh8En+RvIo4y9jBh5WXm6/35sDkZlETkbwz
kLUqYItmrWp32lNPCV6YQcliuS8BAJ8IOUSNdJmNUnF3fRsneq4dJNzYakKW8eg2io4hs2mU7U6v
G79tdGKUa3aEeiAw2w7zQN3kuPXvLyKlf2z0fX1pIzCaJ0Fs+zWktZMCPezJeY4xjTtWk/kRy2wf
To3GeFKoWgfi+YMKLi0nKPK9Q58wRYwHyKEhKYL9IRXqn8OFDqLyVWt6jA4eg7/ZJqupF1mLJg4j
t6kYtxMJ07DtYvq6pTc+7a4JYegqnekGuOH02Yd/JNYmLHAi9ggmueldATHxpz58zngV0zbw3Sry
Ey0zcwCu0RbQYCVREIW+yceH3wQlyUazl1/fK9lhZhd2cFOd17pZVpGZAI9dQPA77PWM7SWm0l6l
TNUMX1zElaY8boQsyS+eLbwsbqMD1MFpvG04Ut9u9kYKz6sPyXTMZET/2roRN2MO5CgladrmQlTm
qGNJ+h4bKcbXh7b2qN/2M6onKdX3TZMY+HTzLBDb+UbjbF2kWUTrNHRfPlKRWs6pMOBfm9Ji3t77
bTrucwQPasnhWvIhK04vaAoH3VL+U60LsG3CZkAaeQpN8QeRNU+zzhJRsYhIXyw++ipwnkvBwdTC
sAHyMcu4pdrHvY3obEoDb56SnUgnxAT7pIfMFgc4Q9qa7be+vpGq6PjPerCiHdspF55Vr4EvXTtR
Wkx80f+PtiqarVrTgoqldmIWsnPcvzmm3wtJModxx0/CAIcmIJVTJ0Qfuw4+hVz0JFVjLJDU0x8d
9TIeoLXqYznB6fpcfYIDs42nWVAN+zpRrwAbZj1T/BQD2/7LL8CbnZ6kqCrYgOkq+lgMFuIyaQlK
1xLRo4Vyan/6tU4a6T60OKQmRJYT0agwKhAPV5MXmJF/0UuEmaZ/OTP62n4fZ0IWZ3hyVWPkSjS9
xZ1UI8IRwMc1u+j+7mt/cR41DUcJbZfTK5Cwl8dFJH6OFN5QERuX1Cq/V3zlu9eH54j/4oQkamDT
lKxhAA4MKh3qog6FZOiDSnb5MqTtqe0Ltq52cuAwrKg6S7BPUFG0iqcfXRs6Ts/OA0uLcDW32Yjl
AKze7WJkOWimn0MfTno2kti0OrBmfxGv1CLMzBBANR0uF6wc1kraHSD4NsPhWAlsVVnahtyA/tuE
W6UIMWj/1GIx6g8qTmOXOfx2/i3ZEq6DTzdJwHpV6oTnYom2ABTVFPOdmSKyHA+Xq0AJz0EMTMQo
Q8G8f6q4gAJTrC9h+N9RrpL1mCPdhJYmN0coud+bkkqxMSiKmbG532DKjfyORXy90N+gMmKVhHpk
qeDhUJ4usiDheRHQ7srgUPp9NqThGkxb4ECLtD/EnnnJl1DdfyIlxq2LCZq5RoRjqscmEud7EbAD
MtQYKbCadQzQItmU05ZNasasvtZE41qN5hLDcWLkUW9AiFnmgmfCHK2LfDOxxAfJ/0YK4r16d7aK
Lblham9kO3YHGHj9RjXGX8nDYC/nHDhhDGt9QcSgPX/SoNtEvvnzMxtRQM4Zm9zSpv/jsvxrGK5+
snOdi7PfdB2ydsXEK+veII9XwKzySu23ruWRiTRQ0sYnHFr0Xg8aqc+Hie94jliQc0Z27+a4+kLB
09WxsZwAC5qOGqi0va07J4zT0OKCbXDMq4nma0Igmmg6n5JEKT+aqKBUB60vHmReaQaWc5JCt4Zq
cxWgjc58IbjbkbKuc+50yGutjzemm9wvRshTOiZFhRJHDGL4rIBqo+cUFD8Gs/xAr1wbZ8/1aPMf
LdtKzPWcI5qTfVzjDi+l8Szt4v2UuL8/2AMjMUb6FB2SxLluKIrtyNYY3c4Bn5Y+gpxXDHHgco+a
ICV06jHQMJc9XLLeMCEF6JKjOjQVQyof0UtVKzso361ERcSq3CjwN8fjm+Glxpv04OT7NGr/3g3A
MNvbM7FDCmKZU9cyJX7n5j6qQ7qp3HOBYuDrC19i6hdrsvwytQQ6zPbUNO3YAhMdbMFtmZA1l26l
huPgvW4ur+df4NZxK7LFV1HCltfP3zSIhnKsgScP+nbFQSVPIczKXjVImEmvB6beT8aCmD2lRmi9
fj0uH38rB6YbHpWgBwtpGw8Xu9LW3HmkFBLWp7LWguZqPSpsidQMKSsCDupG0VM4BGMnu2LF1mZG
NnSIZ+HdNg4GgAiwUvDfA5yyo4yUNSg1iOtxY86NXP28OXB3EhM1rG2q7JdUVCtaR9bJlAoKkVZD
OtwJXCeSQaRXUtwqBkKs937Xyw8TOnANrngOiMaTfSULNcTyI7t4NqeUxpHGJ3oXLOA9RJYhk3eh
3jVIFWgpWyVpSEcYEh7dK8UO4nAiAQFns3kDnyGiOerNgFKF3GT7ZQJgCTvfcwfzvvgxiSsMqMs6
bWgnAVj0PJnKionBd61IQSV54F+cUIQe6oorPoCDCV/MbxhbTFgc3SwuXOggSJOE5F6guWSrzDu8
t7i0Bs8uNiwFdwBaQq+ps9BDWeDo9eWajwNBEgL5sTEpU63CCvzolA0pU4kzGFipI4jh6Pff3CNh
3Sm7uxvZ3rG8r5M7ODzb2YqDIyFYvBZqId5fsdf1t4JxhjwWDb5Qutq7gDW+knQi8J51WGfQhmo5
sIASLoKiqvs+fw3OqjlLzAL+fZMYWPVkMq8vVKoNRIl+TknlJx3gGL9j5ZYmxiQtInA2+CHgnvtA
48JeSeY/trVBcp0rCqsmc7OHrlDLnkOXvPhMf7N1kKFMsh/hL+e7aM25a7uAMerdkKXvvjCTmU25
OrKQUL7Pqn/MIileYqRkQ8skdTefs5jEqBVC3XOvcF7RPRanNi+g9lLrh+m+dPp2oQ9gCM4JLj25
7CJ2UOUYNdx/DBhSTVJUFUhxM6LS/GLLU9ATgPutIIstF1Bs2pqBtPfUxtllW7s+IlI/TBC0sCwF
+QXzwrxhCVudfiuT022TNgaA5800mnImHmtaegB2vzusjaM3x0kdR8uRhWp4rinGsSH/3AlLgzpV
cBEjbsh6sYUZ/DhTiYq7+rKZB4pRG4c7+Yaf81C74cW82DEHH2QIahwy168qebDDdDYSpfUT7ITY
vLTQKfl6tDxuhn1nFuGOSDD4NQGF3TU4h6Wln4prP+uHvqL7FG3K140A/EAIuQ4t3S1KKieX6H8M
s5kob8gx3efqSo49D1y6UsBznjlnQ6kPOqxC40beOJND9FqE40ciATQ0J54ZU3FmeOs+UOxtuwu2
SAbY+SB/mH+s/10pU2s7cJO3pgSQS6H/SoUC2bNsurusjcR2tL2SrBqoTsOFmRx3EglzXiqkYIss
i+WEOGRlxr2k+jsEyF1vXJA162eRswZDTqLoYmn2mxioaCJvnCWLvqcHhcMqL1EFeQbZrqq+WXKw
NVE6ecAMP3I7gGM4d1DRHvUcODo2IiWUcz7kM3o+FCkNHFS9PXlW1AuBUNIPZOSU3hd2PI6wKi75
krAR6Z5vPFfOc/MLYGj6RXXVd3TjJJLYB3OUIW+FkmWy8CbzYlNL8xbow/HzvbjOpioFy6AvPhEk
fWzaXYkdNv22wjgd3pZdkrfpcXd26pwss9eu6naKqsdCAOqpmvMzW7SrrZKch/EAUKpFTfkRisRj
FHEoZzzCcOx79i246inoRY5rSATrAgI5ymdRttD2okLClijWjvRRr8hFl0olSg46Pg39ezC26ftk
hStcBXuUlUwPPgfQzJyy9HsQadqurT2Gmtb+ztOs/o262+Gm3HB29lypDEulG4MlOmJPUumgooCS
da+YX+/s5lJfnccyzk735KzG43zPAexYGy7mkZr9JVILeDeQTUUL2lNG4PxY8MFfvn7pLZjjsrnv
n/1Y6vXhP3PijtF9rjqBigPYf38K4kKMltD8io8WjcXDWrDyjI3hi7U5edC8aBIAqm3MZjZoem2Q
mkqiBWxYhXBbj3q45Np//mPw/nAVaHLFpJfU/CrKDUC9iNB2zxHi3c/DTXfCOwugIYjoEt8cz5jM
jcrSFGwpq6m5AXXuz8z5OyYCACdHmwgvmfF4y6jiB1O+p/21YVWstHfP9pMKJ5yPWVBCvuxLBPpP
0Jrde4tQtpFLDuw/Lg5EpI4GMIxxj4/f3U1RlkHkDqAVaAlsaFWCwaug3KlYHK77yZjDQsfdfau2
wout7HfZO0H9Un0tW0LawNnG1pMVL4Snky1B4UAV44KRp6if2Xdi0jGqaR51GPa6nxfsJ5gRrIVK
BA+IcRTVz2+KB6DqTjjhwXO4mWeCckblFSgXwS4hfYxTZccapB1StqEH+aYC4p+q2gG51GI6RTPG
VzAsNrmtYmPxsaOSgGBsRhkLPtM+WFLRsdXy1rRCPF/QOkFzVuKRpUdlUt9Fp2rrhmk3saqPrJr6
dzTvrcWlqdegi/jjOsXNR5/QXZ2cctMFIgB0Idq+NSkI0lclmo88VY/hskazEu8fDNnflR3d7ueX
1J9R1W5wLEUVESGU+at5YUGhs/6LyZRrh7JEwOP/085sClSX0hXxg0ZzMbISzyFqzmp2mBna/11f
9sawa6RQc3I+TeRWOXvyoERGbtUy+mqYxFYku/dWHDLvIfqs3OS1S1SREWlgJm1VoCHm8yWLjQhm
5iBg4QB0O2cX4xacnCCTqY1Ivr8jhaS4eI9DKRFCgaenntWPCDQErjs9PF4nI4RDX2eI1SGM/4q/
lwCvcB4xGwDACH36ymohc7qnQn7ADYVh0KLSCJFw212vnp3Nm1WOP6egVtiGXPpy2NmWdQvpvQpG
CxO9Wr9QI0eijifM84YCazf9kpEs7BIZauIQVtatMjKT1lauCiu53rmXxo/1tDnUigEpt+sv8lX2
RmaVCoAWcIwh2cQaWXJhGRABhCzyK1gJbkVc8BiS5fCw2duvtyGUtj7A7ROjL7TstN3hEkow3qU0
Gryyg3qiOMyXu1dOjqXGWeJUl9Z/UUq0kkWrCOayIJ65Zeyd4TPS0JmV8ajbxAKRH4QjIl/CbCGr
Be4U5AYXmtFafFJE7/7Jd8/DaPPzg9p21GsusUehG2KP5ZP+mBcSjyzAyMxKV5x8tH2Oz1H1UKF9
AIeLuoVyRSIP/6Q1jqFpJEwVrcGsflDWr9yTyR8bSPKxSUamF5lTHKC6z6zR7y8XsGbbAHGP0M/E
LB5r/gW5r/6gIIiV4t0+fKh69EwAGpaFdRpQRtmr+G6ixrAdUWIVHQBr8wPuX+lP3k4zNlpRzdVY
+csCbp1XrCpEC8myg4Ni/1fEsrqvhhTz1ZYFjRTqUIcKUN4SoDXAbxKfQKzuBJklrgM9VRSO9vuv
b1alVG7IkpCcuJZwhdr7LEHqcjL6od6FR74vBgL3RnB/sL3ORNG4lsxpwn9UgbYgMsamyj6u/gSJ
WvT7lBmvRFpqOhWW3FZBrMjCW74bs7NaprTp4m74aVYeXHlpxTnpD7p4cMOzxk61p4bke7t+mbkm
cJYIan2JbbAygYkGBwASz/6mBnSTXwwwWQg30fK8e0pPWzH7WxaZLJoR2PeN6n0G9EuKa3xulD/x
2IUVZNplA3uj0Tdu+YhnyF4JZUgI+xv3y3rdppQqGPTq/N7ryWQSU56DMi99SSL8RzlFEsxuQ+KS
MQsdnwhfopyNasTAE2ga2E/v7PDpwSt0ptXmY8J133OFAe63MILzGUBhE0stFGMmySkZcwPMnL/x
S5AmC1IH4KULvqIfzstD9gxMzKTVMLjPNEMVIKZU+QYL1l+P+nhH3YiP/aioRu3kCDocmqLiIemm
DFQueeSkflaSYuhVX60LdxA7xqdo+MdOmLqmlO6J9mcHLwu75DwRV8Kn1XUavM7yncdg9V5m/OYg
KmgQQF51PPVb/Jh+DO8bWo64i56DrCNBSI/XasOK4g2SlsorJr1mzGc3o4NVtWmm9ICDodLdXZS6
haASyor2DWhx9ZJ80AZw9KJ4zgkK0bCHSXfrTwTjJOMRnx4UD86nVfgwT61XY1V1acY6VVPacvya
PAKJgZv4+VPVgJqWs9L7DpIZbvKPiK2ot46b47bS7z+SHzQc40E6rddlNYMQavLMNM6CbvLiD6mW
tPVkzqRcudw9aj5M1tWP1v1vE5rAR5QYJRQsDlnjX0U26CDYTzEfeHmWZeuyy9rATVtUQ1MTYM2L
dn2DrCrzndFa3kTekq8xIjCVcQcFeiVjzeDkB13l2I9nwxP2WXgGAgLgaNb9L44qnBEAwX39tmg4
tyGMvQbEkctYH9Gklz98XLE+TpSMdKNChpczu3bzKYSjzMB5p+kZ7wh+JvryIjb/GPQfm1R2Z50Z
90xDZglR/oEOp63MTCiDLkQ4PAHj7hla2uEsLaSWKijeJnQoVzvn25ZZBZznzuiBGV7teS48fvch
lOyMaoFE2GRFit31YT7IliYOE8wc4wK6nY3LgOQBDEFkvwftLGgMnADAUeJ9cU1Uo3V3JTUPikna
/82GZAkQiXLdbivgYjaaW1Lkgez++agRgj9IE43cvabs7v3FOabVPNKamAJrDZXT81jiuyK2uUnR
BABihMeNze3mmm4svYw2WPDVaxQi0UlRM5ccmu1OZ5rwblLy47Oxd8B4PGhGdaAgWZUerdqm0bs2
9f9HWAtpO5pls+k+/T2NHxtOVCqjfHsNnqkBObks23lrKz6RkTyCVwEN8VOG5IPmdcg7ep+yHpRO
JScRwfvWLtLqum+yy1v+qSVolSQvNtsN5rxDJm1KGEZFGcH+kgGlpGW5tXbWIQ4wYBeu7PJKHFXb
+4+z3wWbq4MdJ4Q8ofXfUEbtyqdd8bKPVsJb3Vh4qceEA/i1XqTeVmuCik/pROxbrXx3pfe5ERGE
Aori944vGISVs2lDbBrd/XM08vJYltGyzXfcVueFLNWqbUv4qyN7f7NoFOgx0cck3WxXJXTYq5UO
WWCmHn9lryVMIt8a977L9h2nMVNUmItDqWfCtdJjZZpBHA29ycLzBJyTDJg2wnNj8CRK7yn4UTYE
J2djKdSZoLEBc63jdboOfEJLUBGh4uHfTYUgdp6tschvYVRpQODh+A3x23p0qyKBW8c0PyCT08fF
n+i5Uk6bQ3pFhj/trcAKHlI9tRR1/gCnvMCLihwk1C7kXRwYeuJRECsQgC9LcDUcQugGWrdKQXpd
Um3hKeS9o72Jzolv40si5fRh1rXcuNI9BYL6viAajR1KXo66QmF3ULe9qn3GVOhIeI8C6uPnJF8W
Jvz6M0v8p18acmHBT9GfP5AY3jkSIYzTGZhqJj0msTfy4+26VYRSeGewSsUvytQfypp27OWHIL2o
U58uxpL1gGms3BQYFcAPRsFzpOL40OxvpZiPMQYjstQo/CLQIa7qaQK0DAfVGAB72mH4qIY88Esf
bOSb32OQi4x9+6QvUl2qVan/ccN6GdFVVRiFkYGvCHYl2zED05X+crFzV9jBPJoiCwxRWRN+A85c
C3vT0mLyJhPejbF+HQWix4r3iGVRQPyazoGviUd7L0hxO/ut/T+PR3VZq1hkL4wc6HABXN5rCLjU
CIDtbGAv8bEGEVvuMg81aYBbxsoiLDrexqH8Fjq4g8lxfVA+Jq08OL/E9yte2hxj98T4Ri+1dK25
1fuRx6AxMLi8+CtD7OEaTOQ/6VRWz0PIxGJTiPlr4WdQj32DiReY5GapcipD6tuxl2gsj8LmV3KL
l+O/8oG9ndJLrn1TetGxI2mUM66M3EFqePCYw1ZxT6Ub0GSST46YpX6LmNTTBR9v0lPwzuU4FukQ
QMewmdF/4a1a+L7Zv9qQwA2UQLHbDraBtfXdDw1Xw27fLFUI7ygJ7l529u6i+H8DhgV953ya0TrV
IMXhPx2y5TXlDExW3BpoB5SLL2VpGPJF/e01j4AfEjb2kgt1Y/Ou/aMgfHbujDhuTo6UjHaEOHuV
kUkIaczK7HQ3zSIFRTSllQaLr6wGqclN5J2klkLzccftASTiVc4Fis6BqreH6z+qH0QpqHhO/V7Q
Yceje8pgDZqSN+660T/ZlImVWcB9jwJpDXJn7Hg1wHuYiUlb/akB2pZ2TbKZEhwYezQ/xEZ09nJa
ltdAsltudBT5kEi6uSLSrIizat34PRPwhzifCtpHSv3t/bdLJl/2wllC7+i1+8d6icIz6SogY2Fz
ihUU+VLTDTIiIkE0X8iBLEAc83Wn+jkfjewf0HG5ZCP3KOGn4pIqn6KDhJALjzP2tS4/QPLDTq8r
a1yKCfbYU2Ecbfvzv5YJNnAbMImDiVG2/GMUUGmd76qJm+gwDn9CK4OjvLmKRphg+eUIrMs0Um/y
xkY6KDN4Pi22BLV8QhGp4iGrNqak67vVLqU6qAmUPSOEGy9ePRlT5p9kTOrXrpdfkDvbgF+qviBe
ba3B078qjbwxiyYcFRqn+gidC76BiJEcCcWVUHVjCAT61mV6C59ZCJ7dgeEeLwS6I+ZKGztnv1xV
huI80nA7/BDS17Y/8gI7fpg2tCERCKVHAOvDbSOvLqm+dcl5E0ASoj4iSbGTSLdaR7tL3pSz512J
g1DL2ZR3/hDPsBsScnPT2W9spxqtUX13KM5WIVcdwJ0imrs66gyA4u+abpgLs2WaHULjdrAcytVs
BmFev/R20gtNcITxB/u2dAuPW+cGeDKcVpGECsruixE7dKo/1x629CMSOfc6qTlelN38j4QWGM67
7lNLy47jaQJUBVKDqie0TUZNzm2iFbjK+/ZwDCd/WgLioP484EC/KvEJc3TSiWLFXb9rggo1FrNj
yefkEI3i69oNeo7z+aLqUTuJQbr/T/zoIdNOrVARoe9jYDPAAFmJAwY+zQLAYQpG5od/nmK4Xqxm
sJdwmVfeOTOAfWvz0UAi0oZYBlQfYVZvnYt0KScSliXhPx70VRrlfMpwrIi29Xcki1rwt4miEa1j
n6h6mYQDE4B8Ejr3FT/NxAShYr1LTn9+cssuKSU2K3iJkgp0+PgZkaVvmrmV03GFskd5BFcVTWIi
Fjn6eQEOAtJ4LBK0Fr6yHbmDImYdNf1ZWPvQsAov/kEOTTgTW/qSuJDNLv0rvRrwQPFpBy2ySgwV
1h5E23eVNSNUIcL4XokUA42oxzkTiAtWIhGdikEMZ5VqEh594vyZQMW4Dyw2x1ekaQqolvkrDBmg
vXAUhGohqcUX2XhfanTPfLLVYp7LSFjD3lZ2ucGCky9goKOZ+rN1OxVLu29oKewNirZHGSPBeLMI
yj/zmmnfQPzLP1YRLFehX82tPNZ7xSAY+YQQhWPcQJC+3wA7PP5MfZb1JplWbcgL7cc+qdE0g5/A
haHuXAn3M+ddGtscVeVeVvYrTTFvDypqeIU/pKYvkaj47jm0GWPJXCXtT+q2+1f0+/41wodlWhWc
EbycSmRN0M2bFuK3oLTFTIOGfSJnK52CV1X4OvXZiMMsWVuvrVUgYPL/wY8gzADWGVIkXj0O+cmH
LhZ05kVKePyLRXT+r6VRIVv7WdOJXJ78N7SUuXVjpJzCMEn9IVCy+rPwpsV5KmX7j7crR7VtroJ+
Fjj/fEs/3VxOyFjIH6NRgelyLSl3grQViwaZyNCleFC+MhBRHt3Si2Lj+P6HC2557X0x2JRHrWfL
bp1yT0vbV09xbuwKXPbJ5QeukMxOvNeXTdya5MajyvMmd4A2Dtt5DM8ExGemocKb4KgolZQIPUPn
nLL7BSp8zX2mp3/1pPzaXJtqs5DBLdlNigxnpsT+NCe/C8OAkFJ3X/1GI5pcOU1l88UskLszw7lU
Zam9NXWhupWe5ajbz53elPPHvFBqg7zPLJxwPwLh5DGbjRaXXL9tEUurMyi9Ez1mH08xRXQ6+BYQ
N7Rx7b3wrk7vspvaYJyPZONfZOtVw5BJIxaTYkE86/pvgtV0kvJvBPoKsc83vfkNmVRSvyPVFidh
SPaisieQTxNGfiRlEW5YRwqtmxQLi5+r2J2LNi6AK01Mk4kiiciJ1OZJkEW5MbWZ8wgFfx38Zmfe
5G+D0lcfvFs3izK3ALMvmKksPqCHEzyg6cgqz0EopHMQheaiFCFe63F6pSnfOWB6t8FxFmLJo8SZ
wQPzYqhSKnCMJ5S2AG85F9VPljBV1OBQrNU39UwYegDMbxNWz60bRajz+i3a4rnwZVzSNUrvczX8
EDaRTkO7wD2/e9dJenDreKst3k9p5Tgd8c8Y2w+QSm0qn26ihMQNiDrEvM+U65HOiTRCssbEkp+W
KZyZIyE0DWActQMdNj2AoZ+AZjRX82GTY8sW7JZSo4QLwRAhhDcpoHtMONIrAiWwTxk12tKSAT0s
ypWSGdc78ELfwHJ2MCBOhZ72GJIepS/nqcfFR7w/HD3vGtmnCv87j2RH4Y9XxfcgfEFm3+/GqDvP
spIIVG13BwuNFB+4JO3G8sZv3WMmfPZHulpjazZkjkGCL8qdbywKZdMlYzwk+0/GUCmgJsaFQsTP
+ko8RleaeVRUVTugx+4Bi6Yu6vbqcS2KrroYskON/5W9xfg7hKzLAmgxt7j5X3zlaHvgSObZaX1E
UXtzTzcR1fBvC4xOEKE+kgKXh1Sjrt/ktanZ9GWFz3OhFWPiMvi4GegvoLy7cDY+agmNrJI2Q3Ea
f9syrSYv2HaxYwRWOwSpamTc8Hm7Znu5N+HyLq/XMyTHGGNgoVVm0g7QqdZ/jIXLrLPt6ZG2v8Ls
qkmJ8ds7SAKgcqoddrfhYOLoUFQUDeY8lmLINpn/5b34m+GKtFniDtMWpICLTOUlHgV1RG2Roltd
2uFqZg87vVurgeI8h0GTLVtk5rqbFHhTmq4ZMk8I6GFzdYub8R8+BpN92qosethzCtYjTmxdD56K
WKAgvmoc+w/bQ6eu69nA2uy5vFerfFmMWsn9G4jyCqUtJiTOR9OSOQFECOjtzcvvkb6GmKk6NYqD
u1Eo2t7RW0bwO7IkEME+P7FE4iQaTC8g+EkQ2vsSPXDEV7sWdmLBOcf3bs42xUM+jqo3yk9wTf7b
WYzWxI5lfYlnZ/RaBy53MdPYOkN5BaNXQx0w745FVplrcVL11Fxf5TnME84o4eHBRb61vm9MhTXD
2ubN0Exd+LtTeVOvHKcWz/QAZ/tfyfu0a1zhx1LnFRWMGcin43VILXGmY2j2Z9ApimroMruOj+1A
X2hJKRsZLUB88ydwByQsaG5UDiQI3pwmf10rgsNybUilYuMRPyNgSRH0iqolO18X+yYcQ1i0hDTo
uFXCxdftriKICJ4wPk0BeE17nJlT6+dx2L76jNbVHMDL36pLE6WFq9LAGGXFleSq32xNOS1sqfnL
Q1TzTzZQ3/SFxtNq8LEo9urE7HWdzsiXyBROJk2HNEOGcE24IKcbEmZF6kpzV2djW3ZF6yeE4ISG
TjS3Z25GINIes9TKbO+NnHAfuOBMmwSC5sQPk0MH37mFr+Gc+G6tXBYTAxmOhIUYxLh0f9V9mNuI
hmmnCTXogeYwLAVJMmhy/0oE0EUxC8e3+fmyr4iCdHPxjmcCVaDVmxcoFsy9OwurQi98P03vmSwo
RKV6c7GLueycjZNKlDhEbqI/V4I4h7l0tYKoxLwTcxPss8KmZEJgmZPzDVnBCLfky7dgP23qBXIW
Yfb9XpJPc+0sCqZXyfa8Xu9U8iloUg0gPPJUkBiwnOn4EAAaEssKe5iBh9bVsnT/E8KVmLZvG8/K
RujzHYBm488MRT0jd5tRlZcs+g1Guj4vohlUetlYeIlOC93YiWe3K57+iXaxd7vy7uoNadYxb7G1
tTZ5EA8NX3ufav0tGZfLXfqXlFufGl2g5P2nemUH0ynRSdfEOkcHqKvVqY07mkv+PT/BCgHyPV4m
bqpyZvIzP6w7ui4f1HIQeJUVdUMA9tFHz9ob7pXEeiPZYRZQ9wzLKE8afyZx0bZd0sT9S/2kX6a8
Gyp5TiRmz7bpN9Lqum1vNpRsWShWrX1jhzUpkzaad7YT0yth/HCcfBe4UCzzDK6IGm3AJJ59gKBi
zzYeVtbsfLYlrGRCQMoNpcse0+wFc1MSMJtv5hu2I+MveCHEAxqrKog9l7mixSPMmsa6QrremnOR
4okuVD2t9FAlpQUreDURX1QJqYvot08kgMXUQi2/DUpbEvo3gEt6vhNwfof4PbFbwrlvZZdzJO4N
SqI0ypOOyWoo7Dz96n8iqthjtt8x5mcmKnGrYT0ju7CiWG/dYgbdk5i/Y0CQ6yXMYp5Y9cptxo3L
eOIOsCop4kqB2di8SaRPDV8w2LFvIb89sXYoM6M7O38//HbMyxB6RvuVxPjsOvDlFpRQM/HG9FrT
dF1J3V3vfoa4rCjAvFSmDUGFb6ueY/A9tJpVUWeqzqIgjqBroQipBvaUw9+6aoKNepW0xmKWha2p
4afQvM7DkmAYcgv4IwVkLSuSqBTpa+tKwuO87Ka2uiEKeJIUy+zd8/WzbVxjbhwDOLA7UKr24iCu
lVWLNR5uicBKwuuzJFEb6mwnK4cB07c9Jqe7w39EkYCMVI5R4r0yydOJ5GJtmQUazJPzaIOpCSua
nEOwsuPxOcVViYqu9UY7No7MBUZMTF7oyr7aPoA58yxdEWqOYlYY6419MasMGCMLOqgy6G53g3RD
0RxLK6lWSZoUroyU5cWIH3AFIbgYK6S8ZwxpSZbclZuPEkBFLIwHjwMpdGH1VyF/ycW7ypqPPdNK
xWnTjePDi13TxrgWj1gl4YetQIA5a2rD+k+CV7xS8UWI93/OzMhT1YWNnOnTMiKBG9UWypKWnzeT
qSswVKbdci19kYYgkBf+GM+jUb7A9htMWi0oYdllgRyh10P3Vqd2Oi6x4DH1JASDjOv6hRC++TYL
PTMasVJXOEJXkYbprgbdkOFdVoVu4we0VCgXSI5qpUjX+X2VTMcXOpSlbm4Rm4WIgcGo5XAytnsu
8em+STrnwWgWIiqiHWVlmjWelhpvZ6wtdvDfWYeywcOR0BR7kUCL/grQqT02WI+g4pfRWNlamAs4
XUuYsrmJAQVKZ2GgWKPpJBktElAflEjPRXt15ARtIPx7Jbehj2vawem+/GQtveI/Z1fz5NiCo0vW
w6dwt4aorw89UkocPQs1C7Gxot2b4loka/5Y/NNA80NJ++s2Y25J7KNdPKfpAHGzbko3fpyZTxB4
lBiYZxKUTws9v/fK5UgnWXU/LXOmmH4nPrt3VxobfaAEksNgb/mayvRZEWDdeCywjKJmVeA82Jze
bRVUEmK4jbBPwQ5PZQhHR6mG2YDYTGOBCaf0YshHr2ci94jkyQ+w/crl9adUHtcr1s7tgTe9gZr2
UYiQ0sWoEzYhiBNXDpyHcSYeRBaCl9pw6Cpo7WcsaM/taw78R3FGtnFopimu4Aw8IxLJzunUirgo
1aaQ0rsc8uJjuAXYvtaCP/hrre/Z4x2Y3zkLGCCa9upCKq5lVwrAcBOPX/CZSbwf12Q9c6CDsfTt
IO99YXttX6pJdIlscVO+apLEMG6X0WgU+bG003cciKzk8cMMxVhn8P48a/3kbJ9uxEW9+VChSXem
diwxaXcHT9HkW2hjsmX/v+hsyfapKugVp8p4DNwy4mBZt2Zfq04mbqQnAlaR7H3PlzfsV4eNGPVr
4HY0M/fhvOe9Gm7DDYjtzbpJMU5jMI9n1Dp1773jjjn+CKnPjyhLmPPuSz9HdBLOxGYk86B25vGI
9XiI3JMKGWD90Yq33Htc7+Fewcpm1Y7K0eel/lB5+2UawnpE3JmSxxSxBY4qgFxrXxY8738vscJ5
xNNFT/igdx2dRx9mgCAJaiVtfyCNmUF054/LRHAdWjeX1Xcfh/I9R88jLk4Wfpp22GfE6Rr0FUZ9
pxyEjysWtlEvdbj1G0KyOF8D5Oaz/RyqhSczj5lxqtoSTDy/SQ8fFD+9Bf0OyOzBJ0YCJBDdYoT+
8gVeyeFL/Hc/rUjLmD+2RCrQraJCOKS3TCTiOxFd+ckgYHL2LVSVuVUBybdcrBOcccjwj7s11F1K
vLwo6YAa52/NREH5773cPmcJY/tALtmx8tifA9f25pLxXFsp6aPvrD61kDkJVJg/FiyjRemTMa72
JMZO7hyjSzBQ6KzliN6s/vF+i44ZeV/pkB1x77U0NLEwg8w7e2ycV5U86FIpRWRiBQUh6Ndh/Qad
ECW3WIXgdaDAZmzvXy7yKDJrP7CJ5mDwTRKTlDLxkBmSP+0WW25nlmhOUm2kGDhYJi4J/mEz9hYk
Zom52Iidd4YWI9awrrf6t6s0MuNUUCUDxW5sqeC9vn5DkeXPtjlywpQaCJ+1w3yLBuEw983KZ4ks
3tJY4PN2Aeyu3b5rp40TYwiguEkRHv1Ro36RI1Lsc2xADdv9IS/WL2e7sw2ZmS+qEEe6THGInRXo
Pe7UGcOtSog4eZS0oEV+nnOANdP0d6WeE4aNY/68VqmqA/STL/xe68a1PZ4ipWqj2nQcKnDD0soX
HnAfJJ7BXOCWtjBq9UpPpnB61L9mnW9AjOy/GIlCaJfAh5wir64kI50x5J55er+kPWMTpupcVW3a
Yy8IXaspxGvMnT4532nfRJQoAgupnftBob7p+mmFa7eRuCIxY7OtmRgDoSXXT/hChy9aUbduhN8Y
hO25L/Vz1Z5MJDuvnVJi9G1LrMKh/NKWISBgOF7nGhPAvRGuLx+Kv0CG9EBJtYafMJZCcHDR1x1c
PbF189TAOh9/AklSLQTou55a7LbW4GYwyTvTV1tUjPO/7Tj6gMKIO70PaxttatytAruM+VkZZrm0
1P0opbHgz8R51ZyQmjEWeLI4+3lKh+FLkS9o+7diwqXD+phwock9RqI1Rbb59+4BN+WZIbdy5P5c
xOUz4h4YpheypuYWORe6WriM3xvehrjeR9IYGyLVufiqTpmha+PFDWA/imHkpnMplN1k5KIBcEOl
9EauBzAptHX0BB6+6SxxdggukRylAngOUvl965Lw3HwPOd0H/CejrHdw5tFru7A+mavcDUNw+9SF
FG1A3umY4WE9Ig0oB9lruUzFi4bboiaFNWnLfrvbJlP7mullORs8WfPeVZYSsNXb9qJqx1cQIoB9
JW2D0SReE6qRfF2H0/8vVGtYNG2X/sS9eS4IFvwIUVLmoRr3ZYlwq6kiPpqs7LHEQ+5q02i9JYKt
kPFQbDjYIRRFr7y/VkvFSW97SrwPexO3QTmv5+gk/qLxWe9BfJSvFQJpwbC0j4sjpkNYGb7bMHLE
AwerZwZm1K55jDm8usjJiBfoVZoigJt5Yw2bq4bUNEKVk04UM31n+DSu2SKZfqGTf12MlVEtIyh7
y/JI3t2zdKobG1kflCxyHYb3+SS7s8sKw9idGvrhRKXG4nxLjlwUWaqCNqcaBamXRWC71nUAagk/
ma3fWi6LsASpFtN2EJ8N9WT92lTHZ936YHMgOYd5Qn1zH0puJSn1q+eS3hWaor9CSrivWk/Ve9h0
d9602a+zAjQxjDeUG8HKAO1jgut56EBcNVTaIUo6xeYT5iVuiPQe1hR9/R/GN+9Rk1kW4ws+FRIj
L2i0NPGX/MkdWe15mmYhpc1mYa0/yXHlqcTnbeC1aAircOQ1TiMsNJkUWptwGq9AIhpLRxj9lUei
qIPtnfRyrM3d/ZfaYgIEaZJ7tmDnhnvfV5AJ+//LZTX4AZGozYxA+bftLbeMvuYMKugvjevnWxT4
z/tNGxJiQp2YW7Vt17YFCKsp5ezub9qfMHrypYkoPqdVcYJGJKP0KJLURebt9z3xzHKsCzpLyGgq
tWQ6pIdGdCeMTbRrZzLlAl5+efus+SUXq1OUl+a/1B44QhZ9xf0XAzXELRg+LxQxNqwh7Mf8LZWp
hrkcbCXpSHziSEpPVdGefAujfe6pVL14bpvCeFzwSbnvgJ9pR2OiOKZmuqijr3XubUt1IXGwEqkg
c9j1yUhi4r5BqArkWUxPp9Px/oUNPb4OpI/G8gN/aa4GDV1MT63/5g4wdvF1q+FFzrIK1XYLQJLW
M8J+mEHtSn77g0IiQLeZwWWCzMVUXgj8b5wj6R6cHGWlWwhi7XQlbW9ElHj2BCyy8kfExi+ntd4a
klCKU5Ft2sIiLp4HQzF66IEt91JYLKMRZR+UqUCe/9sWTzHHjTtliFYgYzdT8LMybY41dM2Qk9tF
OGCG/IIBHLs7Cy2hOpJqTG23sCGiyqZuOJo3sgE5ioMMAutk0fWmRi570t9KTELuzDkEIAXS7kaN
EjINMOG76sIFOpShOaXMPHc3YU/xAA0vHdfCr1BZFlkfvkN6EYrJVxH9krFtvcejoYaPMwyZn7q2
TJ3UlSgRPJncNxIW0PeaZY86Cm78X+HYcd5Mv2TJR31tiBdqZlGHbbdxPHLKk/71XRW/RU1csg5Z
bueaYmgYfTZCERRqsGijyYoLBXJB37ONKuvYEJhixmg91YDBrsJeN41GAqfbmsIziwcFeQL6h/TW
BKNl0rKhCc82ilvQ640IIxXXslLLa8MuSXsRPc8Pr4cjLJXIuAkDEud8ZS8UZbQQnD7h4+7LBSC+
EOs4w9Bvd6+vuTqL3gy8EVI7dtZ4MY1Q0MIamwIJaCALTcqvRbpsxL9TQBql9/pznuTrf/o/GG1c
KDgTUdNBY3AMCjtgErZVnvqFS7P+byAF/hNbiqQ1nbjTYb4yY0lrpbpYx4khi4Fq0i2noonm3gI5
cxjolAmO5JYq7BVhJJR5XjuUpBvpfNyx6SfO9dPpaYaYD7TDTKel8IA7m/L9og2jfLnZjFJ1N+gh
BPW2TZvuJyJQ4CWWUcHJjDq7L2AUSvHDqCB04D26C9258+px5WqJm9cTzjpYXJhlJNuRrRltFFp+
vBIZiMFwNFI8zYRlqCtpCsIXdSwETc+L5T5i+sBcP7QpCeGRK0rKM+Fy8qfm3jvXSZbeoZXmtgAX
rkr5Qf4A3t7X+9Oqzi9z+mDa9CMVYQdRri4a0MpHwOBUTYHyjcaKrOvtd4NrKLEJvmoZIt/KPhsN
3t3yrHB01VDJnfU57xvEuW/Ar4sDz4FmrquiVzg2rMuH+7kbonwsyfcEcH/yyaqIcdtP6ocOTFg5
QylZpNM5pQ/fSEmU8L5+Zmzi0zb87PTHyOawONll2mpV1z8LhyfFRRAcR2zMKR/Vgs5BhzYrdKPA
dwqEXurNjorGXt6ghUOOOalGIgu++u1OvkCqliLNWw4OUoLj5dIlfawcpR54DP2vQc5Si1kWiMY7
hlqBJhS529f1FhFMOXPlkcNgg4YBut86iQ8V0qg4SnqTusM9HMZWnWPs+AYA28U9GwrtjqATnPe1
svUGPQzzdxHy617GO0pcKb1RbM4asucsAv6nIjh8+ez0o59T3sLKSVYF2qVKpl5DM8kvO8rlJ+La
5602M6YHmZT6g7C0XqDL4sOaCQYpscSbupVJGscXFQX6x65DKsc96L2BWCL9PRKB/4FQ+Psm+EWE
eiVres84xQ1T0bcwWkD1IBr7yXTt7kYGunPzJNVncGWRnk5QUnPV0Ul7MOhp4VF3MiuQ/xngmZ0J
eur9US7z9WkaEk1hKPOoUZJZh4EXwbjjUTzwMeapQVY13D4qd0+zIWgn9zBLireduno+N1BMWraD
WFYcK827oDlD/pUmRwp4a1OPYfIl4FQgCLZY6AXwDAOxv3qfA7deX61AWGL4A+wyl+ghNqkLMU+r
18Sr55shTtUQ1zutI/J1K34jzwgH0rL46uCGVx/ccXeQ/bemSCAv9aqj1q6sJeN40Z+PA7uuVChc
iTHfG+0aDTgXSviY91lhqYvnLxx179FSbmK4IUtlXqHoLHzpuLSsZn5OB3I4QjouB956Nosw3FMz
RqkJItpWichIsQb7AtRsb3fAIfI4ygXK0/PhsK6h9xLnNAkwJZFcDr1GRfAU701ngsrOD9uXXxrP
FwGa29iWW9qyqvTqmsGA75N3BfYgcEH3g/SbbU5ug4NXgCqx4GLeUIrbs7Qnwf3i7d6e4YFmTMU0
Aw6dBFURDdMtM4QHmo3yFSB67FyrL4gzoaOm3rS/EmFx5qdAuh7uu6l/xuphOtgVVEUF6ZirQLmU
O/TH3X1n7mq3FCuaDkO8kppAoPcQkXC3b/6jfpfYnZg43u6gPI6vIJbI3yp7eNXqY1gJu6Ni5z3j
s1OPnnEOSU1hU7pmfhQnZoQSwwLlDNI2HdTQYgCzApOem6jzcPtTXtlmVB3hLThdmaVY+6Ido9ew
f/2zQBhtzNAZ6Nsiw4YavcGzyqPfDdL8SoTyWyqfTQc9RDR5b0kJdL0PrLtXfU/zB4d+7xsPZF1e
cxWO5pJ4qNEVk4K0MSV+9piuGeT5v/IuRKSyVEWc9u9UcESTJsoL9VT3sfJeT/HEwxkUFYZe/2YW
qIV8zLFVLrg95wuAN+4mxXlVhkeYWNyRtkFL1UYQ3qM8w+i5+gcfo56ujMjOxTULdYDLlxP12nt0
3iNHTF+qNr3FuUkj2+8DX0rCUoUFZFTBuD8/GXCEH7lLDh2rj/+a4prijHXh//QeKjZPPWXA8+Jm
wWOvm8/85cRwTtEMjMqFlupkV51Rch/a15h7VX1KesUfaZSnF3Coofysj9+tqmYI0v90d6fD9nTD
Fm1MqiHWGThJGLAMyLKEb0DqJbYNrv5I0ZIJXda1XFkr3VtWJfgzu/wDO5LJxfGMUgriTVSntV7/
vud+AhyViN8EbviOMjMf9XSUz2zqBzUtW096ft5cKzpgu9sd+ahsE9jhbXFPL4ViIlbHO5xWI4MW
f6bpRBFNRtuu2Kdnjyi62+E4dIEt3DInwusiDL+50Hg9+H3TznKwGYqBcZMOZwrNR3ZVgwHByIze
8ZMkP49BaJjJ7JhcxucNJGXdPoDMkb/HDziZsTLz1dOtpATNxqIj1H9iZcHruFuemuY0YTcALnxD
QNBIzptL9vdJFBP8cuLpATjITfWcz4TWTLNxhw6i7I/V1i73RllQ6PBVrkhSkeQO2fLraY6GoGS+
VT/qFVL5ze+WThM7kj+4kbJvJqoUjV/JyWR8QSCKx36pjv4WZKRUdOQz4O2kLkectzVjRtMbojZ4
DclXFmU3H9wCgfyxlK2c0bciny40+LhLWqdu3rODjzwIoYNynEKEygQJ+Zhxz4SATGOS9EshtgB7
daKvHcjKqGf0CG3cjPciqDSwi8izuiZvqgqdcdVV3lGwYFNw6/+Rz5MWHftia/FJCpAhNpWtUE9A
bnkm057d/XKcqP+rIl/vpNQFK2GIjO86Nd84h5Wd6jDg6R+MUZuDkQd9sAMfEFEdPJmecBhh/4ZD
B8qoWuvlwa98YwU7kwPbRYJFjbdz/qC3RvUgM1SEzO3MKH+cYlw+1Nl1fold/IIZRl/6kOfVJsY6
voE72QsmWa3QxI4wGXqegGjHfwJ3avBghmrNK8vyOqqA84MJ9dkj5+D7kEPXm0+wxnP5JWG9ciud
cTuQ34sMTbmUBCr6AIn2hbd16/syyIE8cRpI3S2LL0TlRFStUu2gmaTlxcYIjEuCqPPKYMG3fEWO
WaYGJiJz3kwuoBiIi/7swRJ+mtNYxF80oaRQeZVP9jR1wzJJBT0g+7rcRy3u0F1Bbz2fBVF6+LA8
tZ7wViwejVjytggyxmniqDmiCoJqThMd+JO+y9TAuUwcfTSrGVNKkEcLEsOkbhOPLAUOAXKVDgeC
OMU5k4Vs0+K3Agpiigz6X5jpUcl5mvrvCF4JAjZny+XsLzYw2rJTFK5Pzv6f8FzO6CI0zolFoAiS
Up4ANWjwLzJ/OAUwgK3dGR9Vi1z/dWatnZe+HbmNOCxqfwthiq7sbA2jnHp1rlJ3keoragWESADw
j+1u14hZzwFDnjgHbnN7OOP6bxw+W3Q/Bw6kZWSyYbQrCD7/6PFWGGnTMxXRjQx4a/E9kc9Ggoxq
/OcsOU/eQnW7P0UyTP/qGNMFy17F1rG1hqVS8oT7xHYOV2PnhNijrS5fa/0wn+8ussvNfQua2veY
XpTfVIOHWMehEEL51x7eAfSOdRsiLaeL3ckVx9mBLxtyUBxG2WMYQ05vgNe/Rxf0CGPr8X0V/l/p
oXGaDTdBJIZfg0eFCL2jNgan3YseVEYc6Q2gzauvoPAb9ofigPTGbQJNdO0hZV9K1/fN4ioZ3ZeC
sPoprQuDTXySLmhgiWApuQqeWtOt5bpSn/gY0NNfqtMDX8PdGA//82x3AfTL+FFn1Gh0GulPJdGp
Cmi7OyURJnceWCF1hzj7IjfcCjtMTHiHsj5jMXNdiSqKHrFmPXfdIj0Om110p/NtdxjfbdJ3dGg4
61guvw2H4R8gRJ2l5yS1ZG1QwlTB+lDckn6zjTfGL2vCjBtoyBT1vJ2EOsbqeIfDQhWbdW+70qyt
p2fNSQn1CN+fSbr1JSAdOsGz4W2XLyXekmaSDQwmmt4oD5RAI3OOeMut0S5xO4Ruhwgc1olQnfkL
7D4ExhidqlKjuwOuu+AnpN/DKrRs44EQEgV3kNKAA3tD742zLx43c0kfCZXieSN3wrrlZHwZRsxd
5aNCpQmfBr+aOrHcMpk/pSJucgnyOrwKEcjACCEW7tehxRHOLCmStdE+gWMqHbCK4W81vn8ftKWv
KbL/jEM9qkF6ctm3ITB0wE+EeYU+5Rz66QUome1tHXiiwb2sonKgJp2UXLAhZPOGsm+FSOehD9I0
+gqig+L+fnDaYS9e5UJeJLg5CUOHgucQoq0whtA4TbH5CVeDgmeQVk6eZObsFeZ6QAso9TCU/ssd
mrzSJqkFjbdko3Zf+5QuJKdZO4YFEQ9JksMh5E2JMacure7jMcwA3wTRegI2o4OFlS6UP+MTHXcm
vArDLHnE2MFa2nGC5X7e8EkbnFSE6I89Oe+CMuH0kxjdJJCBCzd8iBpu5BZ8eXJ85v8/YqSa8ZKr
kp8TC4d+j85AmqwAkLzjdOFbjMbaMBzY994x4emcFbgm1/gChP7647pWJ0wXHdFp1Yjy9zr2gBMv
Rr4Bsbjd2+1HYhvH4dDDAQwy1WF0PA7cz6OpcoMU+UDFlCMT42zTTZwAoAmS/WN8yc23FYIrvPfO
OiU+/EI02uNwIqQlmlhWO4EOMka2dhdfkWFpLAuuhv3lykqs5bpqgxHAaCkn8mQ2y3C38OZtDjj7
QfbOGX3u53a8l0jd3ogQbe8skkr+KaZGKCI6eFKdE7ULPByVyxIpVrvvZYjbBJ8BnD5f8MQPjHw8
+dMytQ5BqIWG9j5BMmFhoiEG6OKWEuB+ZAJmwgm+fbEAn/DqfDx3MEWD15WVOjI4m9jReHDtTWTO
M4B4RMV08z/mykiqc42iInYoftFyVCHep16ws5fQuswXuTLjobsFJEcn8WZtfPerdCWv6AC5kQuC
JLx7tjWiJMNkoxvb3m4d3C38FDE7S7SkCbrQUp+B5HJ3ye+MVSWE3/XC9++JOG4se22Vex0gSqck
yDE312Lri1Ae30cdaZJmiLHh4MNvF3faSs298vFKrqnIimRgpo+EZjoSPFk2Vt8zGoONhhfsl79s
7gay8DhmzjZiUfvILV/QjAeVRY+2+nZf4F5s1CRvKBL1D4+dCLK56cpedwIaojlwUq14FIF8jbFn
Qjc2SI2gOyc6lFdxBYjNC/RVa+RWhD48YQgBX5PAp9L4r++gEp2XAN+dD6Qah/apHMQXnpREyNWs
XyonBbbusb5zyYRNyH6rbJbXfAmzMyto1TaQEyA3A2CRyR6HewZDXQ51SuEf2Gnr/uBL8czw2XFN
za2LmZjXLSebfg5ljuBPkynv3dUvJyeq/o5n+Ue3XkriaysPZbqUvdHDx+HJtZFnQTxxVeLOLOVg
1Ljtv6me/V6VG+N0C4slluTLLbFqhOiSXbLeiAX+6xOgSPKfW3mubY4yR6gj1G4fsg6pT+n8XG5r
tQx6Hzdynz1Q1vWAX23SL08r8exdtpiFiAbnP1Iomq88l5l5SWaKabtWe2EGFejFSXV/pz96ocmH
jsuvuUF+God9GXIfK4/LWWjtPpm5aMEmC8nDDD2tl6weLkxRLijil7MRZjW9W7eGXjfZrjhooxlt
rFywJHMFmBK2l9kLkRM8L6ta4M6wzMqjNsZwx7yviPqqM1ixFaansT1Wu8RBhnBRbuSHCrE7nBx+
3PPX5VF4eWP36bcSC2Iznai4Z3opQhqYDh0CqCHf1FFr0ItveuRamHonggdq6gjLW1ir8kCxpm/Z
X/hTBHpmBJdmieWmGyKRdQyM2dQHXwt33FwbdG29P+fRMGexLwJPzBqsWJYS4cyBsyN9pp/P6VKY
MUhcRWZ1ezehnLO/Lt6hI9sJoGsUx348QxoW4CtTBj7NT24aLcGfzC1HKPS1gdSFRfxYdQcXJMSH
mN3hh58sbe/eTQxjeXCCVLuVvPg1VLiiH8Ymc1IWrFCvUI9mkQYqzAAsB/br7vStI+IamZ70xIRa
5I16tt/K7jExGPisaZDJ6S65Gqwhz47JkogLZYbAwKSWnhT3/3AsHLlB9u+Kqh96jNUhKEPPqphl
RYQ8pk/8j69upn8oqnuK6cqRHY4J7M0gts+lpyIGoxBXMFaDoaTcgWIMuhx5gxderZYfE5rvGTRr
G2R0FTekWTNTTt2nJHl9mifk0+6XdDJVUdVngwO+VxkCw8aJ39TobRe/K0xfhXIcnYonISPAi4fK
XhnJSVd5JY7S1OM+t403eBQ2cwOQMcInNKJjromTvzNSQyskM/3umMBxVQCDuC3ZnmMgkDKzWpnZ
2eoYR2XFrqDyNjG4yiTVePS2VrJ7NkaanHzBKuquGBXKlkA7OwB4gto+CtUt+ia+UML49UilOlnF
hH6P3Fen7ihzQcL9IfL7OcUair9zU9Tb7lgn3Ii4gFkMgEl6zuR22AuMz3V5T4f45hgZcD3KzzgN
M6JMxupb7IOTtQRfR7XENzxAldkPvibGqBWjk5x7orB6W94o64ZRvcQMju21CZhr9gZNOBj8rafO
HiZNaMRUjDSR6UWF7cxxmVGZxQZZcd1kIcOzu2sVzWlN2TQy59HlagbTrpaJCUc+LVuQcRwTMfz6
2FFokgJGV2jq+pwf4P64WMcQsxYvVePkRSIfQIKB92wqCbUySEqWctqxgkXBcJVMjn2ZRM/dM+OO
fTYPRMqgMASNUVUYE5iC55Wx8AaqPgSFWjPWIOW7UnNoJbRxnAnnSw/p2bSVTzcyGWYVswO5L1BK
Re1deI6HyRxYFHLb7AYiNf6+27dKCngF+CiV7Y1Pl+7AtSx/Wbs2njwIdMvCDTEfSM+NJc7V0LzJ
my0VIvtmeiDJLvAf0Bam1xLmN5pPlRns+JovHqK3PjRPIL5B2u48qGKZg7OhltHVAOwHmc/kW0xM
5fpSv8d2+Rw1cooMfr2yiboWQj8hHytLpe3ZQZ9B2jkhvEuW+2hnfH4rwS/51zmtYWKA4ZHEBwyy
kkzZXsBKk2Qf681TInfTuz6Ufaoc7GnS+B03Rag4JWvQI/lRoe2cABjpOlkwBILZdDt4YG9oSQ8F
ENbKDuREZ4abdQTIeHztN4EEpL14qEYK+TV9a8gtbW5E6JbsGNb1Rc+84GheDigcLe1aa7bG60pk
89QJiEGztSsvucttFd+V+LgIZTrTyE3Av1SXVup9i2pql5HlBKo6quqXVgeosfkwogCzkVSigh+3
a9sMXVsl0bDZzxjBFQ8GgS9swxDIGmTMIW+Ysgru3Rq2/CB/tqbxPGzvWBomZPIs2U6S0ntbzZxB
RGbS5I/gIRg6791Qh6A8MlwwG0xsn4HeV34ADtr3Z3pBVYqj7DXI3yNGCFIdmdgnmt5zKcuBKQDZ
Silo7xGnQnKl/uM8lVz1J+E9+K+Ckx/NqvIaDvj9jhU4OaqxoGoBEamlTcmlHQp+assDREWD49On
ibJQ3kv6qM4F2iOKmG2IsPj4hq255VMr9F/KzpWUshapEgY1QBebZMv9oNfzHa2tfSmeNSxsR5lR
iCXaZesubLiPDaNuT5Xm+M/X6in3rW2Upe9vgIZqG2D53kyYkMTclFXcPLNDV6lY4qqEyb9IhMGh
Xr8QbL0faydP2uDI3PhORz9yAiW1m4dA3hfoy+UPfo/9Cp4e6A87M6hw+M6UmfPuWsL3xf9ZZ+tb
94v5IHZzGHZNZUAnbhlw2eCnj6jbWc3SUvgu0W5k5HqcXfKWVJobxr90654/zgyf1VRkkcYOxGSc
Y055cF49E5vuIdbSh5wtmu4cA2hvKyZ+iLgsvcDMkcRigKOItP7VcEH+MJ3a52EGQc8oalWDe4ph
Jf3FOqRnAeaU/nOKseUg0S5xd0SJEjSOxe/z06fqiKYQX1D9T0dsqp3sGMYUQ8SdRCpXssL21rSI
kPoV+7GyNLlqK0rjIbcRBV3JZBT5+/jDWspVP4o2h0aFqkBMr+DG3M4x+9aZNOJSJb+nAMSVh8kp
oEMCHIwcWRILDFW9vB2vd6hIkvxh48Cm4lZ4E8tQp45kcjg3mdX45PkyKH3iW5yGB6oAWKaKWnCt
zrRhVd8Jvet+lUBTqj06psdXgrhjyGLjhK9gxfuC4HOKwqkUf5zQUPLYdgk4VW9wA0X8eFW8tPrr
NU/kvmwlZSwg5q66xi93yYWgAYJ9ksEObbhoPoCtBy5aNLCpUJ0OU+Imn6lPeRbMFsGZvRBsgQ2f
ww72hMkaQZn6VhNdfSujW7CZuVLZupX0nHG+K1Wz24Y0rddXrkev/GA7L53bDrpPZRMvO/kbZIBh
YvIaJR8oYMhTns+EWQZt1KHeyD2yLMXy48WeEeD/vkeVRhL6Zz9fpN0ExHYgt24chcG0GNyAuc/q
Eb7iULXeygRYFzG4nljzysCC9vKPE1FwGLGHeEmUj/kHyqy4sxoa6M3xEfZ77R5eg04oleWwNK2I
XsiJ0J6NSrftEXMr7FeGkZcO5zbAUivMAHIzlnjJpeqcYb4p403wLyzSXqi8EocWRyNcCDyqHCiT
6b7sp571fIoqjaGXU9/9uw5pL5ctyf8I5HV679cbjn+BnTDJLhNJh9u7CVHALGUzpvq+jCe0xfKL
yU1aNzJMYKkgRuGL7rf4t5lXJwLP/NrQLrk4VuzHlH2fJPh12EL3gHS156V6FXUvpHNzFkmexU62
hTSFfDwl1pfZlcy1Gr07yCVmr4vIicfB7cXDCqwDG4ymW25+5M4IeEzvdWiT+9QliRanso2Sxsoh
gBq0XyQxqIs2RgEhDEBNILMuiF909xz781k8OBNt3gaC3kcDHTTWVEwn8zMmPxwdOBVD4PbtaINS
7G3mJFe6hhse9nL1W+y6MD8A5jXpPqCRLNcofutcpoy2Bay/bUop1LdONzoe116KldcBhuRExISt
246V+LLRS44feDWQaGwZQgAuWMwWdXXllCdLSwsDoXGGCWfXHT16Ou4i+yn20ch08HvM9dnnVWIo
FfzfXXt+HH9ezPfnbyWUUthmGkzw+rZ55BPhAXoFoE1K8yB8ED6ppfdUU+p7QlvJp3+VSoBcGAy6
QEcfiWCbs0CVQ73LN3limYp3M8RvR46lLJ3YIpcqWqPLrjGXRbr0mEjxvGu/Gn+0SuHrL14DC7HH
6552K8ceLDREO+vbLnRL8Amm+Qc7spP8aW7VnXgjrCM6RIHwLv2onLt3upvDgbJn3AynCOLS2U+L
aM4TMJtUynlQwhCebKXr/vw/NzsHyAyooZS3YCzVFpecZmLAb9dtDegNUP6rghrb9ZyVU3pi/9+5
D/1WGLPygfzD8+LxVIopQwIrtJQiEWrBXTbWSoCsIkXl0yCsQQjnJvBSZrDMZVkiPhkZuOE+cRXJ
FkUb1kYRbjzB7/FptrwQ8iJn4AKQYf1F2f4wl9sbERDJPqxNMGk3GjEPFIs1KMHwMnXqtyfIBy0Z
+zs8/Nj3ncMuBdjIqT38WsSAd3Jckhg3+d+ObknJjyn3w9ruDcyYKpwsTD4gXt6wrPoqKlZdZvjk
n2Dj5aKwnlqppLj2dyZJnqYeiY7fSH6lKCdXAHMBu8YiGPLcRIHCGNkkgAOHIK2PdszHDrubhWr7
k9owjGLdQ7oq11k7pl+0VnWHkuvlhauNVF6Pj6vNGa/Z/YegvnEyGJ8XEOkFPQTEalZ7rzbxP7bX
NgUqNTrsmYfl0FjuY/hQV0mABTZsvSUR0Op/vj7nPnNZSs7wvzPyxkngyURQYOy7xSW3B2JPpFz+
+mJ4IIPa84twhn1EK9urhsAQ1aU87ocrF+CtuE3ZRN/FDtd3GwBuBQbxPZdMWOP9hcWKjbbXdwXb
DJj8uV5G8uSHJLqSNqCjNiEgTLFrIX6QbENCzuPmRT61pilTYPy+jw//T3lXLsZIf0fJM6GZfIEZ
RjCJ4pgC53rurquZJEkzdpdBE4EdTILD4kZ8d2O27dUzRdbmhz3gZA56uEba11OoPLip1i6MO0G5
w28QVQHCb34LvYr5YKKhYn5Wxqjdi7WaqPu5rAf90RyM16uWZcOHMQWUJnP1gf3RSvgXqaQ2TXSd
LgfWBypxsBP2mQZQsp8K9kzaKD0ac9W4139n2my0CXnZlPH/TCpVGP0aUlQWIUXnJ2XzAAJv9NiQ
SSta30uyqR+xPzOXl06QnpVj0zFReUEokzl/ktXkV4HH8zaKVadS9qHsNbtnpW2/qQc1GbVjLleY
oO9U9L+aHlZ1f3voi+8M2odWnpGt6PXi9yCJaRktEPsRaBWyZRFz7Zi9VYzbD0AtmmDYnojB/qbk
PwngU9eFmYDBupaLNGW+yz3ghdsYQXCS3+4AgfQmXFTbKWHyHp0g8Us//fmwmkqnHx3cYb6EQXsF
e4KEGvV8ZDHIPsoP/j4LZVumzYLpGP5DYMBu71+UfD6jtO6JmvFypkkwq03JboTlP2FbCO44TzCI
w/jL8Zn4lhkcjTvMM1LnyLS55HTm5HrGm6dgEVAdZ7LrfP6vy1aQdyYgDgftMUSKFkzWGBRhK0su
IAI8N9DBvREtb1Rx+OIHb5M5VRfaa/0B4eN5Mq4OmVKg+3ZuJ6ywCivICQk90eFKqE5HJqPrB+86
a6jzB0Wd4xrRYf5eWEgMR7EOfaBcseYX7DNR3yO00u0wPV8JBGOV92dhRUkkLpPi0ROfDmuqWtsb
VaTRst6gGoIA0roFjxdSQmDXuxpU0+poocmovxmhH5q+ZBqBW3aP3BUTELb0lQjB/FXqgMo7Up5n
SXvArIWS1TvImS5WtPMdcKSA4ZsThF4lOcg4dlsKmfW4StCg8uxy5rWsLIJ8awOC44wS/rfrGR/B
fQxBstPadfM3gSqLZ9hvgXkFReoj98MpLAYGA0om0Q1hQwytKR9NHVuHwSJ3MzeICDPoKmJdYp+M
poLRcLLD6XQEa9f0iwdFBCMVxLXT1AIqu3zQoWtRSMByyVJur9OFx03mEjm5Kw+rmIga18gGO3DR
wh59MyDtYuS2iqtKk667RZhnGuUeNeIkAMqHGoGZwakmTd0WTOz7jHWGdWo0TyPA9puE1aGJg+S+
jZVCCLLp/V3MhVpwJd7K4EcSxc8Sq8cqU5J1R4SVOFmX/Vq6Kr64I7fJOy0DA40PaoPtEpoSOJb3
MaRQRz2GNTKCsRXzbdVnDXF+jmwv6q9cR64nU5cllo613RFnkx5tmVdZTkIcuAAJT6GkPG/tib/E
fIdnB+eISQOCu1T6yuSPiUFg9rMn0XCLp0ueebAXCkBLdOB/zD8u10/flzKmyU+T3wCW6X7BecFb
4lLipX0cayBtokFR0bvC1c9w3yG4ZWM/MVaX3i6QW9NC53W9s82PZ/+VI5SAr8ncCniYynfpLNhJ
P03fdE6X0Y9hxgul5h/LSP8qcSSR56sp/2FGnr5NEslAcf7GgdBVRcL3+rtroRDNxOX1Vq4kLva0
f0ZHOtFV6wsq1lRv2IWqzfnLVxxTN04z3cwzgse9gkbuOe2eFBEnekMJ4mZmcnb+rLqtBQd7HdX+
b9J3h6Gafa2/EpA24pxsdZcPa48bjWsqi0sz38dY0fIPyluNPf3XAtQya6DmYQVJmZrMhPzboj89
4+vTf38QmLz6SIow7uY8xSeAjQvWm7w8kY4k04Oc/sb5by5z/KpYIRer/OAO8lVwSQwR7ZNDmJr3
ns6FTJRB1iOMhI3LG4zOL4VjnvVbQngMtapOW3w8TxESgWUU2gFIw7TuHjp5su6MoqKvUVpFzFow
3liT5GRlWWduZe5E7OPSSvC0s669Di0Fu7Rrzuk6UeJOPztLF5Li27wYP+FMMHxHKwDJtPklmPDu
3Gj1133d8IV4RQ9leIM7kWp37FlzdDoR6zA98jGVjO6qM6xurzv+WZyibvYqHhbQ7rRy1mOW/puQ
nfrbqLXpB64pQZ/evJgz8tEdjcf1wqFvLvEOXIqlXY0kciwWZ9JCCwv9flWemxwsozaUa+WEZQlW
HzCH0sXHPP1qIGtA4XxvExnyww7iN9ByeVf+ZofReewwBehm823lMKoL59/GwKOGj5W4og1yY3pV
QFoJfRX+m1oHI3Hl96//i7nzwSu5mVxntjkxRrH1W8YkNVrZGzy+FF64C1zLC7HDwzO7RShKelQm
JCE9hx+IfYshJy+4YiKqr8HEjXDVB2pWpfCcsfUS6qS57M8HiJtkOsuP2HtK32HuYHVofYmCRrSe
4ehDKHED9LCF/ni5TcIXba2IjSKKcWk+CduYtnf16LgFz1sg5b4JmImP0o2vJEhlqV1xR2Lf9uqL
1DCZ4GqGmbrxKJ3XmwK0Z4mxxMS+mUfnR0/YInt8uoXq2LLdWI6kTKB5w1agZvSdmDf5zlXBYohX
z2ESHrEqSoDKd0HjaLZstgWXsNJc1wM1Qv90DIxEiEeknNOIBIMjTclWeRNFXEVLDVM29sto0cPj
LP7LMM8SjtlV9pK/pvh44bvuKS6tVPQEgqTMZjdUfat1iKmlQEm2VIEIBSDy+/jJqh8Ff8st/Q66
4/+TvSw0Q8eoDfjIO1p4a0yYDzTmcHL2D/SMyZ4YO7Rff8NO5JSUtmOdHfIfiN5vWA7Zjq6qDK97
TXaqESspARyyDsLCFtHmFwer4iK29UsagYK7vLdpfXQwxxfpgDScKT7Lqck3MCUGq3AltVn0XnGH
zMU73zMCyoOJ8z9hhkh+9wNLaOBT0G7BxnSm0PWljgjHxmElUjH+dR1Cd/T59mQXAgaG7ODnDF0h
sSHbWFzzx7uk4KwKvda1c1PUIx2xJiVtxSBZi0xZ+E0BeAU/SL4dEH0jsyLh7+WPSPjWM7Km0VCL
0pCP4dSERUJ12462lqmH4rxsfA0mzkJxIo4c036ywbi1ZAeXMFVie1Yao5AlnIRBGH2MxFrxyOwO
7IvT8A/8ihNSBwa+FoLwj9CG8hrgP7WJaS/Njiq2NLeoM0lhmeVdXMOlJJa9poBpaEKunr6I24eC
lynKC9q33Lb5JaXrdr8ADDRV6O8jKLF5gXhV/D5ey2557rKl7qYcJKwOAeTx8fZKInyvjDhyHKR4
LS0mqzV41ctxOKtaQc9h0jubkVRsC5pQ69uvnquVvKNsIwXh+rxgzV3X9tDvqEG5dMKdExxWHaOW
7l0Hi0oQ7fJUbsy5D++r4OgfOTCRziQiJNCAKMZouboECuN+xxIIxsGG/QFCqiJ8WQd6DIc/WRS0
AiWtRngICtyHz3vIKndrcYoy82/djCli5rundYXemHmZRFegR6WM8Qoa7q57DljZI10Xdn84Ox+x
dU+5KnOGjCj+m2HpnYKvggY9GCGGdQkgpQO018P4KP6EaINXt5WSKNwbCrbt0iHvO4pdAsGfnXXu
uPbS9G3GaqN85XQtLa/0hbac0l5xGDOKSuYFQbqAEid4f3xdIiKF9ti1Zqas3ZbBBaOtGFbpcPS7
RtI4I8G9QnC5ws7EfF00Iyc9x1lykaCz4u7Hmk7lRYQkKlzDfok351JRenwhBdG0krShKsC56yXU
A6P2jPzytr36l4JfVaDCcFFv/aJTscIrvXt6Ad1v7jH9ziSsHervArOS1IYLpOHEZkxMtNGlM0dP
Q9JLSz/po93Kyb3pS96zgxUWK6f/bceem09zGNeHg/EVQrY5e/Y1llxs8PEHpwjGPcnyXrCcwgEY
ASolZAdj0nRiQpLyQkTALXF0gySl0jl0IuCzvx+pc/1aiJOqJNaCvgFYWKtl95Kf+Si3+mwy6BHF
utSnyYIgRfXC6Y8mNPPG02sTvRzZ88NgivKh68qjjFoFgBJJsmNMlf4PSWQnPHf73RxyqqgOyOWc
o7E2K6NCiadV2NCIZfHkNNRENxTmkULNX5/OrWZ+N1nXaUGXXO1OLFr8L6Sgx9t/4UMFDF5AXfAI
tE0I/IMExOZfnoODuYnSB0FGLOITuubpwPRNBwzN9rIj3Y/neVzXboOpIy5dMFFi9BtD723Km9T/
pq76Bly6FLAaCdePkw9RDBHC6lUDc6ups/j1KSJr7h8tPQHBjIe3wxjodxk1dxIoLn1AzjrXKz2X
/fYcDW+jZOqkJGVTvv2Fj49EfRIWpN8nRcoX6LVxNl15hpsCH5XhO308meIbTOaDfPbExp5Jc4Im
2ktetHJSrbNofefu7gp/oXsZLrLFcmUDp9kPC9ibU7seLqotzyiAB149E2Sy2ZfMKEOEfP596csi
JF1pSeNmi9gXUldjbIXrO62TH/U8lHr/q2DgJYECCKhpR40A1bLTOBxtU5/iF9Pr2s3REIN/0+jO
X9ETcjO1iIxnIm89J3kAj1qLmMMQp0bGak9fOhJGjWhlWcwZAEJ6FT9NwZwQ2b15yIZnSBuBTdh6
593Ch8eZVMVfL037SRLGmkNbePvFVeEY0fGDBj7LKPk7J7BH/xQkgzSI2aDizChNyiISY0ZxHzC/
Rdt1cRa+fxnPQpV7tR4HFM7iSuNdtUS4zwS7YUuvOmjTtof0NAeH0QPBC1OxQvJQL8HA/1fXVzBF
yf409KQyLFomzpPxNppwJBJTXbvoPmq++Xa60WYUuBPVebabasuKLVyblA+AcY2BIjyPr/+GNzE9
qzQ/hN8yu2k/iJOglqhwKy/vxyd33pBcMsld7FcTaI3bIOemNAOUe2WzOLFd4AyH2xxJdHQ0Kavc
5w28l+RpoETGaFbzrzRPGB8J17KFUUQJ+bPETDXsd72384jOzqC4DEr3Kf5mROR6sepfAvEme9UL
uzDf2/ixFL7IW2Z8kW62QSCqD+HkkGmNYyJEubllyt5eiPlVoh2+ui1NTOGmtUshzcKxIeKhXFzj
6pAydhxt+Q8ss69jjDXbZ82aCQWrbLOUIKVc9HlX2FgzVbbaz5WJ9WhyrlcPX2Cq044TmLJ9J9Zy
0YLZls+wx4yjdnOkBXMbtnSwki80pw9qvy8qBO2CKfvVzrorWYXe6L+o8vp7QbeC9bMB4Q1feeNI
3fPr10nxAmvxl1nyFKV/k/Kv0rmWNfmZUW4R1axF+i639bynD+aMhVE215XKCN0IVG/InrbcfZuF
j4vYLnVOdn1uLJH4wHGjsaRw+88wi7C7YoW02N9OlbTfhmAIrnzIhKTQxz+HAxUv++45YfYPwWrn
+6FeXYR6+8R6ADr+3ohINkrSXxbAobqXjtyU/ddGcbWP8H5UPhdgUzGUl9phKHk02Eblhy2Yxg7T
yfQQiOi37ORAczbBDbK3Ut9t6wDWL0eVgvMHAmrKqy8uh4GiWdRG5Xyj3D8IDtoUgyo0bbnm5LDc
navSa0Yh9DNKUpKWktFYfNy2z5wxKheCA3ItOuOG99wp77AHvTMvfQYZIR3uF/BWa7qXMydXFchm
4tkm2XaFPIdewQJEbtE61aDyRfz88+Kz/8hPPykRpFE6R8JBdDfHO1j4xcz9WSTNJZSFHaxe7Su/
ixVI0p1dwafCrlyLZh3aiVKMPpuG2TPZVPV2eOZ30BvH0/Do/+1UGw7GNFgavTVsGm3faT00nzsd
3+FyzgQR0gPn0ZUljqRgA1an/DUM/nM2fUgMQ7RpUBvnfOQeUk5vBWDIEwqdIAduVyGGJwrHAcJR
98ikzamvJWJGUIrtgzZrdz/c4z/13hgAOPLsGaOSPe96Dc7XwcT4lyQkQ1hQokRB5a78ZyzEHQLb
5BqaqVZb3BN1eICAUdkePQsUOfhb95NsvjF/xKlAyIHF7p1pmK2JPJBDNmdjJaEFvU0YwyU9NTO2
l7FxtEU93HbFhJP0nbukmGlKyB9nLZUDxZhO+LMi8iJbfPsx7RMMHcz+Es24d2CXJ/KCM86a3yAf
r7PmMn1NiyhQFPgKL1NxNl20nf8ISugoMfkH9Ehu9sd9g2Y5RRIdEt9GWUSPxEMBaWjXY+wOJ/4V
J4Uqqrn7EcdJVanEL6ZRpLNQephOmsvEK8qb1N6MspXgkmsSM54kSn0f4je5zlAMkFLIXa5+jk2c
Mwxzq5lYKmOf9Ab24mz/4ltqfQ2c5U6chXpntYQisyuC2XT4mMXAJdyR0pCZMqCwAIHXZKMLyK/S
UKq1fvF/fyFDmuIAtg7cisAsLsTQuiNTRcFnjyTjfdrgxX30dYAoyOPjCHvRp5+dKnAQoIbIa6Hi
kjGNPa3URAdCCciUA/vJNhOpmlFhQ0QUfF/5mkL28TsdSWOkd0bzEMPPxIPVA6koK9mLl9PlXxmx
V2SBECHMU64OvAbw72GtfQx/HwOm2uCg1v1+VYynCXJ8a/YtNRArWuaH6lRsFusDirJtNz3FnD8v
NBFSba47RwLaGsp+kzvhEOx6Am7NzrEucbCiOHYy64QgIdn/GKxCAEdbEVpDatBExscf3nkI7l+O
MEkNkhg9xhGezVavoRdmr7v1ArfhIA1IM80dFhRDH8z95Y0nZXvJNgO2+m/uyDad7o69QTo1JvwV
KJzH11BBMa74GfL4oQyFur4lGf4T5el1JzD7Cug6RtD6nySpJmybrGr5JKahdCsAvcJ/oSRiQdbk
1mXFSRDPJuLcV9WNP4wMQhGLxzuU5uOuqXt/39zxAQ7aJj8ZnizXg0SiSdo7xRis6k6aV3ZttQba
8s75zYjRvr5o/UPgjtQK6TWzGrd0dMNl+AdI0E0uDVs4AGTgFZmiu5EwhQjM5rPQp49Evn4aD5J0
erfjB7jEGe1LoN2GTZk00Up5wbJOzQcTTD1QK+zbnGjI2o915rI38eZhDYIFD9DJnBIogFYO8XOn
bvrmYQq86bzts8v9Oh1Bkt6suD5Q/m/TnGpicbAE06HlLp21SaVtIyae8Pytvkt+b1mtiPfEmJec
H6Zg/bit1mH6LKX+MwYSQvumk38gl77Kgk+cBYY8RtWN1hSlNja3NHiZXu7Y0x1wBQcb5bIPsmZ8
RE2klAeuTv0Glw+4sNGAo79+Olx57T+b1j+Sls/+UGQhflw+eXk2lo7ga86F3Vpsxquzjo59zQBI
bxXG3Ga9jK8/SEeEjSxw8A5frj34NH4jAFOWTjzeYo70uDn+z/KU/Xq7t2V3jFZZM7SwP+ErCyws
LlINkeciRWeBZEP9/HqItbON20cPj7Zoq4DR0QWZjYULIK+btmwPHXovSewo9F9IIVejtFJJ+KbB
XPg3Wbgg+yKCzNq9TW4ABIur96hsRfAKSTJh5WHsmvZ1aWlVPaO2bAwVsRQsd5/i2TPMuyvgdjOa
HIzMkeTZGARjrxUDXN5/ABuSBkjOe0c/IG1mYQFPykM/dBTqDY+DLs6tTL7CPej1UO52nw0D0nwn
+f9Un0FjKBcOB1eF54fiOu7sA4yk+ALzW7wxNDR3m8ejmyf0RgO8QXt7Ibh65uUs7lObefA57cGo
nGHuufF5ARE6qNpGzk013Qn7BsBkKghj0aI594518N3iz+ckpSRvijKaj7lzkWWoh+4APwUz7d7X
0E5zE/UvyynCSVr9JLJwcb7LV4CJAX7QU4zqqO5QB+5L/VU1Gm1btAiibcddsWWJtmFotKjZYJ2a
ZiX5rCDCrdu8kcWLMGQB7dxVtx6tHhDC+bu1ZnMlmg7WutZJqouNKhIj+umnuUPx3RW2AdKQMVik
X8XvmBEGTyTqai7MSQhB2Sx/ASWPus31myh8Lunvp1mruXfXihBzu+TiOMytUwWY3oLYO4N+Oudv
z5nLSm9+YedbbQQCnap7RMHUvPtkB+jKvsvd5gkLVYIH4ImiYpxDIWJZiN8GWyjQZmwXrh1hq3LL
qRR28t55x9CISaETSmnYTGEDDeL38UVZkpwkfvmADfBOYSpY3St59OyWLPRAiPtEAF3574OVFG8X
dp75eeTQLteKpO3usayjjG9Imehlg/W+VfOgcjfvShI4Z8tAa3qtU9mAhEZavPpPv00HruFqRDK8
jbTftoDO/JkFVknE+5qZvzUsdaYBhFYKeWgPODP5kuo6xEXrdNaaP2aH3n4xzqfgv5uZB1vJdAAu
Fw9XSG0tVhHw9S0DBZ9BVaURXb3a9jvydFf84Ap5qm+cA3TL3EcYQ00Q0ZBhlIKGhK1Yr3pTvTU8
OGMvNIvQ4EB2LbQoeW63+SkOq83MMvEweH6dcsvAYCfuyakNX4WTTpzHaqeP9q2PhgEvwc3kBXOS
fQnP19FDrb9g5uxJcvWyAlAyea+vEKmaAYF/z9PoC+utKmYiKDXdxztBGqs5PfiNJnWVdR4lDT68
+kIbAJY5DOZR9SSqbsM8uRvKtY6VPo+SatUMUxHulvEo+bp2Mnc9dDRkU9s+98BqiOb4aVB9+ieV
CJmKeInhiVD804MQRpWPD95BkAun44d9yFEBHiuCKoBhm7kHeVPjEgzx3goKkqrjiRqvxToTLEu0
OToN5fi47FuqaEULEeDTZZnuDK7gBgqgpZcfP9AXj7ieIKvJs1BQIDzLLRYR1BS/Sonc+xtI5paP
Yt5a1FYokAmgbiae7A7ewA+vZ6Fh9NhxnsXedHoThABgqaXgxyQ/ja6Wq4t/7tFi3qJwm+I1Ox3o
AgdWs6IEr3JQdS/RJXH25ZEH46bx5ZiPIZjoqEDfPuh49H4jsQJCY6oTLRwWpQeG6Xgll2NJV33B
cD3/LMWXg9h05zvNZYrrSOlqgc5OgZhJ9VtP7UBpOtZe9BdVkr1oR22KvbBqFFk83D76gUKrMgK5
zXiKCESQ7AZvT3JNxgmDsSrwmn3m87NDCuNncvYsJKlkK60flsazHn49IMBWhBFyB+xL1824+BXq
1ecnwjQGMMvBrgdcegebfhCwGvI/mWuv7w00CjlFLhdYvhXrKfjWLVrF7AwzLzBIOqWYXIK4SJ3E
Ct7TGAU7jskM+E/wlnTdNatYc+ZCRiRvPeqX60SWFHj6dv2cC9zfon9g+l0NdKwrb6Kb55mOBSt+
FHpEbbUPdCURpL3ZSsl2pRGRRjEhly5igNd8HjWlYpbb29dk/Koekirk4Ro4O/bls0WwBGtIh31s
pnLoMNBTQe9Qy5pWd2tFJqOCEIhYFQe+rA6Wz1ldVUWzx++mwuINwq4YlVlcCHYXc44hY5qT7P5A
GSBdaXQTkqFMHidbEdiYYT9I/bOP009f6gWNyV0+du6tfZAdKNBxaW9yxRrX2V5gLRzcO9344eU6
0S3CvM3vlUxdhdU733AkaKhIfniVGiAnwcAs2iqB9WYlZgHt19w9prmmdj9uWM2+iyupoRD0Yl6P
uFHkdYwGD6vO7OwOxegeAiFfmkuWf2vP7I2KR8Fhtl4LROXyonFVuoI0H50AT+JmBPo9TZlSp1F0
X+23QayMn8e83ZaOO0j4LzcHXfn9l2cIpp4uiLKLr0WCV3OCCB9KG/fZNBVW7xu26vXvxmdFJ9Ve
OleHbbtF12BWSetpdPl41egk05VpZxI0xYtLd1zwHoJAaRKdNL9XD+EM49hNR2Vf07+PAkEU4bnn
6PWgC9Dt3t5J91FOgpPfJi5VG7RKG7lbnfd+rhzPBfEB3QiTBCULbrC1qtMwnvvwU4mb3tc3oJso
N6n69j+gUMg1Let4Qqr705L6qBg4L6HqiUDumxPxVumySn5G7/+jBpQGuovL2mZ6bZHIn+OeXRg5
8JMVP3WyzTtqPyMHQKk8kMYKAeevoJKeJajuz6pWEljGAdP61o5brB8C6kuEXS7HLTovAhIEBFh/
N2rrcJgGd+hSpjmwE+vk0WBAsGw7vm4ILZbmF5zhWzORkkVCp+t4wzFnR9tI9LV+bWfP1J9wmU1Q
9KXPQeSvAyVlTiHuQLmGxQtxWC+B8acgL6HJBHH27xaLya1tJQ4xzlh/Ui/Qt78kG21kOIfVRVkS
62nEHqaVhQYeMHAxtALN2dcsLZ9ilnD5H9Xx22YrM664pGzyEvuzLINHNGsHo58wk6UndhEHENgX
e9XIaXDfHaVe8ch+Hsp65fPnQeoBvyMxQcTVJJTPLmIQVB4u6WXDk/VZjXmqow1IZMPsdtNw3gyf
WmIKMyufAE25Z2KCEUEzj8WE4DLi4PwQYz2lftby2lA0ekZAk6a+EbHDPi2J9MPL9VmxzAq7noS4
sXYeCdLFQbbFEBthX9dRaMlknQLKw4pL9czbRYmm9/OQLVuyxeRQveqzXs/euN4FYL510i8CtsCp
M6w07pxvGpic7gNdR3PqSaYjOmq6Y7zP0YP/jzMvwo/aTnkV2RtLShbVCHP4n4iZ9KIjGksxnilM
Qc2pKZByhycczerGioKz9ovNz/FFdnqRWP4ebEGOBhqXUpSGVVbuX84MjHvYf2l9AkuXV1awquYQ
3eUG280u4PyK0ffxYRfkw1NurrIM0XYsvoK5LKWhmybYzpbeuUHiK5fumhCGime2CIWU1rdSIcxX
9jWIkLO+f6uRqa21o9zplYW/4cBK3i6lBR//a5p2Mo6QK2ZSTeeYuSEgLjfvstYYHqu+aX/t/6pD
XCs+sV2Im3z68CQg9q2FFr2YrEioBMVxR77G/FBqirdoy6TanHOANW0NjjT43br+j3CCf93t/O6p
+rkAydQzIBF06SHnCRm3zd2OhTKpfCGWt6dxN6kTe3/W+nzbm7F7FhJlk8epf4RpMkYZetBkTSgJ
5mSAEXFvH27FIbt8LBSt9xC8OEn/dfYsflXeBhtLdEwHBMBAjt9hWf7jKTbKzg0AaDUjVLN+ZK0C
2UPzIz2Qcfdf3MKupiWIepe3dF5/1Nx02SuoSGpiFAmpJlceJ7Ym4JDIlq8ypGuxyxFj7P7FIYHZ
ah4az5QIn2njP5Uil70XYjgnU49yiz1IWM+3hWp5yz/asWXbVeQRsmqTra7eHllfb20B5Sy2WwJK
WcekRGGQC7VWbToyGPWxHw/HVWaQc+9Gu2IeMGZEaQJM89bjOPy5lbRFdvOQzjgKNUO/yZx9xidi
4Gk/RCPQzNFui+IURlr7pkXWwtVFVuhGAG1voHPVe4hxOg7nbl/f2mgiMxi5ue0RCBSM2AIyKjD8
E9TZZg/RIBIGN+UhSCmnpHb2eRJkaexCa0UbhN4RJu73grHmJqdHA8WiuUMHec4wUYqjVp04kxKK
FY9rTyb9mm0wrhiu4Y6haMeCQoxu0/B75D0I6jMjpzDREs9Da+0zOJlxjp+GRR9+aOAJw3KeiMw6
rkrfrsKvs/ASryJt0A42PUDFamA3NPd1D6nHF6N8i3CvBy8ZcL6c5CzABFbXxKdKk9a/qFW4YcbV
WyljiD00bwJgUF18mtDvSzQhGfkDGFHS8t5N6bZL0EOK3KzkcgJRujloYd+N1WrpnJPaE9yI5U7G
rgXPn7aYLMRGkM7+OCPOcMpcobtuQ5ZFplu9cmU4iumwL5J84vwZvu30v2NfErU/vN5TlFr9HzVq
vE6MECI2yLLnD9pcGfeC00N3rXP6nwcjod9qBdkaA6Sz0NWFwcKNpV1WA9inSg0BL4joffPk16Fy
9T/L8XJEMDx0jkd8Mm7sNxoJR87cUrl7UoYYZhD8KhPKgqc7S+UiprmppbHACnQ5pNHEwYk1MRKb
+l7WodC8BaFmiRYjgChLe9G9XdxjRUd+VKlj8pWB+a/uXSjb189CZGDkWyxTQGm09NqOY0BhLYHI
owjAfbSzMFTyb57TL942JrLT01BFyt7DDADFQAN0sPs8OciAzCzEv/J9C9WRRiY08nJpODO51RT8
7mnHuoanm9TxKyaJkuTtYB+JxsiVi4d/XxjfwNbPsFJYaorBCOdFHhyB5wHabJTm880GRpZoKXgK
X7Mhb9ncVD4LAb2iPkiiOcVNZbuUj4pgn5V7eEejcEb3NL6tKRJs8WcTQfPhc/4yJlV1QD6uZBRR
8grsert348mzWGP9bpZICgF8msX6zqK/q2pR7YXqBYMWmcMYZP3cj4hSiu+9fdpP3X8QwM8tytYj
hRhw4QmOhl9wUZK1Lpm4BF3sKbEJ0fPJraOl+xNdblB8bywNCKqCSEez594KE9eE649koTEOctjY
ngOIAD4YKFr1gAGKiB1YzHYbKM21rHvgkTt9n4To73fcKSm5ma1aEGSktqV1IpN9FbvjcumYCi1D
jON1YzJOlF68+6o9049CZ9BxPf8hvDDlLsWMoaCmMjqhTQ+axxbTgDUn4kF6lRUqCVyds/n43J0f
k2ikoRAfRjvL47DH2QLAJPFjDRypFt4NaepHZzZsuixuBqbO+lx74doCdBu5WaNhw85JMDjHojXr
49teSjUBtmVYnMV8u7Pb8hwPRUvfeua8afdovTD5m1k4l/YwNd/9w6bk4ekxTj5tXbwvEl2p9kb1
KdPj/81o/UfI7LFD+APqln2mueh0r9ha/g35YGdaS87juvowLH8D8cLX+y79FaalJuGgS0MgBKlQ
RbtkUExJPqTWOGAxd2TBfXyU4wsWC9K+WGm/oc7G8zJ06FQn8V9uh6YEIPlwNpGmrnDEp6kMC9Eu
i9vBpHoLrK4hZdr/HyVHLRxzN7rZca3XJHZlNYdt79SIYkT5I2hCebM5UK7yw5IZzdum48cQFbal
DkOpR7go0poDWGkgZ78FOmP+RX9rKrAUBTol4xZN1imNWHtxFBj0s1MvY1c1lwlt2LJK/FGW5ctW
RR07F4AJ+Be9o5jzXSL+/lq5FQlddBtwS28x4e6uvLOFYJp9hEjKXvtoM7vlDuv+QjpgGRl5s/tu
D0C+MH2KLukuVKqa12WC8MkpgeXoY6PN5Vw6poMvHUXZcawVi0b1kGWtRR2YhuCikC/0d7Eb5k38
UACjEOInI1yqy6NjqwiEJD4MyqFgKqG/uSlOGhGwQZH0azI3G0AgNfdQ0/iyKY629NT0KrHuVggV
MKQeUXIRmmMj7qLdC1H3OXYePjMwY9RXlS6iMfbpv8n+Q9R0Ys0MBWNq0J09ttuh2r8v7Cot2AtH
FdTZEwBtA5q47sQ/6BZeRw7S7SdM192P0opS4keoZ6XPwFPHuSZyTseL0JOQDlLpmf4GWk1m9fqU
7TDeSGgkzd2OIjkTeSdMBTJiT6brmqyAotHP5q+TMZfL+woFj6dhQIjsdlr8p672w0hnDiFfYb+D
Alc7rULIkOEd/5nekmrTAenb+Ec4NdK8mLBgvBVNx7F1LIf2Z4+JeqlhrnLdE0UJhbNkDuDzFtiM
n/t168EqYx/inlQ5kGSe1NzSe1cvHtrUEILyyMWj7OjuMLuKbP2VFUHYxr+w0kRLxbtJilw0s69n
9rufHIfskpa7mt3IHXEWD4lEc2XvfUpKN1T6X4Iz9u52tigsldfEMwIWwTKcNR0On6L3TDmYQtSz
2mNDrPBGOevH9mqxV4kF6EgvjKmHfEF1B3cvEkbBxOoxp3jcHDhxtFpx8WZ/6c2whprEqxaKwW0P
oc9yUfXA1gaBJMpkrmrvt3r6F0tdMvw0Lsg3k+dpthmn/L6sEQI8YnVIRehsWlTStAN4WOFLL3Uv
2KZSpt1zr5cdWUyzSU3zXy/9iG/CetQhX0GoEsF3pp/V6ecRCRexal7CsLUc/2FT1kENS9RhU6L4
RYgaN+GC/gjjrZyE5Mb7qdnt8OaGM6b2E0UXWpWU+yvJOh4RNHL4/TUcdixeTfco3n8aKh6YDxdf
AXCfnczg9Gfahr1Sj62W82xGJOXRczNJ8AOeOa3Q1+k2opkt8jSfI1Cjr8ontpZPn15c8BndeUJn
9WI81jraGwMZ8pSSTbWoNGaontgzRa44/33V8Fr8WlTVX8cMvLX9auHjNXRPfaeJPCcQnWn4Cwq+
NMz9F6zOafs+1mCUAFg6dvdjjxXeWHTQ3XCimSmZOnQbCyg5nkgX/m/qqV0zbtMiXpJ9ImSLn5zt
P3OHQz/5KO3Gf5VJow3zvhvp+SsHDAFH6EKozkxp38+HM2wuvnQrNn7zAuWcrRcSgp5qTk9mNZuG
cE5Ez8T0KAC7+mqpAqsAOtJT4TU8No3lIOtO3Ixvl9Vlwt3RGTKuEB7Q7g4BtmKJw92oq5JeKeAG
I3MOtjHYO7+il8wr45ox+mGj7k1ReTy62SIln67xm3qmJbrrGSwvN07xh+v80RFR2rndmZsQh/8Q
zu49O3au8fdA7Jfd/V5yT3ojEOOdUcLyO7UaUJ7qH2MRgN1roEcShdU0XeqieMhOjU37WwQXoLWY
o0KHEIembE5+fMZQpuxIz1il2KHTZ1YAueKkEadkQoynyJDn/quBzQQSRsUdAXkq8g9HMeml41Vg
JnRzHK9ZOoeGvmdTD/hLtRxDJstxi43NvkReMvdr1nUF1oIetxYvl4fEYbjuF35XpMPATOCEN0su
kQa4ESWlOEaZ1daxW2/3c8WAq6fYo9S0EhX4AbGfSGUJPWI/g9zdkTmzbN/W01YopTkvzK22SkRp
XDPzRy979W/EBejkIqmokJ7jT73kamFGKKGTNz4JaHvJqqzzP3eux4GjCOPNIAJOQNdIDoLvYnRl
oYEVxOL7cAwo9qEa3HB2lJp9L9mCPd0/gyqRGHOUyQVaX6uAFiVjkhmkXKT/SksPRaok0xm/Zf5S
50dEnP3aBohxry+67zgZr6dTjrUxzWjjZdoF20WbXPXluIq1nRFnDZX8mBXavhEfyixT74Y/NkbC
uOUsd4mPcMtIzc7rlTIhbgrjUkbLB3Vbe76ZO8aS/9lJ7pVGkBDdudDYp99H/Pt7VirXtRWULUbN
GrW382bVzk1JrP/Mek6+sam4DCP8sjwRYdt0RFZe8ABs4d5nPmCfTJTR+XKk5qPVYVdFBmnRrxhd
+RZ6VZd4KuyGodG19GO0ivJavXIHcrSkKjHe5XcW13PQiNeJEq2OaUmCyDQwutL1iuFWGyK7lYnd
9DPGKrB8m7+oz+Lxhp/YUoa2dk3Uebw10/5aZS4Gk5NwfrviJKuOs9EdX0M+t1KtdD27bA4lMYB+
dOPd2rb8DbQdsVEBfU3lYO3yVyAB6HMumxcxgLEh+f5F6o+L9Vdwqa5GSM6Y3TsHx3F3X1Bux6qg
mEdjMu0GAXoFrfSoR03NELzKxRDz0dG7iq8G1MgKBwy1j6e9ly24rbWkVRm9a1T+CJ1wzQlFsUCq
u66FG1mN8ql82hR0RxV4JVsqsx2Y7vKKE5/LRcugaDRm7ZqA2qDOjRVz/5DeeHXEbKvXGBmIo9IW
mOJ4dGztcfhykABLtkYLTIc0WGlT3Mug8deVt76AxB2Z05HeCPLzo3g73OR+r9Yxw/y21kzkM1jo
kpY10+2zlYbbEBYrTLQ2ni7arxHd37JvofQcgRQU59b3iks8QsyzCKywuBwpel3ezGUNglY4XBa+
0DOt2JsR1+DSSb7sZFLkJDktjm9tiL6eCgkAn4vG//82zvLgHE+ZLltx8XVluUg6JSwUTEFd/58r
HNm30YXBJSDuFscnX0QzQOMVIbHpGXHdthC3ZaJRZXM3w0ViAwXWbrJmD4ntZx+3X0cT0lvyebT+
UwlTN77lrQ74RbDehGKkPHxybGTf5UHuEUh3QJaHMq1t9Hee9kl7wCnleQoIkPu2kwfYTUBfelF5
LLKcqBk+gyP2KyQgHwixsqAFs7ytsd4xdTjiqADT9bVIpGPHzQ6QIMv+WOBIUh5miuwCAs0Y6ltx
sjjhFC0HZnLm+8SmzIH27sUF5Qck07YaTN8xnnP3u7WC+a/DU+Nw/Tb1kWbUaijud3padErQoOiv
DeM+rT1KR7zW94BX+RjKs1zbbY0wpYK34JuRATD6Hrua+un570L/w7ga3MFyxlXSCmZEJKFmet56
8ZDV0kBtiwiF18OewMkT5sZDn1CefWrIyT7f4lIh4W5QtU0FUQjSkeKux9gQfLdknoDuKp2UwF1F
qxNKdi/T2pbWnh2p48Bns1WO4146TSZIzUx0d4N5xdTXuKEkJjmnRjjmTy43phffgkSUs8TYZ7ff
WlVRuoiV0CcfjuPdnYZbhdE+3AC1/HwJNTv5INhtyTqXFvqcEvgrEIaUqDNuTs3zb+7BYAeRCULL
0PqYGeDQSK/idp4Ifr9PLhhuoCsIyIXiOPfErK+ix8ziSQNpIsUXt4mm8AF0CIS4Xy7uBe/AnMhV
ofIV23nBwrepmhCeXYQMlKW2cBiFCJnn9pp/n4ONfLngwvEPZm1vMOyQgj5BVNdIyjRQ6GAVywcO
QFPiwg9FDEkYibydtoTri1g5lz/3asAtswUlsruEVXdpTPHor6BLwiHdhbZPES1HySIPpzmMruFr
SeneG1AOsSoJ95Tn96EEUM8loTWyFRT9LYv9CovhLAu3u+30ar1pzQveqtS7cUmZbnHOrvJXx+7n
FGN82y0KqndVSyODeWFMsBYtgJx4FJpB99fYdFKkbdHg1Y9VHUK+kkfTMA6Xx6meT/6GligQJttM
ejM/WvSJFhIlCwbUcb/aUWImy5QDtldIBIqXiQyD+tueibTaud9JOGFIap2SKuBOBVmAnaz1U8U3
ULnwODCuWnHjnY283KzRTf9GbCcB6DM1iCa5DwOmyOKVGaTCdWwvrDdGHOwjcH0gH2a9XFEf6BrL
6T82Y3nQv4ZuD0lIvzX6dbtB7AeV5u41OhoeRGcHQfo1U3HhsLm4sE3/ldffeldKmW6TVZYtJ4xl
2Up7PsgKE0KZmMJfJNHzKHMY4RrMBedXwYYIU7kCnvmfSJtQFSTcLYIeZXvh7HuHEbRTpkg29vv3
Zrvnsm/i9GFN2B3SCjBctcvhzUNADPAJegnBmx41K8/HH2xmBCkt1cWOJ4lbE2ESOmFCxgyBrcOC
ebJ9PrToKRpdsuZ6HB9+QCQ2BGzjV48AEwq7TDW1MY1Tqi6d+AvZ3hSFMvGoJqV+O4NUl65fwBwO
ORc2vpvot5ulpMDVb3c7KHDG0uRYHMHJRAElCa4zV1nj+7mOeUdj88Q2Kbn4ZHgETaalGzMoeFZW
er/yoeezOVICP6YW6l+/VBvffOEmusirbUGPOCSn41U6yAV+CZ7WFK+jwz0fdnmnwrHT/RdPaPbp
3CC0kfQu0bWjf5RjneYp0CJd7xlQyW1BCgrV+sjf8eDPHTLLSPYUxasuC7QzcyhjtjgX8ByjtMK5
wvJTMwciJSfa/Flhz+gPDegHLMqnzhR84TmnVUvXON1DUrPpIMExhNl4vkvd/zRWqgZRo70aKY1k
R4b1lUK72INu77p9is3/EqBJgGQWnfb53FjpRWf2VGOLtw+ugu1BEkoQr5YgxEriNCud9IwdWw9G
tjxebopRItw9XbSt/2iKERRajYsgKKqkN/HzhMrGQtZ5IYQnAS+PpeqSlyvwwpXoeR08Wv88Aazt
DvbxaJfOIYP3l+Fm43ZG6nWAt1f63cXPirDUaI7twtmdtGYw8yQAwkcLSJxsjGueDRVUFierIlAI
W7wBKetG4qqjKWS6an8PLTgPiZYCCoDNofV3xKGpMsJYM/MsIEgEoGrQvsQil8UO0rRMeujIqwTi
XHkeZHhLdOd+tduNWr82wmkmQITsqCrG8hf3L9CEkcmBhf0oZ0KqHOjHxKE/iTp7Vb64ypZLuVdh
6P3GMwgOPP6XiYmr0Q5QsDNlmrYLMaJoV1if0LFXmliKqFI/WAPIIOJcsg+b5+keojSNMkQ+J2ru
39zgAncSTP6gerFu0p//YL1xCuw+bgtU5GsC4zxrnE/Es38A2ZhwMyX7kXgpDdIosoeji1mCcf0R
7ofuSoIlGKAU5hhxTp9xa5bdMkgU3cpU9sPt9mfuv60deZ71tnby9UHdrgkdBzZqrtaWq+iQYEr1
N4hc23FOTSLmTPTM/wHcQPU0VFCJXUCe4kjI4/kUTR8S4LdS0HDKfDAareBFJ2Vh/nFFqQq5zgLW
mVRrKP+1srcfheCq4w5u/L4lBQ62e8Sd24iO72l3k3AG8ub8TSiCmF5DD9xldxXuGlCGbqQtwP7U
FQEj+sYgDu3jz9YAbw17EeQglPGrl8D0Q8H9s9YoxQUScBiXGaDvZCIKh0bX2RqDMZbBD//u7DMt
mtC70/WydxVY2RZYEKp+oSAfaYFbyyoO5PUTAtVOy6RenivYdjt/6fJr166NBlNHwOAHwGLBjUld
GC8ceHJhtJL8+uk+cfQxHzxfLe/+q/EPmnyfzXdw1i+fvjZlSggdZR4IIgUi8uVX8QQZcuBMqkYt
fSKy0B9K6Xk95L4sVrwUq5XCXkqA8qLWJfsFs8C1FVwQgZN+UhkV9get+0/r5HgDqawFSjjQpPtW
QTOZ0/Ibl2BwM51bPptwLfUubjIJnyM5lS+zfjlWg58N7iNcr5fS+uz4h24qxzkwKFB7dtR/Ross
P6uba1u+ganDvCevJ7JXnOIGIi7r4TMkgqiTZOEOdHi46hxSCO91BkLV9Mt4Xf4vAtEc5anqlc/j
oj1X06o8/zYW0iprM/P+g3WIGAsdrsuOWNyt+hP85Z7BUBfwBG+GsxuJXVEbNgl1K38syOy3dgIh
4Vrpu0WV+mNbZp8rEEkSm86MjgDGgV2QAmfVTd6UVA07T1U0ndUi2g3Bp1gpYM7FVEp8Gu2qcE4/
MXOd5wp4JgKNgIPKJaJOTZMXPXZtDvk9uierVJRFEJlJGncg6UbTo/2jAOTEvXg+Rwsjb72iJcoG
Bp+j0QzTM/LaTr/jQlvAWPfrWg1cVf91sr8eTTfPRnwuWfb8N026ccKPU7H5BOsK9m8GEta7vLVK
2PuJt5x2qbuSneWtTw866SGqYiSFYzLznj1iRsjsTdcqpMU2GJN9pY/QGXeK7dhCw5h9qbifSldH
B53AMMZxzAsgFh5qSLP/X9GPpZ0sJjbBRwnF0K0oTe3p5f2vLsEDO1ItFA6N/dnNU9cVjHFLEj6s
UDJHPda5wK+7nGC6HB+K7vhwV5vzzptw7IrH7mjmi0KhU7qbABJyXSNQ/2FjTG3RrL0Wqg3EYgWx
GSBMyg02tQb9vqlygw4PTxjJk94ahivUq6oTPBFlMX2oSnV+/vdYPG5t+LPFTa2hKks3qmpQerP3
5QQB+9wtW1Ti3Y+Pcyn2ndKcbQaNuX1yy7tihpK6iwrqNKlb4tihhvjwxk6cUvSlYODI9v+PxQ5r
6g83VaRAjFKEdl5Kx2nhS0mLv/S5iZdVansEDsuDpVM2KGLn+cBaEE8g/apNHybfYSHiKGOk8Udw
8zytR2HlvT7qaQ6//8qv6X1BWvjDk+cqwf2/NTJLKG2j7h5MQp3VmdSzoJmuc5RJP1tohnODcdZE
lHqm3wR79WcoYZLLVx6pQQ7iTXFpHaPTTBYdEaI6QnWXkK5t7MpwEg+8tDZy5iQk/1xJmwOGxnq8
12x/5Exjn1cFBfIdQd7Wso0D9bj+JetKJwo34rYHmNbECz2exx2yT8G0/JYtv/iRVnB8ppERRBgf
L8ZyXmbfb+pMdaikVE2zawhqX5SSw/oeNqCBjDTcmWcWQnNnMFwc7LUaI+DQCvd1DPLLD+mNw5pH
BOGtAehuZJkyMdYuS4G49t1pIwcqKP+WQZ8phdpNHRbBk07y/w/tKVPgARjU6TZmizw12xFgnnv/
vyoVivJL5uwfECce+5JZlt5uTLiIsdSX18PCfFStdzWu3okl+nBqOfts3vBIWQx0MujB7yiBmhSI
BIiQ+io6W3HJAZqssrYuahLMS4GCyVEStTaXymcq8diFCaYjw6tEh2VTH2nPNHuiM6eytEaibjq7
Q30uNEu6VCfaL/KVaoTaZNWPZhplgkTpIaRXltmKuc/wSZMS9cVxo97sWYh81JVkzRdqjzy5vmWt
4kz5rmpl3jKF6HPQcoZfleCtdQ04o0K6s9Vs0ezbbmc8KHCP3z/viQrWyAhHdPbvSvd3xJ1A5Kpb
LENLfDDEowj8WSm23Frf9K5+yrWU5EqVqAUq3kbnlf1l4TpJ4IGoBBfHVoRBcqW6Plbn0H00zKhj
0nK20u5HFY6BQ8wsOlUh5/zn5KIoqoRZWGJIsUAcgJXEwXlrxy6/XzCh5AGdmViGCq0Gy9FelMKO
9ttd3k/E8GGVPlKe4FATBZaJJY6oXeXh3ZNcFRT36TR5cY+qaUXKOp8ylpdZaGuKfHwXIPNV/i7+
GNzaO/Zk66a7wvgFakcNph2bdwVef0udetbixkKlVGLz2Q42Odjvs7GcQ/NcMR1B/Y9PitoIg/Cj
YD5guW1KkqsMwRDJdemZ6e2+xA8wSye/S+UzNeNDahJTFM/cOSwDfN4/IRLVScmrR/9DYhOJGPeh
uSB3zUKrb6PYwOD30MSEhAbUPcGIFxgOFreEqvDwetQX9Wdbqb3V9ZqXq3hI3z7KIg6CK9nPRhr0
uanwLT4iTaKz1C/R91Tc83pBUGjHVDpfX2aUUDBO5NnC4YFUHECpfIy+BWvOytTlJPbE3b4/v7kc
D+Ihb+Bxf7swus7akDA1ha+Vg0sX9LCiNuUaDX4ioorJ28NGyHtbs8QrYyJj0BmpjzCXYsyvfC2s
g/z6BrETRL3+Qeau87jb5WjZzcwUPjPajUL3kZn1HlMQqiDG2cJo6uj4a/H3LwRA2S8ry/MkUUgT
AI9FCQGl/1qoK5aJJhpOsDD8Jd6A6YG6PV3fll4p+U9TSFlY+0g6Tsbih63Dox2nz3VfCf6nUvVe
+j4s9hhHKw/1H9MpLP92tAU5daE6vv0+OPou9vX64ojpPBoG3B4evot0+eaPj6rzJwQNXw5itqbf
FIVeDbW3x8jGTtCAs+PAaolkqDUPgY6Cforwhe/1Kp8n6N2xCeQTFi0as4mk1713505LtkCHo6XQ
/qeI8A1LAtFfPRZPCYNsqWnV6KSwP41Upb9tGIh85nYNj3n3aIyA1CMwkqbdxg3O/c5hCp/TZqZD
3D4WF0EwXg9V8GJ/Zb7l/2K9OT0/erc0/I28Pn+QWo4X/iSaods+CxAEgISiY4pTeZIYTJuQ3bQV
PUnX3GRVIfzYvs/UD4MNXeRHexpCTk2wL6/8nOKDyOfIHSkiS0Y3Z2p7AoxIA36rZED5d4q/0FCJ
gbNjhNtUCuggsAcz8KtCoW4U7FYqzGo0bzdEilDdureIstEyBEotc+BxXMoyYez49VB1QrtptXAI
A2hiHZ+eEsMWLnUVZCZqqDF9GOpK+gJ2ezshW+XjbGID6TgYd4AQOShQUTI68p6XSqgMEKQs3/IJ
XR8Jy1kFhz0gOHosi1YkU6Rk3Y83ZXXVcYrpG5duCps2qduREXfpAacJgQWETUfAAHMSmC6XTCHn
+xO+Ii5uA3TCh+hV1rflPQ45PwZa9nlQSA5GOGEGhvhdQ4ac/wgRoXOSWIIDswlLprq4cJN8xgiV
bs4cH/EaSI0Tf3a9dyE9j+Lar5PiQAc0+vfeqb5AmYpL+foqU9Q7l3114soD0+010HVPi9NTAngT
jB5To8qaeBdhzRvJOwDSWcWIqcBpWSmWVO7wg9OrTqY6N/FF/tNbr7mKkEKlxhSYfEBpHs8vveNE
Fd+depnI7WXhfZ6wWn/9gOR73mx5EMjD4EbRY6YJQmqtPjohNyPdbF+avqQV5LyMMerM3hfh2KcP
Y+a1dAnqeTMLo3bXsGOahELyisGro6jcrRVQucJpG1fuLeHZARKAQYi3JR7HCq1b9/7F3RuVJD/l
fvG2OOCS0ty6C98l5XWq3MgPkpS4nRkY9eGHwpK27NLLuixbARhqPm74POWdkDEcAzRVoYL5uu7h
W9OurahkEq/9HnWt0sqFExsrHYx/nJMVznsdIkQy8vzwatfVe8Be3NnMKYRu7b0ezpmM2PHMxGyX
Lx+JGOXwjLc7FwZvUHTK3HUl7ZU3obmOnl3D5wVl7HLsvs9O4Ama64iVqxb2kG86WlpGQQ71qbfe
nGBby1kDXjnvT1JplWiE/iSse/tsqwsJFM+rUoPsVW+hwEP+e92dWZQxhlpl6sPnFOKz8mmTijOD
Fq/agcRluK6ccmK+cvvZPmHEicBJKcOXHn4QqmxS9KdygL9zY1or9HfDpNYVtPUr7pUDw+V5tp3n
yxR0XpMLxitPREvsDL+IsdLXTXv9mr2cAO+YJPzo61Rd1O59ikZykfB+9Sg3k7yF8qfOVSZj6KDR
rfcwQnlj2Wbmrn5kb+VidYO5z2/8uk0vnXH70e5O0E2hnSztgS5YzJpbw5oxn8OipoKls78ctdAs
ccQl/Qm1F8XL5aSWifg0/X1tKYK7S3rUPpSTwkUNfi46ZUlK7u5XEFZURx+DTi22d5MQCTSN+R2b
6W9ie677dS1HlIRjcFFikCsirvqzTfTqy65FGWalfy/TM1o83iGx/sa//gHbnARduJaNFN0jAskx
HPSs8njHIefktUtzRl9JEl6A9aXI/ZF7fjxTHJp4DVXqQEWn8Fhr3THli7xpibhBL7OiQpanuri6
yaMwKS5GyuWF1sHN0Zh2fhzV0bbPPuL0pSoKsMPdkEJ0eGB/Cox23AZPP2GaQQDUxfD7FQMkh3wB
MBIk45O7rw3v6iKULU9j1MQZ8DzBocFWd5uGc02RJETtGEMp++/3sc2DZK+imQAJC5aTh8jkBvLS
cnbk/BArKoIwQ56eaOHlUB1GNPdu60/nYjjWvVgnv7HpMuWXPlsmsgGN0wm5ZT2DwScsaGryXMMB
SDu+6rVtvD9/GzPOx9oGi1vfErl53rTC5gWCHuXPzkgozNzs9uGgKdrRKf9cT2hgnMNDOBkMobRf
/Cg2FvWx4NDNunBm+QsBU8PNxID/S0+5RYhMayA6/+KScB+Tpe7Eu0wrDw8IByN2yf6Joly4uQtc
HEfaPvuxnOR/xSfmDKByPAcZgPrzwGmlRrcoEU1bW5ws3EjCaKMoqbM5LfEZoeWiNeme1YKbc8kt
LOoY9rBGU4AnADfqWcZCQagS9e2tVya115hMOb48R5Gc+8QNw/zY7WiNRz6+0rmFLAhh205hI+bp
1bauFkCPqvgx/9J8OWE9wTCZydJeYotvNzxpW9xrwGaAta7EQgvvSEe+KFE+zkwpEQKcU+A82YLd
GuJSJMokGP7pj0uMRLRvSuUoQiU8s281hRvKChopuk4fTzgRB0TddL/XgHog9e/1r+yxIkfd6OBO
FW7ozmW3RUIsOy5MKY4++NlcBWUYGfEjF1dzanqNi1qxLwzQGY+Aed/NWVE560IKvX9m0m1dwvrW
ZUrN7FMxcMU5ZTqQEhrtveokT7wTC3QolVm6737+G0IZBAru4eXZxuKUNHKZ9qNIemZQAQri7jvO
7dhYfHPN8BvIiEfkbWgMEOtbOrvVgKh3/zd8Up59TXF70OLcRRurM6OBdwSlhdXsUS7gruP5CHiz
04woEJszsA23mDd9jozGlBKuq8pgUV491XYb8YQ6keDN1LJCG5zPE2oegNSDqoWfunfFcpBQ2MUL
vTuy3XWjkAzMJ7pyoTns2riX2Se14gbPaK+ueEmIpei8v7aQmUSXcSGthW7veP7kjrET4vZdD8fu
5dlJKLy1NPhOGQ7sedb+ozhoSN7J6f6M70NOJG9211+w5TVDh902CtYaXeFCubO4pTs2lWkOMfIP
0LmtnYSISNV4GwoUtAWncduq0Y7X8p4z8EnCEp7rLm1sR147QWcJYTzijFZnEbdm/UzXCU3jhNtQ
5XQet+dafUpJ7dGWl65YqHXvbVVexD+bbkDeJOfhOROlEPhUfBa1jvWC+H+zR9UH/lgDUPyCGXYq
6OdTYk+xIs4rNNuHS75nWTqqMc0flqm+Fi+e9Yv4Qmuh/WAHjduLmWrCnJDPT1AZ7303WKrqy41K
28zNKmEw3AGT6iMPla5PvWAPdnjl+MHTYWDsHI8pxOTLDxeJcKe3RsIM3PCWaYs2EWa7aRvlMEjf
TpZHnn2SfTY1FTOJMVduN/uCouRMrk5ZgRODBB+WnGUnwKh7fBpXtsZ2SdvglL3yRDSJjWmjpE5u
WP1z02uoD11r1DCqNXMqskW/9HCpC+uX4m3C2onTm0kJenBCRcHWJVaqArQQpNnDk4HKUYlPBBgd
WQdRapJ29KJS58XI73HHWF68sIaDDoZ26M8HDhWxMPaQnJTClTz4osdWmrjRzeTvOjwE+i1jEtUf
it/dTNmfHPW42kkkOH/MVGNRHZfEBvNs1oEkYLkJRvKkKKflR5RiNAirdjST2WyM+eqEX2u9yi2x
lMVdX5DEACCwvlmdiJPZzGJ+IfxzDTuaO1cPKq4mEQ2cExVYOpgoQstqedbf5kwYUO5p2bgCVAHe
Jo5SoMLenHnF/RReh0bl/7YIFIfYeK6HBEGwOob20P5BwG2UNvV6qTMDQo2KAg10mh6P1EbhXhBb
IvRDqQwm9NicBEJuf+7qgASn6MLMsAxy6pSYyhp3Y7EvT0gn9YR3/Nf+2vylvv00bmwhdCvPKTe6
Xkecaw3MlHgjewSJ0FHej984y/oORCm5ADVzVUDNJ4jacD0lW8fI8pbPPMQlroumBSLBbzqqPd9a
MJ3uE2XuA6aiXR7PuMEv53V+R1hsGeWERX6hU6SWJ2nBnrBnxUKUc4KGfbxq64OgdGnMnGGH8K8Q
u7ob5+VZxu76qKvKVsk5/lspFDxcdXbwmLjHPdOWqgMp3z31EDUUZCeWB8cvofCe3YIg02x0XD2e
eriKkLO+PGQeFTptX5KdJ1SsZE1QALIJeYTwsRwdwaz0v3XmQ3VqRRRfggiAv6w3QpUu9XR+98hm
0OFLynfw3hwooiMM+zwENKmJpuPZCo5OfwYp9dLmtOg+8Ji19wEYHEh/7woUVXn2OfFjWC+Y5Vqr
pzICfIXdjUfxc6sFJSxpY5U/e8ImSsmrqUMF1HnFZdgk9yCGx2vFaP80CHUfEyVaf04H0+kV4C5V
tidC144B294xDgZVbNJp974187BKI7S3yllBLo5xiBa0XApmr1AV5iUHc0jCORnRX9MixNyvvVEU
QtyzZr7S+5jQjSS2/pVnFtbInXmr9qXpMcKidFGboNjGAFLmZRV+LWZclTJ0IVIZqS7JerUilwc0
/qrdtljqYdg6RUpnWeIDpwiN2cafHQ5szdECJrdHr5eXrdCMmUt5pRwwbMp3UaG5uIUDFQYHQodO
Zl7w/7MCGPFvbWSQEAV0gl7zi7GiXCRb8wOGUofQFb/leZluVmrEdpWPQ+T1pouyh6r638VJQZSV
hb+ero5j/UYOwSuW25U2krXwg3hjkPeSYXMM/iZmrRjYLsN5zLOoOG8tFjBEI17rWMNi6iL3GUUE
pUwVLslmIxJtan8NpE6wt3S3n82b5iCEANCG8naOp4lO8wU/dofCobfAKwcJYmod07+zn6xAs41a
rw+WqCU8ix6l1qRfrPHWoasy+Ti1AxeR7m7zsDHVbcvOt4C8s1JQ8wlV3xENbeX71KxfcVkJcObz
SzFw2MZlkF2rsEVw1ZS/Ot/ypoftjsdkW/xCX7PprSbg0NFz1PGy7UCZNFWkRQtkta8g2s0y7BqY
2ruixOfzVnVvuHY7JHmFVpCH0IUx3611KfI6JKNVl3mkgJlpp6QkwDu/QT5LVx7Jawcp/H96xX/r
caMuApAq8xQEAYBecKvc4bRkD7kDXFjYXyI4X/Hsj6Gkm4/2pfZ7LK7rQDJ9SzazwD6bRP6kkPDb
d0cqluvHqKt2Fss21xVta4oRF+uWmpYWFqbD0jVRMzQw8yAtwyTjCqBFiDTsyXI/RfX2sCA1Gy25
ml2O133Ny4ZREgy5NIBsVjORU2E6KOYrvn/3deZ+sjKR7yHaz/1pYrTBBKkPhKy+U5LO7VBt3VAp
Wpt3TrCfmj0+pcF6CS7ePCC++regqIiaHJufdeRX6itggDTo7xElVgtHpCdQXCY1ig8bfVBP0xFu
Nr0E9eO0yeMd055kzkQNPYIZJtcv7zxD/zyj6Qu1YQ589o1xJZXzCoD0sYGnaz0XKXtL4SpQVMaQ
thMKzpC2t8ez+FHYEcpC19u0mq6I2fdOUztn1PYBvnp0aI6j/tuCdh3bYt4XlGwWXeqR8I335pzK
tc2j4Iz0pzMRUc2AoCYvUXOrA/Wf6eQ3VIVEn3YUyJH1t7cJi82/5AAXvrK1YfM6zK/+2SHdEI1G
NW9DqVRMGm/ErFFfe5al9CzN9ko+rCU5rYR66BfWdEGrnjiBLERo9l+jzV2qHPgBL8WHdS+oJHbg
RpalBNDe7cU2JNMLZSZO7IxrWwtAPe5dwNk9Ee5l98ZPX7Gc/gUVPSS3+zs5zUpRJUfwrmFFetgG
/UZ4fqnKVel7EKGQ1yzetZQAmWhBh0dtEwNofETmtIrdiDmcE1tgGZMVu0y4rf+RNACvDcsS4yDI
WdWxwYz67c9OiH0yVnsHTvR49l2JDLio5RcN3OLQvovK+6hdCYVP10qoi+fpkzPoZcAWeAbi95Nt
7PqrPY5Dup2RF+LSic80KLWE6z+tVrFDIN6XTk+i+kPtc6aUz4fhCZRLs1hDP1f4szRUwum9KjZo
IPP55nAwx7V0raJLK9eF7ufg1zkA4JX9K/VSB4MxT/HjxkpeuFGCOadGr1X7OUvcUk1RT7LBcpE+
jVhvdiGsKcaGRZRd0V7q31E2lRiLj2GOjdhzP1ESqABp9ePC/MrYOQdppItZCzaSaamCYcEA2uwn
rxDzI9BS0qqpCCT3tlCQafe7/L2Y31p5u3bbYO2TxX5wKUZILACGG5EdBzHYHHb5EyWIQFqT8287
IsPS10FgS5o+MhG0kS3qVNrtt3k7EmUd9d18ZPNWCcm1XE7Hvy8R6bN6fG65j0Bn8IBIllZmQ7jw
JnWu87eJEaeLeIYnPmm3hUyeAxvliY7GhOrkmpzng4K7rmr4MfSnKZuW2pmZXYhWlCXEjmWcedSl
lgJw/d4qbrJyBMg3/1qDgYLCCOUMioaB8Lzfl80n+NoPLdsZb5Lwy2vUF7++DiSXZMk+oAzFPCUu
Tt3RizQiNX8LNRNrlbjk5DScVdjmsfxr3NVYGhM90B+DV6QUZEq7IffJN605kK0qzWIW2cLGTM5f
dX/ak4i215I+JxdOr7QuwRoGoLWZuVwz642PT0KSnk8ZmuGcXwmNQ0UXXUIWyOVD7JkUZDcKF99T
RPRlCNpq3slL6I+DPSBgetmVyksQG/RxEO0N+Wbbv60AnfnuvjuhAkNToY3dGI2aK0k1kr7J2eLS
GqHsm3L0/pt9vYhPL9GvcDD0I7WJhKUTY99H2EJhMsFUlQVgtQ7Ybiucwx/Mr5uDiTa7hf+YNfE4
m5zop9/EXMkiqrx4l1KXTWzCSqZRuMjOk9us62ubGmb3VIBCsP6Pw8sPbZIhIzp/Em22qeDuyGYw
aA0R0VfbEdOIUpts1cw2QWJrw2DNPODB8vQJ6500LA2wBwG+zCB9H6iziqRONg2LvuDjOqkQZ3IF
aHqw5aYyR80eUEUTaYsD4EZp2XmPu2B+CZp3+AzmR3oHLll3Fb8SukMUuoAl3miXzCjkOgde3YWr
dV+RgbZCzC1hOs2lPxIPGvqb/uqbqfxl+wUMVNd/4QJvaeT1QN5WLRyzEzkXUGJRul87kkd1E7w0
5jBhGY7tsNJ0O9nyMSblRG6XxmoRS9CVqMs3kjI6koFZF5wEb2KfmrlaY9XSa0W2FN+pTekSEZow
WeZNhG5ZzoJMj7TYh0rBjVZXidODcoNVdo8d0abn28mPKCxp0VjWyGPm/UsFuk/yNggniXkj3KbM
0xIjscuSGMyCkZ/xz1WKPJTwgNAIthEDXk+DvYzgvT5Wpwr8ZDhDJa3fpDR8tq8QqwJj5tt9uugO
2Lu4CSUfEEvUrvFRR7Do1vUVlJYOiMhvsF70NJWuZkiBxSt37BmEflkhCn2BMNe3ysmiUBx+iHUt
nyMQ177KN/Bh6awQUcbaelW9PmPRqSjWFZvUzXGkKPV/4npS0CWIj5pkZIhCTwpHPUnPvH5euIOd
kg2ow0uXo/lGULlNfSa5mWRST0Cm9zZmPMF1zO/fyvCKboTT+wOMlYVKlxFVEi4wW6phPtVFwJcB
9IzwxDlYogLwpgj7Vjvm3zPfJnIFhJqw+tYXwqnpeA/t8eLXoWFTkY99eNT/P6/pu+apAH22JEm9
qHJcDmeGAPpFGuGvi+JV3ZdrlLqA9L2oP2LMCqAx2HaVLf029flzzS4X3AlCjoArdYQleeBHJO8o
+fpjWeB3yNGK53mP8Vu/hvQTHcHuB7/7XET3FolfrbULANUnaUNNRKEDOMDxGpdjMDPIAIx89Z4Y
4scF8ZMm3EACyTSwj//RPpIZoPtl23QKXOaOLlaqDFFaHxiEET0+XMOI3oMGEWJsSghoeqvePE23
BUqMC5DhcDxPN+cy2Itl+/MFrZpvKZqEU+vxerQeOL3fnpGgmMN2dgltiFgSVtZFe98n0UTdFKuc
OGdLaE5zsCbEbkdQJBES94KYdRmSoFjdfxOuhzEzepvxAxIDb5AjcuTju+PLvCJ/gfFBe7mR3/kX
EABdQCJUKmAmjQ8nQVvMxj7GEjclvRHg2eVvkZGLbpQKNEUVHozo7IA7UYqn9erjv1lGGXI4kGYi
YjXUKGwN+RNGrmFhnal9b+FXgbwaCAi1bMDuH3IEkxu9Uh9LzVZmnt1YElKDln4CsbVlTIdlifsz
RPhNXLiA9Nbe28a0ATleGw5dnJYzvGkskBYv7hD6BEOYxpfGdrBz6av5d/lmSdbeRt/qA3dhDyTd
13BzuLcuM3t5y4X+AhxIDd8cy8AbnPJgvxEJ15HdEFwWEXq4mkEEknl6fXsl6PEcZt+V1JunNO5G
DfLlyOKSNGUU+VbMFAnsYUWD9t9qUMetFWHnWjunAssHJ4Lei7gAbLAosCJRdOjhUbuwifBOLbOk
VjVA7ILdYNO3ng6HTW7uRSmNmGWVtfGHo6yAbMaWIUN4omb/TzEB9R9KN5Nav+1vQkEcb8KnqtYf
pX+lX5rzj8ZgnTotLiy7ZV8GKgdkjImLu6AYGOKjo/X9uha3a9pB1tL6gc3O2prboSdcjGtzbrf3
Tg3p6G0R9Lgk0DQerS6wxFA2aNrdrw2mOE78IdD3SJNix+hvraHQdsZ2ub9krpdaFl1pwokTb1rm
WXqUIOE17XcR1FaBx4jxwvNRVmaf1GbUDjRCMjm6xRp8czK3IoOUCiiB2YxD4x+uJBEe7n/5URYU
C9BZ35gzuB8Ez5tyJV7nq2/mpZYRb9gl2JSUkfFoQnUCakeAQ9w7wtYmHQDqytMLRvLW2SD0kB0M
H3DDPuS1tJYiGP8szy1Nf1WDFZkDYJxow++5LiW5KD3O1JFHaGObm37YdChVUWtP/t2zsSNYV9pr
rv5lVIL7D8iWGcOWnKexpQkJEM1vLchKSESdHXjtGS84ZywAB2Vnmv4Za5kdJ3K2S+q+lfja1hzK
37b1dR2EtS/DRBhiuLI3keQHy8r35Auqtd598H8ZN3MeUbwN3tuyXg+7rQDlzQFDTi3k8xCqAe5E
xDcM/T8EykqZtr+c//87Z8kY4falBVzWpKmVE8Qkxsr9l327IhW1xbaXScqn32/mBJ1dR3SV/vmW
N3JUG9493T4UCHpQbgL7417y0dcyveH92PzgA2pM7lXlJ47kaCR7KHt3hJX6lo7aLoSrOQTC/k6+
O64WXHEnNR2IISKvWLadC4n4qExjOqynC2rdc2orJcIw0SpWaQQRYFXGP3UIzR3C7pCzRIbACTap
dt29Ra4+JxSHBo34XP6oyBpJyuCEQpzliGlBFwNio/caQpxUvJZbxoEGE+Fitp/ztwPJBgr1fJAE
XsTAuSsh265vC/DTaTPhgD0QUGr3ZYUl+YLinHi+18iGn5hsALDdiazeVjIxOTV0FS9KD5jRkAzc
3ds8LgGGFH+iJSEX9XKZhqzVtOZfyDrvLRV9D7bcU+hxiSjJElIRClOIaTY7TOrKLuBx+aWSnSLw
ES3oa7mlCYhRqLfhWgGzFvx6ke76UO52UiDRjDhXX8XC7xM3cxxaZmDK5U+zyb3liSEkWfX70UYK
rHpw1sEki3fVlSVGFvYvTmITVVcA3yEUpmykNVRRs7Sz0ztIGpnuiCJyTCfwturCrjZS61BUlD2s
GnqUZ42E+SMHWMZ9IXeWx22d4IPiZ3OcffEuyiUpLMGIzxRiAHh4L5XRkjnTCq2TlM5SU9wewEWC
2y97pJ7qMijc/fJhwlFmJ37JgPxKa/V7e9r40jCezajpPdIxg9+tSp6jBXWkBIedOJfykdLDS16i
mgZckQvrhn1J9EqWHbPBZA/JgbepqiMwf2A8KW58hXJr6p/bTTqRB1vu9Nb55YLmOaC3R8/Yf5U/
ZiP7M+EQVHI3GnOnGj/tH49kF7v4qWBrHsjGCXLoRnxQj65q24FfeJJS9uNoLC6mQ+1Mox+9kSn1
Nla3c3tCMl6xGb93uzrhCSSHjpL9NpNIgomv84cJqvMmarQlEDZFyz3+pGWFq7JoicxRa1OgfusD
015TBtGm8T/fpWtf36whwr49zigr4lW1/rNqADDfhVI68tkfQaxkNukDWIl5QAgvaxLQJTvXYlDg
+nVmAsgtOwdXHWAQhdsl+utlGEkxbWmCosJjBhl6wHvbILDaRvS6PNB5PCRwqO2eFrpmb/b3LixZ
voLOybzWNrZwyJacMd2YF1tJaP/YPki00EW5SOEdK7FO5rUE2lDV0yZZfTR8dTvQEv06y8NesuOa
RR6plN5x4+TINQp7VraEaYpARqXUa7pqmriG+nOR+WDSm7NnolRHK9QX7O5feQyUiouT+2VeqPcH
e/3GR/JxId8zDqehfoKnvG3xuDTxOiPtxDymM0X9+h7y1ydxkrv1quMc+f9hVn6CvT31wfDeAAE3
y8WCLvh8G0KiWS+YNSNVjuR8+59AI8uukSRbkfC9za6T0CviFqtSwcbC6iRNGaQhpeDWw2q1kGpc
tFpjadEpmmQttWni+9KRCQJ+BaxO2+HDHOGLyPPOvm6TrQx+2wLwqk+y2nWcZce4AMz5xz4Ak1fm
0EsrFDCtFvtq9AwxV3ihUstyYIqDd7l0C4LZMsYcozogOuXojznLPlhLs11usLF6Rqxi7FLZuR2T
zBIk9Yj1MFEO6RbbOfrSArpFDM6WIOco6NItLuIafp29m86Tr88apMl12laZzr3AKp5ALd69xq95
4Tjd9iRkqt4I+Wi6pRsWTd9gv2F+v22taOr2tCwYtthQeja397QfyZhTEtD4cA8SX+6ZsxOK/9Tf
6c0yLeuPcgj85g0tvEd+0ABLCGtxp2kHzemxtbidU29Wjv/iHcSNaNduo7kVSFZh3ClhHZYttvnG
dBo3BuEFYBKIIPM3WfBQUxLMRmovZ/0u2P8mJH1nrJv1bbPW49OwqtSw7grpq3AtqL4/yrYGSirx
1lEs/mfy9gPDSOOQCtTzF8Y48yB49xmVHBp1qtlOCFGYrS4tYR3pmZSbAUEQVn62adkR77EDQ4cS
hQqW2u8wlO36U8zRnF1LtcNJnB7hoZwYm4QNAOkNAj48RLMtvHyhHqscla2RffljqZao/4dmMWl0
5PFI0c8AtJYPCnbg5QqH3x++7soDBIwRSKZaiamxam6GuysbcNFPgPmEGjQ6HjKKQp41g/pJw1zj
Sg9D0D9IJUgkZc4OMEw66dLcZn+bY9rm3RglfMD5UL7xMCzGld+hAtgoqc36uSHr0l2H8EePMtlO
N+nJ0oTmS9GjTkq/TnB+agjM09kelpDccoDEpGU4ANofq41mkMZM2ia0h/I/PfM+F2ms1j2bGu2K
3dxidWtrpUc2f0SewGENMSyhw8h5SzuO+FIr41xxumZSOheqHsHkOk6uQq41S4b34v5UtrAC0Qxs
+M5RoCSzlewohUGLs+yK1z/bsZYU6HuXQr45VAuBIPE++fZwZpIx50+rJDhxsxgAhj3+BCNs6zxv
0qfGM1r7OMfrYTVxpGuY/SP8IZikBI4PBnYVOruYL0HzLF51AptRbBmvJ8k4RGA4F/wyfWgSIZzO
xfdZxXufkXCW99e/N2e1jpYpOaiNYPuhVLHUHYTA5bHC3VZrN9WbJLK9VRWV1JOkyBNCCRVTvEkg
VfMsEgOZnz+7BsH7yNXaaGFC5RERc+Ply5P4fe8sJeWoa+HgiNxkzdt49UEGCIaBp1BdEbWCD0FB
BIxHZu/o32GkqgIajGPhzxJpeUIj5UTrKBsCxGq0QY2IzD4IvtgIsYevZRk+Rf74O7BL3Xxb9VlH
L2CS+4zKOA07IM1LxWm6z94pY3K4m4ATefVmYRyzKf6fJGbiytWg8BVz+Dl/lJRPMxMV9Pz4fofy
CITnU6/r8tTqv4WHrDdQID/5zTPXb4jQHy+P3ynautmHNMNOrY87HUxXEySafPgv/aFjALTSs1r2
cTQ5FLQR1cyY03FDvQkoVJC2av+7nWGelvMwoSpKx1tlxKoT6fw+J8vqbNZoHogJMxSAapvjAREi
a7fk9eHZ23ksxXXMiAAzBUMwN0gkqR9+rFRdEuwy59HI3EACD7kYb8vg2RWocvgMK6NeGbXn6R5o
Iy4y9f5a7afJ2KAPqXczco41bGLinYhkD27oBtVTxzFoWHoqPxDYvJILQpRISveqgrCvjSBP03jy
+M7sFjdcraIynfuMy3P6jLd4kABm2OOBMREi6iP2b7eIVxJ7wSdbtn0KFQfEzpKRqxOyErCeX7p7
5u60oKBnipaPt5UZC+NMnDKZHWwWpVA0qY+MxxHdKcq5Llt3jfOGCPWViG2eYrGa2N4YmjoVgBT6
rQXGpixeqeoJ90XEg33PeUJ2GRUYi51GqoKTftLd/PS5jxZwqP8viaLVpcrexXhCZ9xiuak50t6C
LWsUEjORfZEVBeiNNteSW4y+HuOc+OANpiH0tmc3WNb434/iuJ3/zZSwm03Qy01xndo3dk3nie/E
Zx0f8+K0d1HqLlqIRia8N1HOgv7ql6QJNjU3A8BNY1txQDXPfjw2wbNxWTk1o7m71KW+MUbYO3oL
+5NZnmH2rFhwNW7faKQq6NOP1PKAU8vvbYZbbc96Bhr57P95rSZuB01Wb6WsCoe6tyKtHHqRe65h
DVzSeLsv4NTQl7c/zhg5fyMKZpQh50f7cYar+FhZAJ3xKPKDJKyfFNR+9WJ/3lqK1R+qXAPxsVz9
hrkVeLFdQC8z2HApCV2R+Dz0CDFJAxBTeOWKOfviLxBzdZmRCnEjhs1tTPOsMDeaZ9zQ30SfrZEx
7X4RBH+hlKw+rcO68d7bOUUFX89hDOsyzywKal/fVz45vXqUOG1HPg77Cp/CxiWP6Lc+0dscxEZM
tGBhUbGiFks52xSiHxogVseXX7ttU9cELop/krPLjdq0ODiuhsrnEeFdCAmtTl+jhfvarurwX2XG
IagzuuJ3XVXIKlI0AFcAYiJSuGGOKjLLFhZDVRKEDPffEttdxyGRAdwkp0DqvDEV6qPL7fWjIwzV
CmSEyu14bYoM9WxWXebscqPi5nDInbrAaGmwDY2bzYK5B4aTqLxFRl9NeDP9HmGv2SZxHkgox0Hy
lMx0zrHml5BQV1MhdkE9TgkhYa7RxdoZzuioEQ0Fk7kpsrSiPTJqci66rEriodbQe/YI7utG4iCu
2XEVZHsA4ncOVpGJcHw8oJ1WxTvtQaZgpyont+XbUtKi8hE5Y1c1KEsFyQKIJ08f+scdYitEwei+
NgTKAoUNbIjVAlazOrnGgp/h96GqVqBn+a2UWrkVDZcDsEjI5zrNyorRVY3s8bin5YrTzamuXkNA
4z3U6cFKYxh4C65Ouw+RW0B+GNgALIURrOYbVfhsE3pQybznJPetMWKOY38Qm3ecp8AGP7D1n9Fn
QFzUo7yYVkiurK929RY3zqRzsH/vICsBMUT08nlc0dywvUPgD1qMcnEDh3EPSK+OZVVLu31zHGTz
2eCDFDYRdl86ZpQMkU/NGFg1fk8S5oZfNE7Iv23HR8ORFXlvvNsCmOTQczD1Tb4OZcyof9yD1gDI
RHnnZYmVEyj9Drf0WDl269+4Ws9Tk4hKgCQEQ52PTBOpVxQRPHGNxIllVc7shortWzQqU2jn6W+X
dtHNOgj/q87yCkK00d+recTe6zXUHrhwcsM7NkHSw9ONj26sdiAqHG7rBq5xQ1if2rsXhVw7Y7ks
Z+ddYdjG0k0BhCpvsMllQiFKHSsHAmpO6vNf30uMAZYif1P+3cif6mK+WxfZLM9QbaznbB5hxx1e
CVL1spcKs5KDBgWi2D4kCpkzJLL6uXUNfuEx5qGjmSofx9bCY7AneoEjnlVQRUO71/zZ42Rt8mAf
8uv+xHmkn+I0/vim/sqJFfdErBzn7E/ekoWEwWR7Akw0jy7M5r9rjhinB5CNgZiWNu4zo11cWwOg
pk9CeKg95PT/5xNVI8NEBVbwIh8AiuxWmNi0wyooh/ao3mwDecPckrVFQowJxeJBei5SNW2Qnp0v
kDwxjh5KHkN5HM0/lgj7CleLRR9ZsmRWGuKziN2IAx/siyN6Su2tGF3OtAzen4IXApK3kNojFfTh
1pMX/ghciwlPWbKzNO8/yiiVQbxd5AqBzC8Ce/Un1JVWYHnCqwLoqoJxU1daUzGJ7pxC5OnWrsJf
mb5cPUPGUUm9SNdB4nV9SqJZTKU+gks46Yct+i5wfNo9CcLevNUNCg2+CQCwvdgLhpbsH1yP+SVO
FOeSEGHRSeyXI30xw0Q2DoXt0/u7aWQvqS/EV+CgVX7RMpW0JNJOWnIvhSuTRJ3TQmgal7Kk/vW3
BzgDEgOII23W9y/iplj9yF7erP6oJ38LSOnkCwcDYxcl0yAiHbxWg1bObZ3lMB/wcd+iXzObYFw2
eXj1cg+DKFWEW8EIEjHMZUps4hJ1EPXuJgLYYVVpRh4Sr6AtJnpsie95qzD9IWW3rQQ9cfSlpSJS
YdXsjqTPpjQla47IBmXGHqNOIrQjNAa6YGbiFjOfmj878EiExNcFB3PK4CLfuxOOEsZLoliRFk3h
cmlGFvLLw/R+25H5I1At7l4dW9uhfL5xw1UKGY0ZCgrUSSVuaCT0xzpv0tQqbjlSwaVyl0S3zT0b
M9BiHOYJjo4TyIffKqPm4a92YBImmO80LX05CGwOAU2+W+umqv5IBQaR1WTTL7QZweE9iLM7yR3a
nUxKROYl+ZYuULWnpPk1CPEQHMA90p7mPKPAc+w0CWKUvvMtUOv0f4ggbEa5QOcpRcQ3kgqvQNj6
V6HLw4pOM3vYeIA+WIIKQAHtii6OQjjbnj8/4+JMhCgOCoM0k1LHVHQeVTSxc4dDc56N5Wcgbu4Y
Sajehz7i1iorbQe7okHcRQIwPstlqOfofVJ2umUoB11HoZa+pXW0Taypymcl5EavPdMm5rSL6Wob
wdskMXqmVKiCoeTyTOzsJYQvASxBuMbrkAj5ELfdVVNz6Wuh4oUkYEvvghWUnP9IAWowHrhuVXmP
G9yPMTLQ7jB5dJHvlbf+zSETZouRhUo54u5OJUN2eHV4Uwcgf5/dOSOaBmLiSSO85LWK0yyGEalX
P3QiuUtTfMMqtXhBzsb2pakA0CMI25Na3gQzhfTZ58FDW2Y4Nem32SNfpOXFpdpN+zXz8fmYSqR/
j55n25nGh+LFoV/Bjr00m89Xqw7cOgzHNnvC8D4fq3HxKBsJRrAZaMW1J3Hv95x8aaBb5RghQ1gh
rX6OLS+0USI785c92lWbxnL2EhgnPg/kQzqAAtQahAFck2Wu7TU/JuJV34MyTMrhtFGDqkp50kL8
z/OFG9zHQm3wDg4ONctpWbyrvTCevCswS2XQj49Nf+fHh13St0CPPBlTZj6rXutFfmkoix18RE/W
2f9i6wXE+TaUdHzh/jZD7Tl6qEo8NfzwM3u+KnWL5WQmgHVDsBzHIvFqt49KkgQiKmP47kVnZj9E
UpbkbyHs5GjRou3fCpqoVFyY6q1WsDKt1DauACufPzenQgxRBOf8WOPUmZfhg/xhyPZJBGpnRpv1
XR2bpNUiO2yXuvjZBtBVkH7Lj0i+Z1KKa0atjA2Gm0NV4DblHsPJBVUaXVhI6FpOgSBN9w0ieMZa
pBxRuNW+22abXEq7nUEoBf5FXKC/agtY+pSS6FAAqU8ZZQdPKqv/qxD3+15eWLK4WeAPHFGdMOf1
51VkCgSQHVLJ1iTutfV7hGJuU58z47KrK79j2vnMsGcTPgTnJNk84w8a0nViBvzQ2SiO95pOoAaX
aQSGmbVFOy3KlEhXEcPBHjV4tHhSnWnLjWU3rCKC+22LW3UMX5CZ4qXZasD24w2vdN+owkMWc52C
z5+uBoMsKS6O8NFSg/N4nYj8qTcE0nuqswm7OaR5F5aDQptavktQZcvn4NzDn+4PxQxt6mN1T83H
VYRD85dqNn76X2alSgYBnKrrtsSDx9yh91bVTbuTt8hnVSkcJBcnpJDCAJztA8xRbPlip/kUbs7e
FSAz0ggcjh/77EVGR9fIi4ASSG2HQ2NM+2EwlWTb3QGkidqxDqoaa4FZpRBDaWN6nLdErCxXrZbU
NHEeAdxYmY9W7z9PmPQToDyqpTD+4kIqQ/GRuv0VgS0DP2F9poUHBjVuMlhwVmD7w1twm7yrR3k2
csMFPZ+LobbcgcwunH7VtDeVQEaYdCciR8ZdfT5nB2d5GRBqHz8cfcgV+4jkHN80iPCzRv8uQBFF
NK8Kd4U6gV6NT6l1nihKdIN2mcFVOyDZd5SUnSK6W0UXKmHrdc2lyy0Et0hRYagXHUkmTNXoVgr7
IeceMPLlZ1/yTyQBE0vO835XGGxxcXQisOkdVMNQ385PfHT40JQ/gjI4dY1X8dGdZ7v04GHgvtET
t67FU+Y/BqP3y5OY1jtN5XLRfHXAPrpxspAIDbXxYZPK+mN4AdzGkpcrStDAQ7kKogPzeNVilQ8n
P1Fiiv5FqwUK2s4lyiInUVMJM2y0v7VPwRxeFiGxQ985CheKMCR4qXqCAEH1hcOLiFMEyCiESB54
qUytbBp6FNyPLTgvnfhB9b7gkSskPO1uBkpSTFdIIuYZuDUDLeqVlcfmddL2tMhm0/7nd5KatQ7h
HfE8ZcQ6w4eNpjxmgzvMXwwPmmj8c0mWzDgPXYy+yIOnxoXS6DZ3++Q0b0PF7ioBY25CPBEWRb7C
bz2+GqCTxLrTTTBwrH7rpBvLV0b3mnkJVqKsn8uILPJvYQhSwTFLeMBZXsYY+wzLcu5/sCoxd7kd
7e9lu3MpHl0TD3nRXq2itUQltJ4pn5IkKpNWzEHtxJhLDUeKmVV90E65wCZJlHPHaif7HPFYKDXN
AUbLP2GjnRXfLMNZDBHwXujp58gacAr7uILZJOUM0nQiVljyeH+FJHR22fBxEhQRmT8APameHcPv
9udspPB3n9kEtF5h7hvgopgT+Ul5vhtgFrYlJU+5M2tOhmrQWJL3y4euwbxUDJwZ5f1rZthxbR2E
V/liHoqUKvFFes6K8ZkJzwkICQ3qJHdV5upJdRsBBMwp1XrL5LSytO486KGp+YHc4Ac/a27fjGRK
qLGhWFNddlZc8whXVFL2nYg89SlSCWbKa1b5Nsdta53zgirN4RrvkYGSAQ6GOx3DVAVZDtxb2nc1
z1v1SbcWs8gkUPrksx1MgKFzkFAU0WCM+9+r7TPT+P+uPwBUbPMfaIKOfzM+BvxV+eOpcnn1PrM4
rQ0Km6caoZFtqklHzek2XloiQfQ4S3O2ZbvGUjPZx4dP3QvgBwtN3yzLKbeFWRCIH3dVzT9WnpNy
i51Y28GwCUq+hYxcxpZPFOQk5XHqqc4fXziekN/CsHz/IaGxGC8keMYbAvh1iLUn0Z7llefR3BKd
sc7md1R+9luDrGu1mgCeikL+xKRSUoASy/9A3H1xIUMCFhR+TV1SftMoL79kB6unLZ8583+hKi2t
lBQuGXs0o3YtMsqXa05mXBt1qvvcRGD20HIoToVBcMsSSFAYpFp6Bb99a7dh+t2Pc6lYTqX8jcKe
DiCdIh9l6kcqmQcD0qL03BHOqNuFuJoBWDNYqqt5F/sC4ptwTXrUpoSrEIoYECq6vdPsd6X+BxLY
vYsyENz2vHwOo/5cXkNOwA4uNMRaxyga2Dks3UD2IioS1o+3LI5J5EROPf/2XHEDWq4VpEBTbiuW
yUDVT/ikJRQ++X24BpAU5zX6k7R13eb5e9k/gprVfIGk5GlTDHzYf/nSpSjcojMuERsmSJjgZcw7
hD1mBn5/1++7wDBpIb4DzYc2BlEYA009bGp5W36RoDX1kBA6zQFgV7bEOLWLgNW8Q5MTtg1oKPXo
lcGQxpMeKs7YYXQnYEFpfBXb5j4HKnIH9BI/ak8da0ai5SpLrEc5iktJjFAze2JF92DsxvfZF2Fy
W0QHPcJMQjU9XS+FbuYdKTmpky4a0D8urLiuPuTI7nceu8J11jxBlRY/AnpEVhWbWBGuRVUo8ZaU
16jIfgXkBCFkK5RS0zbrqr2fD4neUhvt5ho2ogB9QnMkgAO0c6lFL1kQMWYmFeJ1II1TYb9ESNSE
19td9b55SiGIAhgOxJRltenwbqfcSRnzaovELn50gjjrzrdnShs0NfShlPcrg+t+P6/dlhpQ8Emz
KniA8vGgoQvm3Nli/I9lqLHjCxknAAsJ7d9ytr338862uuZNA9XHEnYZl59008UKSVmTOND+Gis3
VUYpXXxbc1X8faJ6HpC3My319x913m54n8OLGJrLDQUkXPtSTJac6AG260cXcA3/FSCJLdaZJz1R
lUUR9SZakuve7kc1y1WrrxDh5Fu5ZjbiFONekTWxNiX6pO9L3Yd/Ah7z+1lPRivTb3zT7JN4sf6L
YXB36bnkoFcEV3pCywm0nAsicGI2nlWio2L8A4GbdD8ME8Uzy/N/yfohHgLJJE6lR0YW0+OmgO1I
JuCayEGXkj0ReO0kPb+AbYhPI01NkFqbwoFZytMseol3mkXFyO1uUAFQ/4ONB3wruWtdtmsojXPR
6Z1n5Ijjbfj+z0WQbV98El2ahsVUFyFV039tZPGHhcvYahCgRHBRhWgPOyuiR/wesiuH8m6Q1Stk
q4P15VMjEeKzCfm9im00fHxAKD7Fhl8Q7iE0XYvKHErOexmVeZrzJP49HIKsZXEGJ1KWD7+807mZ
2VrC2vOkLgqG21zv085aQtSlL4sFSHZqB/Vs6q0TNlYwxiyNnxC0DZf5Jxnle/BgKaAJryTq4Imp
e4goG5KNT6pNgLSk90irxEqwuMY8KfNCyhWfuuW/eWwX7Ml+wX7n4dOY853qTOB2UmqAFRM2x0jF
dAUS2QUz+tmrR+UauVWq7u9G+ZQ7rq9AMsj5aMvRJm8pFqRU6wcmPA5uCOa3I5rkYY93J/14A+Hb
0fBEvXeM8W4eeycdbMEui6v4p//jw2RJWmjrMhQV1H0/H9Zh1GVrXmabpZ5vNTm3iyyqpNeWknJM
RImQx2LIKECZQ5U/Px/0lsiO5US35HjxKlS0OIuwkSvLNqC7KwPwcgJFg9WpwNQ1pbz095F+3hAu
oKv38CgG70Xeo0eKFPIr0AQkXP9jnmTPExjO814JR4TXKpJxwaTpO67sOCX4BJyeEZOteh3/L/fI
MZiNB25taK/zrXftJw5VHvp449kmdNWwQiEDw0jFpsZAP0udRQdNjZ5chXZOMWUjgstBN2sHNfN/
+9Uo7kpgz5xy7MZpOTfLjauf3otHKs+Gg/jlO4Eitrw+GRm6psKE2XNE0Jw/WoisNHRAN4pexxby
XWToBsspGBXkxmPNGnORq+Q2eNendNa3mY+j4m7hqUSzBrez+9+MDrWykxwcJ/cAk/UQptxP/peJ
9F4yw+jLLHAQUHFXYjjnR84/JDN+ym1Z0nHBnMUWcpQJGG9hHWD+BdbU+R7G4k2DrMgEwclUfdMy
t9n5+Az8LsYlltjgRidie7T5TtbIkWdOYALsYFkHBVf+MnhaPDZSBdo6Ezoa8GZuz0eYnSHnTyox
Y+jJKdxkgjDnks5KlL0wrImSXVmsCX+6rcuTQctRu4jQtlq0FD7aWKh9SI+9r+P0ShqazqfGjt5E
9ZD8oATqsABG0QJZoBI5bj+VNJYpcRVgsMuUinxXOU9DnMmOO5HJhlYQBGww5kCHuMLgWcEqQZfU
09wOlHihUP6Pskeiq7KyE7K/vxOX87Y0lV+VA/Ipw5l4lv/ktcXGQxupKpbjNGXj3Ow2Iz1MIPZw
D23PDykLZX/4AeViIHcOuXd13SfZHb2kERgbtPQMrUaRx3OY895ICw6KRJJqQgCK2pePlLyAILsh
AU9gMIk5wIzyDV19QdtdXSUkmtp5UJn8p4nZmc5da/OisYalHrPfk+f7wXxM1ShoyvPYu7avdgAz
zyzsGHU5rmLvBgX3qe7CCQurSY8IqD1KRA4tJvdT/81CpSsmcQLj11Qyw/Tyn4UkwlJmvZ8snp10
BhBatg6WGukFhEAN/a9Azsd/sKuJ4vYosAdGIg4s2WlhFiPbn8o2rjsCCc/44Y30p0bYZvTBGwNQ
YUWlkzdzwU2gCvTbhfG5naZHOYctfjBdf9CklWopGYruMtdbtTa7a6GYuCAt8IHJ6j+Lq8U3n0Rf
b3A5DHyin22fGx3WL+0eCRZ8FJ2kV9w36ekyvPHl4h42XD5LwkNW7KmMdhikxwKnCWEppNqr8utf
4G9CuME0AIkO66MMPOk0paevwvg82SxYgCdLmNRpIL+ehBcZlgtPVIv4/0KuhRHe8X9LNJOLqgH0
qoP5QD+MPbbNKqSrfe5JpjCDoJqHL75Oflc4TkLLkNGz5GKJGK2TciIl6VR3lWv+TdevmDyWk0Kt
GKBCY8HzWdrmWXU1SmQSTv7+r88ucPPWcx3J1ODEsCOUZZJfMrH/g9TQawVd5BQLi1I3MTi8eep7
+cAYcV0NDqSr1V2csnV732DPcs2t3MVtFDM1FNG4oWxjGve8jxD+HuLnQexMD6rg9YuAue158p4T
CB2APVEvc+gBLkcgr6+/DBr1Ca4uEaDPLbA8OG4XgUOiJZlAgC6L9hCg42zlbnIhFJKg8ilqEkwj
4HF9SzH0qSN132EAfuOgmpp0V3aCthsRY9+H3afpOC0gNBYkmvTMBJQi0zeWMNB8ihUTYvB6PKNp
TufYnuegiGScreOkROA+cJxzSjj4FFQ0bGHLRbIzcVpbsXsa5x52SK2z65ArTDzNUtfq2z63w4vu
jWDY4hfnmqWwYlTDjujNJcVEgf3llczeV8IjAQO79WEI3kekaN/AntgAHDO7fZlbpA/IH6oH5VB/
Rf8aCfIRjhYddxtW59h/X1dkt8WkFti5vR6QzXLcDTwnsfkw0+5XIi/0QLIBXkh5ofhRQtUEGoWe
sGVM1VpckxeFICQgj+4O0rgkYoHWikvcOaveCHAEkigRhItDsBMWFsdrIFkBDzw2m67vmAdvhDMv
AyFgUCM10+KMz+PZ7aP+yFTN14TS8QTZgEO8LMeNG6DBNGRZXsa2Na7mdDGfnOOTy6/BshM2kd7D
TRe1Ieu/VSwlsM2HMqvRfd5wNvbOubcW/dCWzMJtINH3/tD5+/wsREjBAfmvm3nLFxASVkWY0tQ9
uVxgdG9IeoRz/ek3EFG4EZtrX+68jenwmVkmu9usvcJKufQzIwKmleo78+sHLv7eb/ufncseDPge
gt46OXsIqI7ukohOOc7PUcWxtI3kJqLCpHt1yZoyIIifQaKtALCoFCTEM5jY3Jvtc00LL95h5AXs
/OMJj+7t1iLKSmGCzFWUqZmbiIX8HjAVQGxJ69IBeKIkyWumhjetgWnG1KnVn40olcmSHvpFQ5Qx
RS4P4T4yrQMFuuo7g8Rt1jilTgpQKBksPQwKQY3UPMU5+wxcdO0+Ja/6Dlu4dXpnoe9sc8mMIsIy
mtAyBBZeYrF659IPKyT7Yfp9QOpNeFHR9VPaPj/CxTJpiowY2tSYCCaTHymES/6+0V0lWR9Y+bRj
OItx3dP3YpZE1zagjLhLX40O8kXJPhIsrWLBQJgfOTom8qptwOz3UGgU9jlTShD29kSB1aeTCxmN
G8+67NU4LEg8NqK2shOn/YO2my7PoAS6dahrjGa4v3tki2DGcAlCf80dkjF7vopPAMx37QzfMB7J
cxTej+WvF4Z1GxnHDDkDDgeCFQPFbkCezrhnx+yq9DAWyRkGBPRDsKL0PuY8ufgZQfJ1zh1PTfRp
WokdzsQ/Z+uTpTYDCYsj5SRRz47z+y1zfPZ6OrzbBQLU7FwZ+oplJtDtfAlddOsPNk8Vp9subn1p
x4JZruLjTAOr0DnKvtkdlByX4bZWLCRWmUL2JcnsBLLz6ffYpOokm+Q7HHYlO54+bvJblcCkIaoQ
Ya+O6Zv7M7OttZ1CiVzyUyaLrJwVQXLfCc54myL54q8Tzq+lsquLK2UzcupK9Tp/3WpwtNQlo6Ks
+9JUclTKAXiWJVNNM0C5U9K4V6s2FBgjJf7po9BMhq/C9FOepBmS/MKtzfO17O0PMad44db8vIe8
KCD3YBEZmBOxlHRAZgLIiDLzoKyWO2vmyo4+mOWNYZHhRkkioLlBuy+GZeKyKHXW3qOz4ywsy0Bg
tn41zF2RcLCTaJYV5sBvCT63c+LT/+o2GndmqyakgYo5+LxsA9wmoI0hZB1Uq/VquQGo+qoATvlY
zHP05lH3nOwKZcsqd8eC+asaAFO23hNZupNlokwQhB7LdRnA5NlcNkvQHMoKNL/01isRXwdQO3s3
0dOo85wqtQ7XD9HsLM065swjhFlcH0bBKdASbtH7ZiL5O6H6ktTAS8Rqtn2ZU3QYoJGVHMq4fP4N
f0Glu7JOlWjJCZrfyFsGfIOVaQmyNp7TjOXHgPCOheXhr/BASSIAXAAnrMhDSp8FF1NWUJTqIITf
uZDcoLPBTw/mX6XPjdeew4aTY6nalLfITCk+wRa0jIe/IdxNNDE/y8p+LYWi5H5+0XAnQ/+wHes/
O7juzH8iXl2qrMtFZ2I+QLkncrLmn9HfiZcDcHXeiOZn+ZyRUavWRSwvcxK8WQM1IEhxnCwarKRz
YL37S0XGCNt/a0uyAAUynb/dCptY6vmfSL1q649uMXcGD00Pg/mhLOpirg10OnyD2MX1+W3NQG5k
97g8054bOM7alZLMHJmIAx5By8ArdQ6CzTdedWWmm1EPipUyaDlIYT1tbzC5SAv/XqC9szwJjizl
f5VgGum0htt+z4/aWOYsM5bE8e5RdT6GlvD5GWDWJn55eGNtt5cGDQY3xz1yDr4ZdndWAjuVsYKO
/F9j2xwvhDnd6IHYkNIKFzSOLYRi5sa80JZGy43Nbbb1/zKdGXsvPB4/KbXjQh7MeMKCQdQ5bHCC
YYGq7sA9pKqCmZSFzR0DbtIJj6UJN2gdufVQdlmdmUdj19LSlQlI9JjVTwThd3Z8ooVHlazVgYQx
C7nXqHIRCawmmJgnNSDb1QFqZVbRqPWQwuDL5CUMNjX3RW5rT0Qgwuk9NYsGXh8SL3Vo5msaDz94
K8Ow/qbN0Wo24ZRpX8TCM7sTWb5/uVcWLjetW4v/jLMQRVSMRAhwMuKNsJK0aJXOESmplME8AMGr
BZ57NkKqwpTypMI5hOX8bY2TvQMuggPuS4d/uX7iJvGh640evDB/LMRJF0w3JPayLm6iP51pEtIa
IIBcQTPeWxG8xxZUHVFOnImow5qH3T6o/QaoRpuvWI/KK5dZEeC0XZTX/Su8S/UMgxRNM0owFFDm
SEKvWZ5pzbx1U3ZJKbeHBOVWkXxItiwu8yJQZk7g/VBF6RSlJvTA2BBIo6ILKd8qhCWyZ2gDO4ZJ
t4vKcIg6zgfYiZGAbqlxEbt6ebd81tpYyJ7xk7oDtG+MmW6j7FjlbXU9bw4lB7oPkOHCB0+aixRc
+R/nkunNieadej1OCpuf0qeB+I17OyzZQ/e2PqMmdvDEv78pO+QpT2DOTbdf4xPTSOkSr4G9LLz5
FDMaP4qeCq7r4SyJPuI0cfDMdFw4WOpYTSuBtCakkFOR9ZAZL6ZJhVTdUivvMcXH5FmpwX16X6eS
u7mkgZ/mVFW1sTJBg11F83iX59ytEDypWOGcemRNmm5PtulJO3c0rvkmMi/xTgR72zZb0AddDo5G
xj2w6Xnf5WwzjurQ80Co2kfMfY68cPFgI/OAHHakbgzYABo1wcmP22gNlRFheYQGFFhbIhmjZbt4
NWMN/A6tZNfnMlBdwFja3OzlCDhoobWhvDQgHcg/uZTSe5gF+v4cByoZvFsL8Jr2DWMYYTFJw+pa
dKC/SEokueDMw2wirfiJsGw/Duguvdbeedpgjmw8MBI+d9i2vYI4tTJP6L5IGKbGLn0oE4bXrC2s
53PYO+TzSm/ndSPkUxpXJe5RN3ijnX2znWNmoDGYOS8DVVerh5qoJkg6aLKdm4BVLl7znVwqhuPR
j+aFN7sSHBQ4cw7pGBJcdMT10q6w+JBrudtOK3UtaK4XVl8SSCRT9cekDyew6byIy79OjRjzgHsp
vrRbYbkclPsdNIsnRgxz2GLLGkLJBHnw29vFJvy+PQzfXIOA/IJJUY/Ql3fNF82u5lQzucLlRNnH
/9+T/CZVfYS7+1rD9UB2ORXpqekBTmOlmtwh2jnAvlkKMkrYNcWNto3JHyyRHIcfXqbTzRjGFkXC
hGdMXukfzJP2fQaFpgbIRzCyxkfxbEn2lWlFEIdcu0Q9LIghb1ecYSmtaB+CMz35b1O7Rd7r02i0
4vFUKAUbGyCnTuLC3v7+zTGq6GvEN+f6Guw08HAlploCmIxJAHVOihomb75JNaRd1Dcs7XsCOtXh
b6Z0xFdfqS4sukV7rH0PcqVjOhW0JG0nOUtNBqOmjqJZhHlEkgQILQ99dqCuGxYBJiHC8HByFB7C
30t2K+FKgSdpU9GmabE1GxkwEN1bchsX4fpy0HHQmgEOP52jUDZfLIPWCNpdvavlKeKqijVsd8GG
nTdJVf1cIvYVgl7u6NTzmm9Q0Uqskm0G80+W/HFzyX3tgKpoOAyhZCLflwbzSWyX8eZdT3ZiTpi9
PSGHmL+JkxK45loX2K6MpLypqxUN6SPC0FPEWyVAGwAIsQiR6R0P90TwfmrNQdICf1oJ4q0s7lP3
vWxobuXqvqBeOf1cWptJjL8BQZnU1AzUMraiKwalsZsmBLcnKN0lGgY8oDy0xBS5fDy9xOWC5IBS
XUMYjop7MNG1MOrTPaBWtpO50IaI23wg/uTSJBs42XHTvXAQFNNwBPHCqHSDSxo1E4xOyUZ5DoDY
nmuCUftIst79BG9G9nPzWa+nJrAV9ocScK9EYALJUaDDA/JfkBOeTT8iQmGpvgPiLtweyZGRwGlI
st7m7DcwC61Q1oGJvwEnyFzbjnB1GpLpekH7mP77aSTvwOz7S56/lBCHhje+AHbkfnVO2Swp1iSf
RnHLtsUT8jLF4HpfhzoiVt+gBCh6O/FCr+fVrg1hbwITBl1N5/BFDMyrXOc3sf1Xa0FqqT0vTxCz
tGzzC2/r0Y+0ESBAuBK52KEtoxxgqymmktBinMDw0puTKya+E7zhc9m8ykoIHwZFu2wotE8eEOzs
SJcSFymfaA4Tw2GWJTC9CBIN0VDpmp91wBvTV3EDl+HJvXcWxbMB+zTW8K+S+carru+4LqGoPiWX
QWDJDTZEOoEpShvRDiqIUliiE27lppfjg2nuNdo+yFXlVotVPxhAwF+oheEAzkqrdQ9lDFtGgw4i
2hxCLQX8qAdizMWOCOhIa6EBmo+hWEcraBS5htV+76rr7SKOvzE+KmP+8AaQ166KwW1q+WbUJ7eK
fpEFSF7EBBLRoO8A+e4BqabQye8/gAQEhAN52HfgZSo408XJWVqy9XqFO58FKU+9b9ovgt9n7ozm
3B/hJDm7I+peSoXZfIJ0TXgqpDU5LiSgOdswgJJuffL+/9Ls973oKw94RT4srDuzo5Tn23lZtwVX
pfr1bqxgMDclrNlS0PMmaiok1hUp4LkVO9P6Bm0Nv3ZBSVoOQlqaD+LBczRJNP5yfR/Vl7XexB5z
dv1aHfEOa76/YT4ktC/idEWQBRyWkrKHbjbDd89qoQHJEySJ5yrOeXZ20IU6tsLciZorch8D+qNp
TvXHt/oX7RhOxCffVR+GnSxyVT730HrFM77Ky1Nax+ObWBhBM5qn0AU/EzqQRcQDSg8QTerzgnh9
uUKgVCMKKFlOMJyomT7/VraeIRUpiBCayHvnqqsQx6mc9H3qWARFAaQ/JE7WlNTSJsKqQ7Si0R8K
/Ta6+zjwguJQbYMp0lwR76ZD6ug+/Rrk9x5RyGNiz/UH0GDijLbU+Cm34r5lRgdju6wrEGOlxBhS
RKjVh7kMdB0QJnVtFRz7FjmVK8TmmJ3/ocDxHRrrrONfZ6bqyIZdelaE4zjC5b9kcSz7mQbrJkNp
4DgB7lZLd4+GZY6pdUHBDsTEdeGVBneATb+Tf3QE/NeAygIh8KCls8bcXTyl8G55w7Vd23itlHtl
aWSQXu784araXQgwRb6AlYjLMC59sCNa57TIDirXXkkHVI/SIeMX6e9E6Tb4YhlDdjHffkTCq8eh
c3tuY2SibCs/SpEdqKSqfuQOBV4PyyR8sbrFx+tJb85WQYBeEWIryGDkYLQw6+46LeFnD43C/06y
aeMS3VvHxVGj8S7N/uMYslligHrngXFJhk3/flY+0KLyfLisli+tOD8nUS4eZG+qu90w4aFLNRXG
bHlRj0bnt54LbyxC3F6/1hcH+4G4IMoMWawpcDiJAqhUyHpGQ+V7+9FA++q1jmrfCLOSH+sXuMDM
6aGSnuqnbYymiQsaQzzb0IknlVjCmwrD0wkF2T1B/W0MZtfBrmt47vT9DwRruE6JgHSFUnVve2/G
tdo8SwSASNcyhGgY8Ti8ZkWywJCTYrXouMsr3/T81KHr60jq3+xgvEpKSVefhCVIxbJaifAuT05V
RYdB1M1AZXfe9AMYzJPNNd218Bgcfmux3BY8GvHFuEe+dhs9smCGJfjXCKpX+ktPHHZPKneXbWcz
I+dKuEYUqnG40YuIUXxkzkCCQ87cgVn521VD2r0JrAJU7+1M1IWx0a/5GVZkX4hld7klSZ6E/FXv
EH9XQUm0+SLN6vnvbI1aNu6jUEz9JjRz9e4Zzy//ysNzYJ1E6UboVCuU29Hq3KTupekGaNxF1/If
++n5fIWt8k3jH2iKpaSleRFaM/aHIDpXoTo3edyQ+t00K3mppkX6zbfPRHVCFNofSHvL84yTTMPV
MTNWODbM/V/1n2WRIbFf1NbWYkxQIHFA7xkgIN3+IC1mX+zpK+mT2QKItcp4sL2lWXfdGfB8b3HX
MjAuKRB6HVvUOamcs8LE2xnUmslyzUKrzXekr9ZpL7k5A/Tvqb2oODKeFpM6/xw99kxG2spVgj+q
EzFuGQQwGgqlwG4m8uvdFLuz9n2SgWmRhOgWhk9Hy/ZnLKCnts1sJxZQoLV1GqY8L8h4i6NjHXOW
Maxa+qcnnd5MJ+S3I9yGRJdMXMi4uMay60smBa622uiCThzXyqD+/0x3vd3+qbB/ff2EBnq6tC2N
lavCvpfki5bZgzD7O5MM1ji9FUBOoCYXvtLv0OxpxtIj8BXmuEaPJXuEWln9fv3eOWKALRg8TlQ6
/PDSCnMsodkt9FY7I4LE/bdrEfZQPNuPZcAwBqxCACVXDS6Etj5NIf3eoSZ2KAKIujkZHfOfxISQ
/ylOLnc408ncj3V6anFLkWBLiioAS4o/suDiOo6ubO+5Q36uFl9H5aXnoWDqzZ5b0KHJjtj/Watr
x2zZmCzefVSWXnR7Yy3MgvnjwBSJUSfSwD7tYB+0haFA9yLtVCtrP3rwvZ125pvP6Q6IF78Rh+aj
wK1zFJ0i4csSH2bQwNqMbcRTWrkOByqF/3uJNJXElH9YNjuQsiTSxeV+ra4wdY0Re/v1voFMPcjv
XB7BHaHioL2BaMgeOIRgviWFvWLTb/omuzG0ssg+vO5Ekp/zUIt4Km4Sj14RZV9PPiJjcg6b5G/v
FWx46m2RvkjI6gu8eK9eCVb24D6Wol80GXhO//NAkdJURQEaxkhIIcRAT7C/FBaItw3jyfigzSGX
AlyseV6HXOIaNq9eZVwyaKAT/eEyQWYDtR+RmOuyJw8Is7msTgP96HQ4TPZm6TFFDsocS/F/iXsg
gAcrODv8fs0Ipdn7/+6jJJI+xwG7X2Gl1AR41gMANQgAF8czUybL9As0AQj+c9AYjJ6HOwXglVXD
84oyaXOm363exiFRG1oEtHB4DMkjHBc2brwqqGQGvhnmKz6BnDZeYTU1aVuIPX8yc2lv1duP5Uq4
KnQgf6WILU2SvU+M4cDxvJ81XtFIMr53hnw9aag4y49jn8d4xJ+BRJIPk5M3mjX6dwteIed0w+Z3
C6X8Ed17XUUAXPApIeCNZQVMCl5Szqbw7acASQ+hB4CC4NFfrKEgQqzVLn+dP0fqlvZVYbaccSmM
a37ODldIkjvLvAKWvbo7pB9uorz3G+x6ZskSs+hnQn/LDjz54g68/FfiXI1uMNdRnlTdhmUC8Wzr
ZzdgM5pHm7YzLd3AQFoUB25AhK/+D3gE9qD5ImyhbjgQYGs+/mc6kUbXnar0A6SbYk2DONTCHP8/
uzN+I/osObzFK7gCwkGrQNd+xyvWZIkKftQEZV2yoYfh7N9f2kQRf8sZq/f486jzBCaO5SI6RQNn
857tnN3ZzNYDVYz3g7I1Ha+456k05MsChc+bfJfUDcnq3q0RAb/T7ua1nwZba5MhQtjuZ/p9MeQO
YNDzR7E8x/GoOLFybPLwBzomgujAlKdKirrk62Rs6rKhenO87+dyUketY5AGnS9suEfuPPFq8UTo
zkdU1kj4JdCqbPHknpSVK7HaMHYyf5OjtIcbDw0lvRTf2LvKUigRxEISj++wNIeAvW4FKrHzdA+U
5Oo10CdGm2smzLZHQ2CBFZyPos6X4KL6CCUdt8+bfznY5o5Hn5IFiN4gdQlCwuYv/lWyQETI4QnA
eJWpZAhSZf3yjMkCsNKy5IylRaZOmnkEl3wQ0dhrZ38mqyK5C75pUxPVKQaWz6GS4xUCx7OUPJlW
Y+HwOzujXb5zsxWXPOZHOsxxDB7bp72IIuO7Efx1O+yQtiRtw0MhRbVOIm+wo+MMp/28TjtDzTqr
E0rNGz3RTnE14DqMhMfo3bYvYK/BLEvZzSEwwn4xPu3MFGYrGmYEXmNCYkHb2BXXP+A1UseVuLQ+
f6Bdw8d4AmgiIsWxHEcWKr4jhUmCkOyzCCxKRn4dCzsKWrxrFywaVxuKTBpGyFmpoOVq5htG1IkV
3lEt8k/eKVp6pspykDgkeGDiMoxiaRQuI0rHGDHosXF5Avt8nVyT8PKkMnDjgqv07NX2hT0xhcB7
hl11x3llnqdQEl5QfZhNsAdJhIyxU9yz+7uO0ID1YpsIoPuAn8sBKf8W2UkpzqVjDoX23ldd60Uo
VQkcxzgfiQhqOVbUsnHvQt432ca+hA0nF/9lp5aWAZlY4qPlwEloNhMs8BlXU7Z+QdmERTtX24eR
Aa4LqYsRGPciVBXEmwP8G29biJi+0ZHKVTf5LnQL61jieEO+ynJJDGSCcR7Ski6UGexDGvKrCPEx
QkwqeJ3zBTreAAqIIsTD3UFT6zUSOq1gLTCZIO1hlhuqZk+nEcNfx8gpJWTGSHMuhLl2s0l32dou
2b+TD4ZR1SJraG21jbCSowFdIa1/J4H4bLWdq+284rLYskpalGsSyFfwNEEieOYtkG2HZdCtDmMy
8oakxP0D/AjiDqemlXwoWo8+EPzulmRNF/Itki3Ks5GWl0hDD8ljEsnbYblu5DQ5jIkwnX7bNf79
rBIah/b21L35o+iYY+G06vLP/1Njbpn9lMvvVzL2R9J2YqfDkmxBADMBpmfE9MiduFNYay8+uO+3
LCgrarQPmsOWH7N5RgziDh3rIDoa007SwCaCqa2oHGnh2WfL57wLofwdzMlvHzfDSXXm3F1b0YxZ
mG0s854uX4UFocJpecq/E62HbYxAUGbb5V81EgXM18NER5em1eeilCxYAHN4nOLGwHwo3wOfrePm
BRXOkiEpNGu7uhJ/P8IEyMjsdoVxPaDt0Kp/gkPiUVXQAkTHqCuWqe4X857kWsFV4dxIGC4IYapj
QgmXrq6NLwZLbNoo88POnMUhoCTaZfaxco3k7+sPu5tzuVszxuNtb1qwkppz5d75stMM0g9A90Jh
UGJ07KcYKWwfLlwRYOmTlrtYbL9jItGLmU6sgit/eBh4s4ceVlK6fPtS3cMVGdZe3T90K8WZTysH
CgUungpK9/9RlCnTzxoUC97nXR0QOEEtdl4+KoAg1dSHl3qxw73oN7uFnmAbCYd/1LuW7HYYYA2U
pyP8IbbghkucjEuDMLoITVNOMeE4nqHtWpLEhZ5JS/rB+lQy/919t55R/wXmE2arT/UXhq2oPZHC
K8rw+msMlpTwlVf8nRf+hTSl0GASc3Fi6qOf4OGG4ipHC5nkXnM/1/07MsaNS3Yg3j8Vlj618rLi
+It7HQT7CwkQGNNcCLO/TGvUutTtXwGEyufbNBX/QNC4a1vJgjPupTMUhFNd+BV++kJdu2Rq01Ug
3drkVrPNhdZEmVRnnE6RiBUVwor1Y69rb3elHz+wSVD/w6rP9oDpCxLpCQO1OMyreiFCQRJZY9MY
FgTnTlyf8EJ6VkTCOEw6lqQSKKUSEDQaVC1qQgNM9hgZXBK1adF8uLyZ+v+8LG9QCVsR3Qs4med0
gYSK/4oXaK3/ZQFYXxtz7sJ3Y+AwgdxscaQiXsq+zNovFvLVhXlCtpqseIKJPCPjyGP10rp57dD7
nMHL1wA+P4C4q1sz4wNjTXV+Uq9B2CdzFeWw82D5flL4R1YTTIo8gNwEJ326qJR29AyF3BSfpwB8
lOMd7apu3z+pt/1KdVp8xWuCE0/FMF4NqbPLQ1IvJUaQwidIv29F4fqPVORIu78pxiXQjcRtaXt7
BL51U0WUS9WAiNSXTpkRoA1NzDCs/3ZbSXTFjKTy2tdAbtif89jt4ikqea4Mt7jUPCH62MqMimBs
0BRFSxSGgRN79XyuADz2CfV1sxdCisSE5E4OYb8HgI34FyOsjH/vUrmuykQ+av/mCHqr2S6CidBj
/mrBM6MYM8Hk3Gw1aDoqzgwsdJ4NA42jBL1InB6qpvGZrxsQi8uCnFFR3f6XVdfz+0GkB+b6SNtH
lSNnwqXRf6ygEUbEwK+1JzMvcaIWq+wCuQobcmAnLBqwgefzRaaiS/HzJKR7ATjwL4sEgJEsG0Bh
baWaI03316ZsJl/4/7p7fJ/M+PWrVOdQ92AlHSkl6Cic15pIFldLMba5KJj7uodBOfotiL3EplBk
e6a6YaO1UQDm+Fhu4nr94IT3N/MvQrZwp9kpn0PdTLpoqjY5lORpIBcP7TYKmNZqjTicVF751ii9
VrzMU3PUBi4/rRUh8ekLHgmydf7w65B5cIgMEl2SkOynVai+v4cAvfsolDGsPwyrH7s4msd2Qggb
WPoN1DEQ6u0pzlp1j9sJg0eBfGqiZd/rHwTJg/JXCf8z25A77iL5RHw1t6NIpWbvYFBG3s8CKigb
SW+rO+EhiB6RmAPRX9tuXfViCSZyqDGonB247oAL1m2vlrLWYFC1kCJDklnkmO+eKs8tctxuwHhz
BZfRUlWNwy4bBOC7SwXUSS8C2w9c64fTGuSA/2JilrB7CXGrSAWUKGH1VipYnak66u5mgGwdKpek
H19zGwsGAr4ox+CWs7HAo2QMlflfAOudBR6xF6IX1Vxm3nhvu5Ej/OhIi34Q1X9HPldIzAh5vXXB
vMUnHHdq7dhvM/bfn1xgcM3X96Uh6yVEhuyJMw2A0ItRwCNiHVBp+Eq3vBcqRIkXEiot4NAzWhlW
7FcenlYWinaDD+QqKdXyw1pBpt3xofdoKR3lL6wL7YTZMDgSb3TazLH+GizRuz4j5HEZp8b61azP
PvOkV9o3kQaE0MR9p14i6V3rmsClmwAiiv+1Mfb2HLvpVaZRCNQRwB1aRQEvKWZcCZ17ZQiGibcO
JP1ho7Z8Ae8YibVi+DsYyNX7Z+HcBkVl8MKfeRpYTN6HyIKApQtotjZcNv7MyX+QrQJpg5ymeyNr
DOi2R3v7e2JFgxQ0E3E2h1efKWqOPrQ7hOVlU83wrNakaGMQrvNXKnQPssrdFoi9dTMjQrnpKQ22
ErykNoZHzrvCcDzeAPuRK9UOCe/JTn3hbxVUT6MX1gw1vMx5eEwcOPj7E8ToDFrIt5OAEk1F+kcb
JwMr5O6lKPTf+qe54P37IE0NrL8EtVdoq50EnaLAH27lmwKgokZZF76efz0uP6QkYZ5DcGmF/qCK
zWElT48ltnTKp/J7p+0/adSLeOXXAbmckoxRMhiOQhUwC8jeVVfFJsT1JfnEeSWF48dHVxArrt4r
l8mAFVOaHGzCQNZZgUWIYY5F7gVma1LFmhXC4uKVffB2TmRKR43eKvUjYAYlzxQSR+o0MCHLKCnG
wsSddslR2DU+kLmIca/E6svL3rnrc9+sZkqqf0mh+JIeklqMB9z0jW9fT+7O4SRltFBaDrFj5RnV
XBu3ZWUVw/SmqMu4CU4Q8touFIgXNJ37lfrMAV+IGj+6BGXFoh6fOjFVd5YbuHvL0d5Hti1qCnE2
wjl/UfIlqpDHWm2zmMSnbTQ7y7wZS7wTJFI+KRGxf73H4xb++AC0YdCvPpSX8JtJmDjxhR64RSgS
OlnfmUNN5yJJ6NQASqSKwivGOP8/TQT+OxDUxBctGLVEBpJOocYcACDVCqV1uzRQE5VhamGMk/Mg
2YdqN55Lqr+8E7ihKx/U2LPKkV39OpS/VwS1Y6+bGyByzaG5gvfeRaYQt0dYlH3IL+oO9hqA+Tea
wVT6Ceq491Nwvci0BgX0X58bn+1kVD9t56W+NJGYefh22ZiEhL7zhtGq9c9SrlPqUBN/bkIC2zcH
HOYKr/ZPCX9KLCou4SjL3t+//VaW0bxs6xsQ4AzseVQ7JrVHNmbktX2QrzNDMyP4DIX08odqNi6f
XfNhQqi0HRSlWIHr5UYRtvQENCmjZMJ1MChRwgYBLnU8VornJuy/RWVRiudrtDyA0IxcYcFxD/n2
5IldPmXux//0x/ou9O1xLS6YVCnVWWVaFA+tvLRoEliIKpK7IY1IhaBFh/RRidUPMQAa5VtmLRsQ
j6BcGsmwBSZp8nxXT5rm+hUTN2dYAScL5ktJeCvgk/DpPog9PklK2+0UCI2Q6AqjUUQHoODOdvML
xRkACUofIS53e8GtquggsaP1WKuI48nsgxg9ejfCBcjacTA9aD1tI4Ncr+gD1PHMJ8lE6LQAx1Y/
RkbQ7Qes+FIEC3W3T2/Af2COWIT2/EeygEruRZQDog07ABhBFnmj62H9AXMSXKqOT1h3NdbuoVOg
6FSF6DyiBibpby8an+MNQQMFskG5QRZK+wV8ogUi9eEbg1Q7kDE0wLgtBAp8gGMSU18840KSCOE1
dKrYZXKs/C43pKJQXeXRJujBQGo0fIHDgCrtyP4oe9E6Ky/puLP5A17XCdJnNci5A09ijE7PVQkh
UIIb608FsJQxUCacYRd+nV8hwRgxWxSv2jgTXREQj1VNZH9iuao54FhGW06c29gv2DnYmFVJX+oP
76uqdcpviYvHFBgYpug135Kona8XFNXiwnlAQXPqKTD6axiv2jEz4MIz6y+QC9tWXlaCeoO02dVT
dscdIv9/2sp9tIopupEQe0EIpVjhgc8FlMAt5p7XiQ9GLIFvsKU7usARRQlWZPliq7yslUx8mSKE
dnAxUkSgeS5yzef5Is27vJUqRRTgVM9MjLe6M7546C4wqrclEPPb3RMpDCuDb8a++dejEqt64hgi
ZTh7nDDLtp9nr/vOeov3rGJSqts8iipO4qkGHGxFW0i8Ol4Hf4REXquE9GAy3rsJZr1TfWgUoSfA
qs8AWmoPwyVtp6iYD5Zn+npq3L6UL6aoCz7++35rukGKja9mj2dlt3+GSt2J1Ealz8lq1IUakVqf
rruI3UOGoCq1cpT2lg0kTa5Y9IwoNaw/7vsAIRYs5i5R2He1Go4I/FPyZd2+Txx3/TSlvkVfW+Ao
nvt81/aLhs9IF3mC9mcXe15SNuW/BdUm1eslPTV6e7jLNbShcFl5sMwIOQZm6VGtdyLdyJxN9ar4
MxrJRECo2u/5tVY+p+VutyJbamR4GMSdEDpp0kFyEIYbuoGOJAkue2puenpZwYa+IspCn6HpozFe
IfQQwIiXnG90niDw6VvH4Yf39wY0Uaxrka/gdv0sSbVceSMF6uwgfv03ZOsKnN3u8isGL1JDA4/Y
qIW0DD3vM7j0e/RmFaPklhFxKESTpdAS6Lj9KUcbAGZu94cXgZ2iGAYxP5sZVSNECyhpMH7LHxY6
/PrfyOpY0DH0wjfN+sRyIE5G5zNB4LcseE9b6YyWgxuQj8HDCS1GmCmW3G1nBEgSI2zXXyFmfeUu
lNOLSNGAMyw/ug/73DtWWJ+TJ0+9SddfolsPZvGEN7mquUQbSXvL+KvBYicBRWoNDkMHHhfIoN28
E5WZI7y/U0uVEnyP7eoKZJO6IEKUGkOYb1pzmkboj8ZK0P41OkKJpudhNlyIdpvCxXGrYRWgvWuW
bta2KBO6ALmqFTc1QGwkKWj4RMozkZodGT/p1p/+cDVnTSCrtrzoRA83z1YvY3N+9eFcQNoaHNdU
NvM1Q1ysyTV/0wssKtngcVVhCb+qCj+5rhEmJ/0SoE5MWm6P0tKmzP2JcP74WxAngiA94m2QLkH2
mBWyq+3sZQoRW3WwhysaGELXXfAsMQpE4duY2NV67HzQsRCwFY7cA+hpfJfZQN9eFQpysSL9VUop
lBIbI5AMaX2UP5+31RBby9OPXlgflPB2s5Lvt+OxWtSLf4D9LfSnmd4MnSCH1kqOWPsmpZ/Cwbei
13rpo5IYIXYJocx0QLCdi6fn7OjkfIPwUjE6TnVVci3hjpfB4QVBr/Ygn7OEydyn2V/e3fPK21M2
lu6xyO09lgbf71V2ByytV0/2Na7NPDkaH/+FRlnkrm/qyImHiT5JcFtbXtV6oLwqN+2GjRTtRwEB
nvYzVHsNYRZb1D4FfN9viqHWa/iu8z3kxVLaOjiJn2t2X9mNM69YhPVYTA+7fKGCfG+ElZqwBoXD
TcyeNRvxqSpnGu7XthWrbkCR/+fs6uvyHvMiPLPd5fbD307mlaT2tYMijPRTblp7HmkAXH408zGW
Asi8t8y7zfrhEodpj+cE6Z1PmQ9gzg/XQtAuL/4HoKKTkdzi6BrfnApULhj85fGuxnGouTnE6AQW
P+EvTYCnGtBiCbz2wswq0y4AwmB1ndz96LEkEiTPPHAsZrotF9fBnNlRpMW35fmiQ+abPkKyekjr
0jUNs4Gjb17rnToNo73HK2yIDAiMVE/LcVo/Gs32ArgNm8djkp6XoCk6ixHSQwGb6I0RRPQzz6ed
D56xpv2xvnGcZKlgK4GvzOzwXGjI0zFT/Pgsx/T/5qSwf8kGeaUZly6V+HUMVW5waK4HQtPn8Fa1
VWmo6359XD+pcNq+CbKcJROgeqbyYJjpYrIfQLVewTEZs5wAI9eSslVSbBc2av3emM9TDCtbgzVX
uu+nf+5s1a5hq3HVMVpXs/v24iXcQkFJ83oaVgs7csClTUysmWU2GDwraGsWA1EG+8xsOVKHLCDI
xeLEydKc1IVfW7pe6XiTcDDkj1Rrn2mDFgtn3OSOe/Rn2RSCnqYA6gx0/L0dkGENOwx8AnqlpK25
quz+t5p+Q07M+KC+ICK5RuoLsO+Gk2xBRHMbCa8JaGbY6tmlwnrdTt7brlsja4yzfiAVTjH7bgB9
NwXnyAohTk09e9nBv+00AqGCXw1f+HADvTGWNFqchtjR02vEM0az+5KtwwtkKsJmdIL4feOa32Z2
oKzeKF2fnrPsXvHYdkKAZF3QSf4iS95cC94POnNur2BKloYDYMFJjxkP4LoDa2P2av2QascM7PGa
HAJ9GZtQlY+cl8GBIM5hMXn6tTLLU8GLdn5xV0evIiWtzLSj5i1NiTcmVbr59RdWQq23mlZ8IndK
T94Ueu8x4Hsle6AyxAaEbDJTbj+EWC52qYjtf/CAnmde7ztbk5YdRC7+pMmsOnfcLVduNETrRsiu
sOUXkJHozFWoTB+mr9di9S8iHqFmlHo4Z511HECDcq5Drry5R9vReZ74qIXQzI3EUxGFHD3Hweob
zomONIGQaMjHa9ar3ZwcLnONspexPn2Z1LZZtFOPXJaMbFvsbaqOFxcCCCkygrYz5XQElKP1Hpgz
9HjoXHNcnI/FOM6uTYWxVrJgtfLfF7GRP4rhKanN8Li6EuJhr5rnmXeiusDxEypItZ8LuFbHUZE9
LjxGjOWnRHrGqBs2hy7lq0/E5LCy/1nf+Wo4tSLrvTwDm2GJcNRjXusQYfW0ZHeTIG0hVuk4DG6n
SOrupa9jNMM22tirCuGp/jTtXYnd+LdKcf8GNM8DvCwe41WOPOSEeNUay/S4Rr2IDauaoO/49nmw
D8Bzsti48OrXYa9NW0atbd3bPik304LS6e9ZXgT4hkFDc+M5CXD3J1wROw3yiyGxJJMsn8Z33lI7
HuZvJiC3nrGhL5x2RE3nnHInxbMhyldjxXN+SIHIPipv8ARp+BYSAKwQegDcrLISbVricFshBZXw
ZAKn+6hCdnMQJ7KAxWSFW426zP77AFDVnkRNJoRKmuR6gxj/iEIiera/K9LHv8XWUMmNyrm5nRFF
1xRlOAcj0sumd761Xty/n+zWeqSKXzgPcHiTl9skZrGEiW7C31k2RDpitao7rtYwfopP4VUT3Nm9
D/qrI4Vr0FiED53QtqcL3ealhfgIenJEo9I1nf2YSaSxzIw39NajSm2VyXpik+V6KMsWCJPX9D9e
VvbZ9FuSayR1A+p0wH4iczihSwpj/Y4REzWW31+xqkqxZMkI/IIUNLfV/fL/ORRAjUnoGUE2RsKy
xIFNkn2u46Hd4xIr4wxaVBrnamPbrMBzW9jsQQzV2//62XWF5ncnJ1BN+gATaYyBCgsYHDUECXQh
cjjhP42Z2sv3eDrkzaPGrUn22Q7JiVfGXtDIsTfJH87/vdQDWPL2zyWZ/+1lgO/BwTh326PGS+Zt
mPqg1rm6ROdRVj2XZwSusmZnNMEll9HegEZ7qgjnGzet83Q6FCX+vz7kXGnN08n3Y1JjAoxj6KOw
nFxVWzb2fZ4OpKWInU2sWoORLPn7HV/SMkXboTY+qwEX9kSNmedGB7u2hxQq85Y7jLQJwiypI9wG
w1J6GIPA0EUPN4w67PQFFX8BRonrXb12ypDlY/lzeYDsAxTQQ1run/7qED4RyuyaQIx0ckLcSCRd
ysAjoskeGam3C0IohuxnoYgdc8rIGossuy88sDRJC5ZwOw8P++m55en43D7soJqJ0n3AaR47nnxR
3rtfpCR393UCGSm7rrfvy5t4OfoeEH/P2cLq8SP59B4+280pyKYdfv6qdWh2GsrScjp5t/qRaOco
NBwOxNxV35bM4IVgnkc2F7YFjGRT+mNrAFaKKCrcWErtHZ5tw9GTeAEK/Mlv0rsFUpgnioj29a6l
+tMAA/fJoxlbzrwLRcdl2pi/NvGZ6FBT5PgzgsIAtX36cPCPjLqdrvVf0tgix/3wiV4kuXsTrXt3
lNlOZqJmKoTpWQOQR9UzvB5IjaY9NFyKt9VEHOn/aikZVqfMneweJeyx3VXj5ivPv6xFtUUq+V96
R6ghulTwhMN0aPqCkSZYBCl72OThWoopS9zc94wg7qV6hEpnOyHPtXSpOMiGKX424XZm917aJvli
iul+9kHQ7MVP2er5JcJDT9cFebJ92ErVfpDe93djbzub4KNHdrb11nGCXPqfX1oOyTgdaYG8FG+y
x8bVEbvnOlnMQervjSUt/fH225eaiXxXtit8XvpKQapwk7006LRZjaqfOj43cfHrpUV2qE9lFK1Q
LkpjLxfdILJ8dbRbHNDGsb3KDJ8rIxUkwu4+iL/m9ROLlf8qM6DBMIEQj39UHJqycq+RuXx/Nb0t
bwGLfbDMvcgi6OpifgSMmnkXyO3XNbnXhdX/1WfAm1aqy4CnMRF0+/rpnL9nCdSV5xlIbuVcAKrR
ttilCMnzPJxK6GRTudzPWDvNQeVSa+JvgaPiQ0QxOR3zmT4cSe0m2ox4C1jtFiQo/dlTjgXA+iNF
wWSPMeI1Tc08p4nHc2dhKIMm4o+GOvYdGKsKgUqUtWPH9dsbXzkzJ6vjLmc0ahZNWwG4M14Dg77w
UDFDobYh+GVUayPx8/nM1CjW0Awnqj102nVN/XP/zdxO5hRHO7jobkh4546PCer0qaeqQetciLob
07BGqdMqP2rdSj88PPOj8Ie/3EEj21TdRiW+C5wfS3CLIuJu+WiOh9PC8P9z751gtVdJ8FkfyUIT
PZR63JrqeWTdsiQ6PR5t+l84TRyeYpGFglBHDC5bqcZTETFBjGzG51d0MJuVnZONjVwVLNIyswH0
gA1KexcOdLVvlooUXN4SZk5tMRExTaEvrxVObW9b6PRqnYaJiNcbUOYWUymzeJR3kj+y/mmhunpx
mTUuzktgz2cXnvfNKCnEIKLMsBanKK4WpsLGEyLEidi44zvTN0DDMisy2x/7MFMtGX37oxxEMrFP
Mi0Hz/U3A85nlNqZDpJLPJdEl5KQnkJmfLqagK+JEVs4ooESwNzYvL9I39cYMufLIrAP8d+VQcyk
tbZaOWYM1ioPvLqAph65p+KIQyZmui+lPRSHMaNRnjckjlx/yX74IlUYHKABc512P+ld/e9Ard7a
eM9zNThDp0ElX4BNIQIZjPhIVc1WVVZCjLnxGA6Jb1qvfA5Zi54iPDx3w52Y/aLX29TSCtRChRov
6PW1obDTfje9N2dMgHctWiqqt07bU2xD3Tm4QK3Ow0nweJ4mPy3DZzAlAhWpZQrE9yHVdxo1fTcO
CrmcdX6KggJ3flivYWaviZ83KQJ4RPwrySkR3uyMIqxnSnszktzdyUgL4TELQnIQ76WPtKMmQuIT
F+T30zxMCXHNZna4zbPktXcko3rsTm7xP+YCivVj7Mr8sxKcWbRH8u4pFI0thS7I2ZgwJovffJb/
lGMVHh3EWHpK2Da0hEe0zuFDPgi7rgpGsPCo1wNh3LHj2gAU9unSfhcpkywPPcYXr0kgGT5kOWL+
tFpEaKOovHNV6RKfCuLIRQT5kAWV5C6jiIcuv9cGUEz2Ux7mNLICdRmq17G99b31Rxol1Tcw1zd8
GiDaL0MnAL37NWYlAQoIVDcnMCn6WUxlgmyfLqVs/tCezxLX+PbA69eFJsxYiX/tEvWkGYiXsXhO
Fk3YSs3ftTgUejprCeILPHIs3PvqVdGDxQgP2oFqU/A6EEuddH/VFDR7cdPBIjetxjAwzqy/pJQa
pQUBinlN2WT72BgBX4uJ0M8QeWXm4pOBJoZclNZPr8flCigHeNn7bR7xetca0f9TUEdDc/5T6DZ+
rlGTA5uSh+UNXqbxJJ1ZlwXzOlnc5aUnEC4Hkghx5mrvUK5D7Y8NtOXD71VK705sq0kmHkxu+jEl
6dngMfGX6+bw7HM4lMfZ4bW1JczhX0K8pRRw7ktb3Gh7f2T70KeWBNNetKLEkCQ2fCtg/Twx9ub6
z3ewrscXmOUGKttCv4+mMTsa2NbObOLZMRx3oHJioA3l8zAWVlS4bxNgPwco1CskCrjS0trfsw7a
WZxJqVhbR2fOn6VCjzoOKb+isFJBWLQBPDxYs9lnaYCmxtemsv1GY0U3yp4jiA1yyq4PeF12Almb
ZSNUlFf3IiS326R0AS0qREhQHg6LDYOBl9UQvWxXZNXf+ovIwgqcelp488K2YPSFie1IhdXj3PSk
fPoRHegW2dvFN408VsU/7QlU4jrjmCii8C/YCQOHDoM8qHVWZrx60LKtCxbg/MJeUfTtHjdAJlKt
rveEcRP16xZdLswcRikjjMOEjRWJ94HI6jWKHs3dn42GPrLAvixoQ4O5Y+H8SoBS9QtnIlXuqQd3
QdecXjS0jeH8t/asppbYkxECGtRRHxLZulsTms4bXlnBGPFcEL452CbrZpmHeZzGkUiwfPwMK4H8
wjnvYaRzk1MsIsz7Qm3Cd3aXl2IZKzbL2fK2u/RATUG0nkWizJxrQ7AjTeEykAqKB46YR80EAQLW
Bt1hS4HHv6NLFv9eIO/hmdtwLNDjc5M/gi/kWBaXMpLvZ5Lw8jRkBOu6z5cQVwWfSq5Hitmr5LIH
tvCM5fuxTrRdNX6Z16XaOlMb5NApm22B8DcTQx1klHJyhU1N6mShS4ODQ6EhIu6pecOv1ZjqtNCQ
mwWnQcgqcBi1S7qHdrGST5f6uEehusipqSSxqwQGhhqOKPZylJSUo6GpbmK4rRJI72BxXcuhafDO
NHhL37ivTCuJTrrNP4XBkLIbtoIC+Cwa2701za8cstAnHEKSsiNVmA4U8sUrHlDUuwFVegSitoyh
1/xFq8nGZD+diZQxK84QIiXYs1YF6JxWHpUjqTgTDOXEimgx0+Zw0gSQ6j2Uu/gXa1fe8GJXFQpr
/Mzam0woMdOIczaLqZdW45FYR1NisM2vXVm/lNW5varULmoskaVgHYauhvYkLzxRr1xCTp+3RBwB
tDnz1F1+VKQxqtN9SpP1RUAU5HHGzPsvPJcOV7ky3B5iCB/lobMo9J3+s8+NazFLc/J80iq7g+HQ
+mUJnInY9RaOreXe1/WvudpjUVosCwZ/pfV2JFOjfWQkkoc5p/1svx9qcxO58/oi5P75JUx56Kgg
SgjK5orFtn8kjveyTYdkCNSkQJUo8IJh30JeSB1FvftgiockifkxwL1XkyO7mJTo6x9nFcWMnx+C
BpwtJjy+KZd0069r4QEyGyO76C/lIEJA4niiYLEYPePaQNGbDZCwu+mqbqyhBq/nB8RXOR759fmS
1HuvoA1vqYlqhTuDZbH6kNjBrCd8sipEKI1Xg+dkLUleYQDyBK2mArQvrnwwSVKWrphLu6SBoC4j
4p7I1g6KntrcGfCWPRF0e7A3+WrJKXgeb7rWQNlLGG47n4esGANgxMK/NOrF7lensSiRXbESXMCL
q+3WRGFNH7VvCMyD8sJFmQqpDn9+B9HdYQctWvgWAi/i5kxSy/3TWdoQeeCFsN3agJmcs1IfRqPt
GqG9ZUwVMFsgAUBntYPZwgHuXSbbGCsWLFIi6b1ZznJMC1foeDqB2N6t482w6QjryUW8KS0s8lpV
IsQFndkqPsy6ZG5tYvDbELqy5TnkJJMeOwGHi0mBQWM4p77MDKLaE4nuZZd4PAYS6gSXqh3eX2ID
I9U2JEpHF8DdyMGc6IRngHLPyg+XkA8r308aqpo8teh2QMWZa5QaMDJnKolsbHmgLrITcTxX0NvF
UC78v0ju8q7iLA+kCFzY30G5ydXWw4YK7arJE2jiBoKYuSfEtPZ9Lu+uVyT1eWuOUZH37Zo1bVyG
tEsLi5je2MQw34tNWdjJYJq3ufL8aSawbuIdfUU0BlzimJG6AycGg7X7B+ZeuU2FnbRsTiqjnL1a
nyZyoHuoe5nLEX4q/p76i5pVxitDBHcub/dPPdrNrCBZGoHJLwpOQ23XLGcj2o0grjqra7B36hh4
+BOvuPEhM5nVVlCwBdl5Ub5uYuTTqoa87Lzxy/F4owFtWHdkehKudktFD0cKFaU14HN9JKTazHOw
dRsxrSqPi6yGRHK8Yy+WNT1gkGpkvDit4qH4UJBc0+zLXHhAlHCq4ySKJKhR0PNk2rHlHocGabvM
+YPJ7UAtg9GW6zylvHofQT+v4lNojcFyjXuBKZPBByztQvOVTQJ2m1VmBGC48tqwTdS7wUL0YeEo
xVw+Dj7x2i3dHxt5IhTX1vZKtvfFplRSkUxhzxXfUu5mdX2hJ3OU6Mxo1ye73gQuOZk/MaDdKNTp
YANecxANV92cPLF6LyJruWSQDMOpE9ZZuxZTuwPUIEQST0XcuYvv2X+iN6/p1W94y/zK6cMl267Z
/SuujroznLS4XBgS9VZakc99L8K7mCG0puG0GUYBQZRQse6BQXykDf36Ce2ZxmP8kIBatAkY2CAu
ocG7XBI9hrw/lZlW37Ki7fArs3F70b4DnVU8ZvPCACh6TlZZX/2L0YE4NQ1dCT8c6zQ0/Nh6PGmT
4ww6T6F+IGgm99PJfc4LbBuU1p12KewAqIjcdBjvJBQO0ecqeoltS4yO1jvsnPCyUZ56LeuN7Vf8
i/nPho0C+g5yRivT07parhEm5YQ6m/MdXztwGJCR3/66VfN3CRhrpBSpRGk4KC/FO3JI20nettP/
0PS3bLVeZiQBIY9K4EFvTBxZSy4ntuY+eXgER5M1fiedQb2aF4qmGElOlIu7IB2OktMwiYPdCvIH
vjEfpmj213dV8ye9RRsJppkFpPddT8jtFlOjRj6yxq6VGk57GkJbb/BxAoSaxJWDPp30ZBSL+CeL
T/fpSpxbYU4xJPWytRNeQcNiWFL8MwXltNn6RdmPMt6pCLGCqRpKQn5lF7vqKOvM0bGNCmgzb1PI
+PraLHj7WyAYSgSaesX1iKmvNE5HzSF7eSuc9Fbgdh6HNcM97MKsYHwhcjfZCNNzhhf3dVjJ6lCv
bo+l/XlUvnB+PS2nbl8BuIOGhsVAtlzcAj8eqtAzfZ1goCA+bEFu8MxMJOGWb9zP4vMKMyJoGHkt
GctBqpKSoAky95MYvGFEzCKs+gLhALHZzYofswrWtYHSsMN2W5cCxi9/Dui5Lov0zBO6tmx7RCSh
EaMeSrBpHTlmPuUqCkUWQ/ZVROuZj4WavsFrm9KSwFVPUP66aAHyHtod589Y/Nu4bleujMeGuP9j
RTBfk7z6+Ei6SZ8z+xOTL0yUf6SsmunV2yBzv2FxjB6r34VhrZxjaChahRMNAFtCjwynYZW6++cT
aXSXp370jhDn6Ls5QJGRsAmEzdneTEp3f8UIJOlTHRnvabWb8HvxBr3Mor0fPd2/0I8RxgZelQGQ
YVWmXhkShqzNGpuf2edIMDqFHU+6q9tffyP3TQKblSNyTCQd3kLWr3MKmi40NL9W/cRUs1u5Vnbo
MpxVFlpBKvr8VYaJv6K+ezRjoR6B+QlhT3NSL+mzpeHVavYqb2sOZP8lgfLuzzONZuW174wkxWcn
3kmIV/dJ2AKUgwFLw/UlWyMYRxOj8qarvLzVSKdbNID2w8uL8Owc2+RbnSL0d5s8gN8NwOpCFQ3j
v3mS1B29QRVXPuatLW3Tj7tUmp9fFdOjqUHqOxLhSR4PszSLX8Jhd3qRjkog3t/EXLFpVBx6Bagl
G5LFZAmhREDuj8SF9EmgkIDbV1hbGW2uACbEOyPoMvzt0ugM1lR0fYkfW5jMSfwFQvRupPSS6cZf
Jn15+fs8MEgZSDOiqtUWdTFfWVmwv2vw8+EuoQpvL2qmDY5lIaEmhJ+GQ/6NEEb9MzVakTUccQcw
haiYTQiIWaTgn/ZqtZeOAc/S1k+yWoRXhlNJPuVubStLZpe1PCWjPsRVDYfRxt/glwLVm0yssCp/
B+VqAwPe7FKAVNSUzVQvuGdaPqkY//h0WRv0GxpVdFUb8PMjAB7z9gKO03SJ5NyC6jCGlc6R11+a
VSfU373qLPAPYRH02frGQtenOAmmMO+26sej7GIPfO4JNUrqYg/nQxTK80Nkwkbkibff96qIGQNm
MCfgluXNQ4SwsZBhnXM8u1khH4U6p2Er1/iKAUZzQa+gc/URqAle/VkjNSDHfWfAUiPOxdCaYE26
CE7yS/+0JND8RVC6rtYNk2SbdD2+vNm7+4/rMauPeaDo3hc9yesaMGgYOcD1P6squKE2IJAlXm1f
b1b3r2391a5VQmJCXpHJemoIzbhV2fy6/iW/BpXUQyIxqBZJe0mcihblAvwA1K/CsDrS6nqEmPb6
CmTiGmbRKIkpejN1bjCVsVjHELxTIVKHfKaBgLCrF6txmYY6ckzDXBU335SJYZtNSY5gYbM8mtb6
eWTMikiFXOkI1Ysj/h60Y3Nx1PyLR8YsM3Udu+LZhV65QScIBfPJz5KRdKdCKClmpwPIYMqzGomP
z7veyjectVxwCkpaPAlu5g9uOnZjIbdBtpmipIUrwQ5Y6CEF7vSFupmPmQKCzheqpca5u+ob+6PZ
WgJ2YYXbVbtp9psboPCLrC8eGlxfCBfqQCBlbqHNXZiPASHvJZ6gaJ5w8X8nf5o8YD499lYdBwKg
NXp3OTHGoVcKJ8HhfRUSMjP4mb9TIYxnefF6w/aDfxibd5XwuvhN1qmR9J+4P/CqRqUP6ndMGR6t
xAyyyUEKY0tN2+UZKlcJT2XZiL8ofHYknnIsSOQL4a3HRDxLnrtsxSlcFtwEND8qWlojQeHaBEfz
6byV5K4phoV4YuBAcnek7Yc0a8XY5vXNhl8DfDY2zO6AfRITwBIXp9aEVq+4MJjxTKqnKUi0qpXa
/ht5ayun0rY3TnEQpsHC1Xu28izzkgdMbLrJz3g31Q9+DLjaZ7JpgaYOkh62bup72loMi067gBnK
w8aftSrQrdgey8OqIJaa+ljW+aAkbkyaXvYmzZ/8C6ykyIpRewwIlhhly5EITBQTMBPG2fC8UQsu
TGbPfQEwdxtJrM8gbOoB/+eWJpA3T/p80IKnLhqy1rqauUFN9BSlbwC9D+jw3t6N94hF0qVxRz93
AkP7fB8ETI/8HiDi1KFJtMENeNhcm+VsjVpob4gYkVmiQJ4PMrtSaJJ7eHuaSJftPRdPIuIlQgJa
bHh1PvNQYb8MM/ifhTy/qQkFhh4t9hUWi9xP4T7fF49sSsCX0ljehvOOSrOqPcBAKW5Dbo8vYbVU
f9kKAleTltH6cy/3gIRdgo4XRt8PV7M4PZv7Ib7YMTVWULBrHX2WZidd+w4Azih2CsjhkLTRr4n1
T4GcmiVqeLXm+k7/nU60mFV4xU3IjO/l3EsmV4cSb3xwxgjAHiOv98GUeAl+756qAuKiPfwa7rOi
eH4Wq8ZZxnWbEfF+dBq68mSzIvpcMjFiDKUvRC2CF4SN5xQFqhYrUaJL82FhmdVg7kp6rpkRt3+Q
KklUNHJAWpWc/irbCPdUETtp++qR8AfcbrMpmG5jvk7H+7hkOGj/s4gSFrKk8KVewe6tXgAn5UFC
a6AK1hgmhMaFPMkFCGqlx8Nn3a4la0mhduOUj6S3W2WhbETRgTwquYcNDD7JwYBSAx6za9MVG/cg
ex6eGkL461Fero6Hf6yEP5jJi0wkevc/GDcCX9a7QQebtPTB2O/kGrHsl0UJpt9y2/xamMBGInht
I3FB9siuVSiDmMCEcoOyX0SPGDNbxTdpP6eSZRpv35vQoxlXKDPYuTgymbcCOY05YEXCgFfM75MF
FCp8Cg9z4GH63+lCKd7TcBWCEkVEwPRjlRhVWhl0FNVDpkZszNiE5YoQnlcyeZD/dBHdaFoyLud/
vqyq4Jbit/xaYw9ivIqnU/nI7bumyFETB/Or7srtr+f7GRGu6zMMH98rVC+1QLBsOKLw/KwXF3J2
hdHagGqC1zKiL1Yl49o3/WVPG4ls7mdvmhVVtnFZcT5WHs2zxU3dGyce0LlfNfVe49HXpXYoGN1C
NNeccEV7w0OEQzEiaLU5r8okPzhMtDvZhqlaKsGFuakGYNV85As6FXiZdmfpl+/UsnrmMusLi1WH
tkPSnSQPdRbW6EFBC3ius7LIenMfhJ6P5eOB9ONoYlEeuA6nAvFiYrJvSQo/xlILUuElRzGdpOtF
6+3vB/jk9GEIQZE2K8TwLAQ7qUKm3u+8IbptOSm3j62wScRk5v3QsTIYPwfxbqd8Xn4sZtIJxwKq
8sPVrvQllrtuqYNPpC495vxl0AXYSm/dOVdIWCN5oQwdjuaTYrtUpfYcRltBuJRqPCQJwdWKRYmV
LrTHoIF6AE44VXhk7fkrJyJXaHjg0R8j28XD/ZXv4YQO/W+A+KWaoXS8a8RjbkbbdcHkRGmCRywM
oMG6U1yLh0YeiiC4iPEvjNlTKmui002SSjs/2ZxnxUPNeLy7Q3NKniBajjW9AG/WHQ+ZmYkhhYqf
DS9jIjCY7+R9jXBPXJYvZEctAmMxjw8/Np6ql+9gM0r3sX0Sd45J35P02pzQ+Nqu8+LY0/Ew5iuv
MvWkLi9PCucQaqT4USw4+76roZRG7fT0aDkxiWgLMqZHizHfvl1FsVLhhKvi2DGkG4pA0tDjhqcJ
fKvGmrWpSXJUjs/+XJ93ANcGdK6IC8tDiI3unT5XyAOWzHlanUCCQk7oixmy7S7/5RrQ+n/MlaKM
Nuwh8LRcbmVa17sAZ35jH2DS+NOgqWYKn3UXT/FO6WDzcFIDMn+7rxGrcLgQnsJ+8opNfcBDJf+H
niwMiFJTzLlly1Bd4Z6SiZKHC7wDBEkhapI7JSjp1I3h3whNr62ule/0PhCQ4YXNBeakab3YiQlB
1ia60bpRbrFK+h2yNDqsbzebuZ1i+9fQGL5+DVAlk+Cn1pK42MHFWhuLd3xj6EZ6subI12VDSb/0
rYdeZ+YiTcxYB2EkoGx/qgWThjt3ag8hSxVx3R3OWq1PVfPf+Zm7grt0ti1UsToK1uC1Ef/bmBjK
9d9VMQCXKb/SZgk46oIShiCq7yfJW79GDqz9iKrUZqefA5UCp2JJHLm1/t/hkHY2jzz7GGefr/+l
ydjzwH9vyEVvpoIntEVz5+E68tm0OlEBfdyoBWqdlSn+zrh1zk1FWM05KvwZdm2b8pf9AoNc0RXi
vGT5ELXD4ofsIisXb3ZPaOcP9+JVGwCINc3ZPtm7ifD2dwhcN4f7eAaaQbdHgtaVx7ByF9zcqHYj
MYQtn4VDfHhTvhITty6GX8hG/InOdYBwkGuQvvGDKtTD3QdaAlIseBx0ZcpSmFmQZkO5mix2GwCp
6H2ppwR5pGc1S8+8dBiSWuMQO7+rHW9SbfwdRao374ycDe0AHvqhv5gErlCdKkuEg7posRRpw64A
W5ASm9FEDXjTx6FcMgiGUhoFNPYEEvg+cwHxVUaZ4OAq1bSlwMuhHONJ4kiq/MfLozuNOE6PlPMn
4HqA2uGH9qf32KlDyoEGODOsaO0XQTunS801aLL0UL2KvprSBtranhMuEOTaqH0zUcpB9unUUzRZ
b/wpVet4byjmYpLuDu8zxgBzGN/U1OgOVRu/RU/fUrAWdt1iJ6TY1qA9niGmd6blPoPb7meUV1wH
8soA2toqtbzXgdh7l6QmE4DkiQhCnp6Jfx5g/2F/1yalFCy19cKKiy8wf55QOHrK+bJ291Qes0Ss
2VR/v0fMk2J6yRnGA+4k7IqQXLCMkiH+yleyAKTS8o6n3PjnBOchDJtUq/jQPjoGDCUZ8nhTagug
Egh9ITiYH5EpVWPzp4phZrVuSBKbjeCq2jTy1D0QpY6j3sNkcUf2o+CCDgVuPgIlWNhAWp3oIeRh
GvNxRja5bDS8We91TdFGjoKv+e/QShjwHtczKo10D03GbNjxCUJdcj2au/ez5Aj8UQEOXXe/C2SO
9HdJb7m4aiCddEpuPvEnmIiaW1ijmgni1HY7eMnkSJDRBC8LV8w04WC8To+qewX3TENau1RWzdrY
u/dRc/nWVN+Z6LYN5fEFlyN8uZ5m6iMtqBLEwwokmAYaB4QgnZ33Gt7XpvPs9yw0FiEwuPK+5jYx
faqUKcyLr8njYeT5DeK7hHKXT3ZGjgExF1YK6X/Wmeq6dIyp2Kp1CrGYr0PfO3vMejc34K4dg08K
1eCfoq0Bw9qe5Pj67QGuQVEC60d3c9H3wabl1RcNCfh18rpoQVGDV8Ltb17hOOSEXkw9V3E1QXHr
Q+qWpUtqm8vT90/BAYWteLaChvCqapfXmzE5suKOIfEfxdECqB7NmeI2t3ESDV6hcCtQS/ZZphLO
jMrvHHmuGXaFLMaIsTJaccO7ZHrQchnpqvcxUwd1lPgrpr5Th8xr+8MhRnEoTs8KDMCC3jA/jjG4
Gm+PceOa6lEWyqZNQXkYX8IDeEu8Cjrokx4mwawdbPVJNlaMQSTlgH1xi4r8Mz9ymP030gmzTA+x
Kh9dmFdn5sabgS1HlTu6ZMvkaNaOwmKJ3MYHFBOAY3Vs/ZyCbzRPQ4qI8HEbmMOPlDBke+r9INyu
vnZLvS73rKw77eJQ0mIWkoygLCWE3MYJ49k2SFUaH+CAvQgCtjfjddjtKhprK8QQwOPf5dXjTLiL
TsBXPHl8jKtDRkl9krXadd7zXwrUgzgcgv+yL/DHR8/+YzsgVEU+kPCPBZMgDV54HtYAQEwTD3fa
0wlvTtMDYUSXyX4uZv9yqMWmva2yR0neKBt1ZQZhLNRK6iMGuQRB4/jiPgQnKnuyy9w9aS2FbFqB
zhV3sZrRhOPhjfHb6wfw2pUjqi2kZ54yygA/YlVzOlE79ND0xa819uIVuf50fNh6FbMFoy8epRea
1vAFQlyWGngLP2MXQBLpPSkXdN8rITifwPpvTdlc6suUh/rcztyz6tw7V9mItfaesYmWtnqYf48w
yWVSft7KGaOJGnNIA80MRZ0NGyt4XNZQTPT/ja2zT932WBdUwOMMx2dwjXNVvYP3k+EoH9oMWP1P
sKHViGiWpdqRpElSos9rXspgk3QAdy3Y9PBCU8wJLhpqjdEP9j7E0UFYGNqvGx0ImKfY9T/dTrC5
rsfbCxA7XHAdD/4Am3Dl5X7cl4P1IG6Iew2mhTDi80H+1J2nBfM6/PORuPgCoo+LKe9UJfaOfYxy
W5HClLeycCyBQhcJO8qxJwVaSY+BKh++BHsdiype2kWANY+fcc91UoFnJNNeKFFjT1zAuhzZIndm
M9uFX1yAXeKFLQKm43iw+c1dinhcdR47oKGC4bkGjJZmWdRi2WNrsms+cJJ6D2i6PTFIUiEblrkM
3wd+CixE8fKr0pMYflYhiPBeUPTt7Cud6x/tuVdgZDteiU0bSAd58Kyo6yBd/4XVtFlfOUVSbinO
0m2Nk0nDe4aExtecNQPKAa2IuUGudmq8W0KINLv6sLBMaIBhUfsOq7RdY+Q4nLoWyTDL88j8waR4
03yY3F3kVdOQGCRns7m6Nt3K7Q+S2UZnNHW91Mh3W4Rf6nYsHH4Y9WXkvhR5b5cRGz93TsRCtcaa
GaVMyknAyEOur9iLjcRW+JpF01y5ra3QBewD8Y8tbRFPeJNCRLeQ2gM3mkQkR7iQXtHfPGq9iKkc
lHwRSWEVlNpIiZdS90k0d87KelpfVf8gr1dsBltL7AZ5eOld3PJVEwlJXXmmpXH9XMhCmzHeS9mm
qirTcZe93TpT5zDb3SHxx0xqOcVLb9l6/vv1ZK7FRRdlpgeGIwyLU9PpZrBPMTUgOYZrmEoqyFmc
z9fne1KmeXrcY8af1ozk9pB0qJ/l/EJg2oxbUXxPT79PAVm3tB81wmG2c/DNdvJwsX3WUFqg7EaD
YpWhmmNJJevI5yh2RdlEs+L88swN/RYJPUMLfqdKAwnERVfqUx5Qa2r3JnMl+96NG/ItlDAPDbDg
dOCSWniJPNiBuBZLFzT+T64E8IvelC2Gz4DU1LVhNt96K0stt7vWv3unOsm32N/MFf9wTBCHSFxn
FUP5usOCWggsy7FhUlYUofiPcfbBtyb6X6dBj/CTluMsvu/AFYg90tFwytvMghyah7inaOFSopS5
68TNHDVrgyasyrZzzFXsMbDV1OXrqWBQc9Tjco/bk+G+7E3ALaqDZlEDuaOTr686Tn1RapgOj2D0
Vrux6d0/U7EE3KjAEZj2THvYWUAPerpznUDT03Tom21XtI8MXJg0Ka0D348Q9JrGLSDkXLegCRFK
7c9eeObvvo09SGUUx8pPNUmjhTJf67aRSA+0uDhNy6qI7GBEI3562KyzIgdsMGbBv8sXfVjLS7G0
FtqH9IJ3tQz1SvCfGdTfQY01NQIcgWDi3ubqWj9UQdHW7eCtE/Qxx/nCn6khR+rTXGf2JQczpOOn
hyOH6lERL4c3jjWHz/qFoxvwEbF+6kYpljwJ5aBfO/H5o/WbjYZ54rAYODXUHgzL8fuDKK3RKJkl
ngAKLLvdbtsW2eOU0huf7Y1rZZNbs2NymnJj20G+boslpfkuxlQpw0titJ7pxnkHIK4TNUUYb7QK
3f6bawu/9CKQJEO8QCqSGULmWguHq67I/DbqlIyh+r33hTShRm35vRr3iXx6+Z5yexDSLtOiRXnM
w4gT9b0YFLKtjx8aVVkmI4TcQQvcX+OG6vyjDPeH59qwWQhzu0NXX4FULybiNYaNhftecHREldNx
KDK6nRS0/KYggbNaBcmR7yZ7+2saNsU4M3Cll5l5HOPfnfpaUq4EZ6TRVQbJRVRUAEit4R4AW7B+
CHinQuWGAVDO6324p+WEtw0/XA1PW8JRQRMZOJSRcvJ+3VEa2RMu1cc4fY7QwHYhAAyhIYIl2gh8
zY64GJw9mGGVe1+dAi0pLhubStLgpb5dnP8glg3NyArXNYVFVQblRbgjbCanhKv4PcuUK9GdTGkC
6Buw2Jqh+Az4tiCEXaIqx1H2coWSl1g342liXBcCVwhn/deui60QkLEix5kP2Jm/i5UkEvrUsOIA
JfsV/ZCmO3IPopmroYtxGwU7azcFwhnwOrIt9H2hgoPdq/txDJIQy0nj3WYE7Vb+24cU/sDNyN1M
AxuMs41n/iOkoS1tclOUcNl8qowjlX3epKWaajlaJvzYAWOSTpMUWMThcC9TBKx9oDlIEnZT0hco
I5u47b0GGMXF0hhB8VaU5Dp5pKEs82DHfUDl+vRLFaXwdKgTJKVz0dwlZSu3jwJERqbyLv5ldjs2
IeUPEqWHtmRgI+iJ80u7UcrgL+l/WG9HKkWpbqwZx5eH8QtzwN6e7Mz+7Li8bzsisSYW8iuFewYW
nGzdhYNpElE7K1Swx2moS2gDC/uBRTb/6Gpdyu/Db5F9Dgy10N0S0czCNadgC7neFZk2vGDzZnLK
d1tDrHYPdPyjFzuw3KCysZr4c5ajWkSXGyM0gqMv1zH8rH5QF5rS6ENTrUyOrVfyYRt/megcBhXX
OAOQh0/hAmVfrM3QvB/wfpXR4jAQ7Lni6QpL8jEzFz45NimMUG5Aqq8bC0/GoE8rndPhtL6FMnFs
Sj/HN6r3gR7VpDzYnanO/62UIrVLdCc6y8nEaxbTFngyISJN/Y6i4QWebWBlm/JnH7viR8ADl9Cs
MldJaErbzBN70QhZO+JZ0XjLvQYgx+uiiKrFPdcIV1i/OxDrB/5Nwi6ElgQBdLchX0VOnlYyvyP/
bPGcl20j/X25+R1hzU0s9au0lgysJtfxFsT6U8wnPBXpP7dXw/9/c+Q5RnjBKqyGAoF8u9rizzt2
mZ7pD0e0kwHH+/CnXUjCqyeaMynpZnqYnuym9fD7bwkUQCBTpvy4cGkxYd4bt1s5hLc9X9ExAbZA
L1JHUoBUSi/F2xMTfBSV7M/wExzDj5mjb87YybFar/GFVjmY3l4ulCvGF0TYrsgAcp/ejeP9D2Q+
dyz9neSdUMs10AkGrZuAIZRFLajnQHo0d0tSQEi1KCFv6PHKkqhciSA00mA5H/8ucXu2dBxogEBB
BFeGb2eP/reBNx6JG8uFsljCFDZdqlmWFyTPa+dHs7fyMAObpO1tiLrKE1IU86r50iTdg67ca8Fq
xPBiJe8Aajv2mGAwUAypAJH4ENlyjL/1RVjEVzb37eeUBq/m0DrgSp5acNcb+x5ZDtlowDIR0MTo
K4677uTIvwPaMBu5RhlvPRVgWZklVBS9CXWEdjYfEOstOOT3RjYawyapU6HMoncsU545RpLqh+nb
tUIJ6xdMNPCwvdpkT0LjTAlSvUDazq7h1uw+jf4bzlwWxCJD7IRNmIcR5ekVp5jUGFuyuKHzVuiI
dw+ILOUdZncI+ogGEAD+rP1yuyXOPC0nqwbfr3xScjyj48qgfnnC4ujf1jCKdHZAPf6jfmIg2UN1
uGJiAOsYqN+v49l6TolN0lpbsRUfUtOHP0LbjnsGYanOBeJ39ycmq1BWmIZUjJdTZYtVjwUOMpDu
Ci2g6lywCSQdy/7o+jkCpSbRbBFzr64Y2Z79144txaaOEgo4bSaE6zdx8WiNzvs7fJZUWWKfIP3n
pW6aZjSd28Jfum3iizwr9cvNqKGav3K13uhAMzmBhY/CoV9N0EtBbo8S0BGUKMgWgCu4QnTJp81o
HyUSxps+9ZQFaUWkN7J0uEZjyDs6qC/jyb5p6W5yO5PTzQTUHiZyV5aX7kw9T9y5HQ0gvWoRWrUg
o07QTx1A5Z7ZAT9qYhdi7456sLwGbvzpIMxJa31wB4kpv40oG8ZX2XTc5tt4U4j8YM4mO5zBDIhJ
XQkm2HQ9YPxJxGfaO8YFvbwYSFUqmSDsaO0SiTYPfId5pCEW9EfFWEmkEMB7b+icR0WQH4vh2geB
mCjvpe7amntUQ9awXuQtkPIga4U15bv2xn2fax7TpMJjkOLzJeQmyLgwPZX9bMESJhtuvy4+h/9F
+xP3Ns1ldIpfsOtNc6r3DHI4KcxM25aZO9YYWbcpg+kPEim+NPMDQmJ6eYxV+wzXYAmqy5EWoE4Z
6WCVcph/dhRng1ywvGe+/eqD+ysm+Q40SFeTTUYrxOqgw8hvrd73f6xXC1krWHLhuytswzmB+myA
MKtEyJO13gCrcDzsf0pkKkIa0XLfzFtzZa4C1vmZQ/Rqm6IVASdye/xmEz+LY4UJr+dpyvIS3ZXs
GUItyf5Z650IK8nAQaN9AnTgroltvf6RjEkCZc/lCv5JRqYEIgfRUepogeknv95RSSqHo/A5RUhe
GmLCE1kpHvFy+NpVn5vQLEXbLYJduFSweSmP76IKNVpNDJ8qMt3102TM5ps4/DC4FBv5UyW5oXW0
37gAt/l7b3MeItyhd6yj20kIWdnDw+h4INKvA2A367DPxTtx5tSD+/5dVff+jYt6bMcHN+9Njovw
D3yD6DRxSmlyW0ROfT2em0MNL5qy5jQO3UQO+HYiiseUk1PqBQjY2Z8Oj+yCVoVkRpTnsIW+/lfV
8xg7O2rRcHa2uAbnDyUVrl9pKnFQO6ZrOLwLbBUgL4XUBv/MYKR6qsiRm0RHQDVhEalxHAGlgYmz
fbC7HqjzR72VpT768qo7zAXP8+tpLxiid6GlR/foNkUdMT01lMQHaRjCWjfA1OnBzkJBW+Yl7LCI
oxgioFFluT3/zq/7FU4xV2gGKOaqE+/pRs8EoYIN7o2+5iopO54f/l7flNeC/iDOYlkiSFRf44ro
AMcMTTyz0Ak6aYKzKvbkR0r3K3hckQhSCdO1jql1NC7s5FnXmadinfXRJ4xn9n8AD41DQowBQmGQ
unQWUhwVWtPZhK/1fvML+kN6pNAvORrcyNv6COJ2Jjx1O2y0Kuny9htsw6EfNZpfEZ3R2ui2IqWM
GvJiG1s+tcjwQzwYtHmVyanp51eV1Uh9dBQ+cJLohEb45chnJrUUxXYX6830Rla4tN1gGjkmGmRp
7hbRivgND3V3uJMtYy2eAETUm8D4MuQbl/eSJQMGiQnK+2MycAAUaYFI2z+0XTr9tyXvxT77MGWz
e1XaFBgHS/DhTplZOQrw9H/bUr4P6PYuq1RWn8GFREL+5Eaawnx8VPUF+HPBlihzyYdu/w4wwLL9
yzN/bHg4P5WB8xMtlaZHlifADJQ9H/WDhOVEO/6UCNVN78BvXuPBA4QNdbURv3MqKB/MCzr7RUnj
l+zjzM0VpHCvXuWJljoYO5KFGRJK1rsvlxWkRWYttr4vyYLueF3l+frKZ7ptjLXqRDchvn2/euxe
JUnK+NTNaNtxHPNcRbf2Rnnuq++kggFxl5BsrIe9pY1xPBllM5A8ULZW1bl0yUQ0UcvhZPs+NC1R
T0N+rfPNCnA5oYNTGkIfd56fO2Lk8gxq5qdpaiD7qrhV2Y/cdhTY4ZhCyzbhcmr6gMuuUlvm74mD
s8xKHaodjgqOa/UDMP8EC99XdtFjaBtEURAwJjzi2kI4OdvM8TtDu+5qKI0dTaizH72gWi7g8EYQ
9T+NL1XIXwtHIq8YucY+tm1z5Fb/JfOJ9ThNV5VuE3j9CyN2b6/7HOU7KSd5GsNjYeqamsqv+J58
4BxhG4XaY7ocEDrs869QqJtWkrxlkqnhhwvvIdZdLkbpMdJ/MR+kRDuosMhRERmLIm3P1A70lfH5
GM9bEE1XVbG/8FQU1Y3jeC7kcea3tWMjnWJCOLgTKxdeucDLILRAaG7IoIlb47cjOkyNN6pUQ0X6
ZD0QNg/eg4t9JFdITZgWYJWIIFVr2y/NXnUt9LSf4me/VxmtkjuQQ6o+GcvF//c9hi62np6EjejI
muD+kCUGtauYkTFkJ7GPiAOjUZt0CcesLLMA8igK3MsJVfKc04kydorAIcVnFUWK+q0EJv32AQnN
luN4l2ROt1WJ/g1gBtTrUZTde/GpPS9ZckfWDc2DlBbxgDTeJlU4ocVI2ip1Pt93Fh59M0vdj5dZ
P4KFBKQCuZnCSBq6BeJUL5+LLZx7/PhOGoXckHOCIREjdQTFeNpRm5vi4SE/vRaJXMc7jo21MRMr
fX6ny7XH4qVrp/OIcoclJrOrfZJhZuPNsUzJyCrERis1LB22VvLDrRq1YM4ZvsIWwgBSqy8E00cx
TzEYsjGQFZd+Kn1q+OL52ifk4TgwI+0OKfLPfLgjanfBDIdFydj0XA0PksUTXzwHqDE9UIo+VtMO
dcX+hWROxFGz6GAIHeLcjNH+68j8JCpO3FapK25AbwntvRbaH3bNPyWHjHktMqQ9tw8+fay7oNPS
vq3M3WAUZa9Q/S83EEUQUl+Ye1Z80wztIHJS+j1S4OmI2D/mdlj0xgBeW3egWyV6zfnwV2Pwh+dd
3maPF4cFuUBNu9Yd5Efp8zKimUuDJ+tmPL9+Ug/2mTKIzwMw09mvUNjnbb4POHMQp/A13Sg14qy1
0Oa32VQKtdwE429nz4phiBAdzD8Z0b6XKDbuw3KE9nVTgi6b/VDH2WfFXK9D5cssjza2N7iHbO45
T7Tj1l70qIxiUl0s2v4XCey4CWEa5nqqbD+h5djwgtiF/2jYvgQCygnLJmCnYb8UIbNvSntwODta
P+ko+CSitv+5qZp0O2gk5Hjifc+FZI+NAmcEcqEmHoY1REKeu0Ysn+AHzyg2mpVpQe3zNXjekUFJ
ChhrUtc1EVyOd5BqBKCc5ZeCDETKHM7SZ2wD6bjhjjAUUnSv4Y4KXltPcdUBxMvg+qYP+rG4Qz8K
jC57K9fl8P0NBcJJnyidqrbhJTlyQ4WMUJsBI/1IYHKDhKf5ewcGnYf+hUYjgsMgNEoZ3cxTcBMP
9yvCoLyNca1DyVx/nWbx8M7fh8IuMxCAIfOUo1zbrdcw0wOTMpyTU3o6xK7YNCMLmcjE+mIkaUr2
KIlp3KSthhHnCiabRZAotOL/RWDgGeOF5wqTeBEjtFepA6wCmqu+vE58zkPba6ZDReyrzjPZ3D8m
bCHMvBDqD9NYm4kHe7Ie3rpwyUXPOcDG4BKcfX2f3+91lVXhhB6sBvnG/L+KU9TqY4Dl2uqVy/Zg
Vb/SVbT/f0D7OGm89COwplgzBbIrMDsMJKTxqv/CedSU+BYq5uWHolSPViplzkvyUTYGY+bnxhfQ
2SWzjS52E//VyggzOiFT3cWa+83/digmfJmmCH0diGd/BcPMztLyidyyGBj6wG+xkc9Xg4ZAtujU
yrxvDh/Q1OOkRU1cbI8YxcUSFh/4C4kiN9DasiNdWjKqgQVfR2JmJmnhv7BbnNIExrR8AvVpVjXg
dlhlRX1M1qTKc4lZe9A+FErnNpvk8xn8Eu0AYuNjuijkjj7CBrCn0ZTnjsfNd4ouSzfXvOGyxJUK
cHo+ZPZlmyC1tZBfUiNo30EPgbUotUS+YagABIwvx3eAdn7H19UkeTtn1JcfeBXRhn28T1Gb+0ml
YjStcQRDDOrJ1MZByZTmc68k8W5Y8BHNqsT9gFoj5rmH3XB2MMEjpE9pAGa+Uy4tvUxNVOIpocOC
K9kA7hkUwGsCKL3pw1gbCvQ5GEPcSDyPDDJE+hb7Mb/EoXNFTOOXgE2y+0BYaiFVI4rNLiYm73+g
T1HXJy5IWyh82nI+e1T+EsAKbhWA8M+LWHXKqfC6dw4Lu1ikL/I1MBBShKTDDYWup9ebqqFN+YCo
rqqEZsIGpCyNc830lDpLex5CZsoz3VcCDXEVX3SVPxTj2Dcu1C8Rau6Du+YLgmsXddkWMF+heTT/
fRwIazO4lhVEUmuhboBXpXzKtaN8KqUA1D1hq08hI/mRBUlu7ySUsL/IN94THdwDNyAw7eKxHdRW
W6vOyCaKSquYs66+yCrFkVAPuEJ/1fkSm9Xd9hKj2koxO0OVp25QeTMt1UADyhTVOueTnbaXnUmK
4cQgAix7ykKnsrC9dvrFNKzEfZrH7bv5iQAIjOYvBdZ52aBMx4+bT2CsyV+Zr7AE8D95BgiFktsh
xXMLfvSvqzR4d8u6kNKNT06K3hduac5CHaRLAp8o07tD6cXzFab0w+w4CeOGbsd2JantHOvsSJ1z
JdZfYHUf10arx5WESZ+wiui66VsD7UGTKZq0uy8CVkix7QS79lB2aeeh22JzTdNzozs5ZPUfqhfU
8tFaQu4lfrJfHD3ByOSJrdt0zFpG1HB+A55zpDdGOB8NEieNIRISf3zJPs8QeGzSFgME6QZgNsSG
eBq3CGy8+F3PbBP8wfIoA07RacvMBajCkEoEKvPZ3HXPtV0HrTof4y3Ioq4nQ6VfeAgvC/4U8B1K
6VMNm25wJGWGoVWy0u69z2Ip/Zl6nzx732OkRhQ4dIVw+8OqiSnjymAD3muyfjm7Pvy3129glr2C
oDRyjtHA+PtGEtskXpFWgsfd8uKPMaU0v4KbRkudkMlY88RNA5rL/OlQmyWD98J3JZIDnOu7M8WB
fC8pmd6qcC3C0RJOj6ylHRVXTklMMxIvP0HZnALuI0tv0jkJwT/EvJIAseVlqcKOn8/LaVZYVsPG
mVA0A1kGuQW15scTNnK1njWMVYY1rFL1XD64lUetGTnAZipgAP6KSSmpS0AzSzNGnCRXJsa/HazS
AIxhquuV03GaYT0CC6MufmVt2YCAgSlxKezNAjsw69tv/s+vC9JwtRykC4R4UBPhhLCvzdlNO0hD
97Hfc127qGS7WDE1DeoSSj5CFb2keYh/AiwLQmIWtuzO354wa/0hMbz3abU2Uxty/+JKRQ50v52n
KC3Ozzz0MvsorLAkUAUzT+xvq6wc2gxEXnIa+xcgjCS1zN9PqRaSsQTdNrCgoQA5hIKUl6SJcRWv
m4DUAKPN9sLQuu0K0Bw5ZS1NMwAbB0LfMjP/NAW93ZfjutrjIrgbXG/p6Pzjbf4laldNFohh3oky
sB8qwtZUnxMOizPJa/xviKhlxR3/RbPl4qi2oERmRyZ7JlL3k7fSfIwtEhqmJQ1q200uNFp5aPrI
4+RaoWx9GPrxxI3BUR5ZjL0IfqKOZOAjuLuySOb2dWPmoqsEOZmTQ4wlrKGxls8hgjXB/nakM8e/
vauQ5kH4XMmJaVf8nRn1CFxRJG+naaY29wylz+iGlymvwq5Iyrs+AiEsKIxUzqM/Wx+zTpV/XmC3
5dOelGfdiMmAre8MnxZQ1SFc/+v6Hgub/MK6RMbEBrngcUrZPH8zn4dTDtvmydp2phVvkvlaXOZz
uEG2TSDIyGFGv+GzYq7Iyhe2ZKwXVxK5ViDpYeuS1nSe7n/P16U1ytZDYDOdimZPjZG0Dw4H8rc+
lYwskhnQDenJ1hTyI6wOtCWKczURcCnc5vRZycCgsNt97X+ghdfs1nH0jHd86Xnt4rvzEssKgyU6
H/d7YOyZc+VjMbtFCKLMJKrBzImu5KMX4eS+dsvtW6zfzwtlJKF4ti4hhL7fD6OKFGGzgKrKvEYW
WiWejthfMLZ9aydzxNK72GRDNsgj1CNX0LqgPHu/iPOHV1QaswV3TCaYqa60IhgDfvpdaYv168HF
glY7IrUi0cLV5OVM4ebzy2M1vXZPx7brfsA4shxUHU3wDy3M03js/Lo37ncdCqH/5PJ2Du/4yhAQ
9q7tV5DjplRX593Dho7oE/WsDh7IONB7P3LSQnTcZiukVPgeN9iQkeM/MOnoU4SoLwv5gSeo16PT
h0Nt4wP8pfFNLH3LDLEmV6CgARs04pwh1nOTsMJ+4uNTeqePdc2JQfE/d8awmXqa++/HErEHW9/G
Ni58s+CtKLq8IujyUnv253m6531+AL2pXsTB3eST2q/uqmnPhaAgdQZTXLhlMfYeZ5OJ7EY+UazP
vfqXY3dsM+6hwNUCOI+Cf5qNPAizyTsSl9K+Tmn2FPj/4QcoDuJCi/VtrUC5HeDE5fi/4bBoXV12
13I8KFG5dE/BX+nf3Vzc+CKmZvsjEVgdShqUjhQAxPIRm+VMgZZ2ymt1j+S2wA9UUHP6z9ySAonM
5UcxFr8QgqmT1IJYtTJel/0Wdlau0b6k/H40cAvz08YjXbO24okbX1Q9dfXqrsEQ1VGUD1Fgcxf7
OlldS501Oulqk7M0oaQJe5Y4ehg1FOaR5Fqe+Xlxu7A5SnbfA3qPcB0b1VDTHB1bIgySk89RBvQN
KoiBEwSaHWYJN/7F9nO8T1fFHv6eaSVUsxI+ehuxLNhlb+GTZAl/otBGTXwa60Col5FVEVOukCD1
NCyDdaQUSC3LSi/5cBLqKUjJRwMsM6sBkti9tAFsNCFlPQ0iIW9RyvqnEP8N0EU/MpGHkP3ukEe5
buf1RPwb+4Ui6DdkPAo7Ard6fi9+nopwPRLgWJg9/6MNd59EJKRxQOjjh8aBXviPxT30a1H2pEj4
rGDHv2EkUGrFO6PS7l7WsCPlfu/zAREKllNAUN5guuZL7bOHDhRh9cF6n5Pz2gCQr2SW1S1LPhRm
mZBfT0SFuu99gYymVdajvSkLMkNQufIZ4rM6GGeZK1w1NBZS8nIlPegvefqcGoJUoYEfR0IA4iCH
jXP+29GBg2Co4xCU8oDGXbgjCbz3tWL/BeBhtzFBusMdlWQEAMS1MRZVlSPyX09RV9jkZOJ6/chu
MSFEKDgUSinPE9jPOzO0b1gVh55ofdu+hAQQUShoGCqtGhR4b/GsZqayIiRab1TIqIfIPegH16Cr
GeE7GHU5Qt2GFmutmAC9ANC3bPCYRRWlLVjqjHPf+rhHTC1LQAZWjjWP7rwdmd03mXgtLJDiNltI
+PiTaiu8aeESJ7DaoBaKnLVwoySM8od8btoChOhYwSADtK8088O4v40WaPWdBy3FyHbGWWiJA708
CNdNZgCCCmIfcciWsQ2UpXOw27FeSQBzRMdP0OY3EEJ5HGoUiUeg2WU+A/zmclUSYsc7xcnn0vjs
7zzY40g/V2905HSjZJHHkgwofYB/jcZqXVwF5o30SIu9B4eP3U/zD9k5YcHWxMrR7flDsSE06Gsl
rHKPu1E6wrH092Y9hag/dc2g/aJkMUSzXvgL+WIAaQzYTp14jCrLmbPHZ1yYRXw+ohpty2r4BNWk
oFyYWEuOHigc/KfazuBOKHHTWUeLDgBmixVFOOwwfoEFdqpLEKzeGVHsTP0JAt16XEVZXMCrNUKc
myfcDfFWMLB3jUFIdXGTygKMwZOejAbwVdDRMjng+1hSskpTDO5njeyOAPG5SiFwBKZITvMbsxhI
ydVb25yUK/MUAOYJnRGkaOVAl+jkDDg6CKaH4K3O5J+tI3jr+RvefFMfT4PWOHJu7nwJuqcWYold
KF+qcDsHxe2ETQmden6wrAo9iG38y5i9z3PnL5Pw3vHVmfgCYqlJdUeixbyh9gVCSw7wb5UbeG37
/kYxzkiDKvcqRiRz80AxsEXMemARb0MIQ8Ys6v6qXk0ft+AowhswRUuBumll9NG25K0nzFI+w39E
ZpTTJiqh+8YrJmORXAzXLAlQtDP4heHljp0Oh7uvBpPLEcKgQ+K3DLsAndYlzHI1LtzEdcMuPTZu
qSUXhhYvsk34CKvZXo4ZPE9XDE+bdpwI+q9RU3xDr7TwKkq664X4Hs8QH0iHOVqch8/nKztjhwOL
yGj8mUDWkBMfOzMngzyDt4X+aKnM8zTJKUpR4Wcv6NUqoLQw0Xf0/yJtcjS+7Q30/9qMMWxMxydG
cua4xpobaojuR/5OzPVLwxzuQMYFSjyv279aANYvwYb9fKih7RDNIC3X/Gg3j+1y+jUkS164b6L4
OuYL8Qq6l9S7wVuBSMmzLaO0FCyb8nWUAYpobVVW3vHg17KXVVSGdn8tN2Oh+8lDhgZcbtEbvdrI
ZU1YZu83hQYugy+dPDM4yaGDxtgHE93yEG26pmJXSNnHPOru/NsGspVoTWBii0KmQm+twZmc+lbg
7oBfpZnm5Xx7xTkbV+UF3XGLf1ZzR8YbfkUzYurpLBbtAzr4oem783yY4VvZEoFwDSXSLQMyrGY6
Ov2NqJmREn3E9MvssQDFZn4NBN8SqMNFDBIapk2OViw1y798ETHkWzwL9hzQnpZ65lWYQVSMTheO
RufWn8G1c4/lq8S44YA17oie8TvnSRFKmDR15Yaniyw8WqNEtHQ+PhpKtdq7hrXgZFeZX+fV8an8
Qh7h3RPdqjk449EMA4DQhx4G44+K86cCEdmw5+R2LZ+etGpkwhBoxvosbPaQp3aZm+1W9i1QYO9V
9d7plTZeRjuYLvo+7+oJWG1WYuZsmoec7CzMHiWd6L+Ok9VyIdkcBz6mteqA96t4s7tj3B/PBA0S
GPvr/39FddYysOPLgqKCMAI6jD0d6jhZ7qBQ0JQTovaFfUtmGDvI3movGbv7WfqDKku/TlVW2RZG
HQcCdB6rcE7r4zpvjv8GPyqucjsemW9eQ5uBG7X+KsXah02ipOY0i3vBvyFhsc8GFvceTVhfNgbf
cbzMtTqqHWxLfA2jxmuRCnZqOq7gHe1s2QJcMnyoMBlR+bHXsBRHqvkvoyKfLO4nGkAJPV6u/qih
uRJvf+z2k4+Jbfiddck75fIe9yIJ6ZU9Ws6ZCgc/xq0AZTKjeZopBLiagXz0SRjd2pAfWagFCG10
rjUvpUo/jUKoWuHAn17Iea9wZF9YffnXuEfUVKkJDSkG7gsoPB48ysrOSRW7m4w2bya8Fn25bsNq
8N0sX91RljscE76XvDnftkJV+txz6fJ/3RjU1mzn+46nSx6XOOsKiKYul9uolrGiCzAVIGuDSwyX
cDsNgc4LXAqZohIiBE1kIYKRLdf3TNwPMRWjBelAo8uYKAjHxFW1PaSd5T1QjXuQ1keBd9iXA26D
WoHjsr+z7QbBY8UljzYTB3w5iDESrN5VspR5bVoBKiHdlYmwwA1d7YlLD63+ivgc/7yxok5VUd6m
X3797xA/bekcXneWoh2QE0noZP5hsfMKxt5EfSZZzZEhViFpMhIRYPC7iPrEg3tnJR+Fxxe690AA
fSP6RYDYXu9hxXhXwbGXJg/2/nJrWlIi9o0CIm/ZimURh8EUWgEB3kB1QqUW1cjiEIghJIKwPdHL
e88DA9uLbq1nSoX2KLlIbjkhOxx2wqF0apSnA97CPH0mB7Qfok9gIm2wDLSFk5CsO2FZN49nEAVc
JEMKxRAV+LR6mgEuVm+jaNxCzftxKzeLXv/z2HFPHMo/73f8M9IYJ6VpKVOHkUKYNh/jaCf0nML/
M9xf8gx0fk3WZ+CpyACUrdYF7cUs8GUfJBKpVLmBs+7S1A5xqvnLkNSMADjvCDReOURQ6CykQDrI
9pSmkbzojfdYODhj2257O15RpdT4SY2O0Nu4EDqkqFaWJgaRymzFx+xOATl/M8algdfzRZzVGWL+
QhhpAdkM4Vc6JbwCxQmHcAOK7+DHabHU63e9+uDf5teAvC0lnFKC5ArscbrDEDUSky6my7ujfDcP
H549SVtkj7/PDj1VEw1vF6kSkUw06/mYABQmO/+43UghCUqhmwOfwhUrXB8SfGnHHdrTxe3RjCc3
g7ZQSVKWOtyPYDNZZM2mVX3to8YTWH1YEmzgCXXR1/GjSbDhmWSG1ysENAMoxRzt7n/Jj4Lu6+MX
dngQzTrOzFPz+fhStLjB6FQd9QksN/XnVJ8pZIDnbu6rEThZQOnzynW6Ou32mJ408A2WAWEd81mh
QdEkanTSGLQavEE5UHSvieDnbNCayzFwsghw40DmDxZ0hSQLsEBm61wKnGmbk15lITxnn0kfRPVz
7afoE+XEfs1o7HSqNXhiaYsrO+pmo5lVZd0W/+0/A6Lbh0psBpnS/GH98SHRufcI07punBmwkogQ
LlwfCNXBtrItjb7prWypiXjDutBmNAO1zLO8agFwVxWLQSxBy/Y6p7s1Iz2mUVbjwxX67P5sL9/F
TQcJW6IXnoa9iDLc4AikpBnodPZ4VgHP3osa/lMoAXIwt9rCnVUtnFY/uQME5ul6RWRx7bQSRLYA
BVb48KQS2SVQ9v0H3lM9q9QgjKjdt3MlPCLNcUtuRdrByHuZM7X6xOYpQAvIB6nZeqShrLM8aGt0
/r/aybdKxI3Sh476cRQwEqmhAgJRVSyufeYxDQVz1plqSDGCTaeM81WzD7SPXTkUCqZAO/IoJYEU
R3NLjVzZvNKIxpF09oMZgO0wH0feqmDcECjsBFwaEUfJkmGR4bcUviNMIQAiEohSdv7tUN/a4nad
YY5UE3Op3jBdNb3KAcqB72h2TklhgYRtB7otyxHxgeD+Ai/L94mN1HACHTXX7QkbkKR585WIq5Ck
xW0rbrThSor/bUemNuRPmZ+j57vj0N+Dl6xivgB+OgJZbk26/fSxDvlRYwDlsauQZYG/UCx/nzio
3au/yq3bXHmnZIJJVflXcMLXdtQrIftPlZ6mOjhmCIZvF8YK5JIgz7qsiQkYmUHNl9TNxQSNL8fQ
QtuiD2jl3HJfWmp/iNeg522ANGwPwT4WN5ArDCL2aLBKIew3qSaUZUfjUMQd1pq4wtXXxBnop4rI
RB5r3o2oXUrQJcU7hZIWlXHsSJQkk2clplpYU2hWLBqO9W82nwKSY7AVOknb+P/2I5C9sruB6nLZ
k1o2ti56e7L/kvjoRdA+xlmJ68Nwera/UY6DnLimEkpsGD2Hi5prNZNv2qQibxVzrJwkWNT7kcvw
vYJlz+yrj0MYXoTkbALtrXSSsU5+DSprVqP6KqYQyeeo4ogc0/Wg+l7vzeuh8vfDhZapsVOcYciA
hznqm+x6QvQ64/3FwsMHGwMKH7AahBzmoV193tgjMHPAJMWAZe2LgqPaJg4MIhiYFDt+PCrEnDxq
MMrs32TbwTaKE7lEzGDA8fxR3pSG2PU3dKaYSho2DUeTtpYixD8v0VFN6lwiSux5akZlxGwLslqD
FeDIU2JHpnKZd2+U/G6NGJoUhcyyu0ymSxt7iCbKU6P4rX167mMJCRit553+1kZeF/AhSRNxKWiQ
p0azJHkyhDdQmR7syy97wv4xqMvVEEQ+U8OFH/86j7Ak98e5bacltfmHLnavC1wU8fy8cGrFX1zZ
xaBYeMj68Dgyxq7hwBiXR56O6hbl2Y4JwxUAhf+5f03nq3kvu0Y4BoLomb32rMZzyAOmgyY1TZak
3au60iy1khShOGZPOqORFDhtPLZvQo6EdU8Oi74DFYCdPwa9Sj0M227UBWdExMnlOmpSMHk1Xjrx
yUhbax8u6+dCDKOv7/LvjXY8kxRwQomHP2pOYQz6MnsppUUS+Cy71gka8h6JahjzlDhEePlygUx6
g6ArxEWc0fJ+ZeNW3ohxaQyjrwkWOV860SLiUYmx/pDHXDkOrMqk6KOvPNhxUs7PRMClXoJls2BL
b+Nm3lIYDUtP/WpQ1jAHnRJ0juYK7lqyrMl99hy3gzoKOEPMHCzzuKANcrELgvgYSU5uh+0Vofxn
FewxSbBwljraeFc/3nMJjCWlQJZzBVcoHSgVeoIHiaxOixEtJn1fzfRRohAZz3zHC61Pbrht7zhA
xgxusPMa6NWNoVSWSgFtJiDbVQulCqnoXzeCmnmkbObbGqWxKBz+s4v1DKRNoolpFn7h1PaQTMm/
m//9CYEVvEPQEYLP0fqyipSZtIPl/9gyCd8jvUakBl5eLDBNhZr6sy7rfPKMyOMRt8VnPl/TPaYx
eqJtZsxzuMiVMXrkfTYGo+HOswtEBFd0WJaxn4ju5R2YtuaLP34ToKfRX+BkZzEzH1aTcqzQR3mY
Uu4G9m5veKWyHwHYgf99+Jg9Y9u73hX2ssPeykEtWkdVRw0ikNJbO5JOGeP66cfOFwXMAT77NOee
sLOX9IF4QasIDONcdOwiZ6ka613ZRUcnpdIJLpJy2tE019poIlWVeyipQjbtO75V3RxbzvsgTYTF
2dZaKkvDBEHgX4OvRk7FGnArP9mJpkppp0Y+2V1MpjUqhgNpnSdJ70D6JU3PcQND/VX9UJC6jiDb
6cD8PlKILhdYIXkprrEoifRZ8mF35Gxlmr4mZeh8uKPmnvOLMIfKYy8F/TRjGuDhznmqgAbCmizz
raXuRVKznqEL4nN7PUQ2uMUF9IAPwy0A2LwnvSTIkd9xMTdUtHLttsJc0V3F4wWMd8hcECGZfupI
st46x6urUVb2dPQleeBOKxuHTUysTtnocQ0Vu3rjXglJnfpVHKmqHKd4BhbYn35fO6RpxY+/JM3Z
G+CCyFySd71yUzcEQzheFOjL7PB1yc9GgFJkM+8o4XX0VShqJKLDyx7zw/9DYoMylPYcOCDxsdWK
KDbNcnn1WJocx4Nc0H/wnSi3ksyksfqRrOT6SZeD6D6164vhYr16AlrEOUr+ptilmbc3WxzG3m7G
pZ2awar2S9PFWjZnepmA3i+Ld3STj326pmoCAh0FQV/pYpeJFCdoV9AtSLSsgXMnwN3C5jMrE2O8
0IK3teqw/wwCUcLwJrKrCyb0xl7plVi83bla9Qip3TwlSemp36PqsjG7ZQ9H2gOeIPigOt2mWQk6
w9yVZhT+6ZeM2NhzievvtWQVL1IPQx5lcq87Ny2CE2QACrkJQurHs5TPk+ViKgqutxEeSkBEQcWF
fhw0VRVWPHnGZx0VTfn3DG22uFsCG4ISH1+g3ccGDQNCWiwik1cZW+vH9ob/AHC+jGpijjv9kOCN
Mg4E+Z6rbGFBwJoiMXdb4AFpIsAt7M9M7gvIrEniAdMGJnTMYVG5XvNgCa0pWF0FOsDnSBaJ5ljQ
Jnb/uI9gbKH1Uw8l6WXrZEekE6glaOXkr+QnNQ/9Y7D/xmzASldeb0qDxVGMO6Re03heeOAQT+3k
MsCULOyidO+rXf7Shdf5Y4RNC7ZFpYDUG9hbRAKx/obb10cJkVT1Eae5bOZjTQ5f0X8j6V6sFhPi
faTaZUbYh8qUtLVVoy/0VGIihw+9eIypgKpmU2KjGxQhkEqR9vNrC5ApjjS3WFIgN3gxbvtPfKPp
wfZFuw7ZGL/miCqMAcGibnfbIN2zmZuv4UPaT5mjP3srCIJ65zdO+zPPiSiAum1sEmUE2XimYvmf
TgGTT784Dz+ll1j6HFyygddnmP/IIhKZ7mNmZlA0P58f7lMWDWD1T46/E48YzQIP3tVwIfGPp6NN
LbB6Vqua0DwAG4hQ7CiAk9gp5KAany+blvOyH+rDkePojTkYAK6ugKcTAeVVcezj0M2k+rkxnmOF
2yEFQYE9aAwdzc+A6vMfb5eaSs1O3D0dg0DR+7NDOIoh+fX/kB9mDlOVc9tol36qCyVSANqNle18
zljJ44AJZkC9Q1lo3KchgY8eZX7HxoMMGrAGRXD7Oxs6qJ/B8xRMRIYn71OZVo3zcj6lH/jV9QJS
EBIWaa8h963ZMQ5WqCXnqfZaShOxWHcL2Lt39Y8WTwsFvoy+PxBn5vsXyQ6BV0SJb5rW4FPcQgzH
9wszZo64VrY+WmaJTw+w+VdJd/hoYeePia1TaUul/aeayK/yVje8ww1jrb6AWz8tu5z9/V7vpk51
mMznCKc/R0wYkqb06s3MwKn0cgko6K8Zs/qs3tSiaAJY3dbvieiK09TchN5hHfYT1ImAoluqHFqY
dG8hrEbRTJa6A5++PvEjgWRJOqQXxwIqrQWFgm4OStKTMSXW/A3IxpRuuwqzqZCowUeOIylQxb9c
uIwiJT63Df13FfsQZuWSdi4e36VEjRN9tN9PS8r/3B5IDuGqqt3tek+BoIR+eGNddlf7ho1X1ShF
oNU2B8VUrZJrXp24udzLXH6JJly+HSBeNux7m2lxJrEsVGZi3Lp8Hu0WedkcFKEArDsgyYgDknV2
WXb24dRXdASVg2cdiHDt+1dkJIqHwxPfLw4/F+NZ8btsmoVcdLn8pcb9hfwb70ugMeVH2GaxCrq/
qah7NheC2+67SlEzW7b5P+IlD4sRWJzGHGjTZ90yfHnRxFOmsTTqQX/xva7p30Src9NRJ4UjAGEN
TE8vIc9W1/y4gJ/q4+GT8aB/L5LHok3hslKlQRxk0A8L5JH1bIAZHwUF30BlvDkMng7W5A72kSM9
rtQLUXPS4012fxd+3SbDkSG0NqKpEwicPUoCc03kbQImxOZsbHBceOTe6NMZoX666JVMtAdnWXpo
u21SiimW1S8QazNaX9za5qwQFbqMM9xw55k4mL9pvnWXfXpwMq4feM6W8QkOpq95V2EOLWY+hBUr
GiyB+26vaCa+uGhliJSKLR1Mibv/aIIrnXj2tmsjjl9DG/y2OEjguMS3aJeUdZjx95M5emZUBAgW
XQWAptocxmKOYhGIvqRxKXk8Ke1hXV7GvAqoSTrgJPDKqn47MgfkLdAn/mGVEDu4qnMzJiPNWa90
rQobZIFYRs0GfAUPWNRDw7BDDn13g+kC/ehnYl3AwrdsJWa3oxz7WU3wOXHFEu3Op5CnI7lKB5J4
njMf/ysTsxd9xnyWmHSBWrTbkxjPVVBIG0g2F4O5Wo3Iav0GGG9ha8azw8p+xmcrs3SW22tcW4A3
1RDVZqBtGfXJoqzySOgvtftzmyH0JykOxnosXbQwfeplLdF/6MYV4m/FspJK6HYmz32FEd6s3MLn
5CVdgCjs9arqqa5DHZW7m2/nvcX3224L69+fhDnFdxaPH4Wv/bzzwxGKL7zNB0XDgVGSVokKm8KC
EeEgLD8J3GoJH0YvkQIq29OAD5ba+Q9lU1t0516Tkm6hy7owTXHVThOEHugNlBWL6ZOq02LMVCKl
dFCwzbdN0whFTP6XIlaeAfs2qxPCFGP0xNCBXkhBpWszmN0k6NHBa/68uLgy2DOJPzRL9BrZIKl/
F74zlzYGvnLNLXjhnKPn5ps6h8jAHT4MGX/oL5fFG6LiW1KEoXxW9eZc4PyKDvr7P5Gx3G6U6XhQ
F74yQqokbXK4huPx5/KdL342fl6l5RpmWz5KtdDJ8c+MvVyMqCWcVfoQyYtTw+bNzJIt6F62iIvz
eUJJg86fZsc75OwcLx8hkjft+kOIdx5WsnDZrAYmeI+YSLIKfFtewI9WfGc4daZZIN96xFgzRXSS
aMtF7wuDZpxe8/rRYfZTfWYojlES6h68OCkAmUMWIWF6YAXVj6DGn7pqzKI549jd5irp2gq6hk4h
A0C6QjPERM5E2SiZAVV/pPClA26gpKdYmohcU+a3XoPnK4ERfd5mCAMZkZaiA2aNzcQyMvpBkNlC
L2jXW2R+YlM8X79CUuD6E0FuWSqhQz+L1Ws2goG6Q8yt4gOCscInA0OKcDSCJPOKo3G29x03Rp1+
gVTMjFughLRIRruAUUXOP5XADDoOZwiUvHw3jEfBKeZKcu9M9M6FhQHtgNanabRgstL/dBBjrL7J
1iskLEmYz5mkt+p1H4av4NMErj236905TNGUQbjS2ziIEmtUvSIWmAT/oTi5r3C0ZiEJqCeiJ1k1
wAmDqZ67QNvp+tw2wOW4D3HyFB3/hchIJKtUGr4w4EKHz85DiVSGEmboibifap91I+qXexnd16iM
jtulAW+S3TLYIIXoIDXsWnA7r6sJtjuN3BURYso0EW8PvvRY0P5gGTfXU1WRyuK2my8syJosW/EH
dt+Sy1bbJw9HJ9mRKJst9TV5udBpnSnxO2ptyPujYpJEJUYxhRRsBD4OmxdS7SFZ5GxpesaiyXbn
sADXGMmdnMHMiNnoXXo3Z1VkKyi6VUjwk6/SBJqCXqqX2ytfIt6DoTabd4SjTZes9dBmdoyjih/t
tGcUF0dHI9SozrbeZQTfvUzm7oy9xd6tGm8dT2wm2o7PHLGbjEwGtrl4+NWLJxp6eKNrtsrvn6DH
qekAmJOZTCApTPp8ovs5N/6s9pf4nfsqVfbnP6W/RI7f5DQmS4CWuMv7ZD+Fjnr/4uNaPDulhxqb
r0qQD/NQwo8Tv91/Kt4Jk1zA4aeoVFGj07EFujgpEQriFMjd96J5dbshslcZ+Q3GGOqxfk+vLK3H
4qBY7AyzhR/D1BHU5vqqPCt7Z3YOcaXJMENwxdbntvu6IYhXxu9pPUf3zQ1NnTp128nNZsOcOzML
1vFqMEczjceEjA5E2T4FRGyPv6qVvru3Mng4dIdLxQW3CEolzFR1L7gYvdw8+dSMjNyuX72l9nJp
kvxwc5Ty7Fezf+vmrdDCQb/sRhN670W8ff1zCjuyD8HLghbXc8oL/ROhAhYzv931Bj2CANWSJOEr
S+GnT62VsABrjw9vHVjBh9DawbHGqV/5DZfkFdTDv0Fz7wXDqsurZSBWiR9YmaoX9JXQ6zC3VtUH
ItaquyaNUUepDYEPrpmak3TbmTLKtFoKxhA8u2TkuIlBeovMSnE7Fj/Cj72BXmtp1ttf3KbmU/U/
ZzeBU/iY4lRCuuy3pnk4hXqfz40P3zxo6qsSz8rhJfbD3Vabj1cv4VNa/q3CromhUIio6P+hGiKx
Lx3ZaiV4FOvBxSwoT/yCK9n1qtUrSsK7q7ZmBXYS4pHFx2VmogJ8oX8ela3dprfpxsAIOeXG93q4
xsuJ/EqHMSR6rl1Bs5P6pTanMKbO4zblTOQETQVg8WJrD/s8PBRNYMqKNaMZt9CMFL+Rqo0ljf9V
0nytT14u6hfvcI6T5wIbimQnekHY5vZHIDESgrQm5OoFKnmaoiHjOo7Kt55uVIF3ew/hoHVNd3TK
cLSRP1nvE17go+rbZK2sNWtQxQsV+nDqE2Nbu9mH7BJn9CVffTi7f87h4AZ/P08E6BEhe4poHafv
70NGsPtzRkL8Fq8HDlQQj3p3Xt5diW93PgDQe2NgIlLm+IC0+A14QsGIaKCt19Gx5Q/JfaJjUw0h
xaP3+RJD2JE0syTcj5Wr4mJqoLCbgQPEEaOVWQ5jcwzQbvS8Rs7IAivLGvvMklyb10+9uFYpsXLh
LOYjfG5iy85EPPvIeIEU3PXXBva9Q6k7btT94cJ/JXOfCiiIP8dlvjZajNjq5bIv4hEkljM0NlgC
cyp7dhYVAx2zfHTiSEZy20TCp4kNuvkETXPTM9ZeYlJdtEp/5YuWykSekbHcaXYoy42JxK8Oo6tI
kYWx55e4jD+Q1Ejtu0hEoYl/8dyS7ze5E0hROq17Iol6nPGIChJmsHpxELh6HKYz5GZS49C96tXu
0Dp2yRjwnMKTBy82R/M8kTAw3bFLKjCPHoq7NNwk9AcbdH1DKA/9cPTMxuzli0qNOhDIqUIsP1w5
BM6jyk9XMfi0xoOjeEpDvzag8X0fi8KeUVhsEJ9bJcqSvBeeoS+pLNJuLewFhqrcb63/dBYMfH2F
PhT1Ry5E5chPQHA0VurjnzIcAh3jnDKiK01gmAONeQTN0pfJdyyW8x3t/jV5DoChCzVTizwfz6tT
Qt+XD/0Y1CpzmXO5BPIdE1D9SHXugsqt/v7E4oIvcW7F/dzTiKcuBkCnX6ZTTMXkBZEqmxmep8mU
+5oGvBvab9ZaJOKSmllGo5qwO0phDqQdt/9vm0VVeFZZ1uHzAwzxjh6Ps2gVFnyF1UkNU4Zb5hbf
HFbO144BoaZHh2+Wqo/CIXy4v42d6WAszJ3Nn8QtjfiFE+QqFfAL0KvxeMdZNPRkMKv2MBbiwbUu
o3ku6LsiduXx14QgLFwMeD1UVUSHUHNfHmpUy4SatcVDe+tdxHnAFB7knKLJx5S+juSUtBEOj6To
WXONL3BbjEYAdXfyO+KLn8EcCi3tD2y4uyAwG2hTEVaca7rvuB9sRRnAVSFw2Joa0XdbpvTtqjJS
q4FTGPHdKTbvNjKb09Zg0j5PbnpKQupS1aQOdPa5kAnfd3WGahSgNmqapqu0zRGpZfBKdIh29c0X
7yv3Qw4BgXJxdptqkkZYBaJi9s+CPg/1t7bZ0SIqz88aDvLNyFFvqsrdggbmN/+xOfKZZbcws/j0
vgx9Tc+yQY/il4dHNHLWT6M/VWn6qHN6nuQnFDOUKiTUs/OqRCeMYnTIuGMK9uOBqiO7LmLArxlr
wOFwfmXZU2Or2OX1b66G63e9pQTD2cng7a/SWHEpqhFtd+y57FEqWkGzfrSmk+1fpFjsK+8bEYHh
lM5pYgEgOOhd7dvmgs+YVuANcnB5/BNDM5x7nddmGO8nxJyNoCBIv+fc5HM7Xhh95qR86ryU/4jP
mtcKPuTbYzs1bKOKbWVZYaXFaKGyD8bFPRof8Y7hpQxEathTuP58Egme7LhrCAJtwoUSCQz7u2Qs
VYIzwsAsEl8fONPxdUcxbnrvk/fQvSniyEwDFeb02LP+fQiG48ykM4qTPbB1pLZjsiiEPGbiza/m
A0qlp8/6hfG4vzoIX1zxkt4+Ym2q2Cmw1i3Ro7xFo2LAPBLw0fwxkGL+4VoQ75pUxjfzjPD80ngY
k2dohhgQ7D8ogr+dsnKvbEz/+AB8eP4LEXbBPi0jn8Tb8pPTlqdq5W4bWS/qeQAIEaWiKexFA8Rk
aOy25nOF34ojQcIZWflZXvEG/SNvrk5x1vSCptPpiMzXDQ1S9ryhdfX3OXWmM1QNuy6nzfghC1xV
HsUZQNtYdPXbrhlj0pe1BWpZ2d4FZx/LrGBp7QCKck5flluPe9+JLKfIcx3FBFjwJyfSBUZRM7w1
Yt+jcEk+TOq2pGJ5osNzcRFIwuycrpg7GtR7bO2pbO3RqbOg0hTcU9EXcq1QO/qU7O4aXqLN3UGX
NeM8CCeVhUonQYYEK0cu42lKpgDbYXrI+FKIpuVtkuZKodAJ9JRlI680DXT+7quAw1ODC9rp7Jgn
9kpj8Wo4Wwre9GjAzfTmxhg/zcfhAEmyfsXuUOoFrsOotaYSr7JU6/QoBOX7nsTYAVakrbMPTujU
cjKz1Tbng5MexnlOwDagc4S0P9IrnNtbqbxowvhx3kiWOhBcjwZJNm7Qg9JwPVy03/NrwP8ZGUQe
SZm+jXO9gKvr9CXgsE+4tqJAVqdSbzbBQwZoDCWU+8H4/AHWmJO5AsNjc6rBW0Eqh9lr1fScSzqy
Nl8axSFydgJO/OZzEbzhaQQ1bCwlpgxgNlcmEPSg+Lljg+nX3Sex6FjLgd9KxLl6v9OYzjQl5pGm
PMRJR0Vjj6/Rwls0W0gcTPyW42uERgTZMRN6TptXSJUkzuPMispST4msJRjhD2i9I/pEd48qVgcU
tVuAglFsnjuxoBb7i7adTuJvPKZ7ALzxTEgDjC1T8HG2Yov90nfFgB3MFyYiu2TrS5a/qgSP6CB0
vnNDQUJ3yzttZE5Iw/a8moyySA7IbcadL584yy9s7CefBI4QLgbJK0Mb3Fo8/vDGsM/N7L1vLjlD
JmP4p7lZ+2L6t3yyL6dqovm/UcT1+Qt8umlGVhEdJV7jqYliLKBhs8YpGwmHtiPxjN3GhDwJ+HOl
7i+co9DKecZtVwJGxZwYkuDoya40gihuVOyEU+M0G10qR1p8rivkv9na4dJZx8IEofZjOZ/xzhLu
HFvQf7abSIB7wMN60+OzFmoIDN9SsABD6EaYB2S1R9wlBlu0RGxl3gX5AeX1wPI73kdjSK8thu0K
a6ZOt3L36cOV4kXZskCquOVZuLmTxeHMw6swaCEBOYbZ921/+nGzX/F1DOAvObfMMUNlOhQ13oCY
7ANey6yQvRfnZKDRCdfKOe2qNxtAPMXxyFgI/lkP+qgTX2W0K2fu6x3zOPLpB21sTc8WNc+iqspm
y5F4K1RA90i1KiHAruhp3GuS6X9sxDyw55hZVOh3+EgWyPIV56v3EAJiHwCCqxe7wLDkwQVin+Yt
bhUgEKs1711KF9RBPdGnAEj9dhEKQoxdHb+uaDTUW8b4O/hyzqf68+Qe7WL9WDjMAwBi9Ty279Ip
l2H/0GFc5nMy57+vN5YST5RdmlJqDNNVpxQqw0x/tB6+WWliSSLl0AwmyMbuk3EXU7yP8Cazs+IN
s+hJ+SVoNckghuKVB/CiA7PZozyfXhhwyPTMk26lf/MoUbNtnMDVvNi6Mj4P2V7Jyy/Huns4OVvK
klMKI4sPZnQFwy3kSucE/ehEkK6PV6VOxllaigunaU+3Tj1DO581do797hxhiA8NkzCgylOOLj9u
jh8mqEwI98TDEbEbgrPC3Jo3Y2yqbwGIpFE12quuS4JDdyuH12btJH7FLbG0i1UW6OUAc2LtkouD
at7KaL5hXz8HYk6RUYSAYpzm/Gi0SkciH5iL/qTaIHUYwDtLwSZ8p1pSTTiuq4qTofu9L8o06bf5
ZMbJi0WH4tnbDtCkrwzIffUice1u3ECQRcCWYbN94upNord7CgkRqWg6o1ZG7wTyOxGp8ur1KjGU
G07AaI8XYTXuEUd/7zGlv6YSs/SK+aB4m2rtySxFHJinDtSlqLAxfapgznjAqrEejMm7MAQZOYU/
tUwrrlZBuhp1Q+3zL6m8bPYX9XqrdK94ZjMvfkWWMp6A8iHavg/s4qXwayu83/wTcQw+EX/uhyXN
UIncJxp5QbUelP27dmNWBJyjOEI8WD6+KhTy/wl90gfTtm+WeKwkWzUvTpyExh6Oe5LfiByMHe+f
jeO8uCsMi8pkMS43pB88I7vvojig2WoNiSipJym+8ikctiiGQdxkUYe9dl1tLC5vCqvY5QIyMe1O
t9NrDqi01GpXRUoO6RQBXUsQMMyocILRZvKmo1+vAcFOU1qfrINL5+MjgeT8LAq23MzjqhlwqnlB
kkKk3fho20HA5D0n24p88JYANMpbuPAQG4Av7sSflXS7o1F6X9e+Az3ZSXUUHbi//jEq7rcpJ9D6
7ybMMKyqiejVzWCcSFYpGsPxr4Sj5Dmb7zChbAiy3VPX4OIyNqtq9Gy7KDcmRjUyPHwLd8Cmhg00
/aFkt/mkIKbr3FtYQYtNYc9+OvNY7zd2+l2OwC7m7K/P65EvCyscnv/GFMEvyIsGUObgJ2dyynlq
rM2mijiCNdxkhSxKI9Aw9+f5+smbV7ctx7j0XKNu80aTe4N16gCfzUHnORrU99IA5k+3cU9nSjAN
cF7naPnNZEM35rHXvBCNO3nU7cdbhp3Mos1J1feEQCXXVMruUMtRuiYpLhHUopKI3gwHrej2oGfY
k+h4Ti9r4GKkxgpk5APIhAcusxz1y4X1G9QelESaf7kNoKpBl4wDT6eXVGNWRK8zDdq6dWDTOztp
HcEv8KT+fHXbCOxI9Dgc++/ZuswcOhGZlw/Vles71JVX/FdAOBSPpzAfDlJmSzGRW++wU3Xa6CLR
bT3G+qhLpEkE0zgpWh1P73yUrRMd/nvYVjmG2QWj0ectpnBRUJo6vcKGLl/eQmDNANbCcCyv5Wz1
ZYGqBBTn4FsYepa/wEdQ0XMY1x/LXa/Pa0w0ysclMl4GL7JD9mGSYfZWSsQX5mQskKpgO1wKW5Jd
TSld4vnpNGbuBOwphh+7KLm7wEE1PsSi+ngoakxpfpYKhS5Dv1+RyDVZEWJ/JGcQ3PTHfvB+Plpb
ICvsaIj4nypRTcu+zrBpFs5fPtbvQyFjP+0FC349Q0zDfiMZZeSkS8I+pjuXgv8PlkZb1WHNIMuS
u/TEYggZTJ+IukICKeJYXxLaHVEDd8M2hN1nVa5Laq+X8xu0XO/Mj0lhU0mdLk+SU4LsVrFFlOuX
YIu3QcwXefHPYLkwAS+HnmxtyWokALT70PRvvo4qOWEjJ3dyWvkrKW8Ll7zZJ73Ho3wxxeiCMX+E
YSwd3G2qRV2MpB3GnaCnnrwcId2d7rxoXzmfx7+Xem8G5RPS39b7iBlwJ/LqyDg6p2A5E6B52hLT
aGQioRNpcr3XuIWTB3q+GOfxdI6YCztOUI2EmbkDV8jDKU4D87EISWukX8CQg+smuPyukgu17QuZ
uiu0EG3Jvh/s8GcmL7kgQj7ecboV7kNXLo2KIaTJTtWtqWf4qAAqFR+BezleWBBO2VmNFhpgIfxX
A5ErmjLmfROLZm7g/n1KptFqdcMVOP4VaYLCG7KWq1lP0GJ4bYmjiKxmw6FEXEks4PmcW0dfqo5A
7WlK7OgJf+7qJNmNoXcqkfr68kZs4U9asfOmjn84lO0XdwwjKxwVNS5o1Jpdt9OQq4sqP/uVRWJl
voC/jfvAZseqcWZ62/zU6BMLGXmgYMFXaEVJjYVc/Ky5ofcantDTdtVBUJbSvZo/Feu1CbVQ6EVK
U0bgWs5JlElFxQg168x0Jcif7++tE6x3urHHL/vzZQNk10GE0uOCP4Wi1DZcNFUxzzLDcx9Zkj4I
7F1WjyL2RU+EFYVzL1argLbYkb1focD/5pQsYPSDSAIQmTshXYRdubs1HZeJTs0EMzlYc7wIvqwc
W4LgQtgcKCVx1Zxee0QWjz43IGZPhNZ+JQYSvxgm9ovsgt4yz94+JgZLCaBHNjW1jT+++QD/CoEo
t0Jzlol+vwZg8TfJjQbe+V1GMfQd5Okv5wBOxTAdLh4zHIi9CKBfwt76zAVOUoab05uAWU+yPGms
2MX3GgM4mwToSsqb/XmAQ8jv7de3h59r7GB3pimwXglyFz+j9YR84+cyHrcFDLkxPMZ7oHfTC1xe
0XWvWjfY3Z80zmOebZpjDpG5cjp9kyEK8ukHmNjDuXow5MLR2FMHNH4SzzxXHgxelOZg9u3EKk5i
1Nw9CcSl3FgcX/tn2Es99lSODrDgHHcJVGJwZoHJUlHm+CYTdWaw8ad7hnZc0C87kwJN5nV29qPA
94UbExGvd8m6W46lFbgeu3yWwQfxwgf0uKnL5P3Y0kpXWM5M3jQnStB1jtN+7Ymcp9MKZh2yi/ag
lRuWw8c2RXR1VVJuhastN/pJpjyABIqekNT3KXKZ/KOGj/R20fxMMBIh0d4rvPAulZLYlrm6izi1
nrmfTJyTeOusT/LyNs2qktQKfa8Hcm9+40lw/FRdN21tH3hNJ+5tPhSEM4u3ZDKig4DQVqczn1Tb
IPu6jSRNod4MP6N4X8u448FuwSZuUX5pFf9Ixy4LhmVT6zz4t/Tes6OsPfnl5LkuGort9SqMU6YF
YmEGZQtj1QHc6PIWmW1R33vjfYLOisQhuhlY2pHtk8uEtZbbwpeqO+lm87Gn0WnjWE2QFJ2kj34F
LYAYBqGvwCaFnULyiWL+J1uyAUD1VVjuQ8UqSK6nr6xlqLInRGnss1nwng5ISvLPxwGFwVHRRD5N
9NJ0xHd9JNMAvKl3IIJy/n8t8l8s/m4a/LAzU6pQC7L5kuAGf0ymPGi1c75BalmtIwr5TRnAV1Mi
U5olLZmEDuHJ+4khWVZO+zxzdBuTL5QmwTo+QU2Z2UmiSzJUPeg3cwAruMA0655Lk+qJnYzTbuPY
uzWxGLBrVZ+21DN7qgxCi3H8G0ZJlcfbL3JWUoLlZMRe+iRUQjJ/arMiLYPVO7joFMhUR36iBWmq
CxZ+ZfKECICpeb8WiUusRJUSAfzbOsfZbGRiuB5s5H22VlI1jpZFeS9nE2T9TsbTgTJXm3pNU/vj
OFra3FbFyaYThBn0KdKFcEj8MvhJowHFXv2LLcXQ4HIDbIMqb6w/FUZPDZRTIbcjTmobHS/boP50
MKn38wSIWkeRxItNVg4N9uwk7C3i+VVEnkOULFmN0+eJWK6i/MgJJG6QKPX0htzqSQ66cJ+j9ycm
ryWHSNheZ8rXRkzK5H5/IqhfWJItkd+gGwZXKzkRt3B0g6gwmt5w8PLgXfON5dIoThAeBtwPm2qC
6XDcViTmI9Gl52fizdtIZlXOGDyhpVHxrggwT/L9TzMFf4iXPIfnU8PUG33LJ2PTiVz7GPogvJFR
MjG5T55afvYMRZZrsTzTa6zpbKryOnoE+bXJHuFBNl7tXQPdrOpKpdhdE9oIVc6TA0gtL6Md/f7m
j3lTqlU/bBJjUZeoiILCe4dag+kQO+4bI4V7q8TKpJKlCnhBpYMZ8qEr4XOQp722lOL1WDajswWi
YPdzA3fmNQiBtseqnych0Q07FASu6OhR6T6ASj7YD6hTLL7ZFN7FFofhXG+UZx/Or3tkzV7ASRB9
mbe5zrA2667Jr4CAm3UC8YOcP8XvmFj/FmGk35LFL+yXUMA8BeDi6RQuZOAqLLFYftIeXVCmEW6H
gjK2Hqg2KrWjl82rVL9vAZ3H+5oxIazYaAqi9w6j46rRioQcxPfVvzqvHWrZprtolASyLLnGMsiR
CHX287h2E07+7PEIare+I+o0ICXf44CQ/IW+zHIUV7aYlvUMOLWN9Zt9PTXoEWe3SQBAKgL2SPig
vsZ+2mT+Bc4PjGHGpxnLuWbnlGVmuUZuKmURdedozjpEawSpHy4fQfvdGKOGsZd0DTAb5YHuZ5Oh
UqtS3BoIccOcK4o4NBOshaHpOoSSFxvWu6ydseAEc3dnbFK4sSTW3XVv9WzVUxpVLHsH2d/wdmGl
KK98C2eFekn75HOkyy3CcDKJ4chieMs5TLA61FcZ8+IecXqUWWvVPByqszY3XEnWPlKTvrsZ8tn9
W/f7JIjQvehR1fhJkifuBX06GPU8V6AAAYnw6FATfpeueBexbC6VViWt42qjBBvq3bPx2488q/gT
dW9O1E6s5ySq6wFlNMP6aFW2zz25U9+R+xoe8fgAX29h4K74PJMD5h3ylXu4YLTmmjMRnmaZkwhx
kfuSKDDCLJVQN60ipL2r9Nf/LERHyAo+eouoU4Dxiz6RT2RguAC8tmmLIevBnkEAvtjZRjUkfqEy
MUhvmm3TRwZgKlUvqKDCvvOMBJ2jRuSJT81NfF8iAUDJpxdBlGHGqsZI2EgDrYFKvaq9obmjkkTq
355FjOze3RQXV700yp9J037cCch8+jrtq7pCssO+T4aJ2NBahqfy+EeefcDgi9ymLweIlFNv1Hh8
g2oc1VCYhkkwEyLny1fXJXlwAvbxl+cPxmzN/E5p6NbCcAcd0J9D37YaDAXDONOhaitx2iBP3u0w
zDiEFHUSxD9uAwIxWe0t76eXWvXQwkpFXC160qja9KRqrDhkf/D60WFg4bMEBLZT7SbJPOEA972F
rJwmyNrsZE+jm275RFReMieX4mLyHeNiYVWbMoygpGvJLHgIWKounyuH8226GLSn+JT6s8s9dHtP
8LBjZNub/zK+sdxdzqn8U9wrRwPoJqZZG2IOaVeWjmBrFx/5wfmdgV5AcFA544jobyS+hILWFBPQ
y1QCdjZRNkOwre3Y8V7PYZJbhUziDxmRSXsx6nCUcljm57ZC/q/6YFwZ6a2UJIlpuSho4sF0JtrD
GEP88JcUQYAZzJpJ0IN9BMTsFGbcodiqIbq6b855WP41Oouru0K45hP9vNix46Iv/8wwWK1lkeJQ
X6tDG4+lFpfrS8R/amUAC6JFhpayyiSLg4wEobJls589OGx1u2khGoEr8ZCxsQx7CziHgTlDJdld
V9/xkvIeWXUTqFGm/n/2DhZfMpuheezepKxaULfLsJyJNA7qLGPiy99zDXibJbrmulC7DmHwFkWR
nRQauUTLl17tq5NK4rmrDR3AbBQbB5hS1Zatn0VTI+38Pcy4dJyddVQCLBg2iOVLjxDmYYryQjiR
kUi+DCH3Ckoosra/qI/oS3srymI793HsDGZdv7qwibg0W/zxBVGFXNwRGd76M/WkhFgV89mJhocv
JIRWLVfGnKWOPV2qcf1n9OzsdQgxbly6gihbCLTa3j1OGI3RWQIUjkgK1GzTt9zr4ZYqfKxgahH5
rb4M1b45dENAavnN4OF7JJVBzqEjOEN1QH428W/Dw7mILPZuVwa/DlJkRIxKSsDPl6bYgLEZjCCD
GXr11j5mB+vmHRnoB2UtNYCkvaq0q0mJFnao8mgT97qtZmwxB5gCcvR81ij2Imj6zwSY0aw14qCl
3uFGN5z0Rcn17/Lga8A3RS+728akC79t8Y4iZue+wYLv9SSpr12vvbP2pS1j65unu36LjgGDbHW7
LnwVxDUsrs3YkUrf5bmMDfgyNR8162jliNSFWZJJpnjoCzBmlsOjXuse5ge4I2N+wOHA5YOGepZG
8HeVbCaOVWfbaWuhJ2LpL+iG1GC6/4/hHl3fEDZoc8D1L7ArbOCWXFPrmEtNsEJy/FgXLL/wiOQV
HcFpQcbILxXyyHOsc3D7O4PzjzWl/9GxrZVZtPS47FKNnHyweX9n911ko/FyL81vjBZfyVEyJRfe
b7qHVmIEdXyZ8Dids3+uK/h266OKIo+ttgOfZ5fJNnAX2N9Fbh+1OifDqHxddXgaNFQfhL6uHVvB
eZujBjKKDp1BtvPq+eVyj6Vx4z53IS/h/n45vYPX4gFb8M+cczTGUc9GWBD/rm/fhLWu6HYGv+BW
ZALvw9MhqAOTTUYpcuqgE88eFf0u6F38DHSnN3rztqMpJIeQzVr6osDGn7SFat8bO8YUXJrf51Gi
NoC4kWnj0JY4VOn9JSafCa1bFBYgrm4823Yn1TP1vz/ShBQePvIR8usMFxFmieJV+49IbzD1KkuC
tzRlfOBacGIpVKI0E1AhRdt7xPoy/BIwpVeXgyM2AhUhjCkYcGNcctmpWAHKNyYXz/3qypyRO9Gw
rmZxyCyVNoC6su5RFaHThTe7IYhRqcZ0ajpJufNqXLeHkf8Clj1IUj90lhJHCGfS+5w+Wd5MVA4J
4zvjKVe5pthxazUyrmYlbb2gBinFtTrbaPwSBghKsUeU1Sr/TBekKxAQukHGYzm9JEh9GMa6ne1L
qQL3suHtsrq/YlElwlMK7M3Yv+TvknWC+rsMPImyyMfa5FERqIXVhmu38f79kSaz5Wzb8YU/Wt8a
Ap53i93hPdWsbHW5JQbHSmfvj4pqtpf74uN7gPh5ZtMxFdlCs96whsSW9GMxRQbia5fVIAKQ1Ao5
g8PPizT056SjxqsmdlWuEQWNKxq2z9ZICXcsLnxLGxGx3rQUj0NTLuzFVtwv0Gl2trQmN23l7HzB
r/Y45NURmnMaJnbIi6si7QW79LbpBV7pFbEAO4i8RQ8khZIjUD4zT9KRQmpT+mOlI2kCxsptqKsf
UOwishZUG/TWG6aoDIzTkxg09jf/764pKoC3ft2WIEQ61E6a8OOEQsBVGQ1uD+hnkHNkXWOaS7Vm
StB5fIuDjJb02SovW6UKgDMjGRLjK6FPVNhVQwFZhp5LRKXkdwdDERJdjRT6G7y+Oj0/yZxLlobd
laTZKmqmWDlcPHzYnQZWp3MN++vM9tUN7MSrPkjwCCZzIyCPJZdrCh8pabPnTvAQj6eFL93vKX1g
rmCPLrHZV+vYn0qCYlWACsUIPsAw7U+pqky0wjgPpIzf9Bp0FxLBGdPYU4w9yuERxZImVb6vtQNL
DI3uWz1FQmjHHNuthtXdUGqtTxhWMiPoRaIqikV8gvZgTaMR5ZSC5YZN1+UUwgdphH37x1bcaYz2
heg++rFkYb+o17HUnwbEyVoQpSW79IB0xxCC4X2V2lS34u44XBN5+bjfcPwu03mhhVlXu5AUtZ/Y
sg+JdFi1SUDqP2o8jkXdlzsPJIw+rm+vAPyeqwwAOO5Tlcg4ApfDqnQoGX3R2l4QOi0TqJDt8AQ4
ox82M5tqr9FOXq8QctAmAlVuxLmTNy2Cq1EdZubCWVMeK5PPo20Zg6KBUYmvLb8c05zJ63U3m0xy
IH3h4FXJaTjFNIInNh4nPttsxby0sThkcnT+6rUKJZghCQXzhbf41HguqgN64KO+VEhnNNo0ZM9C
deLyw8Kql5TBx2muZwLsGEDJ6b5YTmqnvpsn9EqpdA3KwMso4PPzNedO31LbYr+Hs33c7HfYNhTz
MYWv1LE70XFF9qdbCeeG/vXGx8q8mSxSEdO01uChO7FWKfvBrlmNqqvhJVvLsby3okD1gDwxwzHk
IMZ+Ear6BtWr6E6iBS70IiQ3GLaXG403HfyYGi+saZTune45+oQAWgEpZSTE6fH76woLF1bf1zbG
Cn1WRcle9aeyEw0HtnEMrC0j3hKJeDt9P94vp+3eOyjMAwxjhs2H98GId4eeToahjOTuuaihXJa9
AM8D0OnkDSVZX//Pph10qzAziHgEmH5spZzqux9G64dEv8YFIm1r2VBCGap4ny/81oEgBTK/yW2l
78H8GSFFWRpO5KMDU4Unn/8VmnQb4RIN6IIgFDZTpO0bXs7oGLwGxroarzJznYp355QHn9V2LDke
9T8sgTCntt3PqVWzilwgSAeERgqwzqCM/HpX0qhnnjqCu0T2ML+Abg5OYQi02uFUMBiT1tFU8xBZ
19Ofvc8siU2KzZOjhEoRO1OtVRMzqoyFQC5iBuKZR//nvyzHBxGWqQio6akon5Ysorbk44pJolqg
cE1ilZwRKSxgFlKouuXAV+RFdGOgpBPSlU7ovmmux0Dp0weEf18BGwbiNgTDj78OadvvMDqkojck
8bPPDgXuPt6TuzwTcS6UwonNGZxbrsBHkCaIm16fT50L6QdkAAeUVOGRWsEcQ+2G2POqDgFMpdU4
OCep685mfh4dzptxDeGflL9jpF9jqsclK61b8sLk7qn+GDLiUNe3zos7xVw5+w4YBuIt0b65WS6S
NPAp6DVwkaQBw0veJphcUoWjBwGsxRy68iZSZICvSYC5zNCc3ExBLLtb365GjrCYS+M/sfZRzR1n
IJJgpaqpXS1tmVsAVeHeDUF41GtqCJTfCevXx63imavaojX5kMbLHC+I7lZLOVE1FiQkP+3oPvAn
AkL7V/jrUaXiX03P9rR2s41rZDST83ohJncjXCVQl25zXL1ttRmX1y4SqF54eytqT6LZAOV5rYC2
+Ggz1dW6dezFje1u3PhRvqZPcl3OPzMBugjvBQEZqJTv8DYRO2Q3XlHm4N5r/5z1mJ3ouZO+EXmI
T48ay+hluzMG7p3x4LFDGdG9VNnyyskto2jIE7EWdNaTv1XDsVHvwgfZBrhauBmg1CrfuJBLrMde
Rg7AYsxNrx0nsY4iiqLNCH8/3j8MuyNnczU0ER7r1lDOu8/+IVVQjwUbuoC9iJbzPwS8PZkyDj7U
qgz8OFdI8N8uSQNuKis2lD4Thh6N75t9aqWmfyhXHgFwxNxcqeBYQVrc+qV04eVdr3hW8Ru0hJmB
pZWbAMGY7i5uUSL823KB8LRQL2geznLCVjaekyu4HkS0dEdtVAjNFooqtmrBuokZ1wJoH1udex6C
OWypxUguTFdDbjnz49kdF3uNIxjRuBRarLMC4TPZ8roFxp77oAHjBlaJEA0GGxIOkTEQ2NrzNiSF
CKONJilW42vM0bErl92mNZlVbVWnSmB4l5uXMaYqhIVnu5AscXB+b0FhjG+4cK/J6kPRhH0181aK
0UcOzZ3OY8oSwtJtxQHW3E6o5068/OoGe/tf9oce3Aar5H6u+LBIX85JOLCvRa5CQsV75nh8ZFcd
WaUcIZTZj2SeLLRurMnWC+3SswVdxCru+gq00bUTJs2Wwbul5dLMu1fX4cvJgEEc3aHjveT0gGuQ
1X54AX5qQMK9lmfNrmHCpO0fD5kveT7SPkdwTmA+9L4tkZAvSZpRPOeY8h0BVQEWiwexw2qKQBcq
AJnwevxLnUmo3DU4hB/Yidk3ml+EqsIBK9CBKQBqmFyqpcoGDG7mJ/+FvrCZO+H5i/4IBYKQ6rSa
Dt1CnaSj7Re0I39WgznBwe6W+x6l+e78oUx/sqz0rwWZxa7J6WDkKK2ooqce+IwaCtdkKTS7fCeI
V/WY6vkYjJ/oTGGFQnJCQVKU3aP1ZM3IGpd3KDKBg754ZiWSN1azQwgJFX7YG3X8LCeTSwq74sr3
U9mzTKyCxxE35+OT8DFr47TC+shOM7CKQk2sMwRYZSHALqOWKKs7QdJqinB41sAQPDAEd0eUTIeH
E2FZbWofZOoy264TgOqkHwkfF6zllXH3QtsQqTD3xK4V4SfUuiypu4NUg4y+kVWETG8R+eH4ckuf
migtvnCzg59RE9jn5B487WeCTkNRaYdTtRBj3vRPDq3UYyO/8HsTN4PldlUKtCOTFKziN2ku+IuQ
FB5qXbWo/yJ1ATQUfoJLyuPtnc+76tRNHGWK36B04Gs99jggY5HEyLO0dAy08fnScrERmLOpHyKl
QhnGGD2mvCbvy4jC5K2+j/3CLVB16yrb/iYaZXSXzgCVlVUH6kYjJJhKTdRM/qd67vB8jL7Org+i
u/BI5dpVoDsW53F+DXmXR8Ang5FcvW7+1Y+dZ5J62cDKvp/KRflWKYasNSGuiegWzQ/ic0FBm1nB
ZCwrVs6dH5PXIFyZbb0XHIMm7I+NS1N3vPddP97bS+opY86s8O3d0biQTkSR1nhvBq6HSYYn5j+4
cZMoHjsXG3KEMGP10eAL/Fa8ibGK3qjo59DO1DKQPgyu2Bpe1/oPh9fJ0MKnU+y9bXd4jydun59Q
nTyfAk3RznClRxudhCghUKWFaoAZBdcae2h3CN4gBUkUzK9trNQE52RtMB2ZD1cVgAwl5Gkr1Tk3
JUQAKQ2uLcjFaSC754Q0TRKvHQwJ81Nl7gegHv1z9gFUY/rSTs7dGtYHrjmgM+gQeVCsY1RjwAyo
rJg2aBE0P+xyMonLM32GSqIdyrkBryneciOyras2Wyf1vfWUAg+wsXBq9hbDna+P8+0pefO3O/FT
ITprqbfRrypFRF/rlxiJHZvJirSP26ZXMj1VPXWMjgPc/YZGbodcwu9aQjBi9ZbLJ9jpugxiUS+H
+VLq2aokJprytl2hUIwg8cGiLyYfaJEKSkFQVJoM9AW6t71XgiQtIvENhMqFF9Gnf05BxrKhXXEY
kumZCzmNhf6omXqOMnE12RMv8pWZR9sAf6Kfy5M+3KqD6de/nI37lSc2UAdbL5lEHYgemADIcw0d
95LbVWnMkYyluX3JBbcOMuyzLDd+HR4vSjixlRcX97tbvU/YUSrm0DbKmZ/hkWs6WPx+PPSzFlCj
howD3wlnqgXoBexADr4bGkFfT1tQ7hu1vNZ4iuYgKdIbqbbV8K+XfJJeeV230FNfC3iZjCdj5Ed6
A2LldOHEluB8LA1mJmfu8J4kSOc7qG2xTfsEyKnn5wS5XBtq9gEM+RUQ023Re1zzsdfQlrdBe3Ti
9Iu5383KM7Hynp4Jb50xeTUMpqi/JHV8yUPmjFcKrSoofiw9+7jZjxaytW6cCkNDlt15GdmCbxvC
34c73cNkBYINKIRUkx6DJTwHZ5V66iybtBgvuNwoibRoC/e94LcD/Fq9SwwQKjVOrcMoZ3DQMNFa
q4fOV9GdyMghoUimsAJH09wXUjZGeiOAaZE92hIKyygvDUG4UB+Ka0ueJ2kSxYedt/7Ec46QWMvz
yLUIqF8/QBPfkEWkyrj84Ki0dxJxbDxe7DPO8TJamutQto7fgNQUJcUvfXLKakLG9LVqBZmrupNO
KBF1+KrMp72TJ81DI8SovWu94k3ufwL19v0Io/y+LtBpfCd9HRYIShYMrJ4lxOAPXuA1VVZu9DES
Vyuv1HMg2CPJUvUHR0chi5VzyTvARf1saAynZLYE86yeoZYKt/7pN6ep9TZCgjR0tqSmN1u6+buZ
MQMQeJ/nTsPHVRTUuW58M031uD/qAu1CamzkyPk/bf63Rk6adG1vsIHNUHSm1l9kMZPNj04XLZhN
psCskkHg468LMoZiYc7rFbL4MEFFUzS8SiYT/MQD90FC/pYrMIQlThljh+ycTJZyvcCYEKZHHHU6
+LwxNt8xZSiVvMQ04ZEhMc+pejhExgN+Q079bCaK95hyEV/uJv05APWSILn/4BkqdvZ0P5VeahBa
5vmM0Hku5ZQJBv5WlG2FexJtsRHdktaQNW7UflsIcKqwbCTeo1gYLK5AhW6IG/PlZb/2se0tZikU
ZGfwg1xsGWVlSbDGkEP4ZLqvrqFstWEFxiET6XciIlmvSdJGJa2NSa/XrxaHyEEW1AgVtvrDBjUS
SWsjQTOA8bi/OXbAR5gHS13NucvAb/wfMNzq0bgTNmCVBnOvyGG0xfhm5W6/cJh9PWNm4ba39Ang
AwXX6RTuzzt8mvVkSgMEWRxv9MHpQ4f0zdiVxkBIegyN2VDW3UBAIatA+S67IizFcaw7vTtjmt47
dNLw9Un0QXX5kWtTsIv0uIO+hDRN5EVDhY53B+m8hLoP/tPF3uKEw2CtCGndepw05hImR9DRiub0
V7YTsUBlwekvsafDWgdHDufLUECpxGCk1KZUxtCOpuF41yHOXz0Jn4TxU689IKF/fMlyVRKAvXki
DVcE6jG247l4hkAvWaqVO0nBM7PSWvaF4mhZFc1TjfNjCHgDC80FzSD9CtDvNHGnLJyfwj9eDr92
KAdhzMQ/voSezl26R1KMn5MV4rTd2PsRt/au+NY0MrtQ1HUiph9I7VzgNzJWYThAm+9ukM2D7q5y
PrZJnth0PVGmLaBul1mwktkYALWxL4esLbu5c//yKKGf3Aurb2jV4QFihklBfXmfXLcMkkmNaZv7
PRSd8dCOQ6qoJNmcHMoJ8aR/TUZReiuMXZflRgZbnQka4K3QS3uAuKa/ZrmzCT3s86t15JY/LYkL
INzwcXMPafVgyEM64aQMCGBiVbHwtFGVOZ0IUezSUy7ce7Ox53jsfOVfSzSaLD1XsPoEWo7nB4GW
LdS+F5s9Rh1cHReDBt4fFWXeI2hcaak8Q4xtbA4wXUs+g4tu7jBgesn7NbPsX1lHzRpsIyDhYDNF
DOIA1UzYjn/+0XJvbVEL5jaRJbzi0faXOW8VG/GlFKsgIECCCdLgSrW6pbbidQDEyEXgLGTKAZ9J
V5pDXmdufTXEBFBVV9PUPscmVMn9r92+IKqdhWNZlTQVCDZZBn9IZijW9yHrfDNV/PTWEokH4dil
tmmSovp5Xe8XO9ydTISLf+cEexTiyStRImZuy0h4CzBVY06NQiHgMRI4Umr7Q6StPnRDZh1aLJ+H
ArfoiBOXo4kRqYK3N8XpPgSLbRJOM/KfoHg8zvV/urb9gieCH1bnhtkYEP4dlxbYaN6xeRpK136V
MGZLGDYG6RkUZIMxdnzf5IrIHxGLsMSDytJqS/8/Nx3jnGp2H3GZNrbU0TJw+GeXnJ/UZP6OGs3w
bfLk//i1p2Yxmfqe9lhS/Xvvha1kbt7MyFzPAiAUW2YMdpq2X70DzehNMoPcGLd65j7dUmc4mXfe
ufT3zZ0jl7cIB8xu/l3EYwk0tlzaDHngHbp9BRLhAVMkNBNuRDKX7ID9lPbWLCeTV/BZ8tdILZv4
oOJlmZjUrQsBectaMOK1HsS217oeQZ1aJG2POCmvmzxRkMo7M4IPHoyX5rtemsw5qhwMWxuS3DNo
t2cjsyiwiAATi/KHoxI6ciygF7tf8hwl2d2/dXg1lB4/gz/rM5DOXjKOXJtV85FxqiJAOKunsAcJ
M0Ai2PUd8yT3XRsau6/cW728VBqbs415Tfzg0hZT6iquE/daO8zE36LgdPJmyZKz07AglBwQt2U1
Nde+w1/kl8+3nhe+s9Nc6MW/3QnXe/IxgZSvrJDxKECLIfukB6x5K33paQV6acebJr1PzS3/QSDN
j6zMWfyP+kWS6KXwltziapS8eFFD0zOJh7p0kMg7j0QlWsxN2Pwr/00bGqUMb0F8fdjFMMLRJziz
EhUr2FZHd6ZzA6FobZp7ch93klf6lHdjkv5ypXrE9fLW0VtxnKJ3fU0D91bPwIJj0ODEmvxLmfwG
Ubp/eB7Rozon1ewiAOI8LopaUOtBCNo1pYQOM8c8464rkUX/mCWsJNdPN028v5K1tWvzwIuDJ9Ui
7jZ/CfobSXKerS0e30R249LaPeBzcM+F8KA2pZxCb0iRB8poHY4P/eDFb/MDcJPe8s4C4tFQ4S9B
1LHNjSaOYluUxr8/ayanwP9KmBIAl6IZ6CDCcoiBXljeX4fkfYI1piaNwzfVmU09FtolRAD97BmQ
jqinX5/2BfQmND6xI234ayVCmNKBQvszdcw5+2VSFiwdjkzpoilMZjLyqMN9fc6lxhmUn8fG83mv
hG88oestSCfpk62prSThOh/WWqepaCmsDYixirTsApuM9qlZNbbMizrkNbaWfr347cURfm7yu/fU
KI/Q06Mv1PNCL2QbNsG5PtReWZctuJIFluZYWLxpsbTZaHEdkNv5IOBcP1Y1kL7x/fUGiGddLcWK
dA6d9VkfQv3h6nSHqfgc5eeg5o1kdiFZt/oGZmdfvrEzVnDQ+gPvUyg42Yflru4Snoo0TllSWPO5
otzxepogwuDR/TBjXahBjH42YawQx5cYt03vPvoKIC6hJUxPThxmXKBSnWBcDE3v9WDVJh8g3Drb
P41z4YM0WljZmxFM6+G5VNtMpFt9woyeu7HaMwHO6rRT4Zl+RSznrpHkRCgq6yBkd5X+isD26bci
+DLF6lfSeT4gvRVpEfFy64Fe+tvwNG5C7bSNZx+BrpyEMz8BMi7uWyTviGvjSnMRHpdHJU4FNX1w
xfNjfm2LyoF5GaREaDc0oQU2y2TBTOCeyhVniv2BjoV2WOwCozxmGmKq/8juUCI0lup1MkoIxFHw
U6p0BxDU/Ft1C6ij/BSXW3eAMhuUDB5zgxjylNFQUoyHSHtEdnisWz66Db2/W24lBDJm+DpYXvUJ
kB8yNiIYFxUO0/wk2cTh6yy682tWt9E3fkj+LcPTbWKBNkidNnKoycZdsxyeDfyl8ntNsHCI4QY3
PmnQcBd0rHFIXj0Z0JwVRJs5gcbs2u25iiyqTOenxKc77mNFFcrRwP4TU3clSSWUvaYBMe5+WG0V
K7BoxcQHIKWboLIz70LnlLBzNTKrbM8dxm3gpPIjXcFkeHkpYwH8UzESAIh+b+fZYVfXhPSCo3cC
8UhFd16xFLf1tIGrvVLhvKhBWQo/X5XS2knZMKmIgGmqquLSIHwSLaC1+Uz+rTNgOg5A7OzQfg+D
Aqz6/IdTS84WZXLwk/E1U4G0ZLRbYbKTDa5YVSjmEwpZNoVHBT5v1bltBSJLsU5mzc1pcvi7nUeU
k0xiwaKVTXSRlFv46p4ENGMfcPjD7b2nQfLfUIETS983imLqTD+tM+sgzXglJsePdqxnGJ/SROyA
P5Y+jN2mknKPtzTwxiT8u8NrnlKNHyU2y4EIgi6s/A4KNRMaHfoWwZkBD2CgBHKthCcQVg+KIxbl
vxkkGyucikIlSr5T5TnMpcEfFVCOSAm1qSQGUiBOHtVUtrLt/zuiJ2AvLcihrxqe9EJ1vkyvl9lx
V0ZowX4TYwwi0xgEMo6QMNN2CR8BnQw+/lzrGQ9TJ3ywJ28xs2fNI2suBa2Lic1/XM9JK+Y4J8+k
rlmLUCbT/8Oywl5/OYoC1G3/JnQs8uBPysGymOB1TTMsP8J2cboJ9wL7oFAfzlgq4hZExmgl/rPF
Yk9VfdoB3/a84A1VinhGKe2HjALdV59vaCN7PnxqJ8M4GLqzaW7nypkVmwM7m0Falq9/ljDiger6
9qMJmWXuRhQROXvIQs4fenkzqvtXdJpMb4Qc648yzKTJtNgmsNQ5/Pfd6qdxfKkVerlnodKVRaDx
l1yEuUu+5eKtYDBVaF+3G703V6gzO/bXlgtpGcR5hfA5R/nfZ6cQujahpjBAk0NC8TZVjl3misUh
VVXV9hzSRn7X73dG9QASl5O1+UIuljuiZEODw5CrFzjnmI+MrqLParrE6Q2raulaOkrImuw4Tyfn
Sj4P2qFmzhZPCS/A3lo6DxdBBQcu1g/txBFgXToKF9BPtQ1kNWnV1GSapx6OJzoheuQccunAQsQE
QVHetyLkKmZmc24+/vbrcWpFFWeXL+T34len5wU8gpOJs1FVGpyJxZBE+7MEkoAs19JwL0HtLTDt
5gtq81iUnl74HNWv14s8FHKQvpYeyaMkBH3L/Ijs1X7XRHMoOUZTa0FK5ut+crz6xNZy3slPS/Y6
9HC2aOoDUr+w8dtsshJS9L6VKYsnVKIbpzuiCMe2zA2baeqNl/a/k3Tc/Azfjw4SiafzagSAJdHd
IoarrOtwdJTX+nfS6kqhLsSY5EnFdYtPJWyblkp1sVaDRtVMEycd8SynypH+WgQfIF0ywGTQPOnV
aLhr6QM8IYMVP0SowUE3OfvKNWIfKYcgISvKATrU/iEfoxiTQap6cco3kQ7+z1j4g6vQJjg564FY
zWTvgyvdZSW+beAQIBdTBo1Bt3IEwE6wskjwc0RWJp3K/nHelgrCu32JVYtSt/n87dIvY9LJAYbh
7f6qCQd3lBFqW+xDDpwhWmNq/YE29eQpUR50FmI3uEuhfYcaENoAjF6exMosOwgm1YFVvSXGvkGn
gT9cfcVVv0Dh0ZDwrgVVBhxJH+jJ14k7lE5UxpHIvwpeDQnDqOOe2FEvBPe+t1yvqwBabydU1Pnv
sPva99q31HUDP1L7fi2tvDFt4DKXM02fyEMesU0gYUWhSH4uBI+ih6G6flaQhHA5J8tReSNsstMf
cFwgSDNlvfm1eUe/hF60BCy6kxfy1+fcwIwyON1zSxxJNXgM77DsyqLBMRh67cKCRJXNtNi4jTRg
7dSZ83KNYDgLSynmCm8reI6wTTUn1lzmfL0sdHBFtwltYiqjCbJqWX+9tRmdh0vzQrpP8KiyeaAd
nerIPVXvFynwR9YcGMc861k5Cjra2Gw3fX/BfY38pltfZ1vC6ZcID3PM3ajUIxyXdfv59MuIktB0
xWpcagP70zwSK8tHqt/R8HuPZqL0sjoexzFXbo93wTbeQIHbW42kdLq5ge16VbJjHn17TgYxiYBu
+rbF6BNhoXYPXLTDxYMKkL+9U34a3gB5tZuBpObBvDZ59NHJJR179wHzdLdo1I8MNgt7PuGuwlnR
WkDdhzwP4nJGb+Hv8YrnHSjKToWSLctjN1DkiFkrV1n53SVfijPjO/43Up1DlAH4nREyD06sVl4r
ICtJzsK0ifsFiaYyJV3D3F+W670lt/9BHmbqAIXrE2fmfZxQfE+HRg1rM1JjDK90HiQeoAsuJ/PW
yF482YQ/sefNuWmS6fgh7tG75S9j2Jqc3bP2KEEhhY/pxoxHLEbO+KEYiE6s1/iUD/PwoKmsl2YS
CRzWMOdfqqr8nMC8jMLgIMnSHEgWy3+JFhozyRkIlkl6grS/omumUvEApJI1gRHuOKkEPLJKlhCB
Hd28uG2nP7lOxtyS19z2SXWk0TnNyP1sS77KgI9xfBK3OTdRbR7fC3P1VrltKF7sMfRDOfV3eacj
j8uBgNZUT+VD+xAc9S/eVSrARp+/Sc2fpEV28xmg3KluOddiynGiFrt7b2d+9zBRqYES+9KAWvps
5WPlU4h0+imkAznTU+Yr5BlmWjBu3nptEJtd2o8xi0+86Ux8fEy/di1/DT3dKxRkMr3aSqqw5KTq
0D+4s5yG5I//JrvH9f1BwVfWN5O+Zh4M+1I09cjCDcHnfJ4XpFtIIC60eeGB8/DHJJW12ZEZoOZN
c5V7clVQLog7yyYPcA6OZbiLQhs1ZMj26AwrYUb78Wy77QaT2tQ0IrC7ZV8Ew5GjbjyP3e9+VIfH
FBncgpFmUJd39qkK8BPl6zkh/4zcalOCCSSOQ7Fea1prTHXGiHYvM2CSuP+flRgsS3MXH/ekiMzV
+g7V43jJK9H1jGNRTeJRiTIliy9QYyClC9/CzY8u/DgyXq27GJ+UPH5lyEhYeflmhqMn+1Q/sc9M
dfGNjj0dbi2ZrFoneCueAzN+Fh36snB2HiKmnFHaW1b76K1HtuIYIKXKazkPla8lFhrPn2qtkHH7
hlSw0+HTP4rKSOFvfQFe3NW6urnQRYGIJ/6I+98dX2sd1OYNWaT3kIwYkq2Gg0Dv3VV1lpR8kf/2
z0meTm7Riw5Q3KJTRIJpQvS02Y/8Ec1ga3wBf1I3W11QmQySDpIpSc4sE9Qu9lV/m33zYlnp9qUI
7hDIfDCND2tVFjiEn47b9ZMad5uSX+lCNEUPrkYOfpo3Jm2SwQmEGsqFAGkOJFHmwpSHbkhYElY3
J4vuF4j2k+GDxJFfaj6FspFGD7cxXB8PHrKJQcFijblBh8z+iRz8xD3B6TmU1BiiSaNGnGrIPAqP
YJ/h4MtUPOghr4UyUehXPYcF2meimqD5/6Qfe6txQPWEq/C64k3lmvuK5bOl3D+OncGNSfb1qFRY
M5oKXtXOxe3u23JQJOiYxYQIjVc2XGBl4JZoz0ojAADJnkUdNRN17EcaaYHEK8uqJD/1XA926yU1
bBaONDyJni6s0BSEOT7PjFCls1SRhXmLS7Q5Mv4Qf2poA02J4459zGeXTBiGVFiyH7+4Vh41zVHb
35jDILgEp09HHlZUfLyp76PCQhpUFEvlJnndqPXauRyvzxWRCgjd58kpjO/BXSQf2ynDc4ia36AS
TKNIt2sH+JCp+1JjxWRgR7lI2xwwowMrJtX7H4eJJ0dkIKMQ9IrUk1bC2TnTjp/l+9H9KZapxbH3
mDqc/4HT2HQNA2q9+uztNU5mwdFCSOTXGnTd6dLZIX8LdWX683Td7XdMtzRU3lk/z+XzaOcueywz
zYWlrCUEywKNsH6GdUH3BbLIAsT8/Eok8p2dyRfdryiEQkvvrHVejLl8U8LMOec0hg9iGLlLlnZb
hdfWflD3XdiDBjaPCY33xDVHtmVIpvSlK6vPmXyiS7M1lg7bHqV+m5uDJIr5mTP675EIdC+W5NR6
7rLi30n/GzHVvaNCNnyqQabjTrjS6UdnlwfyhQeyT2nDhY0xpI4Wsxjnj4CS4I1HIN2aCE4DIAOM
hs2yUOhzuk25vFA+TD2BCpMG8u2RfSRDE2gVSktyX61h+TL6ITNqJHXTsA4XFfbVLbS4ebHaH/gi
SWFOk14zg9aArwDzWcAamBYjs2dAyxAAWA2hFN059Pdwy6XopUJHgoLZpgIMU53xHiLO/tp2MjsO
/82J4fpbD4gV5hpbwcoV0TdjnQ2y8tbH1997kr4eZ06a/SO6oyaJoVGTdhiqZuvnp/lKF32OLAex
e57AgkcE/6/p6adbsf/aITOe+A5CsHSFe3l+1kcI8yWxYyemCptjjiU3DsWxw/cgrW8JZhGc7sk2
2D+qobIhoiP9vx9iwenE/fzoKiaOdTr9UoUzLM+1yQ2Jlajfxi6kwOhi38I1kWViWuD04OpxGcsG
9nvnLtHDYnIqi8nDwibrRkIu/tXwdY2QwgXjSNw7a1d5rX2schh5Ul/KD8dCc2f9N8GIVWyfMbDX
EmRgOW1xGWiOVPvSsTMqC4FUmv3L4qQRv8rlpsTgVlcHp+ErXUMUbI966fq9DqR+OE47W2oYWLX6
zwwP4W+qq9QQm6fPnEiu0nOhwSUchAVwjvYuUJ1Retrnkql0MJmM+2q6TjPiuzWEG2WRwchLZxdK
/MJ2FtzlAyiCvBW/tkxwWIRsJIRJWZBM044kDpRigs7dvCIEejwAgGxxA1JMC+GplY9d6MxojP0m
+9AnI3nYNBkrQoGLiEWK9nfIu0G34Ayos/+pABis8+0xh6PlYCCepsoHd87iGrtMkdZ5onUZaeJ7
E+ATYEhmsyvOQ4Xfcexl+cFEPumjSfDkSphlSUwndTRHotro/CtjUN4NkCuvec4bXtxB/5Z60nsU
jXGy/4d0xAK8nRjicisdRbok+GWGXOZp8mmVqc3KN+MqurPMM+H2T6bnzyCntZsOHMoLR+OvZtYm
/qPssljWLftQfLEvsJIqV9MDd42KHN6mcv7kij6FFU/gifzJi0QqXkz3xxpFcdfAWBlpX1UHc3+v
rSQVhlzKPgq8wjoA9ZCc9TzV5OG2AYKdkhRIr9iTJvhfq+jUtGJq8K4jkkw4GmyZr6uaDxBrAuOm
kLlpxYJQrwNh0uOI1JZbE6soNVPWwp9Edi1BqfkP7ZMx2zKTSnvItuUQZvt1w4Vh+nN9s0aGh869
SF6zehSiJBWj/HSdcvKe/qVJviU3awP/BQvGPp0lVP+afj7eze9ed/OPSdnkSnnnGH7JwjzzUr87
op2rLDsNCG1o0A39cwyblJMpXi4wC3JIH40MC8MZPAFDyUpNbdCzaC/yjdbMsjERaQqij0ppX/c1
hmf2pCUMonPNdt61Yr08WazuZoFPkHQpjZ+/YLKng1rt/xmO71PSO2dkfW8Te0Qa0mORiYWKIQG/
V+8Jee/3o2GiLwKZGxGi4uPfpcwnY/MKG2vG1anD0UJ4lWYL5bEFtYL5oYmW1EbTuFDGvicKWclS
5A+P+TGQg1I3KXLXKqhC9MN/MPgai5u0T+Ddn4uvXzlUS1hgdxTUYP1JoJkPSYUpZjWneFeDTG1B
Lcc6GB8gGWeuWI/n/Z1Uosx7olWj8PI3rGAZxkR1w9abGGtCZUBa8jV+C/sN/y1kt7DJHc3iJ6Bo
3FWgFW/1nrQmdi1HAXo8+z4ksoqimV68ttC9IEoaLo4IjG6tkNPjrLfBGBCFgD6vkf26npbeypoB
5GsDzEMXG7jJjTQrBwBjfyQCOqt2/pFE4WU/g/QkpmEYjyQbjRVnHG6rBSfAi6bOckYqDM28inrR
YVf50RuoDEE0Ysce41dDb42m0OK73LQE81P/NmeVrNf0+oAXiABsmzGrl4rMjJJg4NbaKzgQ18hA
/z+3y6qvdsy9EXUz1eQMCEYDtlqcd9bO2u9Sj6B9qE8WeyJvlnWbx+JsGzmSbOor+ec0pF3YWQBe
uLcCViMbD1T6UbD8muwD9Eb8w0MaAEROlS7/+LMMkFMihQw81TuEtmTKkOuPyowO/ESG/W6M8ZWX
nZJYCxhhFBm/WHQetkRL5CdiPQmxRSRA5iQuDr1jcirWqCaJ/ieNR63JK3R641RxOGKfGmpJ44aH
8bPFQjbaV8jHJCA+FC7+BNZNJW0ST64p9FdyVpKhlQL44QGvvacNYQxXwpxRvsjeEXxviJVjKdFY
FmIGLXWDuij+L8F7b8xhGzOj2zlAg8K5ZSdgJm0UlbBG2wvKg7MVjsQoYVvuzkQKpHalPrKKv3m/
WCFFib1jRVvS2XMeEjxJDmyTnXXBVHa+Ylzr/t04RSFmpWHp4dVb2Yt6SD17INKW/EtpdhtHDvDh
+sPfII6Lh3ZDa0k0+fbQZpvtlzFZ10kU7yVKqs+jTTvMCVsX4AprnI09QTusPXjWXlfDYyMU1xeH
QtSq957OmHmqfDyFovetKzfxJl4gArKVTE8zkxPiKmvraRZcQCw6sAdzwqMABtRKe9afCwUzTktM
qCTwOP4QNa3m0rkEjBOXT6AV4FsEV4BK44hgBwzMOwHk6+oxi2njt3RKaZbM5bzsfnkYFav0q2fC
5K7T6DGJZ4C9XT2zdjMGqJUJUX+33glVxtrClluyiwTpS31rMvXbpMyxHPTzFUorJ/NuF1HWylcL
ZKo9T3qDtpBwMNcskIP++zOhu5zo+pmiONhWZ3jde35BbP+OC1+QUpAr5Whv8gX77gCwaVuHgdpn
5w8ULrIkenHjkEChu0XZzqS/0fLHq4XBo25DdP+ZIRY9CbWcl1vKqpc/wNEbktahTWYsTHWvQBar
cDbw7ydJ0qb+TdaXw+lEBtawZQfVTfWDb3HtTDsPJktFdk1q2u53QCm+PUuHpRXrmm8QPzJT9HOW
YR6Yo23W5e3AWkJycsmSucnNMaZQ0G9YWrynCRwrZBW6tx1+g/eSeS3yu+17u07dV2hoiM+Okysc
fZP0JQR/6jrdLkfY4kIzEjVXs4IAwS/MfMEDDI0Eom8yMfL1nX9uJyr5W9jh3ufkAxE7zhUCCH7S
CkKY9KXY9xHQvEP7Y7TW/0ydOZ5kvgjiXfo9++uv/uCE0wUDBgwQxZ2A5bKqYUREAY2m/o/LzTHb
BR/FA4Wn1PVI7cDjjKnnyC1XSzTcWqBhQMxh5ho6WMPz9AqwEOiOCWBJ2zDSAgSikNhsM89mhkJI
SbqD+reL7NThiiDb59DMwlFZ+N30Ip3OqbMdBJt9ZWcfTvN012g4sgMM3GG13Fv7twfYK+FgOtiL
frAfZBKjBiEpg0+/3r+vSDP+8bPoxBiIMlTlyVuVaE+5at/+yc8FO3/D4gYED6S381imzVBrdHel
SGSYGAYiRYrdgAWVDXgFlWNDDI3WhstKLEN3ytgjcbOK92EtlMSpY57fuGuscW+VYFH4rYajYEft
5teZkQQ/Q74da0/KBsi5A5W5lQizRCzXbb1EKmTImgBP2DDbGMBGY92eH1kiBXvPDuDLpPzGAPzn
P0TNqsHjiRICamT9/p9sQPgwstjleEDzWMiVh1eqaK630WU2oMryhDriDPb7M13ZvvRPcUQOBzhD
EBoHB3uSLhtvBplyNqXmYHP6YLXH4iF1xaKGu0MMysvQhifjoa/rjiEfYXRfv0RdFoKseWNe36/b
FUZAFyOTnm2ApXi0Ezd2pA0XKJjjCSt16pA7xiCqkThGijfcdNrRfXPGXepmvUsHnvLz8oNkaVmZ
A0EfFX9WpWi9dl5OD/9X1m+C054JtKwcFKUszJSHvHcAplnPc19X9XmV7CwHZcBd6zvMzpLn2GzF
XCVI/e5DzsPOH4uYIMOUWi3SEYrb6Jwu8WCnJVoEEZUIO/HcgTqZAIviEHoCDokcubO/HwoRPMJH
aHWrDH1Izhv718m7Z6k5aNtW2XpfWd4z3140V/PPWvouuXc+GyMWgFuITGZcNxWnfdFczF7lag2P
XF8Hzn/GpU4vDva5S/oEyKwF9ZYlOdBe9Z3ZO4H3oLQDbiPZpUuyIpz9o0nbvO0mOhUL0fGdqXCA
HO5WeVxunoRbbDhByoUhoAcC/4tfgvtBtVlLKRFp2IQxzlNO/L5PuXn8A2iqhrMYSmLbZK4ehPuM
VDAvqJ5gYE/kLKCU/VepupfraHNDFxGnIq9jVIPXtZUUnnaUvlqD5SOARNe+I2uNC95z17CdC5I1
PNhgj8z5F2lJfQ7xoUPQir4R+VjBsTz1aRvqvv8jxa8ugaJAj3hg22UWwtKFA3eLeFmS/159Mg8w
RqhZl3uK7ISe5uVZ6f66H0nZ7D5vnaLu8XWRRlIGyARp61ZZy6z/TQ71gCGkCjDH2m/BUhUiB4UP
wf1z4MA0YEySpGpPuaHr6h/qBYyWURNU2i9HWKp4DTPcrFXm8KQmPJ/4BhUKT0ikRRjxFD/bmqHR
nUUVDFvDKCCRD/xRt9+JH9jbGMz3+erylc+Jd60F8CxnO/WbRWXGkjKABy3CPQ9wVRhZSEWfgvtI
YeNokxHjI95d+qB8dcMsqV34tLGo8Uqv66I8fQLONdi8nJevEkuPpQVzpMFVUFH6CkoZ21mbiASs
+Hd9VjjVX/0q5+0AUryVq8vIcQ2kuI6wzYArAZkouNclCOqKsn8Q29YTrPA60bIDNnLEq9LfRNcY
5cOEAi3Qdx6gRfJ6Z40zHIUTUaUoxF/OR8oXL/vmT2ixBoJQJfidR5PHSGyMpy/TEKEaHcKemWFW
n6VH+aM6QiM75EJpkthbTNmrMTwwhmH2rfZiizz/C5bYmqaTSpLlO/dM2hDw5HwFdH9GW++6RJf6
6iOzryrPFNbYBkiV4AfLC7MoxnDaRDxvmJmOQEjrSZ8C0jiw7wF+DxK9f5fcQM5Oy5nj+D/8Au1/
8/FssW/GsWXa38bh2UTy98gPBMNOJKefGZeXqGEBPIZAlL40eA87qNNshZ63gOfvaLaib4PtCEBa
AH6W/gj7Saxq61P2GO93A7qyshQ8ft5RO91duOWinvuqwNs5g/xMlQbJzsVOv1mpb+/FoVk3Alza
WqHj2/IOVx3seR7uByGLEWVvEtOLla08ta2RexVZCcni9RckddWlYFXhSrpWn3ISfjJkwN3Pl1Kb
wODM9jWwIy8isfNbMARX8ZyHYMzIyM1kJIDQwCCHbWlfyMU5DxeyKCLJHkfqT7WsZxn80a7cLbRY
5sdr4cDxwdkOs0U/i+PTX1LemN0tAwo38fDKDOfd4yM+gTEmDH4v4uKf5rud77Y+MU97VOeg0RzZ
9I+HjXlsvdj8CiSSo4Dl41SjSvmfl5/WoE8wGH4cc2pkUs5a2OtflfV7nalpDQsM9tSWP02c0AC8
GgW16M++1DzLEMNiC2rIm/g2IRJOEckxBQKDLcA2Rrs/ZaZVhP9ooP5R135UNHV9b10aMzgwaMUV
2WiE8rBxHJIy4MJ2AuX5HFsoudrI89AlTfCULsW5k/EqUNwsMBMOt6BbgBQCmLhcKvTLt9ZCbnM3
tyTSd+NcwbWfoa5cB7U74mCKSSMJQl2z2G8XgFevN5PbiHCpWrDFjkCc70BZlnKhIcyWtOWoB3ag
RSkV7C7Uw3nQtIuFlvnuoqeRMJKIp2ZrJm3SWLIpoWUN5ftHKLwU3uqxrtRjiWQwgACMHL9m6jUb
kMxdGKe8bn5YOw2LUVuSmcrQ4TCIlSV7VV0sHIdAyM9PtqhbxndKZt/aoOetrX2ztVQJpINSJfF6
XA163+zQkV6pGYeUkq6K4D7ocOKXF9bP066wXxCvq8hL0wPd52nzFWbW0/F0459FEjd30tN4YGZS
0xQ7+f6wQIXEXtdeyT3k3beSw8LK9rFLkYSeurzCCoj8RlOlYT58X9+K7ycqz8tT/oR5kzMhUT1+
JG0JCpjTlMn1TQAbuZP08orXJuHttuCODJBcNnRS9O09DoImKMpgi1rf5t1YPmWCz77VAkLhK/St
QztiuTepyA1ennw2e29MOcIzKfBK04QRYQPwn4FfI/5clXAwST06hMfC6urtBIqf6J5TA6cjR+Bq
U1qrQAoAhNI6LmxphtJ8uof3nW1YoIlALW3W/WTGjPj6+BSBTeQuYRjYxXAvGzKstltUkLbw4OY6
eiy3OVdJHG+2sx/DpeuVpNChyLPfW9dh2mHsUQjP1AZg26BiklMMRR5SwQBffUUF06hBhgPE9+M9
JuubNzMusvu3DwrCf80+nWhyIt6hR0LAC+/Ca+2e7q/lGkQH1yktOXW+ULUIEqYD7aWDEg3LOmKO
mVeV5wziOB00UiGV7jDZ4K6EwlWpT2cB6FZrioWl4LEM/4DGUUHY54hz3t9l6aX1EhlffwnJso58
Z/srpvu14LSsvN0NphwBc121SA9GO7320M33r/OXGlGg2UuxTjkwGiVws7RiElOkxALr8ZSK0ELJ
uDizIRNCkvHeWeVVY1mavd1qXq5QxmQnVeOle4XaWldCiunfH7ar5C8N+XrONyFF4gGihS3OLtQ1
hjONV++6KPWoiNYhMAidm2JkN4SnZpvNSi+Jlc6DDMfChqZQDio4khj7qUZrXZXTgrxoWRZTWQsJ
Qq6TNz4RNfmDIYPdIld2LsZ39/cfWQDC/IKL6+SEEBvhqkxhnn869D8o5jeSv+Zutqpm21PI5K0a
OjxUIA/123CMuAiX9Vrgti0rp5wLKOdjrQrJpbJewtUcgJ0aSMmIphIXpRuRiEjsNtR9u45yxI5X
KxiIk+Cws+yTbYQLxUUskxG+ZTs662XrtYY0oHTLkgO1zRmmQxLptL48k6WVDVuTBu/0R1ZMgHll
VWYxOASrWA2oG6aRFJPNwepvIE3aFF8XCzCpGeq0UKuY76ET14eG+oOKZSVFCQrQPVfIv5C+v8uK
fVmJOjLwqtl2Qpbefnc3v3CXbJhvqBm45xlifn+gQV9sWDM8hzM5MoiQGXEnhIAsuqW/n8WZ2VxZ
/AWp1LUeKbAxxfHqCvl1qu33ZuVvfUS/7+eP7mXHamCiK6mpdOEQ78TjyX89dCxxdR4YdvzxuST1
VuFiH5XCnazZZajxQ4MhmImAeWm2Foyp3HKM0rXN7ZfIzdk1XtoppwICqjiPcB+3UpRAKYvaS5Zo
4EsM4u63LhZ4GytTFM/KVRdbqQwIRuqlqAmmIAM38FGuhG93PbzFHEy5YawOy6j89snE2hq+R3zX
nngkDyN7OHAyI+8a4EDr2FFCVWLW9LrdXMzrC3bH9ufxw7qUrK92eu5UPJ72Og+vuEPk/6zxpd7J
VIpkK9BVAmryitnr//X9G5FZ27G0nvJgtBq/KWjz+/MEwlwucRXYeFwLErZV8kZNPESStTFZZqiE
/7TCubSeKIZyxrS5nbb186Cokt2H/EDBgTw0qC4uOg7JBjyz9yBR3LCF+9gpdhfnoYOhap+yjst3
5QyAIbECSXTJ68+x05+7TK2+80Ymzy0lN1efHrHnns3vwsk1FbLNairIn4wki6J+7HpeKhessGpx
nZ4HOuNGleY02PK0RXP6TxkYF3gzEupIh3MgRZWSgEed8RcpJv8+oAV/xfGTjAsfduoDTu7FUJWu
KnFl7206OrAOuMjAX2dbkADxhMlPA0oEgWXHt6AFHfou1AWBEDbgxz44T4OHxPdp6720pKJurWoR
uyoJ4zlub4VCu390/XARjDJO2qdHhG3J1v6LqVnQOGHXPDQwljnpRu2xQCkmQrGCi/UfoCWpaGU5
k8MVpLL/d1WKi+4EF5hPSM7y6Z/cFQzS2ku1ikQs2jdrX8DW15Wxrre4eAOnj0IXM07mo7MeFKus
DEZGkWTqWZbbNuXBIVMcCrr5On6w078uFTNHNW9I4IS8Uuf9JiK8GwG8Fa+YFAo0nU3Gy5X/slQH
3t908gHhIsxE8hgdM2fidFnffRsU1n3+fORg/3NI8seMCLdHmAbqhVqsFfYOYfFEm1tYLpzMZAMt
DG0GwSksD94y1YOjJTeOuZmZqsuGvObyQySRuMi6xgh8Hzu8pcJg47Wky/BLnm+3D8CBC565XZwG
5K+a19+akwb99ywdaX+S4uu5Jg2+CSnvIoGGjEk+5WyS6PIGCyxzaD5axaY/riT+qUUgh3tD2CXO
85wka2jjqAf+2zAjTZDUEXH8M4SXO49H7GtlHpIsEKXuSiCgA1ObcRucS73xU8FPgcX1YyNkxylq
bpxC5PfxPvsIIwc7hdVaCKfVS7zeb8Pwthnqy2yUOIVkeO/1U6GTx/f6ckykZPwhE2UycoyrkIKw
i1L0yv2uJd6qHOpF2IwJIeSDzQ5LVFKG9DglsS0MRYogbSKfWp/7jHZZ5kyFKMByOcYXB38Dt7tZ
PTQnInLKr3WbH9opwct/FrL0wIGhyq8u2q7iYmc6RlHEfd2HeI6dJf0CI7Yjuc6a73SS7DqM7mEb
5pQc31UFM+744H9BQLCQH1k4kE8L4e33tkEI1EAFLqmhV79iYfmIoHMgsnF4H9K9EpvlJX6x3doH
jzkYs5FgIeGVku76mnWqEC+V05qkST11WjznOgCQh2+QuiWXERnbQ/MX64OUDVo13COMld147FRR
LuVEWyN/RNXtNbv/fach5aK2AKmNSKwhlHiLmzrk0oDN78DEIiGbu79iJGas7zldwcRhagyOyjkp
j6eWa5U07TYhxq4Hw/7X8pFsHIejGGMQcxqNDPUOHIcAti/Q8x4ZWFldo2EXE0I7xyaFsI9iT21Y
e1oaCWVdTfB3J+A0hPzAcH8hn6OBtbRmgV2fqIKGTLv+6rNm4hliunjADnYDaQVqNRsnHZVvmo7K
ZgBBtbOmGoMogDofmknDX6avdACkWd/LPjXNehQj0FEq6lzuAmowGD6lHTuRmH5znKKciJlijU7f
r4Vp4N09AiY1GGAf9rgboy7TmLRZ8BYeWc+fmHiGmnzMxjaYvx8r02K8aLHii94jqPgasDwypfRz
XQfmnZayH/mL8KeaFyaUO12gRBPAAXY9KPN5Zq9PcgkqRmDM/rGx7HO9+7qzjj6bOiOVuqtSu7x/
vPhDLdX5WynMWQWEURB5iqGdAkTn7ophaa1gWNcAGmX2zs8WjlsdaUbOQ1wA35yRVQt4sOhcKG6y
ZjBsqE0OQu4NydbrPThjEg62s7zGYHACqRk6c0zYB1sWRmsDWG/TFfJnZxujW0cfRctUAVLC3lTd
DIHxCRcXJ1QZUo2kwSobsPwYBrUKASngZ1LpYD3YD3q51/xvUoF2Tn0ZGKzEHfmLZnb5tkpX1Ix3
GI5egfPYtcP0S3nxN4jT3hRCO/EG3ep0EPONZh5M6cTN6fdOFS0yp04c/Gmwnm4qAg1yZnRqsRWH
dRCVzZgBUM2KD3M5pfj4x7fr3P20Sbkg4cJjxrF69b+mKGS7RxKzc+Gs4QVOhZnh4HiJwzue/3yH
do+Hy190q425+uxXLr0ECttYlyBuxO8eHlp40022G/7MuEora/rU1KxTJZiMhsbrxa/dp5oZk6vx
A+bU9YfDPib77RvoLOt6uGcPcqP203lQrVc861BSrAFCjEvRp+lorUWmcQz4f+HQyoN5T0/oo9Ue
3rFtPH04/CHlprtCEW2RHRxY3K/ipMNVZi2PPL2YzrkMnmN0IhdktuzYL7hbNu3k3rJLrropUdyU
sd0sinkh9q9+gZFlHGr9/mXdGEOTBt11CKZkouNQ9ukKpBWImTPFeOakdJwJcw8ItJxMjm229fRa
IOPYi2VoAHWHa/nWezsgiR25dI0RO1ACj3sLA/h3rBvX7WrQ2j+luWBQg6oCljU3ixMYJyC/gpzV
UWtqM/m/gAtVyw0qV79QxMCWIw4e7OHHeRFOdBzb9Oba1IJjQhq/STN2MKbU9oQoMN76Wc+w+3sD
y0TqeszV3FC2Tc1d370qVRqduKMCsYwMcVE3heaG99mCFYE28HCH4OtHITlAWK9pIqdBh5BYvC5j
TYwg8ewXmH91b/DdoWm9vndkAaVbRW8y/ftUKd1IeW/iKjr07J0WXBXkPe4JIl9YQDxKk+JFYlB/
f6TUwazhJX7e4m8lFX0u8G+prZHyHxwNha+BpYONtk22qLHfSB8jF/SJrn7ILoKZqTjRg6qVCD3q
nUh9zD8GJcQrGTEbZQyzzNS12r1TxQmQLHIWtVwlWd3pxQuCYXLRbd7vXn4E2A49DHN5Ka5aXNdx
nIjYXZfaviYRW6o0BaSxYnnihUuLBBEFs1Cymm7D31Xp9u5ZKTJ+F6wjNJnPMywDM86ez0/Brdsb
H5rfJrOYF0pWZ35IMZYFU9xDEKrfyDdK9xihf/wSORu97QpKKBmHT5SW62R6wr8l+XUTBfHf6lZv
A44ccN7Bd55PH9TmOcgcgsuZyUZ/K285c4oukBNkio3GZ+i5I4dcWFMJB3tSrbfqsbdRYRe3DvAE
4OA7UT6vUUtnyisbs2e46vGTrKOtURpsxIkf+JLbgqbIUGHkNoSX44wuV/SA+wnoQFB/rNFcXPTK
mdEp6/SdiuhpaE3yL3OlvvVaeDzbHHRVeY7FGDjtpueC1HZGI7lJ8vf+Skao84eSaKpVHLwBn9KK
BpEkLOs/0Yw7q+BJw3TyXygsHWMwSQAQ0eF0hHLAyFWhVBR5b+FNpNjvDNUBAj35M1ISww1az5NE
G80bDDcWwSw2tP2+1v9+OVGd9ZoWYH0osGChBakv0UuLL4m4PvbxlQgA9ffNoRiK919EL/ApiNux
1HSCU577cHSQ/kHtzL4mjB6IC/2DaWxlU3CLb2aum2O8UFSZ1iX6l2YmEa2/NTWAWprPXAvjYbrA
AFLgh8SnQvtjofwoSUAml5m3QJ8XKeHQPhzbbLB4WuUzLYVrHL5rAXjQs+TYjQsKb5QXgiIjjWvz
Fvs3WvdkJwnSpDnXoEhZN9u6lBOhktyfNhnXqSU/F/tQpwL5W+mwI+5VeKJo2Ej03UIVzMyp9uCV
IMyEdSE3V0j1GSxQ9eVjd22lTjY647lsXKuBTnnNs0iWixfRc6g+Og4mS5q5RZ8V71WXv3IkU7sT
4pscDSY7XfVfjhKlAMlSG2y2yV0yYQgqgyu/H7hRRAAoUupBLL33fGEJno6+3zrhdsJsVtDjYGr8
pbOpqm0Py4JG2lj+ilruWM0ysk2CV6JJ7CZRg9n3QEDDNNlYHyHMMbukkkcCVm4WILOuWr1vdYs+
xqHZZefALco3GcJUB3bVCcJCrizVjeQmuxJjTtR2fz0C77y9B36SQ+nU6FrCHVQlWQKlrTWjQq+2
zJ6AaNnjfq6wlUxO1XdbwhjoL1LSCDO3jqADpUaYJf7CUpAh1/hxHQ4YxJwVaPsNMjX4pM5DLFvz
WJVqRTPLPeAzf2tAvB/1Fhe4/hAiNDLQSmMjS9l6WFQQbfRzx/n5f7sgyole3h+aAlTTLCH9mmc5
RpvUr4pDmu2fdF3NgCC5/Bu5lKv21hgrJBCplIoCcGNOlgiDcj6eLQGJd1QW4/Je4izXHowgr0c4
JQttNv6lx4S949XddiZ+87t031w0+HPIy4MW0PHjEAcF/OYD654n40atFt9rpqI8EmL96vQ0FYby
558m6VTeo/wyNBc8AiScqvORe7fYXeFzZErGO5RaEF91s85A3RD52hKsJsuK7LKdtZOnBxSy6cp/
MCUXG4YPOtZmB7u2GsCk9RyLuSIFKbHs9wounXVkr/gXg9/Hg2fDstmudGaPwcHIK2aJpJF7Owdr
rlz+RFN7Arc9/TXax2oMm/oLmEBAqLsbgdQ8xOW8apxVFBwNKwVVD5ogoduFt9DEhSPGwD5rE9Xc
c3T3XVsdvplRjcfT1MDxNx/HiPn8viGY1q64d7jjjlZGa+raL2z+9Kvb9pwLvbELsflYtqTtNUUY
16IUhHCUJtpxWqY+RB8GXdthEvLSTjAtg5r/91VCvre5mp1OjpQZ1W7x3Vh6RvKuPMOI3IeY4An7
DXc5Zf5Ww/n83Ru2H3AoaEMEv9Nh7R8EDiq296FC2vvckCAzooVme+puwEbgOH5U1ansIabScerc
Bvrhx80I5dMnxa3gA8rOO/gPvXCXlbs4unU8GtZ8w+qqOm5qLSjPYBJL0kcJCWrakY8Ql9N+YvD3
FcqoNl9YzW7Vrg/If7RtMTRqPD+iGBPmzv46AunixvWZdKEBEmpe7TOHsuVMRT0CisnhBewT9rVk
s5OqZT4D+uawLiKY6xWOsXPnQg72GphtPyz0yMXmahTSbn6xnbUTK+QaXbF1WYe5DPDiGels5qMo
iVm18FHmGYscBg+gVZlAtaug6lKid+Smb4eB9Gv7NohM+GbNO/plHhEgmNUag9tzSGh9Ow4t/gvs
+9exFr6DA1h1YoOnp7hBTzN9v0dUhj47AfNbJxV1PWWLTKmj9PuFHPOn8vZ5U85itdK2GDHfHg/t
4UMgJEfqqn1wKg92V6Cc8LN1h2phXGLzdO9zuW215X8NgMuY5VcxToUURz+T2wPEoHx1XYro3MT1
rAwEpV0xEpAocw/UyVMXVH3uzSCBrvEg29019BCRvta8EhmVeQ/kio6nCVlUl/2DH15S2NWYmINE
4enYf8sP/OQSmaC03tGNZJKdw/A2d9/eAqab5XBIxyKWx6OdyQpmoGqauYxgI6BnyDmQ5UcXpjqe
lysce1JNdlNDdfNp7F6U+TVRI6I9COaQ2FGkCyXIYDkUlpmzvQN2Mk+GcXu5kJWv/isUDp12DZlr
chJBeHlB89Lj4LYHZ2Gzkdm5O1MxUm1ZwtlscF+KsH4Oq20ks4lWBQbxJ+v/zqYjQCWXw0N8z7+T
di/YmwTjGI4bnJc6r7cDAT1BjA/xeGQEJtvzD68j4TJqWBHtyYvZ3DWK9mCd1lPRqV4uIwcR2C8X
/DWFMhBslMTkW9lpwMz/CUYKtHc3rMMLSC15piQGwMRwtdu0taFlf75FFr2ti+E4gia+0qY7EYyx
Sj7qtE8kWequhywM3GbFeCxr3b9f29BtEPyVL1b0sfXEMyFNKBOlbaVB4QFAY6oWYQBB/d98/xJx
Dmxg9NU8z7oRWNXlgDP1WsG11pry66qegKYNSK7QXYJf3b3MUYZBhzveAWAe2vqhTCE1gfmgbEXR
wgdmSH/WFIuSEbYBIwOpBExmR/DWks/QHshuYCN885b0nfD7f8sSu2656VbW7tV9a89ToOwrpRaC
jCpdcCUkHuiYJpbNlBXSaEAHL9CmsIRKknpxiP/gxU9nRVzvZfD9SDT2zWdIReN7IrZ2jfXbq0Qp
QPA/fo57Bo6E9KnfXk7sgFaK4eTOoJGn1Lp27JXffz65NXbryZG78BERhvvzO3ATrR3CyVgY39Cl
RQYN3St3gxNTHZ551RI8R256wLjETwgvfHLZu2GstjNgTX6MEOGw5UhNewwcTKqeWCvFXFKqRHJN
jFzvdX3iIipv57ZWahoSlxeDTE5ZqZsy1yqqBt5e8fjdlu+rMS+9atE3ZdiNUCQZzfJLM3Bfc5oB
rjzQQKwJpseMJBD5jTdZZCsGQ9/Fx8S7TbRM0+GTkwn5B0VipyfDe2GmCJBmWfzW5coacHq+3D/f
5pBAGwIImAjVtOIkPNVavnUqWVpr6FI3JFC9J2G/PWYuhEB7tWoKAk7tNwuOUSOfoTeM7CTgubXo
3XepGaZXZK5qBItp/8Rt9SCs6KxGtJHzPBJImJFeKfzsuzN9vD3nzVzPb+64/JbpfTCFsfg85WDo
2YVlbeiFfS4ELjyvpyvCyFhXxZ/k2F6HWUwrC75+0VbffHaeGxgCxm5jxfYF4tI90EQ6F79YyoDz
H64KL425VOcmTkK5myu0RrxSZllxTqbP6iAlb+ifz2QwJpbCkijUS3CzI6y41p2Pko9/DJKSbewV
GRRT6Wrc2vFVaJSsTHsgpvWHD2z8IK3FNYmeNEs584ZCTAL0fZJHpjJZjRfyE2TvgFa0bxqO/n/6
oPDEW1NL42l/sDmmYSkIkroImhlRvwDQTdwfuYw3xcow1tLu4LfpoVsbHNwMykF51v95ZUfvWs0t
1tWIJzr/CVE/6mJFSgC3qBgHVLfQ6UT5afC92uBis5juSCQSlP0fvncXfJ1fxBApS4VCvkvaMkHG
qYC7MI/3mc9K0ZwIHX4+JhBQcrrXp3yiMzQGMKgyrKA4L39ZKZ9QdRDmQCgfl6eFlqa61g9M2+DS
KtmJBJoX+VgSAlXYu/RgweKDKcq2NaOePag9q7gasW565KsShWtZ7EmoAFA/L7P+3cd1q5gUPDHw
67JA6Nj5+lTBcVWEU2T7Q7wRmyr4AE71uj9dDRUuyoSrtyhKb2Ryo1yrYDgENVyAzmiHdHNb7M4R
3DIEhIXMUGm/LylDwOafgXB2gPf6GPm+oBbu/BP4eypzpJLPGew1RbjUWncJ7y9cgQj0Z9dSbymW
xSVjfCk5THm4XJLOPNBP3MqQ8fY7NmRNdg0V+1TlEsuXQS4t9tPIyBCPubW6OFstIQzyafGUp3U4
lE/cvQCnF5F2muk+Ke2OaTxf8P3TzNbyi83/npt5lG14/ZUdPB5evWOvdoJfbq5TaKFmWJNWF+HL
PQ3bKmP2rCUiTr0tf48+kM9FzjAcEyPrjM6aIIE1ArhnTVEA7U+C5hFa1bfzVF3O8ERdV1DcOQIj
XmT+9nTOqxwM3qhZbMxISV0YlWqW5pP2tscL/2hlofrQ+4b2NEAyFHxn4B5QET6nwO/9uDwj5IXH
bSRjokn7NBPi1l823Wj04GcZMudoZkOR1z6rl7QzHHtNG8PxWQv5ww9S3mxBjku2Nh3S2cBPVRqf
BCJQJYDJaheZ4lo1naYRNxtC+uuh1k1oHzQ8e95FFk6H0P0HYJfsuoubJ46t7m1Ja4Pos0z6DKcy
6j65ID/K+2WZ1WfWfN1PHJDvyoLn7Fi2d7R14D6lobG8Amba5YoQy4b8srnIu5EBry+m0Gx7TXX/
E2a5038uMeyFoeh1GxlDgjC8R0nAuO/7ZXSYp0sHBpNpZdhpig1rkdSlxN9MjSEYZSke4xkWQY1v
gq0ify+g5aqo1qZJAQVs4DnEglz5sfzrSYstXqpWqPbfqhnSIe1sBqcstt7PRiQBHDfdHTchLRdT
lAtElero0z6aR4Fou7/mL9xyiujg8+wvKelA5l43zmf9zhG9kwyxexAHA8edXa7z4qoV+c8Cb5pr
2LNmlf5GRVVDJvQIDOhdxz96jc5qnONOVQUibAZKsTBd/LyenKOCaUdwJ3tSNMklploqWeqWLRM8
VfFdn258XDxFspSGaCVDfQnEW3jQTMe36W0W69PsLb05WclzOdKXTQt8erAvBcb4eVtrEDky4mph
+Z/IEoG75K7/kiXukj5DYtJY4wKi4fr+OfcAIxPWlhwBCB0eAiYEvJj7brHyn6ABRqviGdQ5NYgR
B3R8dM6oig2ZClaAjqnkr+QwL8nuh339rO7lrQKt8aEDFoJCI2oDDp78lqSd2lTAKLXrCWLG/I+K
NaXkuRflyU08fUQe7baVEFhUnERrwAPH1aE+wQtg79K/xu5Lo9JpJecd2BpMaZqH0JOI3X9avR9i
f9nykJ8M1EMXIpI+b0LRbfL07CDNl14qskbfsOFDhUh25JjxUaGz8T6mBpVSyWRkSVvS9Wl2V9y5
dkuEbWLk/zXx272s2RCNhuCb0lUZB6LQTM5tyER9mYeTFnUFrcO25khSI2Ng5osxoe1xEt9twD0w
RRQ2PF7g4LKM12eJWMZW4K/2KB7lFU7e/eYn50Zu10oWS0js1dDCjITS919rcd9zVYdhNvLThH3T
BQ8zKm6q/72m1U97yE4uSd3xSbnhLqDGEdLWFxqZn/j7xrSfLoSTC2hi1xrK91l/NLS1tj+TBuLd
seeCkiv1Ll684/G8O9Pbtg99kpEbV1dOa0rjfYpPna3e0vwafdAgXydr2sxXIrVXjCvoESLtFKzL
A0c9qZGXCL+FBL9O1eLagNgluqlPwOhmGIsxz0ihvx0owAXlDZ7WeEbgGZ8BzQQctm0bv8pgK2k+
GIXAs4LBkVLjQ9tOoTRzPKcTM9SwoPfRdJhxcEg6pCBrTR7b/n+EPuJaGktvg69SMSRBR19F+4y+
zzsp1bgdbFIMIaqn867nMu2ZcEoZqyb0c5DsPVpz0idcGU3TJDqhPeZHv69tOdAig33VhtkH9/Gl
54zTT/3NuExj4iVMGA7Yjv1Seb69ZGjQluxAtV1AfHbwyCbvgEUg4kPSg1HFyNv9vlOK5P8tTiSt
VD12s9tLTzgK/yPW9xcDrEAOBh1hh1MnjSu5UUcs2BIiJqcOKVVKc7wj7P0D20QWjccpZzZeNQKU
9YE1mWbjrgyZE/ptMcS7voz+lTz8Km+5kcbsafmL02IQ+XsBHMOyrI5aOlemclzrC84rjCUxhPCy
ZR9aeeRsslLopSPwJ2IhQAwycjf21lg5xGr0++8zVo22flOWxmAmLmbGgGz1OH5TAq7AljHgPtU9
KlsA7OzwNPcUSi1lLzhs0xjTQnONe9O8CfiIXEhMBw4IgdV8BGxcWpTvDH62Xy/JYS9OeE+YMAOr
M76/6IEDAgNgB0GtehBhv9cI9kbixGqndUgEDzMPnE13yQD+4ijqODY85XpsYBT1ANsGPCM1JL8M
Q8dRyXIXCQEzuuDMLmfOeCQ3qbC+VCZ5Eu9ApTn1VMn3nfCe0UtybaPI1ccWf62UhZZdcsZnS+Da
3OAOMklXurxsOGu1pRLtFvfW/Jl4pEBpkHKUkLL8x+Ws+GwtZ2bAumFhysfeEy4mVc/qGGQIFSHh
Pu5llSA3GzTkQSZ2q9XcAh8NpndVNClxmsocunU41xBqvhrYXDVY4VrR+u/hs87BXK+6g5NJkOxx
72OXm5YJAExbXNaqCIXWQvrOSNe+du7/+ryKgXdmyIwPb4TOFm6hfXA3gq5jPmiW7KFLQspk44uE
0UKuBtOlKi9KAWIHsHt0AQKzihNPaUlPAL5WTdZI/kG6hfbk0Azym5gi1ENYVlM6KejV4kCa3ay9
8/HhXqpK+g1t6UwKMdsrfnkMR8/3lJvJUmTFTSaXbb2b3Qtzl+TfXxzI9Phc9XQBxKzCUS26wEZS
PsKNfaaXM9lvDuV5GJBkJhLEEcHjOPmazz5LxvvYxra3r1PnNcsJfUQvehH1XXmQarfppnhPpj3S
2B9CrCBuHhnZCXMzZXVIOBhNopLEH83PmGbRIEE3foP82XrUA/Sgq4hOPkFuvpPy99IrIob+Qe7J
dcprvivjACHidSzwb97flJ7+/UnxB4xuWlaiF4lVc2zPoLounEECzJeD4ZEPOmBkDaAdf2jNaOI/
Jef2QWr4obeZcB3qqIvKex1zjguklOxoZnfa7NCzpCLsU3QeGQRZZJVKijSo0l6rzeblLmzeYu0g
M33AXurdCxu+P/wbExJqEuia6lSLXPbheEo2bbWyT8ZOtjksBZWhJHPrTKkld35764BvUqdY267Q
NbacvLBIPbcS/U4y0qm+H/28R3Vv7m7JFeaTh1jnZTeBdp0JBSXmh9psS0vH9/ph1u2gP6hwhSTq
qQhBlkkZk1VVahCSEy1Rcs7OAXonvDRL+77Bzuh7Ig3U4s2zNbBkt4tD5hYSuYtinNgQebx41FT4
diSH7NnLF61IiWiDpdzCYPDpUcr3tXcWLO6VdyAgjjd0YWoWZskyJEhqPTpGp9RIhZ5qMlEpy1UW
5O9ds674wjM8nKJ0LGuw1iX+igF0J4jOcTseq9aMTgXWFvnsG76Esj0ifBejhaCARfxQ6z+hT3RY
v3kGOrsQ37gUt26DXs8dobWd7duSg80myiY0c7h+PwM13sTHtOHJFiIC7zd5kq3ri0QadY3eBFR+
K8XC43l6F92Eh7cYgnnveNSnzOnU7wRcDIwuxaT9/0VFQvjJp9ofLEExwyD8C7p7vnV6D0q3d7q3
LEKflxxq3f/H4Op6ga1h1m9nX06gnjZN2rnKkX3c9F3c/r5/880AexW/5qDvnZqbhYDYdGzGWXef
C7xfiXIglxDGTrDlxtmEew28vX2s6ZOBpP+g1IHo7QJR1ifE0ywzhS45P4DXkWWjZv2c8qsMHv2c
0zAPddV7fNaSWrPIhO1sd/NWs9ZTXtzs17avuevzxCPp6qP1czh6MOi2fTqKMQDZBFWgaJKRdhyy
dXE+PlV3m6g2zz4vmF/gHww1pLpC5v2JOmx0ZLGzFGyvAJ/iMB1YdRar7ddJRGafn98beB6C/xXA
sY0Wk/yBCtAnF1K/kvExhNqEJxXS5S3nnaTJ9vQzNEAMcpWxhB6impguHQzkQOpYV/0KkN/V+OrK
t1Rkk80FP9Z+pRbAM/yfegZCJGU5DwpmkPawFnWF1MA16/ELU05ECKToV7pZEY9ndKBASIB8j33T
D9ThRLkbgm9MJCl5Syuy3kvnZLeRQ8DEMbAj6bWVQCLFbsCksF0eVBTJXtSh7LOEaIIgfjnVWYXa
kBS0cT1lJioo+bh2CJXOlbf38L2574h4xT17x/QR4YEVW/cm/WxPtBArJ4ksdJwRusLJfUGjsbpM
wPVlIg9NzlaiUBQaISskEG8iyM22PfoduCq7YE524G9UmqZ9jB9fktTsBlBGuRjyiL1toWiWtw3J
Lj+4ak/xN6U8EaZawo4ew60UUQExKVQtQxswR41t5d0WBqgfYvUzCTT+dxUlby22CtcCqbZPpjAL
U1Zo/nnEND4PShwLU1O2/0nd4iU09FKmDDtNvkkdLgFrBjySsChHMOSOEPKFm4GiqLrcErYJ5U5v
d3Mnfd3KNmdHfwCsnwyhuzHWzlc5+UosJP69Q+2y1/YjO5q0cXrHaQYXpkKcEnJWtipr5CfNcGg7
vHKqGP59DoRR9hozqOiZvkTmOTtg4AXIzBwR+7/RfwHyxTiAAT3GTVB6gWOG0Yrxnk3LmKdguwtU
c78ecVd88eI0NqzMG4mlq0jihRvKkS8wW1GXn8ZYY61NHtzbYFvFHuaF03aW1i9Ar560JXwMYUF9
R4Y88ZAFBeQU6F1m4moBXWjjubGBS9GfgA5PEDm3g+QYAKjTUa3t+AjcM4k5amBeHB4AYbTvpj4f
7GZVpRJnvgNfcyt31O2PsYYs1/p6knLRq7izCrBUOq3wrXKuArm0FgwUGI7OwGlsqIRetTPn1m6w
AgQ2kDUc2wDZb3RtNB0wVoddy5Z+5/ptSB9G42TevfnF+dfs0kYe17nEB3DZ/+u2WiTxnZoEFdEl
RAz0qiDLPYULRjDW5Ro1Wt+/5RER+6PY3xMQ7pyYwJ8xn/Y/3/yELJSGDsGRE++YkiZkydU9diRE
D1TldlAv58tTd4/fvYlZ76I5/r2YyG6f1LMK2BaESFhRfJU+XGJohV/2ejXj08o2X9OunlpeMq6p
8PAi15f85Hr4giC4lZapEVrQSapQnPxvVUoyGOmWauRUhwnguIckDozA8JVCtonQLgtQ2PJ40Svm
61eacmjyAZxSAiWqbdMm05H9NTcmbELX3S5zcRFRYagPM0iOp6Ez51pCQ1ufrmIcvBsDiTw//nYR
eftJfmlTwtjboifwb9M58m9Sh0TR3nezavugg9fhdDjFBoYA3vR3ae8SKYpppiLb3UtHfV1m0z5m
+abG3/m4lCBTBLZ5WMcEh+ri8+5BYd5yNzVLF3sA+YxPBtI5OuLgAPMc3e2ai59lLhGBELWfrjHA
bta3rwWguek1ANCPVvyUfXXKa8jnAQ3FfufN39YaOxYAUaNUrbAD0zyzgcNstu3e8meFnIAJPN6/
kpUQ1w0Kn56prTPmmvZuO/p4pcc70gdb8qa1k1b7CR8EA4P+lpp7RLdHbn9INMTlwMFV/fJdA0ze
rP8HmnIq8WJjA4S15kJJFFn/JHbX64oVpPhDZH/ovzbpOtWQOWMJTk06B7EhYpXlZqReHBMyNdsz
3Sd8kZBYoAtoNiIn3X1suGHHh4DCXZ55EEXZydrHx781J3vDOrZrsSTtoUlO8zt9foKywbUQjvgw
xdkF2mjHGVHmi4Lzn+7FSKoTVD+G8fd+82sQggoD4zD+nYK7zKK42FUtWKFN4SCU0xiuxE4rVPWt
9XCDu5OQwbS5jkFjmSN7120NGKf2eZyx9TA0FQCTrAUARfSXTAHIWP80URHKDwM4ubeXOlXFi8T9
zjUpJFjvzPBIIdYfYFCH+Wvwfy0+w5+RYpSYdo4wGdkqlH5Ez6FTpgtjKIs18lCtzVbHH3GTxUM9
+jMnyEv17G+jqqCx2HQRJWdubuQQPqJfhPpTeKpyHjXI/bMzct+2s5LWxXAVr01E9JBlpEZeoUI2
quIfyNmEBg4RgKS1i3OELV7MEy6itHRwjHGqdzo8iMIsBJChsyAsEpeidevYwxTZ2ix3A0/zhxLR
IpN5AvXnDoVcpSWg+9bfCAieGEZ8rjmXRjLeRJtc6whWKgtgOEkBLxF5FdTWQfi24W9BSrrggxvB
NarDVqJybODGTnfSpD2525pU2jBow/7ld5nRqB18mvRZ+ysf2BGzATjjK0toD8p1kVWu6ii4xWVY
0MrLkuVN2I1a7UDsY6a7pfwwg5SjhXKeUwUf2C2cyjcGuEd8fnTgw43BSJqxyhfRf8kCn6icayyA
m6CBPelIaN99SQels4vvobhyZugXLQ5HS4XUOUdq/NCDWRJFvofpfplR4rw9CgNvanTnlmS/NTgw
ZlvuxqWoCjIiSw7LZoeoLUk3M4VJtAcgh+NIF0TqhSBqWty7p/uqrVAQRhEHqj7sw5q2N9p8nr42
W4GK6ahuV/EggTcfsjoxUrn70xgvTbjK8rDhUqm3r8ECL3riWq8SnMYzZ7ZggQj7iz+3DUfvNczT
pXDhnDcYGiGhZZf1AO8QA94dYPgPN9ab+1up5y3OBBVwbqnpw7myUEkP5Wm1cifDqfuO+r+G7IQC
aBL4PbKQF1ngb0Om4i7oklMO9h93rqcffmOyJeaYLR4lk4Qfe24IGb+H+vIkAEXYXLGx0vFyPBNG
/S2YdcHBjKjXONOHYapE4j4KVxaPlREqAcQffASA4YK5S3owE2310/idGu6mxC/v2/nTPtUK4b+p
RUXmRkF8BMoTPQ7k5IIzFbM2XMIP9HplzU8jEAbuA60thBmY2r32pYDTg8OAC/LAz2UUWYDu13Or
6cv/g4u3f/nYB2wjwQBMJomwzRfa493p3jL8KpJfhkiOZjXU0tufFoFUsjEIShvE1V3b3Apzs8rR
oHhIGjhGnkqsbT14EF1IAOD9UtrumBmnCrTgFHW1+5Q/xI50o1Jh6751zafVlPCLwlEmpOef8t+g
yi0Pbo30sd7PZgaL6SC+PQtGJ9rXviNjeIo1qMhhMn6ghcBErZdKlN4CVuKZ5qLJ6/PFRTb0ytiT
yfcn1zJH8Y9bFUu5NlXo7NGFu8cqKBD7swE3x2hx6EXrqxHzfdC/b1PhNoM/smKI52gwJ+VeJgSe
G90HDCI/zZ4tENogSkE8pO/DRMgJQvKv58drsSsqVZk439YUenIQ+qfwWKX+JVzg/jXZb0dGTvhS
DeEj/NXsW+Z+tVAqabumVZ535ouhXLgcKUj2gkXKe0iStZqv7frymQ9jQTvlCv+NJf4SXMTwFu2C
du+m+Vz/Hzn0AT/0oJsLBvwym6mnKsfEZa5WPMsjTcvghJ40YZApAN6pi6i3s1Yy1TgWDyJ+nuNC
g5iKmGqCG5QJsvVbIYDtY7IkHsih5MZp+zIFOUWG6dJYVyDWIvYoq42x9D4boKZoA6uY1/QT5Bxe
B+tYKHFGs2tMxmex5ky/SHPAyA4aCS1NQmfnYZu7EDYmcTyDmS78pdzqcmLJujnc1Ibbiwj9hK9m
N11lnhP2FG9JLsfsQQn1U6BNJ1+jsm44SBKyW0M26NfFJ9INcIW2RAnMSZNJ4AAtIuCwMiHsDZVQ
Ap3/XILSMSENJ5fxSRdCtfSWMXtBysGP3Lr2RUvjgZv5E7aDmM9nmqnkAhJm0wsQqeb6GDoKilXB
jUsAOidvt3upew86PXGEGZo/6UFA/tAhMZJARpPOx/ykwHIWlPvLTf2JAETM7JzbJfPnSwZiesLC
jBJc0MbsjFG/TDsUXcco5PmB7MBdy/BnaSJsOqnSSJW/4Rs8FqlYAlA1KezUiLWmYQnk4eEIdpki
rWDCJufHYaeW1Ha1BLzcqF06Dtj9yzzim2yQXX3pla1738iI4oxbeoH93laJwalAc7p+0DltLH7/
qVN1VhcwAdJXlJx5/SceDnvyG6vaNtYcy0uMrFvOKd75xsEFWcz7PjXvJVKrFZb5nnj/539thhY3
n+uHQ2nfDCWFN814VrIlH0NQpvXb1fdEn7srGU9/qm4RqEWkfCBEhTYaA+uLjsepoRRbVX0s0Bvp
woG+dMfhkWaKFhGMm/IGkjiWfovpb/6P7no39mpLXfiptHg209AnDMPWEiHVrn6AtJ3uwn1c4ri5
c8dMNdGeQST22DP3jR1lor3wxzMOkNk3+ahCSUDBsclDtaZ2R3K6esssgRNtjVqR5qiV5dt5MVDy
YznqamI9QA1kb72YSnqNIFaB2vRfVE0q+KfAV7KlUf73BE4naqbyF7iJgSvQoqhDvJChCOMIkAlW
hOSDe6twZYW3JCGFdb2mMeyiiaYASpmWhYdzZ4DS2pNLdW993bw/lsGaLeR2eak38RGq+uWW4d1y
oZNvjfh44FloGRtLXShbnJ1YwSv+XyNbw5ILsMNMz/5ntBYnOO4+vKCr2t9zv9aSOFxekosHBXJA
3NNkQcBg7wJuuBXKb2jri2g3Av1tiu9dcov+mvFANsTYV1FXrSkHfctmcfN4GPXLXfe/0afy4KPv
rOCgyUhu1fpwSUjN4bnJTNcb0Ay9nJBfNHQiHs/XIelLCbtV5llCzp1zwG/Jjy6FbM3d692kxvHc
1QVCQ9dFd3Jyno9GSkb3XqGSHT6MSdzrXyJl0UyZJB/2RAuIR5s4Q+jsYUuVWLJuRJaVtxtOLSkO
GSfxadOuFqI7LSsYMnv1nWIaPyz2Bnx8kaJwcxmPKUOy3vMOIKjpg7dwI+ySzbMFOdG8AFh5qA6N
RojQ3xrmosnCFOKBItfmXMPEB3AJ+FLa0Ms0WMcoIf8Ot7a3whLiCA/b1BRKe2eHzayWfliBS8/S
KRcxaVpzEY1TCIP8qgeZ4+S/Ppu5HyDno2EFAlYjDU6OZiIG8XPxIX1CUu2Mw8X7GiozkmIcM6nR
F4usPNfhJ+i0xQPnd/mC1HLjQNs3sAN77heREddbVvt3tA5qqZvE8TXE00EIDVtk1N3L/IclieSi
pf+cEOa2Giq8UROtaIFVeTb6+DFl3hT/Gjz7MyP4TAeblbfC58W9Br8cCB1ufyMEr/6V5aWjg64J
3JcvEZO51M0RUXOcKAFzWsA4pjAtWrfwzQ4msTev7zu5tMUejEKYh/rGS/h4KddxZjIeZ4RIxCN9
h6hXncyZK3Urr6RC312pN+bpmyv+U66x501LM1rTEINJyqGamkULtaMyOLe8jsijVApEdsJP+aVt
nnheh8xoZpTcsB/FzjPcIDgICLk8vWXA/YnYPxH/BgqMQkeS+8Qpvejni1qNMBpsSe6RvFo1GqjV
KDMiGfuQxcbcpVrTivV7wSAXs0Yfpj8p0nlq840ZLd8dhVo+Ynicr1+n010Cz3Rn+Vo5MQ/Fpc0q
be+fo0KQvzAWsoeQZ2miwxgr/oD7k79moHrSBUGSqgSibOwIMaNTOiOMvTY2QPpu0s7kcqi0ocWT
R3+ofFjvUDCbG8gAzu+anEKh2gGpYRbnAdzm+eH+MxcN2aQ8NBmmph1P4Hfy1VRroEpezqDUe0LG
/qlGfQWZJx60P1Ghf5f8tTdeJ9sudJ2u7qRin6KpI7bnJBzL2mIPCgsfR+QMEUJTWH6hX+XTNslD
8uV6KKPh8Ggos85ofta6ekE65Fx1M0iDVsxCdzcKEWNRfoFi1x0lsInM9M6d3jyVxhLH3S75gmGy
trbWI59qvEnliOfpIz99yTs0lGeSA6AsY303Y5CFmkSpwLSz+ZikSPGTINlOxJhzl+hFFQ5vuuCB
Ctg3Fy+LosxLnzlsIX/t8zyDUqBeNNHe1gZ7bwpl81V75pLa4Xfu2otB9wEh49bFJIxCQ0zJ1X1H
b1Mue6DrxCEC+OjNWz1rxaJagRDtde/kaXTI3kQxzIbOBLc09ndI13YrTRbOhCi9fdoXkdtNn3s+
4Qw3lceIgyz28N7ylp6yaEqEokKjLG/XcTNkhivlRWY/UANOLZMpsuPLZo/QIgVU3kaQUxJ5Gj3K
yeHRhqNEhrUv6hz8VrltSMs91EpWIR34SN6OIzpaQ3Lfc7bk1TgkvVpO05RejMY1yHyKuFnxNHfh
hM/W/I3UsnnGpgZ7KDUCttuiVo8UMs9AhxsGvooJn9MDF0Wo1fSDOVH77MXvTdqCyGa9T83txrqv
EmhxJTHjzIzZtB3MVedMwsfuQGopojLtskS8PGRIIsrHUIfEvvvzue73L6XMUOSkXkrvg8s/YmoE
OVc1NB4SMHVi3vmdlbK4s8WF6Hq8GSyb8tuo+U1QksOyzh6HsnWGJlvCCEal4fCv26/Dlmj0If1u
ng1Pnr/4sKPFO3NNOEjTkfwKIulD8rZ/pm8+tcJNEihWqwrjw/EuYZlCqk4pgug8XgXWA2YbYsLm
++tWHm1T+qPPbG3e1la7GpYWaA1//ifH5NnXWKMzVi6St2aD1NMEWTug51l6a/Zt1y7dxBCiHX24
KWan+rqcYIJJo1ARaIHXZmZsN0BdLu3UUU8aWX6iG/3MtD2DCCN2iYphUDL4hYB4GbGxrsFa5MOW
LVU+g7I+o3xTchpuUMrRAO0oSh6gwTON6UyzJ+UhzFbIiRN8POP/RddK0q4MfpA2aL5fF1daqAI3
BJIIM5cHi8cFRBh7Ek5Nb+kdEm36YNy45lXl1vWc6ZFrXRLg2pMBaXaJYftk1KvyF7k88tI/JxtP
qSV6A7T0CyzFQwO7z7/wjHKcVFTlXHwtBEulvMKA/9G6j0G7PZ0zNb7dC/MD2eohsAFzsKzGp1zQ
268Fm/HZa+MazvZMT2IPUVpNqSUXxlbkHODuFXVLscnxUzQqUdEQ8x6Wm5T81Oww73f4B1oTFcEJ
tCqanRwueB4EQuush6JqclCvVp8LWdTqee+cfDE6bA+17IbObLXRgxRh5d9vIHsWW2S5NP9tQjhW
SvDjBCg4tw2SQusQdzaTQtv2TbYZLkRbW4k75tRUGq8TOVdxay3thfiMOI66TMfsh2e6vq25WWxr
zw2/fYommdYikOqUkDlYc3Y5vniV5pekSWbEC37wxyxx1eiCrSFdtvSpzkXBr/zig2BoTs/QjvoW
vl+hi0aCt+GatbMGUEh4qcOprIxoWGETlb6VueK0mff2eAPsWikXZvEuaXcieoE6G/6N/pFafyx3
NaSUg5F5RtHahy3S3rV2ZU3bR2IZFKefv+vo+eUOaySdRTqH6lN6H8fkMfebBIGkgQuycjlVJxsp
pk47JdOSEGfAmvS3KTeuBmAnMjLVePrx0nDdDDBtKnB3r9Bq0Sb8l9aWgfFU8cVTy8BRwoqnRwn8
2lDht9WcRmBxvlCFBE/HyN4QXzPb72pgrzu06GtH/fGRZkYZD1mqWkD+FikkY5mughjO8QM1cVE3
ssnO2FcGd09cTvsCtN0WVkamoA69QaQhrKdw+AFEDkf/yTVzqT+rw5bWVUXqR78eTdOM4AD6W96V
x/x0ItVD3vNg2pbTHQOynoo7Mb3Q43LSMzGRlNpJk7eyuMZgHgEnV4rpSkGsUuAHhGpRsfhD7Wrp
3v/GmkYA9FoQ8XXBAsh8lMhL42scYy7OYeSbOPZ7ymTQOC+iXypNXrNHSSywJAKKQkAA4jn3yOqx
zy2eHJtpV8rSmzwcfyZLA6rMtdF7sIv6Kkc+em0QlayTqEhkIqhftnev+pxDOmxyd58oM6El94tY
eqmvlv5mCJ1nqyIaV/YeBdy2KbainIR9Raxy1/kteX8MdMzsWI15lqtjlR1Q51omFxMoHut+c56I
P6BwXD7t3u3RXxYv10khNJYULggGSN6SzwBx1hwhMrKHXzMFMJThQFoJ07yCsTAGveCOaBdIUogs
3Wpg2+dG6T7yO6EnoVvqC/vpz84NI0me8TF27LBDRGEwlagBTMtE/AWXcwZ7FEkWjkV1DlZWBQaH
VOLcj/v5EJdXjIPKttRuDPiHX3PI62nltdewIdkLSdG+zydf6F9BcedmXwjD/+839lidq7seDJqz
KzTKQCvM//kbU/gbRZ7/HTdiJOMeHpgBK4zQk1Gpr5jr3Y7ZV8T/V20Lhl4P0FSDaouVvi38uCdy
qtAnGto8xnlxx7wn5gnvsl1c+/WY7m0S8SsHLC08i1eAcmC+VK77uwCV7WdHYz1/DtIEB+4DC+Vs
jw0bFMLSG0q0espKUG+S3SwoKYp4AKkEWK8hdVVVOSqNm5JA3x+aBq1U4ZJ8GWustT0HNSH3GYgW
9MQpUdsfqUN/VLRsTbYSPDgRpJjo3onWDpejaH3axCSjfpDqrxV56FswFAfvPo2SQ6XJEyZW5yqz
uMH6XPKLjcW77zZidjfM6PuYxj1JLLaA1DLCDc/Mg2yfM+CsEfJr1J0SjBOrvwj5tSj/opmKfTjD
wUgKx0b8TAD1H4+3+XaM4HjtPEa7BTjtq0gGlT2uX3L5hJpieCZk1ZJmk1s1ex2orOvNotkx3HNk
8x6kzkxco2pYnaCLOQuSwVA58DseHFh6ZM8eTcya0o51Sj3kU5E2OST3FGw5+wc5X3gkopzQhYR+
ECphHyOb7+8641RpUV6YCvnsC2obFWr10rL0TBvapRELR8V7kcAvK+oy3EivyXMR3qYOUQRIkBab
8YDu7hZ1Po1isc9YmTWYEdsgPPM+pmCgX3sdbBCBZlrRst5lfzErs/G8gj6t8wurB7ns9hs06a+f
WHnrKXDU9cTLbFaOtqIxGD4fbr5hRFUA/aOn9gxjMfGAL/geAX+F623weratXDq3EbM3kC1Bwm/+
9e+Sct6ivaW06i4HP3FrW2szre05NpFWESfJ1fHSUE4uUw811Xci2n4M+4kIr5wHROp4N25y7/5z
Yu8s2t23JoK1BPMuyAoFcGYZhkI9LshAmpyzE+M2zA6NfrAaUWJhmFL5R3AhjicdN/aC0PSDQbi9
J+XJwiYGpfp+1eGPlSLROwmIflPHHWF3VZXmkJoWTTsz3pgqgghL2vTDQmLfWOQcyX6tv44ka9ay
K0NeFn/JO6+YOzpDpP+Op3UdNluBZUJObT46qgBOS1v70Y8wyNSs/K7MHwCtCRhPPxHIXWqGNblv
VInO3mayLPcaFTd2Xx7BK6E/vdTgMUnmgvoGVRC6PsjnRyBPib+Ywv+gx/9HDHWl++KByRLCZOZP
9saG80eJw2XjgzqilAd3pK+E+NlnrMS8Yp7nqfLWIMKT8M4+ZrkNYpD89++7rcq2U2LR+K1YHDeS
SQ2VXf3n8AODkPoKTCB/aozMHLgDlPkfpwoYnIrLF8c5wEql2UGZlFB8bdNhbjoDRbnLLldjbzjI
GukWBHskd2971q7mSjmnJYKeqBooXkM02/YFQRk3KObYbPbCJv4a+xw3x9TMIEzszDjSiXY9/JCm
Ja7wS8S2SGFccxe02TtPGccPsBcUKUjpmLIPlqxmI3RfIi4sHqndRk3KDr0mNINL8fbG7hdxSiy0
FJCcjju+RbBKSpsCvqYVMC/oI6yFsHUuJ4HeHsMaT7JTSew87nijEMBUYSKaIC7DfuJLwmOKuE9j
ph/PLil87x9oQ31NXnqLzak7nVtVQAgGTKNduDsFjoyCOTISWPWBiOH/nKoQRTV/RTmc7LFxrcYx
NVizjRJV05Asu2xErG1vhV52B3iDGzGA6odd33/aoFJWct3jqI9ao9zE4cSUIoaeRzet8YDTLsLV
ULCni5szDjxRdLFQWwicRqfH7JPoXmLGaQFmJv30rTghZTmPAdOeCrsLqZXHbJ8dXrjCRVbum7Pw
5vg6LjBWcXFjG04zn+r95xHpbMGAz3/A+/r2ZQUqzXu3oJu7wAP5gFEjE9K3C4PEXrgyxuLstqbR
W1UHZXmDpGKAFu2B60eGm4qHR0rar5Nja83PPFVVEUheoHWFxUv1cVaVfUTCZBjyCdBgEA8sDRCp
uAhPkG6yRfq04vRXB44BelrLJs8KmPvGyG0gVNUP4t3NPcRi2hzVeilmbCh8wdn8kD5pOnVQChJt
BDB9MCc1fyMAxLn5vRbA29tFUX+0sGGhUFcWewaNrwimnmaTagYrVhcrfgs2cKLsev4MUD+n0an9
mixvpOnCj5CAhQICvqIo9M5tUbQ8F4vU2L+Dblf1CG1xuroKgAn7xZpm1t5CWdy/qTHLHQV7Ywb4
8yEelsvqvr808IAbALSXk3KR4rPI86ISfITiuJq/9uoymSGXKLvsC9DSn/aouK3ajYegb1SZsOuz
6b8xWBsx/uMBWEZLvLspWVyoLrnIJTcn5UvY8gYrD8fQmTnT0iowWwKHDXpEbCEe7uTjSAvEloyJ
HPnc0OtXUKUIIe2jeHV/CCMVqj6muDwwpwzWniJkIDK/DjKgRRAn1P7helyj0heT1lT0rHq0JYWi
CcQFnLPu3a4V5aTvM/4y1cNZ6yIviUQY3dSVWAR7opH6a/g/TMVw/31o7pXNnp8mqHEXo9o/KuWS
FlWdAww2rSM0sDvQJ1R8GHkChGrFqrdQPaEq49BPpHOHaq+6jdyBgOvEW9lFCm85/FNUiAs3xbHA
5CTaQv78a9hhAblV+ESnA9Rl9R9Rf5+w39muJqsNnOgiXhIgzyvrVyiGFDA75JXeWb1i5Hnoi5lx
c/aVZRBIHKdhtYBv52d50AjNi4xz1uRjHWLbJaRIhurWcB3t6PT6VzOf558oazqGwK4VxJaksyYD
wSMFNz4gmSCQ22IeHg17Wx8X3T1v5cXwxZ3jYwC+i5Pfld6iJj5m6flOfSqw2KfGlYsf3KlNunxJ
dUVJPiuYO3DyeW7eszBriqFiu5r/kxL4kTNasawjS6WdpbkzmFky/L0C/YDZRF2FiJVYDlGE3o4s
7fhXn6549S5c4cGBfcA7fWsuf1RLSwIvQyY+HeATt5wTopV6nqz0/z3P3dlsnAARuuTReQQiMl0M
hkS9bk6M2tTEJ+8bxi4EFtyH4TpoJB7djVzqpnpdfSHpsHEt48dr9JgstRb7tT+MTOMhL2WYHFd9
QF8fOeFWLVPdeOEA7GDW0EWrti597vcLGuBmFrFbyfpJ1g53BqpFnvcQKFXaCe1mIp/I1FN2Ssep
T6w7+CqKVqMlF7wBwCrKIGp8XmsgT6/vZWtiGBV4TZ0P4pOIGh5VxAMpdnAtUr5HSCQPadLEKIrg
So5zpJroAoZAIIJ1jgei5D6+476E9Sd8xnEo30gjIuMC8HkmdGfvuo85CSPXxOkHW1/AkGIKcMLI
wNsS5GteqbIEf5A0ulLWE9zGys6hfAIY7jxwIyfnDhI+iMyaI1K1n3T5RJSd01J6CS3/lmzGBT9k
nvu9UT7tRU8yXvXSXeSSLAzCwMrxe4Z7veZ2liUDojpdEEPhh0X1vH71WVpa+oztAa2Vx9wASw2z
jQd65uiupcltuxF9ml1Yv5DcN7BUBYiGjI88SOW+c1mZoELNEw+H/T2+ndzvJS9ixvcNQ3v2pbAa
rClIgCUeBmb1Pm3oyx4clGiuOaJAHxySN62S+Gant06UHs5xonWJOZC+lG4LvajvCB9uMRNKW5Nm
SxKChgqpNz3NAaAYagwBMyY5XdzOM0wvuO0GMRe2KLoNkIEvR5Sup19/foYBVz5LedEJejCExCbY
e5QgIPPTujr7VH25WO8DjpI3wzyTuaEHcXZ9UJbepT1uNnZCeibmYKaEPfWSMJ8yzYpqqheZKW8Y
1swMKqMPTVlyYDe57NLRqYcohjaoZRs480/mgHxGi2pCaFt/lF2OWdChlShovcZ8aPJLu+Pv4dea
+cCZmVW9c3Qx+u96CgnJrimFS+PUPUEQqijHtcWWkkzaiwwSm+vL/xZlpGfQTI7XpHlfudIjHEmq
3ycRJHTzTSXi4aMVoczcY0tejt2ralHFEh2nX+NdB/+gxq5JBpiv5tWZ2l+VFN3Eu4S9pJbGwvq5
NwVY5patHY5McRbq8Vb9Ou/NZlmeSAhFz8reqcvRWtJRANPkN8I+Euuv5di4aKLoFGGl0MSazjfR
tHChnWtDnPKTX4nXPzvh0Dwdq3BTCLnqxdXs9bF2PRrt4ZfPghZ6XyMJfMPE6Eb/KLVuyaxEYNel
xWW5Zv6YahIij7vGgXZ5M7HkG8HICvckO3N6COQqni+BJnQNCx6XctF4lvpwgV29IqsFOA/X9MNM
WBprbI8prioCNLKDKA0ZGRBloaRTnXiDpE6NfSoTKO7XcoW09joewfos0GkWGhjamHMBT/n9G8Sb
k1PmqM2xur7OX9LSKzVneuZwymlbYvmO0aF/0Y38tY5LxoNQzU/MWiJ+YLsmdno02banpO0a0V5Y
rI70u+rPulnV/mQfllkIrgGeDdQfcVssqFOo40YJYARunfVitQVlJ/obN7TsOXOXCmcomuXZUvzC
7tqZgqsbduaim4VhlNh6fqBKfNQ7Q/TgP362kuMBnbYGac65PwxDjHeFOhDJRZapqI+DxV6VhzDl
iJrkOiSGY3BZTLu0AXEOrdvhMHtgsYH8xFWcliaXCzp9eWtRUcMHeF1rHh7IYWNpvHAgIbE+iGZW
unDbf4HaVe6fD3OzziFZjVqq6nDJM6I4DicChAMMO+AipWDeMvYRM2RlYKy/eEtatoNB6Tv9KNsu
JMzzjaBbHNW0lD6aSQTIr8ltWeAV2JfNIk4ASe67wKSeCgQbFG6a/3JZP2zghRUKcWYMAulCnM/3
nVbWgYgaS1w2LRXWMfUez1Q8UfAYAKB9LZnCoUW8O7GfdJxjSOb3GgwgxvQrlSwDbW3PKDNa2x1c
Wl/bMSnoyX9Ny+xW2dSNoRxarKPc7QxomudzPwHShF1Z2ggUWqGNAm7yILfIYwRF3vyicvfrhQcP
nc3esXYyee4SuFgF9MFuih5rDnxatBkD/8uyTcKZxAHyV+Q+DMlKJrPyknc2rC8ZhbV/MbYENYjN
g/YCpK/lKX/crKEnOov9wUciYCCe0a2CVJZYfmrbA2OGu+pjAJfnaP/TUBShQUHuKpxro8oq5kcN
CXtVP7ga1rGY3nErwcb0lskGsTC7PqOVVGrWnOi7S5m6siIIH3wMULyEjTRRzBuLRKYLQYNVy0hp
O9hAK0kONn0Ga1tfq4/Y663idSKk2HvLcTQEj4waeVCWprTD4AeJAEgXDR+/9JmDmPv9c4rY1S/F
QlfTGEDq3DXzpXLajJs1wGJFBCysEM2KhKZbj/17Q/RgTGfL1R71mzMta5J2x5dNr9dWe8TUsQW7
RHLiQI82b9J/vQEGnEN+MIzuQH6b4ZBWhMgCsnOX6azIzmKp1cGreRecKUSpMlWAzkRLEUgJjRZP
37uPZo5ziv2Kpk1uZZdkarGKBkh+i0LWTSHuLOmWO21rZWQjF28J/H8UM9sZGvKqkDu2rINyOezW
Q1rD8qUHUUB3rHOepX6fGHFvDe9dIK9+zE8Gb57+BPdl84tuoDSdk+7YolWZuXrDMCxNq3pDCX7D
P70SfKpZ1NVByD5/I1KOrovBHcE8d+KHryzYIhAR4HfQZ39DuMf0jhTwqIB14Aft/gpU4zqASJCr
cLuvwE3Vgy3foYdTaLPVg8jnlaqIgTfKB4ETWf6mwvddrXKxn5gom3yXhJ1F8rghUsrgScwB8ibd
ogqgBlTyQHKtf8gRL1ZwhIie0MaSzq+R7fqtSB+FX7+kxC4uC0TzPsJn1dEWVftwihBCmZW6iZ2n
J4wa5bFhstgsumD2uts3s7DRF9fFRZKK4Nqu+z6dB2acP0e7F2Ew8sXRxKafF7+gyiAYXEeZ1oZ9
FyqkvnMe9lKxFkRlPPCEeETbiH1LccgJBFcwdDv+HvTLJ6HmwTTcjaX6QAw+2zSMq0Uai7XxKl6S
QJfe9rV3BMPoiXAt3Cr2tOfkXoVfrfm+p3Tt6T+c/YzvPbxQ4H/Z/KGNoGXv7uJYcbrWVHAsUNku
0LoS5wKZva5m6/0g1oCHAasHusSwfq2D50j7gDKIVIDV1kNTtGYGY48/BaUnEgo5Dt8z+ofiVHL7
HQx+XjOODejXqSOS44bVb/ujqSjLcOmkO3rhfnrMtaWg3AHezk23EbLMiYKYDjhllEwaZUZgJiV/
xB5Cj2V0yHLrM65ZOESzyAp/NdVwzjqbP7+hb6q1CG2ZcL0K2cJuKN6XfapN2+wC24z2+kTHVbcz
Q7xMDBxQmIEiOY57sV3F0XDWeBcDXySNi7T3wIAZRDDoDWI+H0oaS1IGgWzaMjcsczWGlo1QFul/
z7e4vbvss7dE2qt+iHVMxrpsmJ1x6jjZBmMEPavinbszJ4MuGa8z5YR84sAmO3zluPBgwWp4wJ9W
3e+JWtXiAC+HWjwclpN+SVByvI/jM+yXVUSccUnd1ejZUxBr+aExgBSm+u/GxBv3zII7zvYARZDj
A4Q7MKPJHlVgeoBP5uWp+A0K8OmI43f6Va6MbS7ybHLWNKkpWwz/sZBiqate47r8jsCdwE36ebfK
mxyQ0s80k4G3XI70d+g84fPmOXadJ00WZcCp24BSo4vg003heDXKyOwXXafGMh5ClZQyzSV9rmsf
kbU/6gOENGVCBk3vmM+6nEkllj2SnwKsoFOs6aLhCqGYIyA1RHZLJ1jvbU0r/Lz9MVwwsW9Intbj
9WzuBYr2CF0P/Pl2KgsutuI3Lp3jnCDHWBywxuZfCkLfufgPb+kRkqdnFJ7s6hAiu73z4WS9FFDj
JsN4yDouGfErEbORHWKBFgUyILbqwc+2gGBY2+n2LHc3R1Hp+NvFcJ+/AFjiD+37zUvK5Dr9VWmk
pFKIQDnraWpziriWXgv9iQKT4hwCXly6gUfgHziabLZjjTme/K4fBa/pwCLc+FHsm/GzKI7G1k8D
5iLyitIxiGXryqMXtz0e5ljjgViuL5SME/ZprVt/Z5oMh5s0KqTkBgEPNn3V+eO8NTuFDoYweTa4
CRDeIvnt+WG4NxeCvIbrCzMoE9SJIyZ9oZIdniswaOUAc3zGHEsjz0EztfcKrLR2hTtMH5u0syz3
RzZMoX8f6v3XuXOMP5GhnVv720PSuD+waJ10b2omKCVUpEay/BDEj3uMBF+2oTHq/1XqU4MvWmDD
VjMfzQNrhyq+pnKANCowZLmgjuipIiC/sguZ3Jv9JIQZMnT/ObLNcem03d8NYTZs8g+cI20SeQjH
V2F8nIc2hPlIaqSVUJdSv2GzLuTI3o2hPQaHupXBp8rkKvpzgNXWb4Wj1tngc9+T9r+d63w+3gwt
Y2T2tCTk1kVlMHTkSY+IyIduH9vvX2X2b9xFX61EFMfg2NhW78KZH12HneUbt8oCyWuaadnlZDny
T1cQVRMpWQBl6hQEjY/BRgYNOiKPFC4aD8EVHSGb3+js2vdy3xrrYbdoveA7t2aqAZU3ubWZohbB
w8Ck1CcF7v0xoH7kWS+ooe4Ts5Z8o5ItwjlHj4bnXvX6Ki7ImwgDHwMw9NjtJGI0u2bcTNr0qrYz
qRXJ5ioC1mNs9hz87gA5K8Cetp01xa7fAOrShSHbr4zottQjQbKojHk2KGgnsecX1croQlzT3bG5
rUVzWPTo8dDKMWtD2PeBX07/YrqlPb21VjFXqFgZW4KDKN/+t/3KdVu9q6lahT/anmyI06LhCWWu
KWfjbeA1kCWees/EPFJcZf7VZTKJ7RxHzCXSpLdtcmDMgxQTZ51qzuW0hJBtOUllWJZXQQpYKLoa
YCVOyLe0sAVqJh/GHb42VRboCxoCh/xb0liqCZ6DKxaT/b6sw3JUxDPIE4eGAiBz50ZGkKep+Eut
QHE4+U3EJxIUXynQivMwQw1LdIS9JsifZ8R7kLct5JIzJQ4VP4Qv3ccfp8XxtZ53KUbZRpp7yID4
wNT3fOl/xV80zLFUywsf45Jc+wpuCBETB66YhEbh9VCyugHaOcdzNOj/osLgrGXi/adGyqtSJQ7+
Kt4g2aEca9cjgTUgWLclrNYV4vacKdOeSgALEYzYXOg6E+CBBPXWwzJAolLD7RczTqljgsilHN6b
k6etd6y6YjFlLSCom8l4jIjhGAOt0KDNU/7Sc0h/GEGF3OhGxmL+H+VQ8LUfdYzu5M/w2R3cpsnk
XwnzVYfgy9w6/nMJKPOVBxdnCpCrnmApXDzY7cogdVy7oFw8si1+ZAGaGu3LqbYK/5vTb/JqvrW0
XSGT5A99GJ3csWwbNOD3p9d9WgoBtYF7sWRlNKEsDCSgbRLtEJP5JMcSqz10nW0puoLMxv9kLDGh
hBrwfeA1/XkSIrdCXSTKrIBsTTCzyyAwID1X+C74ZbpT48IR9V7Kn3NHMBiBzq4SRUWkQQW2XVcI
Ngg+7vPCcd6OFkZVEM9tYuPre9VL5Vce5ZHTavGsFn0zwrcKKQCkq4q6EnXWWfM4A7/3vTgCAqy+
0sBu3zCyMryiqgBBAzjzJtreX1woc2oD0UT5XupYHthvfZcVBrP8WPVLtBU4vu6CJvtgNyf6HDoL
oYxZkE1TqO3j79FYVl7fOrtajz61Se5wLoDN0kUYOjgJG2yuPXycfQUe51rDCSmi1Ri/t54/Vjn2
SOaQxZoeFiZ3QJIlfSccQppyVzrFuTvaBuj49mS7c8RK9jAEFD5P6TpshmHiWBgZOEKG6TnV+zo7
O1GGtJGFoS6czwkGQTI5BuXL4jBVhcQp/m5McEBFa7nlJleWaDYr/nOyU/1eByVTYrkC9bPmvOyc
j+UgLCoPGtn8FWNYTImx9Eswk5tHu5tmSKV0D2m3KoP8QklTqxhVVHptHm3gLPxyyrCm0YGgqNc/
LwKy0rxJ0CnUVnxBfMGXLo2iC0tlRstPZ0HBEBhURozKZZ0sXO2kjraqnsHts+1TLSjP99VTvOoi
dkDlrXMkmz2YWmeTCLTTIYqyBRCLpWGefGUy/nnHNzTX78rPfhJRLhSU2Jt06mgb0WPzTOekVY/F
M7pPoBnyHXYXRSuyOsN26EVwyiUZAvxNu0wRCM0SYRkMBFnlVqFPGC8kBgQJ+buh94lgLb/MU+Pw
IAGXZva9RAvU/BYeFmmQb/9hoL/fWEAj/1YAzMvIHoDgx/zcoBfeU6ZnSNLZrN4BuMgjEvvBF54D
lob7eYfkma5Ez+XwfzoMufBsIPxmOT00BNrIFQDw8eyvNuFuVBASHlTpAwlApmBQD1XFQFEmSobn
SdcW+83fHVHYUaFTQTSB9mr6KOKFvTmRDM688De0BhTQLYA1OUGjiXiY0IO94TXdORcwWgDjREd6
xWliYRdQBAheibHuKHb5Zro49Ems1/rx6zDJr6vMSdIjw4ZQdWO1ISFMyucYdOFjfdU9bVP/WSHU
hTZ4n+4li8GRIal9iJHEK1tJczF4QDxk0xHosfACOahK923WdawanqgPfKL2oV8SLMMuNL1JHWbH
HQXJogjoUwi3/ENC1+dmYfRgb/0ykrkxaen+qnRiJ0Dl/ZDxXENQ8u1O5b9KYG6cN/MX6nzqpF6U
nPvwhifQ8TkCda7R6Rtrs3wT7JBl15P8Am0eAXAVpRAoG0MSNZoHnCLcXebpEaSanYbasIlYB3kN
ZbLdMjypz2AI1Yry7hC0uLLK93qPTY87T+VdrHcfO5G4wMpqLFAQldyocMBpufga10/OAc3BJKlY
cZZYni38KUKlXfwLx1NYl/0jWqfzxqdlLLA5t2NnMejR3Ctr29zsqZtOBih9q9RVxW6X4CSzOIPY
r8/hsWYc9IlNimEbTNNNNiB2mwzYf8rSl/rvdmP669fQXizNkkfearXHeRXqDTIP5wp08P4wocCv
eAJIUEMdM7q8S5DlMV/hvP1LZxlGYTcw3CnTK8ZMywp/8b/KN9k/SWzKn6fCPckVUL16pEAXd2JP
/1DIamcBwin1sB39Pzx/2+rYdN+ywME4fZFTMjo01FXMKVYa7bTM+0aqtR+fZJOpOBHNmqK2RGri
OvbB+Z8+Y1twJ2QvwgZT4DMd79UAH8jGjfiS5z2vuVlu4FHD6cxD7aiHql1xzy8q0MpVEinXgP7a
w6w7ACgtxLKL7KzaQHoZjT6KA2nUq6ycdOLR5d2kkdRB3dU0GvoE7AAZQmj3fMlp/jvBoiS1v/Es
Cvy1fytr/JKwpekbRpeZYqR+MjJ+khKNZyHv/3NkyrW/MDq7ChHvHdquXfbLylpQbRqZSk0EwgHW
utFReg47UzYnBNY680ar5oNXA1RrANvDOxNwrIKljaJsLNvXZTg6x78Yol8qQ2u9tcyj2RHFAPiu
9+5PQIuoPqM1qsuEzQwsaBVaa/zoy+kExHvDx7G68BEpEk7MxCbFTTNDVNGBQv0jgDziaafzrBC3
0ECgYUofN45IsV9FWdO2+L4o5IpotC5D20pIahU6Co5QqLTAfXcDfZWoEQCv6H1pjbY4Ui+EFKWv
4vTHE/b7uRLSCk3Ck4+kpnX8DwZJ97UdVGG2QaT2Dys6iQt43Lj1p3xs8upiOXOJbK33AEm0qqcG
9lbcAx1axPYsEquGZwSp0cnWR+i0rzAKbo1vXxFCrb16T7lvapd/dqsk4GCdxAiA3edgiCdkcfYQ
UqHZAjKGkaepHOyMLnVvLGgOyiprSarq95MFB/z1nL+008yq5tHZScw7A1BSwlvonxzKKzQpN/RN
7A9itLLkVISHRaP58+OOs/YHFoiw5cjute7dGVWzJUWPzeC187R90uasGPH5V5DbReB7gRHKsZpX
gcjAi0prcNDOpbqCkcpf7bqDGzNyPPNhD7MSPj6Xs1KnbX4mOUEP4naDls3BJ8futKR0KSmXYrGT
AmemsqLUHIwuOewrVF+DLen9lzDfVvfgJmxTy9+H4G5W7ODNkmUCfU5oD0vqpseBq+dr/57BvszX
MSpeErO2uzv4zlsSS+y+1aLt+AnBmmmzB6dITpLpP+kRFzRWUzEhA+8i9aFGnNJknO+6l4n6CtK/
1GlqxzQkFX1vtQPwHuzPEH9pL5yWW3n3JFeh5lPVFhyeykza52xEDUJ5BgWsOVr8GPp+dtmeIwgK
G9s2YYKzbH9HVrrd1z6quB9P71ry7NwhsZxWZD/+FkZZhqK2q3ql8gQpdiWlihgpky7wrx/zCEcy
Nn8sbeHOnPK36Ci022xdjk9YR4lFuqMDpl/Ki3StHeSGIBZifqsqIypMQNVDOHZXCtBOfi1yR4kv
GR4sCmCy4JIWrlU5wEdbxw5kTPGf3dyYPbFWg7P4LK4dfeKANV/R+rOSe5SqJ06MxTwEyd4WZLgN
0gWJ2S4SClUwMPk1d7gZ1umH9/yTRjEyOdn0RKZnYadXNsbKFR1wZiH+qwpQRlBaRkN4VZhiLy9u
M4Nh4XpKDx+0wpm/SmjLMDuqKbUqa0PZO9qTfDyPDdiZ1gn12QtH2PPp0pA6WMtf7N7dTZTlTwd9
u4RPjO1hHw0WLdWZRKM8vprnTuHqgbvSnHMJyHXZpiO+nB0B57s0XFVAJuHwnGrZ9Znryjw7/hm+
RqftXTdAMDZ1cySEVfc2elsqPP2ybxcyYymL+DcTw5XMnWXeoTGbaJBeMr1KFsQxTZn440fPKclA
ETwUOulgZ1u1XiJ+eG2tez16JcGz5EmfUeUk0mdCkwfiXlbI6K2zNUzLZdMw4DfhCjE9YqIL922C
q3d/9KjLdmPOPecv9J3+FSJayRonrf4MD/XlrGyBujT2YHY7FTXD90loa5a+OPr11V3wSHnic5J3
vxIahR0HsNBmt0Af9L30urWnT34+1aG8L9E997Ms/Nk0XMi9+aXBOfT2u3lsfFDDACrNcFnUxOaU
K/cFZaMX4A26z9ZD5kseF8vFAl0SYVR4sgMC5cVXv5JNng/Ne3Z53c86uNlyeR/TBZ5MfXR9IOKk
Tq0xD5wl8x9ddlkekukaDh8Z2I8Y3VDFfZaWrlZuquq/o92hARpf7SOAWH/nOAryRVRCQYJQkxkc
Kf0hAo9MHx/THRVhnXSrn9DLTFmoQCHMgUhHFK0CEDJYSLzuQj5GKX2Bym6N4DsIjYq4wKFRxIa9
271PuQf36KnAUoxTXBPRGEyaNiIn6GBefotd04o4X0m+llCqoQKT0zUdo4+JeluJ0NnbIG/sLLMo
hQ7aexvnkklduKHD6gdhvIaw3OElj3k4iRGDCyTW7ZESIGtR6tTDBsR/v7ZXLp/nIIdHLR5Fc43a
rxR6P9xSMo5ltR0sb49K68ivsnBt7WGa5pWakk0bRTl6eCej5jgO6ApMPCi81y52v54EUULmm03H
+fXjIW1DtF2qX29tGCOXhbgDUDwmjm+r2CkgvP3SLmXFC6VYykADkWqG7Sg3UbAvz8i463H8RvGR
qjZkBeZmbO2EextaWeo+s8Qe5qXzfS656r/GUSLHOwR9A5HsI6pAkeEiCtol7CoPsL13enkAXF1e
dYfxgo0j8KuCVBUkVnjHbF6ettOl29OGMYT93iTrXLvBw/DZQa2KUA1TvdFmc//dRysnwYT6rDGC
ufodscDBTN1NWqzc10wdxM2FDreocVOD/WejNKviRfidoyDTZwbdsxJIuDmcgJVh2u8OXi1jdcfi
WrrRoujIdIh27lAEmk/xi9VCbnNKsBS1fpqaPl+dFKe1N6SGF5anwwQoQY2ujj3wk/aQWeg6oIMH
nCG573OjMcyBJzjqYCCpYp5W5f8uk0Z4wpzQr1BeLnNfrmDuqkcSSzEYvrwCBgMexM2mOeRx80rf
x94mwt9KQKG/kSe5r9WkK8pW1B3SdtBypqcMHZFOBYKr6bmkuGi7H/INXo2mozxmGlIz9CRBZHwI
gzw5SvyRuTDknKnft6WtoO1NXXkkDFbSBwj96ji6UefGD1mq+Ijj/7ExXXQvsoWc+UhmjNoDkfgu
sq1HgR60f1CbRyuHhrhHX1QMOpip4Af7DeghwNo0aS/WE2vNMcKPlv6H610ZZWGMq54ORRXKi2qe
8lJS37bzLm0gaq7ItO7KRixPXpY+UUYG2ye9SuhKXCTptwBi1PHkaHQXYCAOu7z1F1NNRMKrpy8U
yP9TghRCxk/pEVat100uVdYxQjOxkTOgpNGRY2H52zW6BhdyzXgMhjDcvL7RlIW4yk8gnJp0VvOI
oliGvNG8G0rRO1owVRrxvrJQ9nq3bEnSPmlHCIhEQYgIgazPjFkmBtBrv+iSxgeDQqaeqpwIACoH
ysE6DKgNEVaRHu02Qt2W68ySIn+4J3ci1XC/OfpiiR0Dgk+CX3K2mq1cXZ1WNoEPbLiPT27aZqnw
E3RDZ/ttx6pZ2j8UYXorHhVEoCP8aRTBaoYRvRT03YNOoByY5iMsKe2FCjNEx39Tj4Zp6Omhu5gm
CDJpGw2rQrMNV2XTBK/6t+KN0p92pLV/U6VkfPSg9nYq3MO1d396VUNm+gUrEZx4DmBJUJO2mS8B
UzDXCum2syfwrx23uTuostoYw7wksqJ8XPSMKcBFCivQqPIExojSEsiU5TY1GDnRj/P3eGe/r5dy
xOS40iNa7OSPvu7ozy5rgfwk0RLHAm/xa6sATdaIXue8LpOF7suEGQ05OaQ9qbj6wL4jIEOWhHAX
snSwQDT6Ke8ryz0ZDBcL6U4HgzIR51jTgWXU6tAU5J67p/KK3o1y5kTaaeCCzjoK2nVQLqT+TD4z
XtSViprC7Rl+I/tf/oI4rNT4SZDJI293lyynbUmBeHoslx5FQ8FIo/2DNEJ6t/FswPuXGk9Ywjxd
TzseIWVhMue+boEOTSFZlHocml2H5SW4rHoEPh78vg04QfITuxlsC7B8vnrFLiVsr4sgfH7TH5F+
wcHNgZdcy9Dpvjb0QkakpxSREHmRl6QTUTtF1eMpUjXdIRCR30B0DDmL1sjecaDwipA3YUZjrivO
V7a5EtW8spxfAujz7barLMNPThOqfpJrlNYz/0nRSzgn9mOCiBwERkIBWDSHbLsUd4jW4lmDjoWX
LoDJC6VIuLmZHJbj97JOFVEBTVVbbWqUpISIAz4lFTMyhQfdAyI3GkJ5pTtle1BsHR6Jf85yfF9E
hP8rMv7BkW4ILerLhoe0CAwFYKG/5cwA/xpMrOKZdC8qhPhmZSYu0PVhCJg2Grpe4tUlOeYTiWzj
p/rOWnl0MCFswlZfpHYSI1jveTV2jVNJ6FHaoivoIUtqVgQMGPK6wtity0XjY6WZb+93vveWF6E0
+gyoJYYA02ZpnOwyXvOjLdbDl02IpRnWc980jo0E7bPla0pt2qjoyTG/DbtWO5BhdIqAevDTPR2F
Hmg5S8/fo/5ZOkGNmK0ltRjSUewuGmt5LGJkikXXgDA/vg3aJIaqrrjdp3uCIEZSXBAXkc25Gsor
U/SftPvZrX8ef6x8nANHfJVMBvlBUo+P8Z1Ha0/OXoTZOqZgwOuHvDr43psZQlOJoiRbkM3jarJG
Pnc6FxLikZUudC9GN9bxuDtqzCgzQ44WGpwkLiMYSGtfDgxSuMLzxbFp6YMoc6YG1vW7fjFm4lJX
j3nxBO1EWk1UR1fIFC4FwSQXUJDDU0Bz+N1PGfOJ3+K5T7r7IvfhMa9d9dBWxGGXOjxKv+TBHZSD
qARoU+MC8GsiZfyq4AG1MeFT9rkVpTGp0UTVGaE+c8cQMm1/cxDiz6N17EZc+L01DphhPszLfHJO
9Pw6UNdVSArwxa1IomXyht/4v083hyJnYpVfSLULfLkRO6KAvXkW0C8YeeXL/zh9humOaYNMhpdf
/dgxewQdyndtEAgyzCEy8HuisBS3BbCmAsnfakHER+lhdoMd6n5WY96KPizhCAaOLnyR2T/5GfmS
9RJJFPXMkwJW6dPxihlhcdtx0rYOQU1DslXVBuEarvfhpBDCv4nKLoNmLfI274ciByuJWTn2yZOi
eXhrKJMTLpxYaNIu7Bq0CylhRl+WuEE2UDWlX1cHow+l65tPR1L1y4e2ImLsifehdRu0/EwUsp7s
HNv1Ri+DtoVbpNdIbbj1rMPUbJi15vrtrm7WD0F+20FiQguCjanttxxNwSewMFHcamHB8+NwHdhJ
+3VQYzPMLLE8np1FJ+Q4+Ry9gpi2sNnAP4GQYU2Ao2KdTn/jA8WRlb0qinPJUgryFbA8HGFvbXib
hg/nRgcvp5Ses9YQF3gOJX/URr/oXRZszFIyjGvx27stTMMrMoY5MTRgCOc6A7Mf+3mT8PBFvKRq
TdfGNpVGS3MXgdnx+GeQxKiLC16Tq0cf8RjT5kfUw+iHd07IyQct8ebYXhEGau/ZxZZDaDEsfzJm
pZEgXMOZzDZcVxDFjdTRpF7tb3vbvBN2sTuck55wSz8r4vKKagXnrKdZh1WjZJCH67kmAHiP/Sst
5c9dTx1Ti3IiwqJ7VcNRv42i+xIgfk99ycqmCpJA4ucxzKUgT4NbGgCKRg7Ja89z0jsNET8GZ2hX
08I/a4sND/8qk/3BL2qa4A050ZHl6slnmXoXgLS7OwoqBbJ0ODoCj49cne1hghrgPQF82c6LHWJj
6/95wMFWZO47hwcXac0kiFvX6oFYED7P6xM/Qlv7m3359GAxVNUc6UdrJJFUqcUy54DOgV9gR1NL
9WaFqVkHp9E7iDGSQdWHF0E08jwAbeIfzru2yCDf1gh5zArpHrCLYOpa1JEr5pyscyjJFcm3JAOW
7OsgcZM2LcgWEgDtCf3S9TlkGaJoIzK5/O4jDRGuADpFpfNyqLFa9EVu7d35F2q1wfvbaUyM/gDp
Eiivplz31gK4zswSxpEn/YMCX2x6DhCw7ASYi68InFFDTLWvzyU4Ve7KDR+Rylnhg6f5Q5dhlTL2
coIYizIy7+GRNvpsC0gS51wnPgPRNi8/lRkhliIBwrA70t8VYstyQkYdeqrMwV04p8RVEYawaR9V
bKOEddMfoUYBFypp+zyjJQ8FbfOVr8JugY56jLzKDD3sPHjeEY8hLxgB5a2L3rm00Qzd1dqfEtO3
BN7V/JRLCC51WrVpQdRzeekMtz7z7IFh8rUNkXvLZ9heJdxvWiOzRMllmebjR2Skh6R0ns4b9cSX
vOZYJIftlo4HYxJcttsN/F7M1NdsTZNmvfcjW1lys246G1cidZ4BdQBTUaAy8oG++uR/Mp3rwXRK
zxqN6cKevNF9cUM3VoQySZw342W8vaVQGHOz2gwPn+Igw7ryOcoZ8RfPgRvRSfwYp72NAhKAzRBx
cN11MtbAXt79n0QizG48TywqjCv00btYw7MYMC92dSUo1nkiAGfv+kRNt/RpR8t0pmxR6rVntQIY
8EluW7nfdQuqI5ItzwMIOEfBDTFm/fNXlrg4+rAxYUnp4+nANFrvTnt8IuUUYi1T3UOBzjxIThRk
MThyakrOCTW8rRywJxR9Z86W/QxNz3VkDeP0EE7gNSDyobMGHfhbfM6k6lfQJ4IKeAV2NemKkGqg
25lAlH+kqbzZYH48NrJYMHCDO5czJ2gfENiE6GXs8jGNztPmm0yxqKhvf2UTym8g4Oc5kvlWGFYk
sPQ7lDnvIh8Xka2NYnlcvqTRjjKFCeq5nOZS/OCLc+vEfUCUDFYlZSP0hjuZVDuURAhUv3Mbrj4/
eaLQvnell5QgYTFxcMxGeY11JfXfdhjS+Ne/Bp7a7L3zB1kuaWzKu9G/c3MUnnMTh7MFqeYR1tJy
Hh3mpglkxOkcKIwMuuQP35/dmOGQpMU6tH3gx8Ky18N0Ljp3VL5LOOWdiJW0DZzIo+wnuFL0hOIx
65Fq5YkvpOpUWIP6TaZgbTpu9eJhkjZtllTfvlAG/plDVo4OqOtw/WbAhZhbWz5prDz4z122lCcD
gVSiEPOeUn/VhIAlG4kf3py+KMruSmDKxjln4hi7LPOWeWqkwuq9hKqauNrP3mfT74qGvViEOWfv
urBG9CeHPdq1j22plcdCErGE0zDmv3unJUoqvNh8BgdjoQEopq3L05OWdos0uyVn/MA0Y/1zXYoJ
Kc4U62bYZ16elExQVcldbLnhmmmHm89a0VHKN+2pDl0cSNyryMzE301VxDSu37MCEc9/9rBCG3LE
y2MF4n3X/BkROsAXYG32WMfxuq+kbMB7Dl5yhu5aTg7OyBJmJ42YWbrKKrLhRTo1k/bYujH2pPt9
+CQTlnKZ6LklN67GWhwgO+p56I7WaAzrd5LSIv5j7LKISoLe3lpbLNtf95zRpPrRYBGERmPpRILH
W2TPTEEY/ip+7ggElzAc4RJpic/2OCcB7jY71U3uXVQudE00/fXBl+bqzc1pyus+4W5kM/9vTSHo
KtDQpSy2+WnlThriEzRsyhuWSpMZAkbK5rkDwEwJRmLpaHsNkYRXNaP4c2iMXSyEBeh83pk1PJww
sWoULnqzf3LLwHoBUlX5elCWJgPALZcp6xRUGqroOMPqibPMxpqtv5x3xHNWvttxVMEVdIIWP73Z
x//TxINmAwLgJKJhU19p4hLsBfcixcmiL66vyu44OhhC0rKmzeNohblNlIM197PnTKkrvNZJZL8i
M2tkvvNHgYxmLmYN8tMGYJUtVW/2hEQ5CnpbErnHEDaV5hSnsXu7EuNP8PeYPexk9wyHWK2+xJzq
Z3Cym0C9u1VIUPkS2j3cdgkwTrIhckqKZ9p0D96VObsMcR2P3l7T6zdNVdIsM+uHRw2mnRnUIcNq
gshe06gwHtnlfNC8gQ+1yj50Dy67daUgalPmIGaKSOrQSpBzDVkhTZvhT3Wucv6v8Dvoc1L+t/9N
z+dopfoul01vH3uinbDp/JdJApHDSnKpfrockQwZ9MvNy4zofwq1MPHOmErOZXCLIOYnoEWQPHMY
F9feXNQJXUoabhfMPvvP6KT1t1+uefpweeCQaPH4odC+aRfTue9+sAXt3RHRiqKBVG6XsaklyTlX
YcbX/nQDUhs30z2N1opyO+7WqLYkSaAB8Kg9Z2FgS9dpiUgyMTFsxr2d36vGm6No7nPYQEHmxe2o
HSvJWTknOemCCRplKWJcUgsF+FNpXzGImSrsPR5zcPV2eWdF2IpVEUDVimv6LJqCrxm62PdgTxmg
+D7RPlp+FyNwq3pl7KbnYRBOtyelFGf8atQ5eWtnVqZnT691zwtuq0hC4QOM9OM50sh7UxN+IfNk
FCJSLb7EsXmSF7k/kchAalngaVxcx8GusaczSA2/vTRt0eCndfYC3RWSFx2sYMs9Qfqib6LAi69n
U+Hx3XesKZenot+GK73FNGzEcTKr3UKP3oMB9CnR39GBiGFoOighAl2EnIYd+rAsP/wIVuJvs8KR
qpIwxueXu9vJ/55CgIQFFBqv/apHC8znfHSzptWET+7JgMAfJKXkgqVZerzk36ZX97/fCJLWNMDn
ybLna/0PYldPK+J8u3DljBItmN1v7a1kRaaZwzdFuvUuGw+7PTSNq0x537YNPViq9edU4kMRu3vY
4PNMS40PW02tV6SNomf8R3CkR8qyoQ5gWddO7c00SCIZa6GaYxs4joegku8CxrYGcn25dtFgvHjC
CTr7gIDjfI8J8+dtIAEkzq9d++GA45sjgLu9+IHCqqMEkuY1HudTEE9lxPBvgQA5Mc1JHf4+bvAg
x1kxjGzt1s/+hbrqoaKA/HGcbu5bnfELZis87kGTuhNbqrHu9OPtQJq108A7dIPu7lu5jLs0+9GB
1Qpy4S5l+3kzPM1V+reBdj9Q5MN0JQQy7AY1nGYIqT7DYRJPmKNlbNGqERIdKnYuLp1DTjHWX0w0
RalPQGr2u2yed2ga1D/v/fwwHF5/BWivMFUd8EWihQemvLI/RbVF+tTdkyXUGK6qEILeHPYCGESk
eGyfp1CEIWtPIWhpWJlk4YeK+PdmHmLL/mhRTk8GMXItR8cXfLaid28axmUAGFEKSG7htS+ZtU9m
gwvE5CuEnhBGN5s55+sy4RV/T8QU9TghGNxNREP/P/gIYup3hdtWd3w+7GWrKv3xqAUkc/1o26eW
68V5Hz0VlbtiAV02IPeyXqgMJqq9u4lDaKxw5Ml6suRatzoaIuqzCBgCmUzsUkxDhDRBUHYAI3fM
ZyHfjcC86HdDEn3WX5POKnmBN87VBRNQUuQttxLofeYPLruifkkeiWvfhPwTZlJRBZ9SdETwBb57
bgQy/V+yxdiHB3lGK+EJMatnC2mLILT4G22jve8aqm5EpAOO2KX0OirHto82IZ5I4Y9fINI8AdXy
qhhj2kFi0bfLgPjkuGTsFdn8rR8UibYRwl7nYKIjgoGTWLtBRVdEHqMAtcq37Xn9Q08Eqy6f8Kxp
dkOuROBmjQmGtDR+jXUVpTWflhrj1KsS4fW/rF1ToofT+npTlPoLf/w2bbNKF+pmPnzZ1RkyohMr
TuE3SFK7v27Plu1e+MbQPvgrI7agXOXFINLbgcCufxpaUkHMFYUnkr9OISusbn41zmhk70ur/wvd
TFM2X6+c0ywG+f9a9HW7OXZEEAprc0Gps93NHeBgdAIbEZqN8n1iZL6aBlOk6Xijcb2TPhtR+3YI
HQ9eFPlpugmReIzUOYk8cJmO2tgqlrEo2fzkIMWFqAZ2uMbLcieWxjBcge8RNIoVXgO8Y/t2cPjI
hIybos4BBWeTZnXJfi7Rqhynf9AT2cdfDmn/3eHpeEDqSdcZS4OeYVlgcj9NBhrog60X4wMa0g1T
0HMhbh7r0I+zW8Xo3MYSRj/vIsCYtRQI+n6SEfZgMrMwXbnNXBH0gbG4RkFUHnrxcIQNCfcCg1wc
s+EZNENQTX/4XP6FIqvfKdUrRJya3lO8zR7OFhz1s/SyFkCr3F2EWUudOGvYBgD/x7X89gJDLOJK
gwhZinD+31GR2IO6G6AMy1yP2c5sion8HnSSIJvq9O7jzlyePCuFbHtQLxlVsntL6yNk5DtrCVNG
854bc4i+3xaihXa+dqYq1MC4B8dgNNVs8vcP9/DYxapqVjcxxdBUTJDg5vXJKFlmQgJcNtGO6EY8
rZnMzEtJ/nHwljRzJOa27cNpEttZbMQQUhjlX9EqOc/8wr/ezAn2PThWM9xMeoS87wCHaTkkMIjZ
4qiZo3V9GvHURAWy0a19qvvLHurSj/Un3vNbwZd+9iwfBCw1IWaPMsRCOPeP1s2Y50yzcqXhQo27
K9XlQm5kmrJ2PmyxJ16xSQqht1JOeLh7s7/XzH/GXU8MiD54krnw2PH6Ae78Bwqu/Yh4uccQCmw0
cBJ0e0pfVvqiUqZlpJ17OJElaPhuv6BXXyQzT9Chdw2ukHvajupquoxqaoHubnZGJieY+gEzXz1Y
hXnJqMqJ2szQyGOgNxKNdJTYjXhUVlVasMTsgdP91y6JRafC6l5SCZr2+EfrtCWZduWggIWIbu8J
zugOeS4FGkV06V52UNjDl1uGNIoGdv8Ka8IfojQCyzuOd0OshOwdKD4efxPb6D18zmGrhPeEjrpK
h6tjNk/1G3oPM1zxRWdvaxa/KsEdVEqZ3kOAco14Zi3uxb8U56rI0VOWzem0V1hSxsOySewZXSwH
+GsDXJA7u7M2RNeSGb0N+hVgX+QvULATcC41M7dJsiS4VhLmpqiBNv6yvjodXtdZJ8oVJuN31/sg
wX5ckb6ORNE2+w13crWNhNGjn71DfWT/TBlHcJ266V7UWgUbwei8/nss1F3oWZUHhKp8zQvUQ2Lb
S0o6PZzNfa8H0Rr6wmCN/HVAc5GdWxSsH2bd9htLj3BEyBJ7eQBBCGpa3iYAK7j5BPa4uiB4Rd0K
PxVqqginWmF991CxEjsB0B8AQRA5qnEXkJo4BPtGF4BLju/DdxKTGT4twNro3BDrjCtAUflc/I2X
MRS+IHIxz+eHxLLWwylC22vQDNpFodSfxd/3DogZ26qgtmb3A5Ug+pHMl9UCZmhwdh9SamOPnyqk
ZeeFPd6qGEBndIceenro51ctBeyFJVJfhPSpcoCBRAq3Zf+S+cLLf77XRYlM7EDwmngYYsluwIHR
9yFyioSZvgDF9crgF1emRg02hLJuNah+ljzbvbJp0v8iH46KNbsP549nNyx18JdUJuqSfVVTLHNx
umhihZmhZ3zjVr3fmoN0AwnWJld/765JfFQyR6ZTBroy22i5hTB4ha9EktlOWQdLH6LYRRLtcpz9
YeiDBBHN+sXyotHPdIdAGf3ym6M0YPYfDyP5dirVkl7PYy8+Qjfir1wOs3rswtAsVkLUTx+6egTR
WzqkjcTsAmPPVzeIlOxsYNwdbT9vsQ7kMUVgFpD2l7nfhKNw9yeD9abAn2NImAfLMF5iypDuTuc0
cF7nQPgClgEaXqMZ1cQwOh5J+4igjm7Dw2rFpFMpjfM6XfkEXA0ujjQrl35tjfQ9D/Z4Rgb9WSbR
L7YEcNLx1TEUlzLC8uluqmVih17vR4rCMzCpUMJHJRMA+14n6LbcgMYl5EghvwoFSGYWw+y1QpIz
g93PNDG182YhsU1gjmngsGIGyXLvlKWFw6QeFXrqaXJpCky5BIlNx2mHU2ZmXaGNf7yeAIjD5KV6
b75CNAEq0Ld/HmsDrfukylq5l6XEX0pv6N+wYuHcbU8IOxPz8cl68diHdp+vfWByTs/Pe8rAq54v
id/q56Y9Lrgopc8kXCFO+VUpK3jEJ0YbvnU5JBdjgk6KBgWWh8atpLKe7nALiN7fCA4oUVsumZu0
hEG7YRykvUzxhW9G74+TY853shAaNBm90/hi93tirrO1lwjIZJxI4reCmsoCiam4L1fQKOeqhThD
NgygOqelwFSZWuPuf08ueva6ZZcurxtxt+1r0ISuohP98vsvFyKJSWzPrYXM8Puia25Q/N24j+fs
QBjYZwIjq5tVnUvdNQt8GvwIFxnIsoF47toTsLC6eQTFQVeIB6/13mSkPd6UKt4F9VPPxVav78ke
KfGJ/OSuPzjqnQ+EgC9SAiRfR/D2PjYCZiMyKhCMd89D0vLNM3seiSn2BCWI0UP9/lqV0w41aAfr
r+sur1t5qEhsQAQwCoFPyqvVYtQUX8X3YKaWTU2/n4mWptUDXv49i0M3vJFVmsuWYF+31yZaXV3m
Gugpc3lHLgW1vhDSsU2PBWM/hk0EeRnoRvnKOd8GPiE+BTouBzHkYE6wzjtuZFtrOjsswVkwFZ4k
ryuEoisSEMIl/qaFbLzUZZMxb8rSHxLvLPNW4XuN5fwI6CQ8qqLr0/DC8Qz7gkbIP9qGnvsNpsZn
qv9o4IsiG3am9bQae7mLxRCkN1GlThc8Yu+22JWaGgAT7FDFGukSKU/N8HRych24IXJ1AO7ZYkqI
dg5bst7FhkAD1XcWOKhiCgMDs9hM+Rj3WWm2bTqJCVb6Kl555QH3TteGflgr09M6mb8nmlNYOrAr
f5yGNnCFlVrB5YCBoM4xruPSqUfeH3Kase1LywUrjeKfQB5Tnh9J4K8Gv2noNzyPnNRceZqmUaIF
numrlExPK94bxd4iv0ABYzYcgpYjJ8KStbxdJkVrbSC/3Q7L0LAaRDYoJpl8I/2lcbvaombpPfxx
j88bjhAApSqE1RNdxhH4pTud1U0sU6paveqceHl7SVkG+frsuPFgvyV0o6LAwicHJYX3jU2X6Rj4
WVsylYDPs8cFWLINaz4RHnk538ociaEkBMJYVmoVZfYOqdEwu8RFTgTVUjkKRTNCDlOgF754Db44
c+/32MCXJVrV5cBKNjWFUz2jd9jIvqaO60Pb1GsiwZQwIXH7vQgIta2e4uU4ohCS8/EQulEJxBa1
9hQX9kpj7oTgfsUgib3hX15RU8VgrTiEfY38m5T1PGL657EC/SHON+/jICJdLDlst2AP5mTQMKn1
he3p0lo4CRKKam6DUOk8X5UExplC8tg8pqjy1l79ZiOJBoH5LiGfncAHG7B4VRlzcS44yj+2TOlT
XB5hC6oiPtHvNw9dTToVV9HBjuLQgcQqYz+AfYbltcE1L/sDm4zZFZK3yM4TB+TpU/voOYeV4wrX
hlg0DlqoSJYdR+UYVBEmMMHlPKeKUayzdyGbTpZrxNwcQ04BSlDUsAvuBG0wIbax3/JlGKjihk+k
8AkYGT2z/UAoBlM80ONC8UuTYMisPbeNTvhINmpMd4JghmxbcK3iqqwrfQ/UIq7TeNHILcykdPly
5hZcu/z81vR4jQFzkSFWW/r2UQjHprl5X6qX/fvUOIi4kaU60Uq5ao+Qn2yZhUytIXYyPL1UQyTV
RkL8exesmokjvecdEzj2Y38czbvhIKRBHXm1+GeLorfxa/n9/Y1zrzj12XXuEOWOkqMO18f8bpBM
f6lHgjRDrqyu/9GbZg37BYP8tZi6vMfXOpJ0muoPzm6iFThrnEp1rc2U+Ny+yPlpk0h9hycN9qtt
SYpDU6+Eg2tqA1wWj88Zd5xzqsmocV52Z1SvUMdWSrFvjJZ1wZMA9Ftz6rF6T+yt8W+GDj0N+6uJ
DtxEszi0yvPfrerx+OFBvH/D8C/EV5aH9EvHFjdKSGhha+5fZwLSJTkjYCEvpm7WR4kSO0rTZMY1
TgTqMUv8dZSo3no+8Z98Pff+v/ijiJbVVNC54DAHrIAhaMveTRHDfh3U8LbIx70cfLkSM2n2s+pF
/PgLoJvPFHgOI3hJ6KOBo1yrzLnlfkmwR42iB8MJPWNy8CzEwBMYK+U0VPkbWMifgsWigLTFEE10
k9CaT+N30zWJaw4vZbDlqA8viJtfsaGz8l1NTL5GirKVUHxEZbGf/QFzZJjbu3+T+ZqfQ5Pclmur
gxutuq8byJtukketEycT64AHTPXsX8RKpcghIHBAdAPQAXJcDE+dThQR19bpg/0MzD/sQe2k0Xz5
8G03e1oZ3hXh41fN5aZsELKWEgaz8Zz0K7GhSUfS99/nsF2KAPc+AE8ueh+cOfVhRFSDudRJTLem
torX+vY7adrwboH5G2NIS8ata3b8XqxG4hTGXmXesCH2HMcGDJMIseGceMITUIdDeXUsDHdgvkwk
WtRECcUAI6reHnU/nrwPGfN86eP6BFR+/VntrOHPw4bKYXcFyYGl52U6AyGrwNRydQn83xtrczJs
lJ0QelqmceIJRNMAb5DGxDH5Ia0lSuNVsDwl3DGvdpTkpHVQCCVhmn03+GGN/F7hhJMGytOuo+Ro
rEwXY4zGwDHGVHCgQF29mDVPm05HfkXIt198px1KsxnskzyKdFCGqb8cthCquTJLq0EUxjpSaI80
1eV/H5KX1FpwzXFaFBUECV7+ieRiKtSpp6ztS0g3omXaK7AEWaUTjBI+pLP3FRnomgrcQkb1xE7y
bBWHrKZn09keGM5NmLxd2T4QYeci+XFi5y8lASz4ugYne1nckXtrOoj5Nrr9ar0rsnuL0wEPDCT6
V8dW3sCnetZNact+3t5TquogfO+HaWVhgZ2w21jTkNjHCh6TJQ5AlHNMYv6MUKejsfwU5shGEt1W
67gEuYsRLqyHr6JG5DUofFmFqsWD167Mgf0RkpjDO+Eact+bAJM8Fw5li075bCQCPDhY1yUaAEyG
Tkf3gLHutJn9Tn8umjGkkg28efq/AJngHBHDaz9qowsQMxBVahJtaAsU2/3mPoJCIdvktjr6llJ4
1FtCRBknoe9IPCsDI9z2t+JIlcEMXUtUg8/raG5DpImSjCBZo+VfCIHTq1COyT9gXs80yskKxJx6
snpyzrrQHADrrb1zdfIBuPbOBrQeQpyQGxaHTQ6x3SAfkD6HI1sdd2rfeWfLh2dxZthRJksKP9HA
DT3gnchdDNDNjgScTnvWeLFRg8dbR5WoBR5RJN6MptRPjYMJW7bH2diCdO1ig6w1HQU/QwctJ3Rr
AnOQNBumAqO/IiVLcIgHfiGDh9kao/tpvCNBC+J/J5WAe7h2EQr+FMPNJK0/bSKim8RPm9tsLDH/
pUAAsLzDdPDpxff2NYdejfsr8CaWUT3e92GjIQ3MfqZJ0bEIkuqzqcqTSbhUYg5++sy86bQxp3jA
pjD3g5+aPA3bnYadcGagcgoLu0vYYufgdbTNvCKwSguzcZ1TmguHk4Bi92g+e4MtUMniSnipFTfs
uIS4+wHZ1ScABwOSAmigyC+jGcCrEqHTEGKUKQuFs96YzMom4+oO/hKUUdkKSW34DN5M7aksZ7za
5vie1TDM2g4FppKPZPmkWUDwzaOBsHxtkPmjlQwRlxN/iTiC9h8veE39ZGKiB4TEWUER/djo68RO
lMLDVlytrVk1sfnHRaHxqS01E+LChqoJ9B1z2GxzYd2QZ3w+/cGiFRcNARsJaUS6+dFsUiPTA4I0
eeQV5yHB7Ij+qLcdgKbe2A4AMRmAMOp4o7xtxHsqclhocev1/ID4JrAXv8CzUH4Y/1grjJbo3bVL
l7z82iFID3Wu5d1bDTXNb9MlgdEBimu7Q0nQn7bxvXzblX4hlorKj8pw5XmxrKLoyboYqjz5YhYC
jvVCdH7MFaEZS1tZDIlMnQmMPbBbL4kbm/lwnO5HKgmaN+90ELMoHyajjNQdJsMCmVouuYQGijMN
Ry2L681rKhIu1jF9xtl4yrGX3a/jOMRyJ1rXnyt+xZBAsyUasEYXjnzm+XJ65/p91HdVVt3MoPKx
YV+TOBAesIzW16S2jMrSdt0gbDkT0Mh5JshGj1CP5RSj8JvaJFXRTjWDINjJcBXq3Da7YcB8Mb2D
xu4L2O3aivtAwcpLIjYa7XNhcnYnuKUx2gDJcOQUu7CyKNDmyeCyofeYbTh6iFPhd8aNIpd0ScXf
GU8WAoCUOWHZWxj6C32cdZXuQixtsGuLjxsgQjta5fIv2HD8aFRmaMvJImXhMTn0HdZlHOZ0jfty
4vNqi4DfGDVdQEKhkpjoJ8zpSEyJkgrW6acH/0aOVf4seOQAOGbJsrcxvN65xXeuigA7wnr87Vsr
HWeNmYGfXMdmZwaZbRIB8RTCVs/gJhvhJbhy86hzxdpeIt1IbFtmNloymay3Ya6TE/rhusKqlLbT
oo5IaPwwv9Nt7ZqIU0YDbopgrK+2DqyYrdxEVcG5dhuNFbcHUcbDJAtTEnCipnRZIpCy9XTeaFzJ
oE5yAzsk/LM4YjLncqa3DN0h3PT263AEYtQ2EXhxhA93et39p0E9GGtxHkvZrI//n7e72jVwLQm4
tNiLHOcq/hxvMivTq7UQaaqCnrtWjrpa8Aj5BW6nqWNzBkOA/8Y0WKlvsr/gTqYtYuZ0Dyei8qt2
W8K9cDNBbTjaGx4f61fGC4PoPOCmOvSqypHaQH1wkAgXrLTlJdNg27ocFb50JIRTUYX7pK+GPa1u
4gQAQFSEEiBPD1fb+eWmlXiBRUnTNf6R6Lv+Dewm/fVjUq5uTpldLk+p92VbwPXn71nsKeH9FBUg
143QG5IwllN5i8O4Ox/6lffQC+aejhk+V6aIRuGusrAo+isrbDgOlO1+jEcoByj0dF0gUIIiFJR7
6qltri8nsKSOw4Z7+W2j3pz1HmoWYce5eVf1oRT2qqkOj8k6pLzXk05jfzG0dy1EHdHqaPJQnSGu
icU1oAj+kSuj34NhYgYNWrW9eUU9wx4fxWU+HDjkEZt4JKtpxSDFLbO3pK2uiNzTWLImC3CNUEZF
T3oPaORLl/KaheBB56h7XwrF8SUbK3ErjEKnbCMJwVKXzWXExYSC80RumcCUpBzOFQKy/+qQty7O
dZwLMPnt1H0YpvZkhf5/cpOcaKEBUNJcWO0FVO1o3//cGtrUY53i3JWRKYQQR0La1QPboIm+d81a
g10FUV4GQdUzk7Y2NebOOeqB/KgTnUUFjaGl1JaCeOR/IGvmwc9uC0SBDsQKKTe3W9d5PKb5uGek
+7uobxXmGFqiA+8Pkvc3Q8mwcGEJN5RJD3qrX+OKOhaSSUbfX89fBxbVckN37ZmjnvrgJrTwMU8b
2aiOLkjBikjZZIDqZcwbs3XUqWHAZ9sCQlMgZWY+2v0k790w3tBBKsN/A5FKyeowb8Yc6wnArEh0
G/40mRHjpPUBP2nSuGpbzR1XaIpiK4opGMAc+66Q/OREwScFKWDLfGHUoz4x41a0V5ZiV/VzDEfS
cCEclDAaax6DrSl9W4CYch/OqHgAYNlANBY9gkxbC4NGE9I/OrJpkITulSwzYwoEdiThOWSe40wQ
RAymfJpOGNOC4Jl7inMqiYl1W69cdvPytbtTdwZvVOxkZEIMNaALrnNEHWfviw6PAeAnYMxLt38M
D3hJkLKQZJ19YSaPrHtwcNDEYwJ+jMCAF42wC7sKawohg4MvOrxxk7eMyoIX94LosjMnyiMYlTh7
Kd4/SKlmi+2pX73Q6ggXqKy5YNdqgvQPVsw3OeNfyHqGPY/o4rqmlfuhHZTEn0RJjHEAPCQaMlXm
MUr9SqDQPMJ1AMoJy1G98NMgV+rrLjTNBQpIjeieC/k6EY6REc3ZjGRnFDnSjW4Ldiz3DTTX/g1f
6hcMUwSfGMkyGrnD8IdpyhZkJBNPE8+79I6F76K4NxsiBH1cp63MSrfxq9Ka0DPutT2z5WWPxZW6
vdrpQEY5XG0AecjSshGIljLzTWMpVN7rjwy84ikH1VChG7NBy/uJJnw86hd7pCZ+iblFCsmmrWrG
82J2qAzZ45xEMimBfghz4qvTC/dAlJoFbMpXn67mKvFBVGKvEYe1B+wbXvEA2JDV6AJn9SQaRanl
KtyFq6qiLK6mdUJvE1EnahLSOhQcMVt/xGZeYAAHfrjRzO7iF0/XbucojaV5/xdKBENqfcPjz3lO
1k+o653l0UxVyEMeeBx6Ae/CL/jAY77IPEjnplomoVFdBeCualX3cMvSWGliDLRFFdVlhaFvwV3F
qmtNTbVx7hur0MghA/Q2j/PIcWDxWZ8D/3153Kxe/lnwOLAyVGr/nYosjrKW+1NwKhESbUC22cmy
PAhQEkviYhVcOCkg5stZgm8PVRmFhJEfUg9uy0quEx965D05ApsIItWppXit+PIuo2shdgUDxIe3
65Mri1kzvAGNPflRss6CZYXVIBGcrSx3xk3rDHMg3+1qqzeYZFg2xfQu5YGhifIkzt8z9K+syPvk
IUMvKPVe+gOipKIvqx4++hOrom0z7ZskH0nMBLL4G+5jDvnTJo02vU691cqvzBDUQyJpGvetWdF3
NeAxAHnHIm86559nlXPt0gn9OWUNEFVl+ZLOtYikvRBhQIxAmM+AvUdW45HA8CxvkvP/33bqC9bE
EGeYkuzG60XAuHktI94hfwOTTU9ZZFFIbQJ8SaqXsdzAI/gZpqvPzqIN7zBnB3L/t2MEAZ1R3eB6
x6FISV0bcsJxa/Ud5SKYjQiXtELxqyNcaQ+kTSw9KLi2rDLTaKuOS8MoDGCeiOoArdFD4kEP5eC/
9MY1TvTaADKFyspIEmcU228xLGuugFe+IrFgu2m6uXpx9dJh1HG/+OaeTjnI1IhwXo+6mSczoM5D
23pw7L/YIolv8D5AaHW6wQUUeszkdHEO799q8RVFaV4v2+zq2bqWBfuPZ5Vip7cgAy/SCg+FcC8/
avc4RBRzFBYZ7PMh4N4goY0cKg5Gm0J48PWaNv9Bpx0ivalcKFzBXTQcbfUwrridSv1cc3qg4ZoK
mTST6jlS7DEGGbSJ2PLj11kFHsb57jTo2I8+X9PxKByWywOuwnSzNV/w/QJUt35euKlOZkMF1GsB
EU+QQvGBRN9DwYlHYXBN+djQhfx70eFqFHlJXg6PkRF7Y1BmYskH4hQki0sTGcJFMwgtAYKCjOUQ
UMWLpDFbIEqj/YeUygVUkc2Tm/731M8wBJpzv/XyAfjs7ifCfVGxQPxdzD0ZKTxCQEMcZSn9a1yr
X/5AspHx+mKBH7sTyRUTcI56b9JLmbUgp7VX+zbCB60TMVYEqoS4ako56ixNlrf+1/80niJ44vWH
ny04jTl8VhXJaXsvpAV4tCGh7rf4TGlRAzw5R0eGzTdJSgSEqZJ4/bptr9Ih3qXMPkKjuqWWY/ZR
rGimu3PztPbb0G2GV3aeg4D/PQ7LXPA1W9ofyBwBqL+CSabpMeCWPlNg7B0u7+P/3cGEl1WCC9DF
AOYXkNBJ/IbeEnSyxTIOL7m3NiInWOFw3sqxK6eIBIUkmryhAqvR24/JbNnMcQZrH/NmhvbPyvSa
R9WXkDfuoCYxSiR02nYxCEK6KG7UGUHRMon50gNwipZdQWcpXq1+wdK6jx/rOxNpOhs31T1YsOqy
nF3jsubcm4sV34o44p6++oxe7yAgzmWkAo0bBnkTCIuYYQ47RilOuEZdPC/Mruq3kYkRy02aMMHd
Nxc33vcYhZls/WhGkxpYKBUpJxy/QnckRyKnCUrwsWL6BN/BvkkXhOtwfn9O4CRku/UajlFqJnMW
rxqy2HiJlrYgEjtSd37vFvmluSiTuC7DnYAqZiapa5RNAdCWizWvLt1xWeytTZl0nNOsUe6ObyiJ
QYHMA6vrWc0wP184NwGD6riqLXr39tCsCmB6zfn8oSGQTDinmyuY/jAdo6/37XvF0lnzfBALTqfd
mX1nbDOL18INP+vYC8b1wkqKVcfkFvjYXqnZPJFosqDBm5zd9QS22XVSx4ITPkVRPZ0AciIhUNEN
B5JXtUHqINdJr7XsLzxfd0UXN+B/vj/P4Y2u6h0iBkACT5kcXbMU/iHdjKpflGdUDIm9wi6kAi5p
/xyigMYeE87ZCzUMhGTsIbRBr/L1SSRw9rR7hMs1furjwiYGv/P5t6C89WT0kiFyTIKPYM1MmvJf
7bX9mx5WTCt9c0DHgntash1QgREyV8qV6YeIsmEAE7mopO6ngncOonIsN2vhEDNyt7PJtNwEJfjm
YfYJyNcgyHDFngv3SXNTUxSfTvr/SN5gbhket4JgIbqXV1sno3pdmwifdG7kY/G0vDe/fyGQO1sb
i8SK72o/DsTqS6q4HEedkIT87/Q07E30JOjj3q2fsEcGD3LJDiLY+VEYNgzOyhUfS3zUI2jSNPv5
zkhAjPzZaUKXiEe9oNYU+27uel2fvdufbwPZX2rDF1y7hyp21qBgzJVB5oLt6e/HOCCbnKD5i1h5
z2F3s+Vg4S+Q6Ojtuh39Dwe8co/kOoRQc7UtZbjbodkmNBkD/ZyLEwDSW17Rv2l3PMOvfzSQ51gv
Ci0Ad7UCQcu6MYmZIovyAozNAUEKscKDzcTUyNWrUC6Z/OAEGtUUnxE4apY79mmNZIyw4JEQpuv0
U04wX13P22GrlNrphnEGhthab1OJS9zDy+eIQy7sUpbEV7KBobmPFqQg/Fv/B2V6H4vt7sXsXgJz
nlSd1EGo4fiIjsQtdLMOm7cWbxknlnlaBSoMDo4K5uVyMMNwyEk6pa2v3liyHr2h1vYQVB1kYlkJ
26n16T6Ofvth6L2+L2AtcdAY/JLagpogOqI/TAnKowYi0h+gYsq++IuSg0HFZ3EesOilJHib8/JE
4ZL+E4T8pu9c+ECAU9JnASHuIMOPZTmZiolai+kzJEVPHfDXOQIzqdKS0aIEZyYC5JO1ZrE/O8fK
XvSMO9dYb/w2JSEHg/u/K0nttskK3g8/ZrZpt0l09EsZKD0uuszJ0Isb28fo3W8szmMRaIr7Z22v
SbxakGHloekXDM+fdAbEJxgP2hbvk0PeBmC/onF/8gGBWSz4aQzrYNGcFLOfkohiAT1s6oIBJgLN
Yzt7CgoBkZ60qV/S4g4vFlR9LFPpaD230VyxpGkap+vGB7cv8EwIlXLh/3FNaqz1Sh8ICRItaMje
BZVYQq9c4FjtItVz6iBTCo4X9IGTB9oY/RpPpxih+LZxckESKMIaiuLLdwKXNiVXupLEDyrj05FP
waOZe8HwyCsdYUD5TefHSf9uCwFofdLHiH9udc0FDcxNCPdDXGNe3ZefcHJNhdsLCW8C8TGkMACL
WWNfwmjKBa7W8Y+XKpUttK41hlJy9n08Qp+MOGaquVVcCd0l3DfvChMZnDTXFqnWmSZAaMTMAs5+
WLLUipdpk8KS6yObAlTESSwF76mYq0n8QvRvdTXMMDTfUu8rPppXhVjmPEKGkbw2F5g2Tp5aPvGg
9SjE4Ww9gVbvMfYTFeC4G2VeuXBmirgLBAroTSWqGBqjSJbB2C1xJ/0V7WXUjb0ssk39i4q93/TX
IkSJPo+dDxYO6ciyUWyrmOik69h7JcTPtG1JM4uruuLXMrtaxdxTSOBJwsjgr7lt2qErYCgbtuxP
1k4N0P67XS+qTBntBjmie/ca2vXOJ1GaoieZF5EHpDZo9OKmHQ0yEuyT7eTDBuUsqJqSjAjvH/ej
zqs+ttRD/kFKWcD4vua/LBcz0OXTALTkTnuTu5VMeiNQT9dodhVj3ltuUbpFQhlIlKVGL8N0Hxoq
SeSRinuKUB8xZ/lX0zBHYTPoktgLO4sNa60wmj8lVkk4uRrouEGFL+ly8ZHxuiG6VoTsD3IuwxY3
E/zM01P5+c3hMzhyQNztxztvpZDzhJd/SMR5CUoEE6FTZ+cVh2wnJjBredJIi2YxOPnSApfm7Som
MzL/nlRTtA3weJg0aJbduHzRLaq72ihrouXs5x8G6A/4WEnEg+Ut+AJc1bOP7e4CIj+bOt0LpkTR
A/7DfJVPc20Dr8SD5lMuY6OGlmKm7LuJEP2a7BCb/Lm+uD0Qyo9H1puDpiEZLrC/rgNnPBDu/zhQ
5/vYZPs2A9u3Uvhy1znrTGkuBR8L4PC3vvvBbwtwcccYLqVUCFB/q7Er9qbTMsxJj+LoRNp3c2t7
jSlu9V7ucaoSPQBVU8wAti2g4ay4qt5FCGx7nktG0OlbthqhFpK2svC9/8jWRkgAM6YauodomvCJ
+f2RJ+QZ4kzvwqNWAe7kUj9Y2f4x3yAFtXDxSx7QBBA1iN/M5KELpOKqGfHanhEXeexj2ANwC24d
W4EkD4dxVBl5qUQYBi6G52UjTfAPsRuPF/XbArolsrsz9VB773wdXnKUgbt46QiJsdgzSDurrDO8
E6VJQ4ZDjkem+9m+WffEUTJDty5jX6YZYlUa8UT4vO51tRnRfKLHoqvIWHDywefqnNuyoBc5/LVn
CK9Zr2PMeHrKZRS2BvRDSqwC/YtKvxqaBqKMWq3IvCoMs+lPAxNa7kY3RXkwzLJKKC5buecJNKKl
ivP8DacjL5Yh21+uW/VK3or97Bknly/sfuqbxxRANdOyGt1wxANSrNS27HF3HyqLCFkclqYMPhGt
fXwBKlszZa1YwhFEixfb+tmqF1jAUmB3EUvAFfdMHz1juROp02GnCRyBh2mrIYgJ4IfnPSiv62HS
F7Is1Ih2ISjR2CDxllotdykcxik4Mmhajsf621qMtXbJcJPSbIWdzrK6ajePa16Cyr50TPm5gBff
EFVJTGCNnbMCZ44kQ1wLcRm9meFJXmJhw63X4+a3kXaIhDVs4u6fNbFIQCdx/Tu9SnP6IMQ5Ko85
nl4XTCy+BUjTucnm/MkN3aKX7dLaY/aWwQJr1AuIdjcrX856WiUIOwQBInrwn+X5NwYpKE7vByHI
8EIkbFjJi4pErrzaLUB+jnHC23XFk/7Gd8DMoVJ5XvwhvjBzl0Zzc5H6MxNg503o33HbpWq+u7Dt
lTfJC2FSW8Ll7wgiT0JQ5O8eYsy88VHQJnT6j1IG2DrMQckAS9TvL20+AvB/hBK/KqtKjcshUXHP
56pqEpRUKDgwTl20d76KGUnEafgjBcMROqQolBpNp2Zr8vQt0AJAJx5KFdXoHmokR1l3JAjos0qE
dmts9OV+912zcIrFxwRkiLFgF7U3L8lTIUgvJGze15FUO3DYTnoaLaJYcmOW7nw+abU+8C0y8RZh
CJ7B7JyPWCd6Uqx3bzntRQkdYpwPBwfMR/wWh7wIErq5cypstPkyUQYN7kP2o6lyvAK4cYDicB3l
EiTi9IxlqMZFCrsRUCTd9IBkC42SoPkpDHpd5FFCzOFnzQyoUGxCtvm4+KqmXI5vCPh+JvYS70Yf
nqQ8FXzsRRDkylrC/ATkubUJu9QqPgvnSynePNShcSJLnF5zyO9di6a/zyV2MdJHZF0DcKk7huLa
jNoJxyuc/ZN6cJnO3op52sOOkG9TgGriRqUeqJLV/wCHJi4o59hOFOQdTyWwvtImHEsbwj6NBOZe
qZ+u4KCCYDMDnxtmWA4hjQrHSUJi8iRIryReXCTzx+a5lpDkjANIqxTGEso3tA7Q3kIhpo6oNnFv
0VsgSvCCHX2ielLQZ3S3h1aE8CI4BB0KvgjZTh2H5e/pLHK7JKnBMpd0ZxV0ggnSBqUso0kAixJo
GNSagzqCaWIbaMHqRmutFoGgoUctKQBk4pB9wO0cYffz15ssh9sBbqPiTnvwJoJUTktZSHEkc6UL
vgcTuPypaqRaOlYaeatvORB1wuv40YmsvMLsJaCN1ZOQoLt1JoRGtKUnVRspcCd0BBk5iHTex99Y
fOOPpvVZDSNEhWo9n2uGKR3M7wBrIB0esc6D2AlNe8vn+MGYbXI5F4j987PMq9rKJEswPyUtGze/
xn2uSpQ/TYIH4mHyuILVQ2yF+CvAIvPEvsgDrOeOTZeeORjSYswiyfoSBb4+UQONI3m40IYDKvQf
VKtP4KzeeZiAe4vfSSRK3UbEnng5X4vEanJMG/4mmm21yfVS7Boy+FUYCBqNoKSGQTSKA4u652Ta
0nYWreex3VOtpqErYQ0qaene0q0nZb3eoCrLJvuTl19jkp2Iq9yaAo9LcBsjP0KvlWRR3QM7LLdx
X27Y6b6WR07/KCv/IlyvRVCRa3MhC000TbB9+/EhgBgVRwP5WzTwl+CDBOWyBh/7CoLQ5sksHqgz
+NvDBfszuH2LmK1ReFxaB94cuI4oairT9w+ZTksxOfUndbbRNFbKpFPRcAqUmvW7wvlheY7WuJJK
5v6WaPkcpVD5viNHfIH5Mj1WLoqrmhDSg56GyjU+fR6NZzBCOEab2kSDObANHFDXwEZ0v30WfJlI
Wss39jmDoG0TO23DGrHtTmvlkABzbaL5CfavMqf2nQOciTnG6gtkm9Jw05yqjzJMHgjlyt3UlKUE
B57ISUZq5Y2QnQpWCanElBE4rqPS31VFYciolNl9Q2b0/6Mu9ZkF7x+MijfWOgpiDMtAknQDooFT
SeuPrvsRMQYWXnRU3WMSdeSWJDBbDE1NxArYhP14DEJNTBU1GqX9yMlS8sSsuBmXXAWWrOCwZ5ci
VbkFG2ULJjN1sp9sgzDZOGO4n01vbSsg1r5nrX9BjT0Hwl8/pnmi8Tqbd7n/6PXvY44m9nGI5mTy
F1aSOOBe7LIdGrLKuOsET9jIAt57b+0MqZDaoxH7c9PBGEZFFgUB+jBM+AkJe41hCH/y4drci3fG
0sHQo/M61T1dbBMc/h1torGvd5AYwlIgY+QrS7gHk0KwcNT82lLX70cI11VF+RbBJY9Z5Krek17o
B3AuweJLrU6lfrvUrlmIOnoHyoF68HucNAjqAn3tZy1CLLo59I2aiM5kXfbEpLHvuFQ0ENwAD7EE
XKIy9QzGRjxz4cqFsRbf2i9WB5tZ7AUparYQuRyN13AlYeEyWI1WGLYV/ZPOrFFTsBW3fTVPlOeC
BW+W9r6bki1hrx/9ilk0Mm5FfMnNTWSwTRrgFp0jyViQ5SHO8/V5PU26Hq7X9+v4Gjk/iAm0Dn5N
7831TVTYnnYL0KAggNZNkUP4S5hKXzwxuEd4rqBdIA+Yr7E7OU4WYsOd4C59mWsVJnLdmlB8LQHS
YYP0Vcw7hRzI/COFqwW+33AOy9CQcED1qf4acHkWu3L49NkPrpo0zruEWXTOT5sRmBNOmLJIN+hk
FUS3qiGjW7UW1sXha+NBr99ewsrVB3u+n3lGAGvNjTHMoPuirTWX6VKvbJ6MAWw8esMfR+NKT61m
AFkvFX6Y0U1lVURYQNYQ2fraotCpmH6s6UvexfuPn9oM1rt7XPk8YEgVRCR1fPgmXKcCKfDn06f4
tPLyG6FK4gcQW36riDhH3N8USOvBj7tZ7k6fYO3m8gNAeNJgNk41kKV9kYFGYHa9uVd+F2toxme2
g8p5XUUYu7G/u35v4GNMlyonHHZu3p0qex+qMS9DGK8STRy6KMLZCXB/+uHAK1hJclLRxsgi2g3v
eqX/8dMuXgxraIDtD708yaDLZkYnhj5BxghNRV2vagiVd3MdmHOsi1EcqPVIjzc3jmlDNN++XQpk
m/tY9epk/UmCYVnRxy8GfLU4IHa8YM7oVEoqOzjUA71Ddm2SXLmoWdK0MUePG8LE0aPklS4uuPu/
PLpr8DK4ZDk6d3O12EpXuvuTAZV9EXGlWKcyGPo0PiCbPhomKxjZpTny6p5wEwO+X6LOXbhEIs87
iLgdq7HXs40SCPjGbT3zt1xzXr/m0oodU0UkeI4GcpLEqJQWm0z/Ad8RVynH1Yu+av/rH+MDjzdq
3Kr5T/dI4G/vPnJpwEK8jJB5nF3GxQpfoD9Fz6NTYmTfr9nI14qKzN4WnRPRl76zCk7yuhzMcJ5I
keh6lmtophst2fbfb45heqQG+u42cmxVPOGzUAhaiSwqOjeVewbFvEE+oAWjcmBZQEMa20w54SiV
TtKm8K8eWOsvfTSAl1SxtcViCET4VPZd+qN65YM4a2TW67Ddqes5fuvM89U9B6rP59m6EfEZkpgG
3TheuVI5BxmW/6pCL4pTd3fjExn1XwZlU991bkiXYw4f9+1g8N+LQx2uiMGlu1ppKZDMoZ79E30Y
IS21HrUPFWlNutKKwqAS3lE3I638K6z7EZmSiqZ4GujozC9efFyElmq7Jvl+DvUj3IZ6eSoBS72v
pN5avJCjLqxumWtg4y1+LWqqauzK4DD21OsjGfrmmnDfIjnAyiMj44KI1qTkyeztODxhvkcLvOb0
QqeoqeTWgLu1Zt0XJ+fBm4SA9yLb/HieYeysekH60wXUXlIJ5ZtRXWGcEfs2+8fcqM64cIzaEwnm
PDdevXaOLMOk4i50n231sME/3hVGvV1lQ5FkfKLqX49QcyOlk+o1dL6aFWaxt3QmBdfQV2xaUNvQ
YoIVB3e2nthTwUk0dTqz8p7alZrNSv0/Hg13d67rkZNRSLqyZZVI0gXFU22H1SrJVhHSfsPu/B8k
DPoOQLV8DuKkAHAPeI5GWtM37ijRZbXeCmsRmpkY2+LRvVT4ftEB3+sELi9PfS/tCudZ3pjRUFI7
k+7yFIGCgjFdrRiiORXdBDCrp5iZ0Bko9tH2PKL9WF9SDOU5PjvITyZsYH/jUaHoQhUaYICNjbh8
8hbKHiy+ltpbv4GHZ9Z/4cnoelK3oAa3E5ZwFn7MuFhqxOtsFAdWySZlrDLzManJjbedMx6v9r8/
lFCn3jHWB7SL4AWYry+fOyvZSnayDBfgz+iZ4lbh9YlycZGY8lzfzN25M6AaK0Mod0b/EcVScLZ2
Azncyn9Vu9JBfsS3Ab0MNT+nIB0JjcXOsQCno4oRi6XPofqPCQiy39xfcmTYCD6YSzY5BOdzSLRQ
zU/rEl8RQimPMhYLL2bJ+zYxwupwBYzmIuIcY9hB0U7hxGKPV0Ravoc8pJbErzKPbDEGfOBO+xrs
/Gep1JlOftbzOs8ZJdh3Sm5FNwr6NVU3QR+FIhc32GAMMKdhCOtr+trVLkBRIwDLx5ECGBqUE18f
CbuKqmQwP6RpZ50WKKEXwO1Omv8cI+QH8YzW+IJNGSNlP697rmaALZ5WEcYMb/Rk2t8N5f9xgzSf
1fJQkfDzH1RyuDq0S9TePvmxRBbKzOW2TPx0r3EE0KHzVNaeqW98uT7JWw1wnAyRX1O94XkRfmDm
2i3kp4Wl/H5Mf2BV02jlDL8mUUZ4aNS11vuABvjCtxET8pa/e7An6a7VV0URqS+oKBoc5L8jJOuz
W6ibwVtWE/jVr3YsRZII4C1WrQmT1/W1N+ByvD+/XdGvzo1GlmvEzHxmZ4Qf3sULTX1qhZzBPj1K
ErUOjXX5IK17DJR84V+Xj9XZJYAavSwj/bt44CwwmU7IVK/PTP8ueB1PPlbss8HPAezt2xSENrvH
mFCnG6E+721nd1W0gwGcfF5BN38uzWHngNWpFkdwPr3+uls75YIiNkRyCZPu/w2w2r9cn4uvU2do
onmMVIiTe6b8D/gQV4bqsali8c/52kfl8bHVt0z+62IerzJXsRRWvzVwsplwYqkgqwLQX8/Ga26M
/ICykWjzbWiCdunRyWONvWPBuhI2ZmLNRsCSa4vzvxukXu48KlIITiWS2Fm8j1TgoeY+9X8HAENF
yi1dkWnDY1UJrcum0j0lynZ1nKxE9Gxf7yF1weDqySYTAdDDf7xTv0J12aQ2JcAsBJ6ABPXarFMb
qx2D+Z6Ce4xseDlOX7c2gwr9wR5IWwnNw/9J/p5d3TTcMtlEBumwvvsEQ69O+y9qnTFPAvy3HRN7
xpwDA1Y1Lu4JN6hGmp6W62mawFy/EmMfq2x6RnD9UMEZREry8MMEI5zrso2wcvPLpYi8erPWIiJ/
od6KkBiZx3vo+Q7tirZBXEkWbRvMe+R9abvyzDLH8HFAuFcK7igKzR4TSVVFXgP17DuObDfWtBM3
94Q/LfhsRxR0Mz1aQZR49HzR4qYfjT9rBJyskYsHMUybBm6IsE7eokZjEVP+t+brV4RPGTaYiB4E
oCq6++O71QRyBEMGJni1IVj5UdRp6Bjbr3v0WIAAOK7TLboV9/djHWk2aqIcFMBmWb2BljIuMu70
HfDevf4fizrSmc5TTYUyixiLqVFcpvNnmMpLQorooYmkH6ZHEUrT9coJSeXyGeEtcA2OKvDxAQ3C
vLFPRQ4fp6XKHnvmZi+Ff1TViOIMNHfZTDrlkbhKXoV34nZiZRGqMNYZ8c7WCkcINbgPu1CC3OmO
XDOLnku9i7BNAhrrTlsdlKVr0j6Hn0RncSrxoc7GiTPY+uDpf4H3lzOM5e3g4PzF9Vze6jyf3K0V
T5uKAXpB2unfAA0tNs4W5w1VDXQZM8yjy25xdN0zXwZtVOUwmugcqx75W03aX5i/sZNc2pbiP201
efQtEe2rM2jEVF5NYO7dd1CAuyowu/f/GqvUIVViIciQ/jBTcCYTbYOebjh39/EtFjKWTpmItzla
eMzRpEAUAsc/5n92HqmT24aTJFVf9emw1vF578HAaP5Q7qSr4xMfnb/BtmRvhiylAIOfVXpMzUGG
fcXB3zQ6flx+4m/G/NyKfJj0ISTZkaMm1H/7Cu5/EbE5xuYwqzzyvZHfduul3um5Rla8n5yYmeKf
oqUmtAMBbCeeCeY3j2Eg4mhRS3aC8tjqwD90FjgGik1o3e8HaGJ4GF+I4g6AODEG0AXArAiGAcCy
YmTljlClfPESTsVACB155xKuNxr6O2zPnt1Gjp1npRPXd0TISGlsoPHh4AqxTcJUCuFr9hBQJ0e0
lVHBDtyAy/Tylx0MTv5OpOxmtcDFOTdWNarSwfmapbo52VWMDV8ruk9CzRt0LKQZX3F0OVN+s2Ti
jnqxm7q1YNmUlJzQIPQPoIvNB+S1JfMfwnceEzFPlSuBzi5MkaGle6PLJthbXToOrnaBdTqha/PY
96NR5GZ7d5iyCnfbMUYTREO7uaUMQBN8FMd3EicRFtFwyTRZ8I9qSBYi81duVsdkMNdlnRTXk3Dy
/Qr6bExT0JQv6lsdZDnLqs+U3aI7vSceYn3s9k1WTS/46l2ZPIV7Lrj9FwxlJGJwf3syWfWgqx5M
wgWjqS6MbID6/ItzBKw+/rrAZ7xLNFfXyEplyoz5ChrsiVGPrEzAeT29xHq16BSzQtQOH1y4l57Y
zkIsneeRDL4yBAysYlvJ9i9oc6H7nziimXj3QUMu/C6i2nbx+7ITm+RiURdzTsHAhmO1INFcHAZn
DCOPRGmxZsazLJaTFDAc8FT7zjDS+kQ8wgTDQuwq0+Cd3QvIvOf4ugQafhjzkB8kYUyXvZNgIurt
sdzrTVfrw7UFnV8R/M7CtBSMnTBp9TuY2UHQsWOr3TrfEOkpx/prP8cB2DDOjxyXvENhNLOrdkA+
6i5Jt47pbdge06L89XT6WTUdmrgEDOSYGd4ubSJrzHRTmmJXuzrQJfQgffmAxKpl5E7cIjC8ntKB
pyST1K5yCfVBzR6mtVXPFVs+IB0cjP2iNl4m3OLG4nXdAT2xVcHlPw+Ikx18nocPGadxTG/votiK
gVi6YIwqGMJknmRz2ZSdC72XOxeI4rYezhG51jIWh5HuawKF/npc8JPIFfD2Wd/JLWnvQOQTWd3D
IMnQCyiX1jWx47HaMDYPHrghRL9eGoozsUT3jqWLTxYS+NlE7eHalyo8/kkeo7MaGFhqHQEtQNYc
n1LCPEiUyPL2/8Jq7rFoaupkt3DeLZwpmeHBturYAgv8eK0exH9tLxOm2h8xztXjwkh/DcmnxT5g
SxV6d5SMK2G15S9MEWuy26zHvgmPFuMRHpZbQ99CmfspNjTGD03WvIoCpZ4ukvNeMoTkUaksWjd6
P3N0TiJyNnYurP5f2Sjm6i30GZy6Rgi8rvswSLZ+u+vIyxuEZI90n1fkkjOuagBfOqHhwcSxBo27
gYEVorL8aoTyewfLi7kYfaxvKQ/6KchLkl33JbIr755EcpzME64RPw4BWGN24WBJ42Kr91psi87E
fLPbVzgrsG8evXyMZtL1QZrFi2E7O+yks8zYFCQEtC/NRlLCxlS9KEHeSckDWYThIwfHlubay9yt
KWVvSpF0HY8NWvK7u/7Li7egKFhIWm31RQZYcK1QSlX/IHsMVLEEAFOXxIql/mg/+JIa85UIMagg
NvYQYqX5GIWQKMR6AkyLi0pDHtcZYwbc5aDiMzp4jmd6nENi7yR60hnI+t7/TwUvDgaTJA9amms4
C84Cm9KLBO5SlS8bkZ6pkg8KgyY4dB9J7C6nS5DsPSiNQJEN0l+aDghSFqd/8qXq/GNmWiO7oc3Y
Cbp4sTr2QAWWjlcWx2R479EAEC6+TkJp0UaP1j6QNRfcgcdKnLwt68cT1Ed/4obG9+XQ5Kl52aWW
bjgQH9Tzgfbt4FPgdRY5sRxXfnS6vukk9Q0MYnnpts+VGrT/J2dGCoNjGFyPxuqo/tcdupGBAPDu
XQP1VQlDetiTNOPslu0K0GOmK9ebEJ+GBfduEM2cCFubJI5OybKT2MSjka6RxwcPFGe/zRYdmhpc
k+kZ6KRTLdL0J5T64X/uiGAzWITqipE3D2ZFEDDN5nJtHuyRb7QGDm801WQbeMh7Mmtl/CcBi1Xh
Cf4o7v8+irVDLrycA8Hul9tdY4DWdAeKVZ9b6JQ19kZJuqWaMfzYWbMPTgdwpyQPWCQZDCHjGYUE
Tq2SUGX63b8u7pPWsWR3rBfnTaqJvW+OPlbrROpprHrH+lEqe1f0VMsaqXTMNl62QvFaL+5UwTPy
ZogvYn5gWRWwJwxH4W8O5C5SKNxJceMxz0Vkqs0wSadVFiVAOD5/UFlSLsG3rNqOWoxu/JGFdOmn
lyFOnmS7QARzqzg7Oy+H1NkmdgxQ0vFW3WEvXWPKTwJz6gNnsSP+sGSdJdendGQM+ltC9cZ9r9nd
Be7Xj5OGHn1DRy7AapHv5W/YLhrtAbvBsCSIjwCqSG1xbaBU9O6yKwPBqvJQqdALEKwA+Nrfm8Ur
Ptog1NfIdIvX9Vxu0ViP9/PYfxi/ZaawHPP9vU6aMo7uqzVqPIcqxRi2byH//cR5CHAw5+ZqoqDz
o79WjM/DLJ4+CbwIeFI+aur4Fto69QDfetBuqBRPt8vnxsqfjVmiI7lRGyut7A91ZRu7YH7XHOgu
ULDh8SsvBIu3zHA7rhP8lEkOBOM0Jrb01z6OZj4AKF5mJmNWLPOgNWGMi+5gj8xK+BDoRJxh1sOO
D4JqMN0LeTsyjS8T9D1tWaYp02XhEH+fIab0GoEhSrJMpxi/X1IxMRvZz1Cf5JRTPvjbA7vOcIId
eX4NNawDT6Z1KW+Da7Onqr53Gv7OPT4kOfOlNMfw1dwqKORVNP+fNvzBsTi735Kra56raw5c9HfR
+UUzsGOtsmsgESs2BAs7sZN7ZX9FNJaq2ByU3yyK9jbO6lvgn5On8p/cnVmNddDgAM61F8Iy5sYh
j6T9vgLrSPdwFjSiB9bkFgQclMZ/deNyb79W3QrUrV2Xm8RZ9nas6VYPoQqa0fWNZcKZMEpktFzU
q2iZuh9olOIerL2fLsRoZsytTQe49xulDtzvhaAYI+pCdw1LCqi4mzqTqQEZnnqKaWhsRMU7GECL
aFdbDcFwCETkJg++py4OCY0uG/ON1sgIFpwE2U06dKtBF8SydXCRQsI/3xlZYSAEBtJe5DbXkLF0
zi3tzSmU3YeqgFOuTTQmn+5Nwf9Cq0QDa5s851gtipTBrkcTT8K6VWV26ZfKtT/TvohPq1pAKtyg
lxJr7WOrXcRwkq6RRRQVBgRxvSNdz9E+6Adm4M0kzZZzPb6Zef4/y0lDFw6j53rCLnD9rLFU65LH
R9M6Yeaz0k1U/BJWWr91f5Rbr492+35c3wqI2J280u7YyckHLtv8YypnBcFESM3b3J2w/sfd+wvB
bfMNd3w++SmgcLtogQ8S9jwj4esrx8cYuYs7bpQquxv/0PmbAFzApQQh1b1eufYCPOC7z24JcxN7
sqWAnfoO0tZCCYDNLPSzZI8kySM59DJybj/xuatVor3FUgsQv5Uxa9KrflFh/zQGn6VmTpC6w1sD
paUUpbHpEJ4/9K32wkfauZh4D0hmJVwHfkVJo1rDFkpaMC0w3LZHaiyn3pwDgP6w9wq0TyBG4QPv
lE0Mr8idIVTqyW0L0MBUEa5ojsT15V39h8xYskkxA0v7MQfFjVMX+44GoxAio4uva5nx9JR9dxmX
lRkWZVO1XZgj19+dWRlPFR74r3goqEtu+T3Ul8bg21Wb4FIcaN758Zsfr66TrzoSTG5rvpJwS8yW
HxeEcovDo+2Q7zZ2qOUHg3EicuNgsvZGuIsISlS2+Bkmvp7VMurA1X2mV1mdqA7SStAk1+yAEKUX
2hDWyTtPJu5pqSJlFBNA24U5F3Rydtn4dr/o3diH5s/MaDIURp/uZtbAEOHdwYvdYRSTdUiINDFO
/K4bmO0VwL8OD/HsViOwMXox88zAUR2CGQWVi/PWNs6QauOJXJkHOvd6sELy9XtuK7Wuq10mXy+R
hEYZvUsBlZ75nf1ngo2+YKWoUG+0Uv5Ga1ERagzubMJ84jV50LwKDW2Hw8VwkPTwnUGmDyea5bGz
UPFFj7Ofy5Bcy+m38Aa7uD/imA+6Gb7IfkqkuDhXx2MK377HkUk7Hi8ueCaYA1/lbRCGssG5U875
G7vahn44aEsBYDD2xgLUyXi6Riw0LvnCYUfgkwo/gSRRy2AYs27WN6T6OZHoISl/Vu6QXmb2pHPR
aZ+od11k89WaIrZOlKXh9akQG7ImhG/NqRnI4YMKydeBcOFZAafocC1MN+DjKbHsrTBzVEksRm6y
Cxwd0S1GxnRvhpNVCYtPVYhf1wPs7vPUXdZrqfvitUUw4Ii9R3ls2z2dbyHLYVuxv5cm4xfd/6Fn
T9yfTCrfsAvRab1ys8JfMrzNNQxNwr/bBxywqWxxgeBXkiT/HsSA7l9Q/qBDVqwwk/CBCIVxeU6n
Idv06fsxMp35aZj7alxZzFoixy9Yyw/B913ga/w6NAITQKm/VrZuB8/IiP0teGzowjv1W9WBnZhz
wcjmB9fSO3zIpcXgwVC5LnEuS97+9QkxabLFcre/Qyzr8E+1cCIjkqetMqDxTgqkRHMcbwvDPka8
0LKdpJJ+2+W+Q+05DgNOm23M6760Pey3YPSAesliHwtr+O/O9HtGywJn/N4qLgQSPFL+hBUbZJtg
6cW0QDlCpQPeGjTrMPkcgqyA0x1OBN1BTAjYC4dBIawLx30JrLTBnxqU8rM4kNylH0KsotQXwyod
qrnKCj6Rcg7y9L5SOEGljCwfQRBgGeW6Iw6tPGvQ3PlQjfs/wF8wKIWEIAuxNTs8w/5G/XBdwpkb
Ejy/x8DkmkUIIJtBZAT26sXz+40wCdmShXI1CrvWZ7tgvpexJUdUpsLHE/59+YlYgmMNthaESNSN
bsTlEFDE17BILg/rCSsgvlmcV/A12xxcEQnyW9rCu0Z8VmfJQUInJqKSiShmMzV94eftzBYjGrA2
mp+8I/IVT8IDUzWrOwZWglDtlzx3Sopb4z8RiTRYWAr6xDCwdvpxZL1/Dhx/PZ9ULiodJ02eZyl8
RVjDw7QtGQQYbnsbOHULxFycKF/uuHWHIF7c3AcGJrcxCQ5uHuwlITx4W6xo32JnePe2/cRVsxNX
B6NAfmY3KFWUbMnW/p5KEcXGq0wZ62kdRN4ChSEO8D2Bkgdz9cl8HAHHVvBl5mZN2R221mojQGjU
AI+wFzEdzr4gdP2Ffj0CwFkLf75VJhkdDbYKjx+eVM+OjFdoG2PP9mRxt+0JGbvFinmFaLJ4HKv4
TPrGMJuByF5LomBtQSs9uTih+5pkY67GP0/6iI6o2K+GGbdlakYRVxkQtNoBx3FlpC3b5QxwIW3W
P6e/tm5tQOC0VJl+SIn0tuilyFrcKeHgnvWp3l463YrIi3GfkEky/4gye1bC755irLmLB5h/zS7C
YYNRSSRKkHF14G5mMEWo1J7TOBbDBMyp/OUJOJjJyq1KzDxeMExZNjnRh1TOe+0EPn01i77YgjmV
nRAsgAVUkrR4VP+tTupKeauPGMg0QjSzQry9j4WLG7L08JffcZkYljKb4FCDCTx3+F+/XpSzc/GT
5ls6YlEriKezc/lSiWSBFb30Tb5F/EOVw3OWK/e9DqB8soRhgm/K+siV9tzQOwIGxZ0NAaYz2ewL
fGU2nP+h4f69N7uOPNObpoo1IRgzRH5/Mma1fZotUa4x+k9UUV0lgfd+dBECMMcsPTZidH+JFGqm
DeEMtq/+0oLSmEM9q4WWia4ioqQ+gQRSnGkd7vZ2eMpuXwqo0v4tM3FTOgLjxKg3KLCAmqvyHi7F
ZhoM1FGT6tdJgUusdjjby8t1oUw1FMeom0hXGanECa0jPltBvQ32/v3evaY0qcoeHrEJo7o33GDV
o4jMoTTUwSVRGHr1S2CK7qf46jHc8svrFYR/WYxOAeIP48mOFJplYXcVGLqfm6eUcsmMA5OHXuH2
jtt9LDBheWaqCvcNI59tRgoa6CG01jy5yEbpz73UvTmjs44+pOOIsXIWgsdJeZPJxFZMEUiQVJWa
w/yJhfVJMYxwH6xx8m1FDowg17K2Qcm3cddpoInZfOS68BrTFdjZdzVVDIu/T1eI5YKr+Z7lcL5R
cxvKyPdmC6/AjxndWyD1PWAtAp97IsrTKBfgOzr349FchnsWMAowp5fX/dRdgZgNUSMxBvYRnVQt
QrThyogkmbYxTCHa9uSDQbZLsc1oTnGKNeadZqG80NvGpoS9z3yKqZvHw/very6uVKfta5UF0X/D
C1i50EgRW0dTlSDzbYb63gTvXtCjuCat6wIniy4SMmt5Sb87rq4G1/y5UfMuFSx0YO3uvoE1PP3D
kZ7287sm/1wGM1+K5DtRTl33cu/7vbv/M3aLBuhkHioZ8P0VfydzdSZY5+Q2qhdjVvHPTefhYMjM
0RIAK/phFyEAWOdNM70S2P+Pg2SHzN0ltTaJZu48vw9P+lOC63t/j47qf9Ial328wo+PV7J6Oo9P
nzcXFHuRyWJEXQ5FKotmmzxd8rgHMXuHt5BDh7g0h0B6Ax8CCLEwoMN06522n9cCBpQJCSOBVzr6
Dk9Vr3uMEp3XFzFKBtx7XDY72etoKzF4SKL4GcrlZeb7ODOYHdlroV4GeeMNxhkouSWTOgjQSKpv
Oj8nNuiJ221Hh7n4nyvx1IV/QVsF9aDh/s7YAgCL0l1uMzeFROyxTkafLLQ+UEo/+F0lmFc2VQv1
pQ3otNgc1o/AxiRveHUkd4pfDPw931B3prHEGOVDIxjG7+5l09wOD39zL48txXmkCeGF6ZMputR9
tTeH2b1N3rPkKEU385Mc/XD38FsL2qP9CfZMH5hxMRmkUuAYvgzlXBMjsLiqqUKKPXQy966VcV5e
PcliuckL96V3aGYjjRV4L4OA77urm5lHqC4XqFaOi/gdQLwDsF+8nxWLgm3tcHCClYLZF3s4GQiU
LF9uTtIu1iPhMxLhYhj01XDcTv31HcW5ZTHTezTXl1zegu9PgF7/2U3gJ1yctbO09m0pM7MVEWPs
KGGwW29XZ9YHo97mJ/FlzvPhD6ZJI+W9p1+OTiNZkOZQJt34UkYxz55U+EOMUHV90dnH2HlP3Tj4
IVqyn7z7bTMOjJ6zlX3qBGWfDOPPCneJ5lh33GFKYHpooZW6HHOAw4daVa1+fTUHO18UBbokqr8k
6MMvdILO456X+fonwnB3kujpBOe+suCdfvDF9GrfwLw/hH7OUPZsaOZOGuuZUacJNS0nJ2g5BPsz
1BrisNdcCWtF8Gn4nyqdypzCu58NWq3ySi4P5W0xWkSxhP+wY1900rzrygFL/wzaiobDxS5wgQ5N
iQmYUr58cjdE6ekts9jduNcMLEbHjB2VKudsWU2kCIybXPnFrfyAJgbjaCoTcI5e7tXkhLX+9+eN
3k6r1DqT6+Xri5H9fL1SYIk6W3BZGDWWb4++AOUFba/qQn8CsY/RKiamvyx31dUlN/4jtkOyjr+a
jjdr9E23nMLVo4giMBJMQfCJGzaTtc4CqVcqPKRzGG8u6/cVVVQu+GgJk2yGOzTks0jigRrnhtSU
4NUTAqLV6Eabi64fWAhYWGQuieZ0CunyHkaj1cls8e4+e0o4Nxeq8no7866hIwclaRHHts1FXybs
h6+Rol/RAf/TqNdZSLuNkuDMYkXadawGhlo0Bq+vNSeutOBULXeH24TVI7Q+luZGdMt2KnDK4WNQ
CLQM11iyjVNkDDcp1YsPWy5CGdhKi+ctthiA//x6IRla+AbNrGCNtoQsp6UjiKpF870Ud+avOdX5
S1T2dGwqD1G2CS+h4rSlzMdiyL4RLF2n37lR1LUkuVzeNuRSlYxMT3sOxwlLPXuBB9mFsVp7inTr
wkoCpdA6uoY5+FW3ISFVZUIDSis7wGatWm0uReyl29Ry16oadE6bPGrQsfLqldLqsmO/Aq8IcFEt
4BrC90LgY9Zd3i/LEprgb799v9DFQN/zu6/kUEo+gBxjFzYH09dRY1ynpEBaE6slOs4G0w2bo9f4
D/8d/KLBTVEC6VjiQ+Wf4VdePcPpKVE2ezYAJG6S21t0GEqKYVU5QOAhf6zcud+18rQ4hVVZTlp1
bTlxv91LH8UB/3R32mSc7zMPdUPnOGZ9qFbCV992EF+lYLrfjnU/cWhI7TuNOaKJYzNOWMLoSgok
SWObRbdcOwfKQzxSseB62HFucnfgcp+VlbsObzvBb+r1ZvvGb8jiTnfLw9p/bXh6LmK5yJHN/gYH
aENmsMPUJ9MOye9TYF3Uey8Fe5WHnHFbzbgKWV3h+rPNKEzkflo4gcPUK6sk0b08IdBK8HeQMSCr
4cf8GAEeBzWOgoK8m1gGQkObTv5l2kDTzPY4lC11bWw3YTBjkCLn+WLZXCmk/ocudiuDtFIM7rej
Rj9DJJ5g08Z1NbKVy0yzFR/usSR+l6NaplGUbuWjehxckVoW47+DbCdRPWm9YsE+nm3Pmen4bhbE
dOPy2bqb0TIW84W6PVIFbUW0aYP2n7aUobXcoLfkRGDWJwZjNUSgJvL6cA4vBPlgl08srvjr/inK
1ieWlB+1WfTTzkCScnszDeonuEpAaG4/raNNTROh6fhyvYu0S6DZgVsdN5Kwt85aRf//UpmVhBex
hSPVVHBVgkz3yr+dG6wabX3zcr1QwswjglIYlkxjAOj/e16iUPgd/tmnDS+v1Pcw5TUiKSlfZR0Z
+srbDLqJIgDzimHY8YsPpgFgPCHrYDzVXF2MdNHTnTQFm9bLeUyfEp91/vtbFK3VNzS7jPZd5OFN
krlJM7y9iY8LPjYC20o/JlaMCqYOe/4M+CSQxQQEYDfMGYZybTe+j4sVIFBw6AE/Z+wjmP3QkJ2G
qe0IP9AcKjDOupHnR+9XxtDdMEAJqQ4xuylEpohJ4qAbzfWxSwAV+OWUS6fiXMG4fzS6HB9sI8J5
XXYrGQZb5+yVpfw0I/j7tMW69uctZOPZTTGfEBLrhmE1Cy7T1Q/amxhBaqiJtlC7Lf1GgzNUxy5D
UajiOUfQ8O+7E9W9Y79rbfegCWBdBQxA7gDLp0ZeQN3JRc/AnQlBNH9nrthHRMuVRt6qj/6MUCsd
V3IhJBxtxBK5ewaoyH4c/tvGqc9c96E1JL+n8hWJohjV27jSYdfUXylYtkM/a7qp+B+sN24OiNZc
/TjRjpI25n35X8+W5qMI9nEjtXEcmheNHCfxnPzmDs2u/jdIK2aYPbonIGFUflnHwIFCIyYZbgAu
Dm1jlQid8BRm24owkZHs5gV8Fe3pIdauVOuyusy7vjmazQNuIl4nsWun82tRF2pY0s9kyMSI1cI9
wE8dpYCTv0YLgJFSsGbN+Z/dauI0KpxaEmp8Q3pDW3vOx+0DzKF5RY233M/2uacAi8Y0TKXS9GIz
lDKNclQISVPCLgaOZyStkWrYrefSZ5SgMPR1fwhjq2kywj4BG8D+vzva4Y3X5vrUyG1lpZobDyqd
vdCaaq9npNSC996MR6yXizUGA98H70lY1L5DZQ5aedZkYYot2Q5/S4S2BKt+NoIjAuuz2IZihWcP
GRrpYCee/G0DY2yk071gH3LTNrFn4XK1wjmwlHtqVE5bGGktrNIr4h37krFlCOXkMTA8VYO4/6eH
3EROTyuymAD2n8xAgZB6c8Mbyg98B0Q3YYEZP1capeyAaQuybx77x9uqUUF66Fa+Q+wXmV+zZzQ8
7S1SHgKb+fSyUQxeoZhsgh58+5ZJe11GFullKtWclPqv5TbeMcKw7xTyeB00/LUlsWWPKf3XsLWH
Y6JRByATainDBvri9kMiArt3toj96NyCJM32mGVt5rblKeJsrUfqJwabPweNSz+bxJlpt0O03v1t
E2sDFLTUJycaOtQOju2BYbycOUDv4CiN14pBQ+Qo2rBHSDr+/SVnZ6/rD54ruQuwZI3zr7FhjUpm
2PCxd2idQB5b54BVHEP2aBDPXMNy5h7n1Vva4YFR0AJPqrvhXbVRew2R1EuV4feCS1hRL3d0yiw/
0lsOSriexsUWgNWpue/AVFJNLb7Ofugl5aV+rqZhU5xmZJZg+GHLCj0FpVbbXDSqy76GXDo4eedi
8vm3GaQA+rbZXteJnCVGafdYck5LdnnrWRMVIVKDkVNxSlR7BBIakGHS7ZwXLer4iYlOiK+x89VO
GrtrqrG7cpbDdVmSrDXEyPTEieRNxB7qKbUUvrGiS77NMdx3OdcmdAWvUz/tEEfcpFc0FOewnY9Q
S4Hda2dM/R3jrGitL+bxqgy/3c6SfwYIXeHj9L5Kq4Ki2CJwNccSSFTQsdXSEtBAeSuqtwNPrEXj
raF9AXybSFMfAaxeMMOK7uERqBazinh/OkhalKF/DomoVY+DJZlMbJGrLZBWJ9I0FL7OMNcScQnm
hJShQ5/U0857TuwKAVFvY3eIOVEfWypdivqwD3NeQAuOXCFv43CtAnw5QpsiGzJllGVbmnIwUtmm
Rw1OtYz0IntwNJ2nkoANI+z8+/YSvvTy8J4lBr8Cg+wjTs9X+n9J/pztJQMLwJI4Wy0FHXB7qYM6
RaJDB6NTnKUsXct51fNLC9hIteoWtW2cCAhwdgK4kQYufUHnmQM+F6l0kksYiIcNvlle0Bf4nKHC
osk6S+/y7ipfoSKkviYtaTNsaXqClWIDwBg994M1MbZaPAt4qyo6ujVonHh9e97bld40XsW0Mwk0
wgGq957nwI5o+wMfmmYT2PZN3Cx4vd5XDBdkdq55XeOTVT/6NkVIO2OBLKzdew3Jr8BUPGvx3Vsj
pmA2vQBfPhrNQp18Mxcqnz99H1jHu/NJRtFp4ll2cfz1Q+ldWF4zYXNczZSNCAsptDuWMEy2DWH3
nKs1NovnSdXA/PI81TgdvqlwMCvzmlqpHIAe2tPTdrKgXJOiPTM2msunhpckq/y6FDadHc0xXiep
k80WW77bfFuhIZXhQj9RvYX9ZwJbOSDzeq00A/yPbZC9ENhkdrL6d9en4/li70pyl8IzPfAGcUYt
PER6w86E99hG6Tfj2w1VcVnAVnl4o1TkJvI2kGT1AE8FhQM102fENgDXfYYzM8Dp9hYiM3yo+R/g
7E+VdONA4SogJWLqj/EXEpNjbT1G7SbO6HoZpbm7pWU0zFdcMT+UOpa9EOKYuy5/yDm2oq2Bto9R
GGVZFTO+V8z06mTDNj/JJBpzei/Ax7p0SA8VPqFjh/1Su6I1oDhHwilpvQiE2zj3FvYtyz9U1HNf
QP5CkVsf/x4zVPynoZaO5sEVzARZToDGa0zb5jHkYoLT9+OaMOZCqmyHJ44hJFZDucuqiT0jGMs2
6UVt2aXR1QAiQB1HJ0Xlgoidxx0qFZIxbvmHPQyplTkqUVCzkZA2XTlHcOwIYH1yLmdXwkOtfvEv
Hy53g/i0bgeb2qe5GFErcy2DqBTZPEfCCRbMX4QrCHlr9eTGcteU/yDNH8PEeyI3ZVDGm3zLvSgE
fHaciLK1uhehXgqx4dezYCqOTiPCjN5pMAf0jNGIHwKmeiZb02AwIR2UdjZNyzrW2OXR0IWM/9Mp
yhH0jrCI5vLZRf/gPv1QCyFtzH/fqmYGQYuAmhSh8VRBpQikWRxlxjiH1H0NB12otj7ptVneQP4n
gzVnrT67j1zADATFTDn7XjJlGkzZUQf9XVpeNzD2Iz4qJ8Ob1KSSkg2ilJqfjsHDD1LDNxRGMlEa
ae4Mrq3vX0UridYRvv1V0D7ri6hxFCPiFVAchMXu38wnlD6uLmbrdmvv+y40B1Py7B4kmkidgnfq
Pchpu6M08DX7obSUM/STD0tmzrATeahbn+zUFZX7ISU5F66D/Sl0s2dlteyu9E8hcFNDnjTm4WkC
V6VQoQ4DdqEDUXV1wC90/UXzT7yfKXgpLR2eGtVUriVwLlwa1qf9Espe4VilTjbTPvmianJtDOMB
V5pQQzpsIZGsqCgAic3fd4nG/x7R4O7N6K5SHFAtcngDgMl3UMKU1jMkwt/fBdMPDhpCU+v7Hc2f
BvvX3DCSsa8D6cHKInqIaq0GW1IxeG6fqHffq5DEtoDyUuSfpFBZOIvSYglP/Isu+8wwvQUpyH9e
K6Wfsip0Qa/QzKoOoVMGCuQJ7ljH74ko5e5SZmlFocXekA27ox0LPDseGXX6PO2zxEdKZSU8pDDZ
0RwNIX2HLyicoHSq1aQuDJDjwCRytsW/2YB4DqrprLOxIAdgKzJU5tsd25/oONedYrrAQDzIlW4J
N30rZPPTcb/HKbjCyChS5+9nLs8M+LQqpAEcyF1zg7NxV+XsqK95maoyEl9EICn3B5Nt0+jTM3G1
KbAkCqmUJRr/T7G/zGyupo/XdNUET6HE6W8p2BhDtM23IResg1+rn70WwygdJR9MgbiulUAS/OP0
wYpDnD0t/EWKocCnjWzBbos1mPCAH+aaQxzbTgXLI/tXlAYu+e3BTkhoeqkEVpNKys60M0JuDCdP
uSpfM1s+8dybd39Gqkj/Gb57E0djbrWWk03IbNoxVrawqYdmY9mH78PmVV9vZpVaNpOvncrrV4Nq
vGUKrpmHTkFHiRX8q81VqjurXIcQ+v+1WoHlsbuQgzWs85G/65eARlwSbdT9b1vUzHecy012Wpje
5quETBjnIz7kqaK0R+TuuoBqK81afK60WKbK1iEAbzU/+pRw4rUZkqBw2XS51Kg1W4SQxSBUXsu7
0bRqEJCu5bThon4HjrlQ8/vHv1obrilLQBQhtGF14jSkaV4m8zCZIyiXHS64Sb4RHD2rdPnO2Tgx
CM7F+VFJZhlX6G38D1DNbDuE9yAOmYGoXfoidkrVtyMjtcw38XiKk7zG1Te3v0gpjPeYgH7GBCU9
bZ7EEc5+f8ubH00i4hjQDGISdmqc1vJLj3bke8jKe7NAYS3l9WNel76mcaubu7ejMG3C3F/KXklE
1ysCa5A+0vZXf9rmnnabIH3NApIdlpsphd370E2PmiOWJj01VpB33rxGbC6ilAqdCHo7bt9iKKNA
faaw7L34RG4oQO4HCC+0VUR+4Bx+su7drUb5giPrxVgFoxwyJ9oJka9XltFODK94OidLpdAWVl/F
4xxd7PWexAO7YaGMUBnBLXJQnhCqv65iaUWdAZf9mqc0MCu+wH3JniKoru0rME0xzz+lUKiwhshY
raI9jaW3Q2KkzOJOovcDRC+LX7QRLgpUnd6y8rPWOKz5BubNH9DG3CerPklt9NmTB5t1kZcjTXvL
ERKozc8FttIZ5f4quqfW1+MhkW5IUT7jJd10pZ29LTP8SMNVFdh5nNTIXdI/2emktrd5w2buT9qt
XQTSrhi/o3APnJ3a3HxRfUap8fBXLvAnci7y9LjoC+f6DcwSpKmQnNcyLTFtEj5vcYvFolh+lFYW
1BRSPylWTtCw757g+JYCfMMUCJB3wj0N9wbTQbxYb4tOB0P7Nj6yAfx3GxbzmOyod8xvJODKvpD+
cS4D1oFo9HCkcDFcojuRaOAwB8mnKwCBs5bhVZTZfHVq0Cml9ssFJXX4v8Gdcd8gumu8qGgNXr4+
+ydI1D0GOlCdDz/5C7YjAeXfIhcAlj8iMfbthoYZt+sMZCphmu30P7+af/AZBQ6tzXC8W+UDYVtY
1+33a3FEym5S9A/kjyu/ZtAHG+I1FqEFWuBaAz/jpRL1FQswd3PhIMDR8WKhNBX3b9FfYQuPRFUF
hx2B8viM5QMzGTsWguPSoW++zMevmAEeTG/6D3DsU/pRbJPeWbuHVjdqHEXylwH9yKUCBkxtygUM
PCCuIPwpLdg5hbrFhfQVVovPhGt4XBzrM9M10sgxc4gH7OZiScFJKS29O3/YNaL09ZEyQ6+CaHot
fKi3g4V8qJqF+IwUgwHvQ3x7zXrjXLkwpK39d34/FEvJQ7BvQ9cXHkXNgF6OqAPhshPv65rae0me
Ow0WLXo7KJG87qdu+IXs/Su2oVpaiazMRFe0ve5tUEOyxbQzHZoTdsoOPd3eQZlvO5FObVyyUn9O
C/Up5WflojOdXg4WNG/2fN9dOEwbNou8S7WurT0lvJUKJiSmji4p6dMsfzKEeVPpEGMIFOA0V6/S
MV2oup1SMgldfYhVoeSJ0YFSWvJYqXMtilD70X0BslVDoQFDHkdry10Gm5q/3x1GD5RworEZ2VuJ
ZFhGxQJ6MDE56pvte98vinhvOA8E8KAKpX+UPqvwHUmInqgc12b15cxLkzWJjl1Ea5sahPGyFwYo
4FTnstKAL93l51pO8RMIZFT6CJHjwj8FHUe3mMzpN6MQ8LR0mfiiLsTto0aATwrx3/qdn2WEqtKU
TTuRiPPR9ZKgy1tjPiFT3JCWVPHKGwuKaV7pSHAjeyAyNS8U3MthvNKKAhMQc97QuDgRZazjSxyp
UUMltD9R/bmjA2/thaMAXASrtq3mxk7BiLOVxL2mxvDT3Ys9bTqS/Bqejkq9y/aU+MfL6NiKkHZT
RHnW7lAgoc0KqZr9MbZNQvOPThzAfB+e3jA7ew5nMFsJOkRksTRyRfljx20rIQSA51pNwIOgU84G
kyfME/OFUgX/nW8dqy+0PaTBl9RIgLTS03oUAnVRLtIE4vx8uPAZrLPdN46PzBni/ANwxxv5raZM
uC7ReSiVgqmWyYR1Xw8evmiyV8EZ2nOlVkJS/NOd9V7nIHQ78QlUXir2lW4FvuPznwA9F3mgToeC
gm9WgaJau/DGRH5Gav3gIjyqFUOkQzJR/bGhLeRI9TSuqYR924VWnhGrPKJxVIo+yXznQF3XaWzg
kBKCCeM8gEu1c8lDb6xMNMZFIz8C9RrK6+j9uVX8xctx6gRF4z6+iFBJQYuq9V5J7p997/6DUD6H
KVq78FWkyo8CVqAcZ69EO9RBZu/wbRhcdepEsX/n76QSe//uOndDEwu5Hd0JKS92rE9qjRaF89m4
lrpb8YkGFG7y01ESkyK0P4Nb7oWGVdhScG5LvLhc0bnSlRrfij46P9616M3+K0+Rd50gq3E3P8ye
wixkqz6HWLzS5HDajkaJQsONDA9gADi6tmUFLS2s/gSrrY3+w7KLVNFbbM55oL9jDKC3er/swAkW
i9sFLWw0d6qQEJXawRIsC9yA0gdu8QQPGyZ++yDA3P6vaHOjQFzowj6t5yu7RPle0ZYjK7gq1d8j
Da4iGtd0w/xqy+yTbWm0L/m4+g15XJTywt2BZXsdGVlMJsJ2N1NNlCcgZz+gzpLx2cZVBzHQbAv9
vDtGEgVWySYy0Fqr0xrAQoX/jCrkRhrY0e53tnmVynjqQw31gSUujEpme9obLHYnU3FxOLzzJRbF
HAjUoCajReebkehgq+aMsfKq566+X/mYxXuD74T3TQYrLKH2x5Hj4bFig660GudxfcdgyUlVTqsk
21z2AqN7SzDb/JsZwEZ7R8ryB6sIvJyYsB0tIm4u8VrqzhiUWiGQ/TQhOgqbFy69m34SJ4iZYGxR
KIuQSTdqar0lI2QD5Mrm86Y5jiK3GX4BOEMsViPKPICii//gysj8a1uPOlv8ecMnzh42e8Rj8u9t
9gCYAAllhQJlHVVZ0N6JQyvLREMk6WQttVfc/71BvOMwPK4PrTZr9HG9FO/+m8AmBGx/cz7ysIUr
Dew2u5YGxUdbsbivtEWQjkMHyDW+uQtgRe+h2BJ3t7A4ccbze8XWdNXr1DwxBmK3nWErhJTieGsE
ZrFKRMjDVPeFdnTaXpdbM+XlXzHcLYxvroo0V7XBrWM1f1LPxTxFvyAesYbbulWOui22xsUEXQH5
hwaLAzL0ESKkdS/STWKBavWh4yptlsUfxgJC9NDDi5bApAO+FQfvcWeRsgJOh0EHMDpGnfGplFvm
Uji3c33gWg61H8DL0JnplsRCLkGHGG1og8KK7YjZ9yqjL2kTAWzJI3qMik4X7IZD9QfpVgs6bDmz
8WzIyXRvt3NkMCLRULrPw/mUqqpNJPsQEso5ltj1FvtXCa2DFBj6hnU3Qed99iz1xcGZSf+T+58f
FEoWBhDsqz3IVoGf+hpAMQo7gkqWB90iwmvppBKokMBCQ6ujF8xKFcFo1821GiLYojembE0ZWiwn
CtxMuTi4H+MLsa5fKD1Uivv47oLJRrPslZ2gXH92M8yIpqJBEh5u7L1PsifAJIuswIE4xA1jjEhy
DIRLLn9q+oR7KwHrcu0cgc9WuMdkY4UKg0HcFGF3lljRNewhMCX6ahlEfC6JWH4VPngZYeiBS/b6
Vm9+UwbmjK/6dtXKx/IZmjkzmP37n7sycFW0ZXYwvZJomRR5KsjbUUA2ijhmQ+9PkXleSwzELxlB
ukr8A+i7h4DpBk3n4x7lREJ9VoaJpjKFRgvL6U93NUCs+ccWR5Ml4RHr9FWSTBKTn2qF/xTL9ZjV
/aRmKVYYDKEPOj4GIDLOmBydN+nqv8yZmPSf/RhOvhF99HQsXzDv5a+OamaR8w1aqFLWh49+OhOc
9mWnl2ffRfbx1qi5sDjXcPaijEESB2uCuQ1lL+D6kYhVwrmQt/3wSR3Rbe9rd5wqBzTixNzBlsNj
mg3zt1HuQGJp7ZePlXFep2fGBOq1bfrdyxz21ueYrLS83Zo/Ko/H2kQTgbepLuopRQoO9X3H5di3
CYPCIlOv5m2tze77c44iiuF7Al3tqwmCTu43wkBVEVw24Lr0PiBjhXkovEUqScxe2sXD00itRcUP
3orUyiWmP9PZytTZLqebpTZXROcEo3poZODj7TjwqhlfsET6ro4Xg63ANEIs+wjOZGzMrq1ifh6W
wPoIaSB34CUsYPPxVuJqyJIlfntYDSHa6QreY2mOwmgXoZKd+By1SzpdkNiQxftKz0Odj6sI7YBV
VX0g1i7AS7FtDD03/0QZgQVANqsrvNZiG+4LiGYU+Zi4EwvAxI3jvtlO7ratBPCvIiYZ0WWy5f84
YeB2bfFnE/L1qV/pMdPxP69hrXLhkFbVYMi+CFRkThtteOtVpXogxhsCdrnvhZZkz7MsSu+qaLo2
ACNjdr4azANcQ5y/6ELZIL29IBjiHwspqLuagBy7I7WOx/g1dOV+tDlqd+BdkfM6FMpAR0lM3fGr
0f/eO2WUiwLao/suxn7Sl2mVMjX6D+XOj84wx3S5yV50252Joh8kUEXfTnFU55Ytha3b+VQN1Qc4
yFCpYQEXkiTNt2hsubzldG+2kcSkeODLBadPV/JgCXGolXfor47mtanSaZFx8OQ3mH2gwR8l1dLK
AhcyUE2ezcoaB6l1Kx/mcJtVMZHiCb92PTSc32zsBVRrknBN0bTTsT3FSswN5OesAY096inRwu57
X7xh2kKGQXFxaBPKEPh1OpVfLX1vHCPFiNplGt0iGA6Oqzs/ZRsFFu17BBymLHjHQZukRwIL1NNb
b5jO4fmzv/Rfb/HtKxJRs3ErM1zcpCglVMIDm+5DSuiQHI2cc0cb9sKGdpt7XwCD2MAmRQgkojK4
gs7+3h7bHMR0eS2ykINWWZX8VUMSJZtattrHC8uo8Nlwha8muLoRP1+bp3r5hmFGiPgJPEr+Lo9X
MENz2xycqTfCG5pGbKvUfeAYWrbPe+cTJSZBdznLrPjGmjEJCL1avsq2d1R6G1YFdV1sFNC2BH3D
VpuIHAKiNDzJ5J3a1KrPjzcMFb8Zm/3erRZyuSgTRSWgGxcp6TZ3VdJ8FImHzpFeWzGp6MqtkDLd
K4ytkRwiZ0aDwpBAZ/WKH2gUeEhGzPLa6cyMX6r1UgvRC+HdAjNrpKer+zkk3zeNEXo7IVJ+pLYd
JV4hmqxWeOckutneRWSgZcjirCu1uXvAGkWneMLdcXYN5YcPqJLrnZj6kEKNqA8nXW/kL8HHh0YW
0sc1pzvR6urec2ZxMh2OYw0fn3YsBxICzMDRTm2KqqpHomPi6wsND4+bM9gAeiIjzf0XgpVqaj+H
DwFe6LNHrwq8SjRY+OTqhTCt9VRrlkCcALPx0P9/7FUNMfT8qb6yccE0r6DDfc1PQIT/0yGUp9rS
rGGF2RrJG2EdNDq2qlU9yUOe69N0XgyW+4oOJYtU7Z7oDjOtyzHIH3eR5UepmBggrbflk42PdhEr
cebdERhAbydW7OPyfhlHn8/UMYCh3gDYFs68iEQoioDnl1pmXG9UKM7y3JuKEn4JWoowSP0dXLNu
WEeVCCIFvOQ+zaS3MGBP8oggJdQmhXF4tENywYw+6tf+HEO0yNO02nlOk8MOlBwx8jJE9JD0dL/s
Qm29aWd3Z72BS0892fJ4CoRS5VNPpc6z2odCapIzah/2LBRItvWJ8CYQilS2q+6UvEWYgVGPXJcz
GzqWGJ+LBI2dEUs8JTkVmgT6yNNPp8xSEp0vfbx88tyyPcaTgAM8/qhuyHFvAsFyemo0Ajzf+Xmw
qlyHo0ncZV2z4v23xfiRwAfnLfLhzVLWfj0Fh9CJKPLHOQ2HNFlq4JOf0es6WkhvXeG/cxnfeeMD
xqTsB/pEGjjMecTfNji4UjuaoJy/0FGOdrAOw8cGF15DQL+6BL1b6yfuNh1NMU92XyKel7FAJuGZ
/bPzRF16WdCYYxBqYvfn4PK07TH5ZT3hsnboMfzPiZ94Cx8Fetj2j4JptnJ37w1YfMl8ZER1WMhg
AXqrn/mnfm5mrfN53/8JcLxrYoeGx/1d2mLq82Si0ofKg5iArzKWtAxHxes65A9JIjmXD3m6haOY
WPMyZMUarM7+BEgRn0Xq1M5w8Vk1CFJ2VXEE44hsGAAX6rha7uthKw2yLfAnd92HJDYPBLLhWTGA
SnPH5BOgnbXsMxXGMPQ5xZHclDXpFbz5PAnIGF1u0QEVV1AlUkkeeRkXZecgfsJTz8mdWcnHQSu7
8H8LAc/pNVkOgzH+2FJqgK/Ihr5VEsviQ1Ts5RUgmFn/9itS68NW5flEYdFjIsCwccn8i0vjY9QG
BwyhzJvuVRtTV4aT12/B3y1os1gta4aYIg7AZmD2ZlN6kF057Vt26kJwqrYA6CzLxbR1sKP4q7qS
JWyJw5jrSP+Z5CjMvWwnhBO8CXjt2JZKnKeJ/0W8qWG2BnR/LoTI3T79tMKN+Hjr59Y3u3YZapYo
vb8PAQBoJrfjCTyfM9AXcFr/anPAyW1BvUGRjaUf6dP82yh0r5JLoMvaJJaKmSlr8iqTxF9oh+NS
fxKMvW/dUjEHQRErPkLmod9N9k8+xMBay/+Mee27z1YO4N8b8vyk0k8AnbFN7cOJYuz7QVe02B9l
MQSc49ZL+GP4gAxTLjUPnd3qmXFH2r6CZFBvRTIr1qodkGwSzQOooXBqUgoZPgWQA/qJ7hB+tg88
0+zaehJx3cBJ50POyY9wmeHU6Nk3ZcxeARefLiqVN4Jt7CQUGZk5i6lkleXDindibBsILM7ySdLS
Y1FPeXD13MRJAzXFxY2XBbNwLSXxPmkEJbpK3hTxtEMM9lZJ4TLUVJ3kklqm232vT64n51jWBFiC
ZYqRuHvnUUHU85Yf5hmaXBIATQYJjVPWvXSNb2ZNnpqFdl6GqgHC6+5lQ0jddg9huwa8x+Odbeh2
XjKmOvU4kupK15U9o1mMY33G2g+uABon/zkJL5nfHY1++ThfcEBvwKN7pTnbO9YSvv1jKN6W68AD
+IYrn9Kb5zYeMWmzxQvAI5f7iE81/r8e83A14MwhcNNoBJqXlZfqhszQZbUzWQ0/PUSbi48VIPnx
+9fQQuJkCWHBNCC5qJoCUXOUhSXsjIy0mXNteC6naN0dt5OclmGmWr/Gesyt25yR4sPEyVF5sUrQ
uF5WGsBhNLPz23T7Dsyb51AT2/e0lCWsICo6/T+7KZpHo3bUSDb+H3aRRX2Pe64Z0lUcSAm/1qNo
KTP+mFuIZlFGu0lvn/DXq79SjLRguXBn9tO0QaELzdkbaEz7qo24Laj3lVcymmNpFgy/El0G1Wxy
AgXrwMU7YUTl4j3zyxOP6pIWzs4Y0KFrZjQUM7QyV903O89GgYO1dEjO6827L05MfpVPnEW5q6T/
wMOVnAn1yb0SXUJq+zoIgkOkj96dz5Qk7X3u54y4QvzK/M9wfKwQS1+rW3Hl8jR0gIpDBkKwos0S
EY7LvEijCNThn2ci0em9pi4jaGXDaQo1y/RTTJmVkzwssdEjU2qJatco9bz521TOesEEr9cMmJFX
shbmntkrUfVICiqlrH8LrIfk1pX+Kx9u9YmyReStw5C1nofXk2QHL/f4wZGOHB/3X09osksaoDo9
GsiKiod5jgDs+tmumZLDLYONKHQLkhDosiYcgibCA3zDp/NTezjK4ByLbKxwWmsUBvzuDZkTAScZ
hIYYkhFUWrY1eXdM40/ZpUGWFDa3Lj97Xj7cGJdHU32IxIr2nekishn2zuySe9Y3zbvTB9ytYyre
/E9hzAQyppTaEboloCFc6dJShIwPGB6yNV4YhkrclxiBlD6/1NN8gpWVLBoJ0QrfaBmW25K0aBWC
oOGhEzQX0DrV6mEX+THC5P9nBMo4mLIzpHSqQCf+EFu3RvKxiU1ZWr8oEecZQMiNKQWLYV4rQEBv
KX15SwBsxioKF+Lxkgewn54s95HL3lEevf3hene0Lhub65H6ZzdN+6vHU1+SQfb1bW4fXduAxt4y
zrO0Sf+TgKsnY/emQPZKeE8aa/X3TG3H4UtgXLVNxzigcT+3PpXBtWSyNdkNEMFUJ94t4MNcXbzz
Ne1JRddJQvB4+GOIKDC+7gK+/6XTC0EIG/Hp2vkaa/HSVuSjdAMQ4jx84ZszFST9HX1SCgDktJVn
JIoiVZg6I+dSfNbaiPckbUayIG0+n+lZ9QoIj/e/TOhVVIyt+JwXAmsKuoHQu24+4YeWAk24P+s8
ci2FztYKDSeDssnRjg4wAY8wsIXrSTjFCC6QClU9J8Qz9P0Ia33ypx7lTXrAy1heL36rtXK9Q7eq
S67SY6ztDm3F0OQ6EPd5G5X1pLJCKtpjd0Ou3kAvRok1v9IfcatnDPabTdudp/BUL6vYA7SH/k/x
eCNdyjV9E0C21lJnSCgGJSB/vJjP6bkNWB6+GNdo1lRIYmq4hJl3VqkHTTgp/0oEF8fs37aFB6Dp
Ca6KnM9nM5rAvYWvez0I3NqBzkQHBnn6HefQa+r9gNq8gEuu/+t9FNSq/3hd1JOXCcaoMQvbi+n6
esLs347fEbI3S8GwHsJJF0T8j0m7TrKh4idj5n/PibRmXfG4Umm8AlvfXuDzHhlo3guksPxMdxEb
ant60li0O3ef9ZQqNJ43+w4W9W5o39f0n/W4BoGP1zEFBy7sr8fm0AYmO0RU7VHEOGWYJmhshWWk
JbXZK7inqX7vvuBgN38ATsO0/fPVA6WgRuvhZgC8UnU83sxiQzIYinhJplk0mp9YBNwjSVtwRIg2
jHK3VvTDhyI2ZW3eRhqMnqazKfSdq3sy2hrv0wePKEZQhUSIVMO+1O6m7eLO0EmepSjNuS/8kBnb
yQ/V2xTVf8tXkxksH56swQbaMVbZWEmBflZd9RnrUOEwpKQTucRqoPrGILFlCVBPIO69LclNpnjp
Bgk+QdfHH2egEbzbcQaZ94NGOccNR0Mj1Dwo7iDg9JQhfAy6mFBCYWo/F3TWWk33c+i3EtbppOWT
M7n+fbwRgEHerAomn1ad1BlrV1h6kIT7QqCImR7AI8+r8qi4FeSUSXUIoaCc3jjiezRxOdXOed42
dZajSE1uxJFSpKKK8q8iL7B2YZcmVOMIn3WQ8Du97MNGrTkCjTNTm1ihML3nnB0nO96GyTZOzGqx
u62aZiaeLbhV80fr6iwKE9czjVSOkvm6I6iCTsgXMKwxF7YAGMW0y8UaS+eyiI9GBhiqZWbB6xqQ
UkQ/+qqC3zkrPIzkvNvfMoiBDPjfhSaNXKNGmwjhxJbkAE3CIi8UwIku+yOF/p8l1RvrLNFtm603
1n32YEN7oYpTtH5/MmuAqPpIJ1961/+Q4Fw8LoYyLa5rvze8XvO6qXhDLJ1XS4naVFAuwJTG76C+
c9G0bI5313AK2VFGi3qdigjhy6a3SD4fA/IhA3alFQ1o1cxlkUG9u4JSXPtLErgsyNavAO5Pn+2L
v6bTlFgKYX4q6kjfMZxldrpwvt868KfSMG4p9pHlWt51/a0zLR8L0rpbH0SUFo++odev376xtb38
VFcnCWBxIMS8chTa4MDfajZWYOBxQcZITZV/S1XzmFZeydVmdsFgOHhtNMzjQP97uRpN1Unv846+
PQeaMmE0vQUDlEt4nVmV28s1dpSjlJznM0IoQf9nTh1ahsyjoK4b5fNtLdxU54bKc+uc3B9oTaVj
jx/3kWURfK1AFZIy/gjVC+xrI2nYQTm8DtPZbR3ygUgh90HHlIS+DOnQobMRrQA/aU1rbPBGb3OK
SNplYlRyRKFy67GiuMxGshjGjPovI6zu8yetox7vvOyBOlN3uOntWt/JjkTLSqrzRYR4Lzx/7jkr
gFqqOXkO/gXSSwYO6L7Lxcc1Th+0m3N11ulqZXxdyr3TIxXZ9NNwgPAO6t69VPULLs+UIK5rZ8pm
pPtGTLaQNmUHc9A/+lEL1fi7QYtvU4w3pf/nlelWPdUFAYgAUOvsWZUjRT7Oi/ebtuycCLQROE4s
Hmard5IOXbDTyKxZQ/QhzRsOQi/aGa4T79sTiOoQH4FZiv2VtvPfn3P9Yo2oL5D6cRpGXQDtJirh
rQYqcfBEUGlRC3+rK8nyX1RC2P8AAAs76exhT+mhUj4KJH8205I3A2jbzMKNwTDbg5/UF+T2l0Gz
Upn0fC0eoZqoEEtZVjkMjSZ4P+bQNhq/4AvzKDH5HRMbO7psVDMepZ+nuCeHLBHHg5NP06p4ABiC
cx4X0X0t7liHvj8NNzzZ01OqrZ07FAmFDQ4SlAZtm/OSwaIGieEZJ8UVgM5JtKOesHj/gFb+dbHz
1U5V9F53s9k/VslrkxgMS2c3fK6yp7jZ0+a71VrLW8SV8HvhUvxQQaGynPG2Knt49relq1H0W5P7
p3XJFa9HotyXwPfIWMRzzMKrC4+heDxGcXHaB6cYu0QrL+asGaLYfP6+D+WX0dFZ94sQ17Eol9eB
QpmcFDqlzJLK3tvv1fp2qI1le7Z8fVibu2uHdv4t+qayzNqGdBV44csiZY1iqlKHUWsAQCm0EBK9
KV91UemiDAUhA2KSsu6lMHsK7uLO3dFabN961MjNSMaEgxmTgrjqsOvEOS7XO8zI7V+1GaAmTfHA
gl7p9R7oa1/1HX9Uy3lwoTnBJ8DFWZTQlVB8TVgqgW9T86Y5OVUA790vZA8SHrykZ4G5JVaObOAe
lmyFqDYD+PK3mPnuk7MJMoiBTCa6NRdwaRcBDuTIoDvvXsAR+jnjTvcf3sNyXuS375zq6zt38+j3
RjHM5hA1ecQYyxLLkLPDkHGE60MggzWDNOdV2Wcvw2tC8YkVWbXrC0yyFeTjeRz5ftlvxVARD8bj
WVFLVUzzPNtIJL/AVU/5T8W7Bzm80yXgR+OKWZHGUHLafRkUK7mgjCuHhBJqDoZTlQG7HmvJSsNg
5Yt0ujtxCh810cK+2JyIACukBpJolnjsIDIpzPLE+0vB2edghKRKCuXQ+4qgO/PBuucmUHyNzAc9
DoINHPab8lAQbL/orGaIEzAikOIjmaTB3GOxMSPVyvh/ii0JZ2F8/BBOxPMN6J2p7sYOeSWD5A7i
LhjmuHuAJxVxpayLouO6xxRrqXD/P5QQelWpj1J6QjAEDF4Na8Hw4TZAwvfCH1pBpxWq4yU4fdoZ
Ka2LEiD18ona1Wit1lol/QQWQJC4+G5rIug8rVB4I5zulPBqF0XErwPJif+w9Lvl6U/0c5VDQhB2
4gSQcehjiG1TIikRrcDNpZl8RY9k2K98h/PEA837QNbL3yWaEcNin4ZBk53GPWsNcRSnDkEyirdR
MWyTsRP+QFlOTnJ1LtjgkqLNQdHexg5jsyeAm0hn0kKqlEBvqiczZIGInKUungXHTHnTjNMzWHJ6
7BcquOxA4FnjfICuBXPgLGzYiCxGkzHVwhkItGLnoiE+Vk8Ejs4LsXss+RiIm+54BcXNngIIlsPK
q7znso08SakKR7WxfXRYotPH7otM2katbOVNe1Iks7bzVcgS2fHgBGpQIF5yZUpLd9JEF3PWVHCT
IcWGjNHCU0/0cueqSS/T0i7BEy0ndoZ6KnG2P/Wy2fMhoK3m/Ww/SZF6VO3wh2OecBzcv+0ns1h+
sKtmSlFEPxLDKp89zs5RflfzAIHBIcw4kbm6pJHmigL7GpQrgInngBUZ6LhdLWapRcv2BVYMkozq
myT1w0TvqZFxfnA+to3Jil6y2H8bjFWQdl08Utvf4BOGfUiu+0RCmpYwy/a2pUXpBbTzThxMXeFf
ehkFVGbhIwTV6A3MP6yCm3OyaJFLaarCrtk2+b5tPjvYCir5M8Ais7pgW34WO8YaahNwcvOgFrho
gVofjj0LL/OMv8jAxBMkcgPIAH2lzC8eYuWJPy6PrxejfNepN7SICAi+L4Rc741jvLN2tFAE7PrM
G1rsYp5vvn0kCtOdyXUz3NWRhsJoYXu8gY9QbKqmzrcKN+0CqIk5HYdqi+KXyJA7P1wdNfws/0N0
mC4s8ucV4lBT49UzsS2Zd7Nmd2rGMf8ysK4Jd6fkyb7byMU+e7CEVwHF916uNFFZ+XIL8hvcQMVs
7UdBZ36SY3mgp2BHEGrQUm/7SWPgO6g++6oaJQILcy31YYUVuMJQV2RInnDhG4ahk8yfsgAfU8Oy
Hv9emLk2iwDfirwDxhR2emjDfBLz5bqkmbjy0xCuiYEMqc4ga4psWwGfY6T+8aHBRCmNN6DWAKv2
HHg9Vw2Br+Cv2kI5Y8yvxbi3KUUg7LsU9Pvndlj3saFtM5aMYYypO5LfcIMbWnJmQg56mIlqT+dv
rztqohoGYKNsQlBBxTLenteq0U3SyTdq2OhbRz2fGMm/GEKsrDtKplXK+4lMuEPS5N00r2OwJ859
f1PBq7gMbkGcudPT8D7b8k7DCnEtfYWJIr4uLAGbRgM9RxJnJnrqbhVANSbSxCO5Ipp5h0daSbQs
6/j7Bf7CRDayq8cluYuzHfiCa1reYuVVIQOgqA800hskU9UsWGRJzB8kmqeQBiqncJsXgfFz5pZ2
/khDuVKmh0ErDPcwtFd8ILp601gjhZ/bEkWfghxmtZjBpEDJ2xqjUTASXmhHJDZ/LhQt1hvP3KE2
aQdUaFB5/fIpZiRCoTJjHwlOYHc/8roSIhcT9+n1D2gAdTEzmoUTMUu3zw4vJck775ZPIPFvzOy6
QvYx6zuBVBVx6MFdaCVovL09rU3jbB0u5i8YyZbe/AYD9Oeo6lEm6A85QQ1tUWylb2LPOcWKSsuZ
Cr5eQBPaNLnFfOeKUtyJxmkgAQjTivNzz+qaMCQ65Kq3jKHaVcYydyZHBEmL9aANh5pda1D3TrBT
gRAfq2nbv47HW9JMVeBbQZWf8C0vD1RecN1KlnmHkPqsA96ib58A7ZyzDcn1mETpiX1oSZa47CAQ
VMDQAzEgQLq9jdzeMmgmpdaYpdhrzJ/jd0ROE/LR6gNDCfdUXn3XbXl9vcdShPt2mVRAMLWUpqdO
vzsBLvLjdMQFqyLX12NrpPpbXbEGPF0LbNh0CFrHqz1CCQIYk7uWC3DOlwF54GWpVSlsnWBM8VEG
UCCcZaTVpemC6BQEtv8YMbTGUD+GKqhwulaaMEgG0i/rKwVWwy7KBv1G+KINHeRLosvUKHu4ulWi
hMSpNE+xII0hFwYrr9ihMsh7w6sLTqKHejzII+PY2MzvgcxiCF6p6ot4LEAOY+dvZbN5QuWm0sfB
fltH6A4PFr3FzlayABxCOqIklXN2/MT4xJeMBKlFD4sXIPoRlVF6YglcQ5KJfrS/PidpXGCKJsmp
yl63u6uaw3O1Mpznlp10PIhfEZoXc96kuPlT5clXIEttkr73kI7KMkzkVJydTfgqfG5vz6i87pAN
oNDW31K0ZwLi/xOHZS3Bep1lVKLQITA/wAUaqOdzpj4PLMhvb9DDMawBpYIoyWX8PUfpNW8QhSbr
js2MzP/erewBi+2281UGwZyg3XeUBGEzynS6H02Y/WRkdAhXhOzGLeuG3wElGotF+KegBzg9gqg7
Ai1xIBRAeET4maOGGo3m4X/GPgMVLEDPVe6nZZuSAK4OpfOh7246gT6Y0Eur4hP6AqaPuNkCpD7I
n/lcU0Jog33VyiyH1gSyyCTZ3cGUew+qWvJzEtlPNeX2u5VPGu9WdVfcnS4kyei3KV88JaH0zzUA
kpqAC0t+738lZ7dL2FkWMO/0Kgyq/vo8BzyPKP9S1fYyUzT/ZgxfKFOovkBkydkLM0ahmKbtcJLC
k9Dw4chnVKeJ4lZM3fDmGpYFld0Mr5JM4rO3gQUCugH4RBRpNGYgI6IH79e9unQ2Hhvsmz4hRzC0
2RBL7fuSnLillZDB6QM+lqw1hGsW+W1IBg9s9k8UfmKxSRZ/8kjJQjor6oRNJRrqSVROWize6ygx
y+f/JBJtgjVpVQUp5/s6z9H+CnRgupgJK6WhDlaC9+NlqDmlQzQUbpjOl6VW9JC/ahnW3UZikjsh
IDDXEcV+PO5SCAoThYMZkGPfMhRHOIYvNMtHfNcEQtf9VqeRBC+sHfEpmoynzwjwX93txLdchIbg
73Qa3s7zBSR2f84h5OsAF+dc3G7tn2hGIGgTsf4vIXJ5fW6l+LlaTn6CEOAbmelK6LI+7xU54y9O
t8GKyx5hVscvbSzi9TE9JaZjcYucXTUHzxCZppay4INPgeDNdaWVQFswhy/WoSXqHfSUjiWWzm9M
rWcfATs5mQsaOLD4rUM3S/tJ2y/pH+mGT/YGgSJcj311X+jxiZ5RfYqLPUVUAT8FF8zMw5uVEqDQ
pTK1ia+V7T4WB3DN+rM9fjM7JR58sXNdOZtmj8aMC5Leqnv8TotW7A7E1db8QfUyFhE8SLVfHp94
hRT/Y71Kpwl33vB8MC482KzLDQzZluEhXU9Apq9nKotGSMe5UQvTos3ne/5nkaGYFSZ6xNK98S0E
epzwj4ky2Mqe9wYcrvYthuG9CM4hLxmbuo7O6gH0parXufM/DJchJuu0myFszHnnxK6cHbdRL8nz
f5U69uJow0A7p+HT4lkxi/qFwqSogXqKGXY/du0id0Kok8C/VgnXMIBf2LQrlRWLWI4JcNtBMPCI
CpJHGchY0INmJd7rEhPEQJdY6XikqtICWpPs38t9wDO3VKwAdO3bN5T8iEk++LfhGRHqITB8HlSF
QRen+RqLzC026vr8GgPCZlSRQnmV+8OTlzKlFrM/P/j8KNDAUN7T6AzgkofPmq28cQ+UDrh9fwcT
VA+BHdZLJH1cXxnk5oAf/Cv/I9J7W6G/Vd60lPp9Q81Ng/g2Lcjf4MLwRG1Y+aEGoooXx7axXCTa
UfAAwXq+JRHJHQ8l0o2NrcDHMvNgw7L8HdFiqYwzvT+cJblPiX6gTSnBzx8KEYTNX5LLZMD9z438
wXWunyNCZqpmTp4mMwx+WKOLDQUKgj2J9v7KttWE0RZtv7q/Lx01q84rK0bWgaCkzY64fZp8x3F3
GfTPHCIp7Gku4cOyJMx8PqS1tTW/vnKMe91NsK1RqKN7k66t/KSG0d0TFyMb9dnSuiHI272Obgyn
4eOV4IGzVwLUlMJy0cWPyoyJxTY03/Ipbpi0PhVqBtyD0UuZPg+M20Oa9qkyaiqQJPsOEF8b1Hhz
+nJZCrrO+BDS5vl6NjT8aT6l+eHtIiDu6gl/0BmlHsgbD6kc/iIxuqeQWPzeNDsfqz+ScrXEnGy2
izw/B2eHhYjAvI2tHa+B7pwx2uyyUrAmkPzwhT09f5fzqgVT19pTCpB74rYz9mr07UqxZSufGzXP
OTD2q66WXyghLt53pAbOAQVWSBFnuxiev4wZpirLxd6XMgoZet4zhfwJdTFKOYnIEHSSYUl7Ll8u
IWPULOFp3JLqcAZewr9woRiyuyeD8CJoeo3QM029Gjo0oy+AGo+3IWu+pw3jIwG2m/lnnE/N3eIU
bPZZmhSxccVRlHU9eZ0Ue/UvE5WnJzqDau9kFsvdYbAqfbftGxjuhzRmfjoljf7kUCaK3tWV35H9
uRA/1fzdAKTBTNJZirG5ZbtlLKcL6OsPQTHUL0sJHxdEwLeWIM3tlX6DinKUa4qkwwQKbOVPpeHS
WF71RgaRUN2f5EWtBcournSCkNxHhuKpBHu6IHSHw+3fRlhqop9LOcD5CvQOUsMaUWp2GkoP1FHN
NrsJuy7LkZ/bvt2WKBBqkOhYbeplSIScV+f05GNJqxZn4AUB8+LsFXqIRRkd11PSGmFRXhG1icIP
zx/5rZwnKkRMXCzz6cYCHlxZFXOCI5cP1w8YfB1OFCluAlsOSJ9VGlvglhf26RKxbQZVhzfJgoV7
qCHzXm9qIFu9E7K0NY755wDdyA2V3jW+G70X9jAdFb0kFUUOA1p5wWJAVXeaxAR9i1OJ0QLMzZC1
nH3RLJZXQPX6NThkJYsFU/lq1U81OzCEeMvLULftXWW1d/b2sGsde2Dh+GaEHVPPO6rBK1Qy+Zfk
R8XUj+Q+JkQUEU1qBlMUMFlPPBaJZuseqVhCygFdb8dGa1i8U4CkRV/8Zg2N9pXQ3RZfNLJnunW0
sjKMXmlJqVXePJxvclGoZVLMrvmRD1PkQaT1DOkYQUxuhr3mawjAILOWQO2Ml38HbJHhCcFG43VV
Uz5xSdc1GQtH2ErrXOjU5gXqEClN52RiWS23qI1jjxQF2kBm4XA/AwSHY9KclCWRK4abWrNuZW6Y
hHOjp1i7SxQtVVC3nZPrmPQq081v3l2Z0Lr68y4NX19DDQKVbnTcA1WLCseB6rQRzGQjE8L0PaVU
MbNCTdD8r1QBX0/1kNlYozIZRLbN1mPHY0C1D23xamleoiXlAxh2tgto/xcpEz75QZH+dhQzQ8Jm
GqtLOlvHrg0hjhpIkhi1dAc7ctS5SA0GI9WyZss0rUs9KKwwj8Mr4bT7OHCrrTXSt/Lx5N7TveS2
b9QQnoebR1OspG22gcp/MdrrSF8wzKFsCGwxXx7llh/Qjg5YEY0FjcSb2yTyVxT3nce9jfB5Ovwj
FtrRGimrpXF/A1pcprgAoKV/gP1TwQaRxpXQZjRO1uV6CrkgjS2G24bRSnyqrOV0Wjq5s/OIlwe9
Tvce/Pwxv5YAdheSqcSAmb/3++YYHvJt/SDJS1WH2Oq99jdh+LA0aYPQQv3z0gP1nVEc0xCLYCRf
83PSCF1j7wfR99Ms/0MIrZW/mRjvenLUW516gXarHqNIYm+cIZ+SaO6bEqSZ6Dxcl+KEteyTLQBs
TcxoW834Ur+nOnlNVwJh7AOgpq5aG8MXFocvmJNC3oG5OULVCWVkY0gNsbtHhEz8Ek/05rwNtdiv
RpRp03oytfveX65PnwqArxko2j82cK4U8zB6qzzb8tFlufS7TNiuPlUuDk67YUMeVOC8Mu+Yu+e5
UQkIZ2MZjP8ofykNSrQsMFF/7d9x7Jg3E2qKgSKrf1Uz2kzGRIzxYq0Nc9ng+cmUO4U/RkbwoAK/
/KiKc72in347SOURW2W4J5Eh1kBldYHA9L1/BOdRo68/QJBHdNDgUos3hFMxgnTIMwgcQeG5nwkT
LQvLZqKFdBzaTZ6JxLyqgoAaEnH8Lh3CSeikmLipJgPpz3BCsTbtbgkPCj4jEk8nT0zak7OOO93Y
awjO+0cIxZ2M+RM2pFYYIpGP8gJwrzVXcyyDR1yfOvRwppbV+wGDmiN8rEvpjxlwR691H8kHh053
nwkir0xyN5Tjck4szeYD9YFsh4k1qqxfCrlTnRPa9oY5MqAnr1w9sygBC88v+fuNyWs1U2KpP1IK
cn48hfmF57QjquPKom/mqaEWzU7xeHMTKfJ1vzVEnC4HZPTaLDmtz+ylV4kuzwluhZfvvqpXcIbC
kXDgDifk+RYpeKDzlVyYjnDLRTr3uFWR3+Y0ZfOBjh5HOIUgc0ePM8lhNfMcAVIoWH4AgeIkPeCD
RSo8bsOvqEW6RHHCk6PDWZSKzBHkZImubM1gdBqwtv+FE3meUC96dOgOlHhHq6JXaUReK6Bx3+mX
qsjHp4UwksO5mkcWEhLSTsyupYQxwrcuHE6aRklGp0nWXup0hoF8zCj/jq0XDDvoPPJbzR3E0HxO
pwW+/warOUmxsoTPZ7Ke0QPWAdOWOKg4pvw+5rt/XE8jUPiDog3v7ptKbDp60oKgjFlAIpVEeoER
hzwhe4PJ/POVD7/Ym5zAiyZsjg8g16fENIwqQNptSLciMqAVTaAF5wnIiNE2+I9xkgCAjuXPWuGS
TP/D5VUi4+4DgJZYixA8odY4ei7uvZverYvXoP0JaQwd3mISqlWYlS4gG5xFa8Jcbz/amYFgZUL/
xIJkpHJ8elq2oW9xvp4zoIzd1vUkt7doSlQ3uOds7jh1Lrd7bTHp3tyfcPe8GtnONSUnwzIK8j3F
OKnqgFcJkaXQpDxA8bTOcIy0eh+uKurEFu31qZh0T0YCk1do9Tk7FJtRm2CcpSdCFyDAzC2KNwPx
sB9MtS8yYCvz1YV9DzeD5bsKpVG5qdWHHwG3xHXKvkfV2kndILtKKLeg6plmD3zBYf2r53HZTtmU
6d9prHUnIIKe5ea3PZP/SagvwyZV9f3EI4PoIZ5pCkfc04qdnNKLvv8XAs2uaaRZyUf2OPD4GxNU
BsRTMTOdrligeI/IlpXaEQx4BHsR9E98Kh2k2uRQQl92lHn/fEgmTCY5mvRLF2kaBnnTPOHE3a0R
mt3+PLf3M0qknjr4Uge5naeauRCC5tGIgyVjt3KWeJBRNbuthwsM8Oau2fmIKqYv/Iz9KpMZTm8y
7ojQXxaei40MGnCmm4/dmIKvPu2ECYYR/0VYRNxy+Hr40kzpP854OYqLEzeHh2Ue+sFtzRn8jhZt
n+5L8eLoYO9nm4drw2nZ5CuyfogfAUS2uYk48ypeDWvcvvEQF9z3i6sto0l/sYrCeIoBc8hHyRPu
1A596okMf7GgHnMdGwfP8BfJU3SsHrZLfjqNjLMdEuju8g6Aev+fXrZf/wE0bemTEzKwi/YT9Jqv
1NmEYLzjniXzDh8hu+hRE/M51Kme+FeSZjHKjxm+Y3OHGhpieUhYp4lZrw3mgqkOGqkTyC9pdiIj
bzI9OQHNTK+zDOvuw3SBQddLYp1f6HBN3Pdh8DEMlQa7M2Tk6nwQPswSEAZKcok/5fozdPAXPkuk
hZiU2apv2yQOqbUkuhLyVca4t3FYJEPqurCtLTJvIP69sb+aeoGpLTuUUXC5mPW+cjKEQUcmElA+
qeJeCDLZOfqOkFA/B35cTAP3tCRS3cVFn5BeKp1nE11Y7K6T/jHCB7Kw3TlKa5NCfiLwm0otN4QH
gCqMrJr3CNOUOozFXKO62qqzDmQKTM4DAiz5DwqeS4w7xCeRSCxfURSswQAbzOLGSlYvwcnjd5Lc
9zhDUUgev7SDV25bM2qQa+6kbBweqDbViADr6H0/5kLxKjVX0ZscyI03/HPXExSgYB1AogGS3E1A
Hae6mrO4qFcNMRn7UryqP7vuuG7gOHz5nZ/BvlHODhcvv+kqmehb3bprelj1Iq9eOGse/zkC8GlD
ics1mF+MXF4/Pam1ZP/SLetKvaOeNZdzApm3Z7Dvx/PBKM+jehyKpXiDQHZO6qzvGGsP1ehnKSjF
rkxxcEVdmiJqlpXF6544IdCLV+z+E5rw/HWtMbNU4q1o4V6v6HNzKjZQxbFBEa9pFf4WZfMwGDHg
jIu9Y4+NO31HiDYzuihkqYji+69djq5lvCBveqr1pczPC0Ud+v9k2/vl9mddcAGUOpCeoIqZiA3W
zluqbhMVrskAXi7GG7qRE4y80eXXCxHqU6KYPDGViptAvqJ/wIDg/zzt0feK+gbnCfbWMNISD3su
cJQb1r7BwlhFSkB4M9OtdZ3eZTrPvAt7hxu9QaeMQo8V4Qnsiwjld7iBoXoxUT6BkM/CJ70IMYw0
HeeJzMPfvx0BkyCIoGnXfUKjbuDfKJwYc0khewobikk1SRc6OEWvr64ZCT77dJ968vH3WMfUo/39
oZ2eYUpFiO04mqu9bYdqOgN8P5GPBRPOyhfTV2Odr6YFp/F5lDKAmctrIFOB2qVyzw3pICy4jWT4
d0PqLy/SZvFmXJAOO2TMNLBMBjABYLffQKPnTWjnYdin5NcW9vRv+8SqTMe6Ok5zsEz7s+CNZJV5
Px69+TkZhn3uUy4N7emHq8jmcSh4gTHXawU3/oxBzwFsTa5iQ1TRJTu6tCxhJeo+NVdwdGW3FHCa
AQUIb9gkyCzBvQZdoIDtIPwuwh+o5rPTu05VHcbr4aOSOn5VArwDP6Pe7CutFLAXWK4z+IDI1oFo
OXMf6gq3wFAs3Gsd6J3CDwPGmNNadWVAE7qxWOf2TTpWm/M7o3o7q9G8VqxN2xN9YjWzMl+OehWf
4ORg1lUEpV0CZlzYhj3udykYWrrPo78ztNBeIPitV+mxm4qZwVdToz3qNK+cdME5aF26yG2yiMWd
v9fwCSzPbzz3/pYlXXtulblF3rSXfaiFIxiu5VKmO728hYGBHPlQ+0Plu6a/gqj3y8oLdgPwE3O0
dUckYgpsPzANJdosIcZZr8a42e23/0m0H7mWF1SLDoJeweI96wdh6hQHzOp9pHjy+v3+9OSjEmIA
LJpkKXG2cOmb1mlooGcAHHuw7bar8u32gHuX9hEPrzqJbADExLBWSfX2z7/VjmeLfvosR2O1Gy43
+itidPOG+j8s5Vk2JzuSlxgQzi67tZ/2G0x0e3KA4M7/VDFPPDLh+nPAY1iq9kcH/CoPIB0+EgyC
vgvEJPI8n6w95zZ+xT1cLm3yEZhVvELHcgin8F21nETr8wCE82PN1iaziU/uUZ16D1jjz730ttV0
YfxpU7UgVMTihOPhzvUIR423X6NHwXuwwIEoCNA6LjvoQuJz95unhsveQNrUNAHibz0+cVYJNqO7
GbtdwUriNUCXCGm9jPzWvQyeyYk8pRXfgCYspfuqMTy/OENmruOvSPP0NHuMXtwtAyqxd+QqEVHz
IqKW7IwW/YI/Ph8pHCdLuDfvmFczJWJRfgucDzYOYng62knjRpYQUZJRmsQR6b/A/p6+0tRcB4Ft
WIpgT9Tued0pP6h35/M0N0rj13tA8gB+ykrEzsu+8q1ohcPPL5BR4boNA5IcBahUgQyEaIZi6tuM
1HvMgexkfuSCn+WATfmRCd1+pQJsylG3nfW0Ai/mXQR0Lf4ByzrGfwksfFGoYRIk4OvsXPJFzZsf
eRfkC+aWBqY/r5lXqfZ3rCrZik7OIW+yECsRg/Q6gq72KlVIqQo6RMvDWwdIrAXnhWmAJtf+u75o
xlrskwHEZUSULKG1h/RltI0ufxNjP9ZU3Pf8eJqw2uaoXmZcupSs3LITOrXhfUvpUpKyqF7KHfWe
rZG3BcQWODW+5u7YcTaGTMGHjMyK3uNFsr0ewNjoFxWeqOpRWjgHzuKBbH++m9UC8zSBdkEoJSpW
qGIxFV9qOvO9RbH5ch9SXBT755kios3lCUfESKpULVN1+6qt573TlspFJDx5tsotnv66wrjCPvOI
bhkEpx+jDikWw7YSguPkMaEkkaNtiJ4PiWs+/2b8fUhytBya0Na6116kG+X1VMTclI20fo/IopBR
qilbfT66AIsx850JyRWCMQN+s01RLKE8KAmQKbT8s8RRRwfoNWkh+Yc6zbdL99UQFSlwbLrFxpf5
jI9Gxv7ctikjyNYJZv4FxqhVdO/a5IMMWo0ZBNVcDZkYj+VHH6xgM6kPyqa8oB4S+QzIs197GGug
lQSVADYcFiHrNGpfyJATTIZQSReWSv/e67eL03j/YnZOjRnOItrjwBwx8ogd8GmVVYIPYtkoj4Qy
YukpBJLaGzfE5QDKTPtsUiscRBQtq9+M2me6pntEOkL5jnvTu7Lj7zPMc0KQq3TLBFnhMZ7giOb6
0EfxG5Zv6tn2asxnnugLIu2oCn7Gm1oWU+5zFO3jAHKzA2JGhmY3azSHzF9SOr/gewP9HsR96lk9
dXPYbPvgWQvJKAq6M61fU9gwde8iXawjAaZ0i2G0gM9LdWgekbwB1KjoTNTfI2uK+iXxuA5T8ToL
+YdpWuayEMHK1faWdiyRJ+wKMbmwzAjEgI9szIALF5VU/0ngUV8oIcRLbO908tTy9NfHt0PagUKz
RxqAvVUrFDLpDqf2pSX2skR7Rz2JAwNZIpvFqx/2C9iZiEQiHmMxE/ey+WliTlBrbrqp4GF0oF7+
gWXgE2hqvk22EHX7s8OLDvczL6BjXH4smEvFe16IF5FoF1bXJiihW39Z20pelaca2PYqlv7erBgx
LacKit7Lpxpa6FGo2V1bnTYyM/L9Egatp0e3wB1cHLkXhdQ0MhPRwhq5wb7NClzNIEM02ZxnhzXa
VNXDdDhrStPskyxhnOrnYf/3kQTx6K+tY+wJSTmFjkQjjrbK0vv2yMeyOU7ES7iHKSBEp2tSbuNz
RSpmm4cIJzAPUX9TZWFYmfn3Zluv6Qvw8rAwixCC2FZsAyH8XuyIWK14ShJNAamK3EsAI+3DKHDI
G94hWeVzwDnUeYIViJA+Adg6wArhiscZXktnYtI4eIX3bJO3EdTrDKKyumL9gvsynnztXjurGzjs
WVuTYB1d5kZSuOYeYobU+SLwPpl9gS4cJDBpSNne/VTUlxqi1gjTQpfBz4+nBGiirJj9cwue1Vza
/EB6+n+IPp/pCLT88DO+Du8RlDaM1/zX/qpQQQBZQFNb89wxvq5fmRhj0TLmBgHTLc4mf0EaOQKz
pa9IczM6REkx4Px2ZApeIoNO0xUH24cWU5N5UluxT+CD5ch+tziwpSA/q2unhzDuryzxc+e/55Po
iM1vLANk+Fj9/JivwL3fqVXDFxIvM95GoNnx/p/yiqpsUfSyTfYDGbPfONrcvOSo7QhtWrepJ+DW
/ozLBQgP8PBDz6XGeMK7gP6kUEbv42z7OVNUzX0Zvweila+AUNAm7SShDbN0RPVETTHT0wmv6qVq
2ZqIZT3w7AaQEmlh9XnckCngVV2VcX6xgQMcF6zTvW1pq+NuyTQfg2b0gIU6WEUVn2vyEQ/XfRdA
gLzYs+yfweryzkHey8pimJOCr22ECPUi2nyh8mfD8i7/7a2FTO6VYSr91F6Ix9SP3Qd3b0Qzm1CW
KfSMKdo5MTNMZOSegXe7FniikxLU+j2/9WWa6I01u3bM92IEJMFhQ+9F9rzXUqPVgp5N+gis1dLk
CAV34vAGgSVQ7hsuR6IbGuopp2N5sJo5rlqkih3kTK2dmjfo7WTWNDnwd0aRMAxKF0N1avdBx9Dh
v6GXW0AcbC+hWWJh3uPWFnDX4zwXhq3rjgzBAUtkKnnhQjpXidr1hZW1/6r0T75XFCDZNoaPdppj
Eov+TbfCNI0n/VEeVl1KrGnKx4hpSUeicau5L6D0lQKBxeIsR2m/2m3IGG4GBIbrLo3U/WiTeTmV
QCEnOqcFeKHFD7apjtvFNPKwlSGX6W9lDURPPvZirU+FNqVL3rRbtGgqWc+3cKkexQOiYxucBP11
anj84Sp0LsZcNQTmbkizjga8sAmhZr2ahVY7Z6oLDvfFxL6Y4ajm4qCAHu04WQpkVgRqVttCnVOB
Her1Qs9RkKNXT3e2fRXFOPWgFMXa+xTjZgiwavsvAt4OK5hCQZHsEGTjymth38WvbT+HNpGKRZmI
oMzAimv6qEge/iJnkHPg+4AGeW8VYf8bPenS6RV2vvrDN65PvLWKt4ZvPyY0bLVbYBGeuh6Dhkw7
e5pTROOUM63mdjz36e4FuAdZf5tlFHu+s1dxYivQIRBKL7hqHh0UmKX5k5ctWTxxymd/crQlsWWx
fVURbC9Te1dgbdGkskSA7fYj/GDG7tDoBT7nNKm0nJRnQx0n4scPAB3x6Tght9I8TtrtIdrd+Sti
kriMIRS66r/qoRZcUdIjDGe9SGNFc/rFUXSirYldT4INGdrwKOcBEWpY7Mtlw+TnzBLmNyIqgowE
1s+QD0jUmKcTAuOohG+HiTEzGpAOeAql+FQTHrDXOOJgyrd9sDnLQpl3LO7nYLkXvkGKN/Gb5jB1
qzfPJ92yFKIuefgU65ubS9IrTDRP90vfTO2PsUE7kLiKsrhl55m7S1DwrN085ahRUqA3ETzQ4nw4
flMQGcu0Txhfqd4CPUIrB425g0x6rTkbEN+Y6qQu6WuDbtFBWtGKTvk86moH2u3L1bDvc+nMtgnp
UzqEYGisDoCdLKEl0FGlW7S/+VUEMZvc0tLIoUxZ/aMPb5tLp/rrmI95ugDocoXSjd//p+LOFfg5
SzDT6UIX0XXotZxzvTsKwhGuN1nqkEBtJGbw/IyMuTlYWUuQqg8/DJSyoR+Rz/2HCXtXyo4mYNbH
8zNxdntRkGSS9GAomeV8fdHH4EfMjzSmv5zBB8FEDsDcvlFr1cJLCq4eeGfVQ9p+XVKy0k8WcioV
Okuz1F8iXSlAC0x0EYn+wrucEoWI5oFEZOf5bn3hcz5NjJx18/fjUIVoxQ4doDIsMFESpFdCyna5
ezWRuljWGJy5pT1qFVujslLJGyRGUn8tTupn+e+HKslzf4LIHLXNTDitm3VTaZ3K8DYdRn+S+Hwu
cXotbUOAJkwf5leQQ0mZ1/X1I7+dmu0Iuu56gZ/kzPhQylF/HnvMi03P6wmQcfvtd1bwiOO5d/6f
RZxjyqToNXQf2eE0NPg+zR/7A35DEyLRc7tX+Bh8Rm4a62AsZPGAUreIoGq7Lk2MbSEW2lRgATNJ
yRAr9Dgeqk6ZKrDCV4US7Zsx81mxUU3nMPYeeWV/lpcU7agvtBvR86a5iCtnrsujOz6uIxOdT9Iv
1MP09oXFRU+fmh5rpFOmYxYqoaXJeaWfQRvhEd3FrnqUdVXHxiSTVEJOkilEBwR3La/Ze61crlds
A3KK5ThAg+XhMlBlLnSAjldyO29qbQ6FbsI+Gm6NS5y/qSPphdMlrOY4+5r+SF0pc10paQ2k/vuW
nqJZtIg0kM3nDNyI+Lbvtc2ACerDEdakWZfB8RvaOqbb5pD+Vk3YtGKH9wfHfZ521Y36YRN6DWVU
pECU6avb9jqYMIcLlatfAnYcFmiEYmfB5T+Kcu6w8OzXgewQzmq+3MZPRRds2rIfagm/YhqUkqO1
YPkoorksEksoFXmQAxnemLUKSJWjdkQ8xFdfQec4ZmAXH1VFFU8DpIIeBsoTV7hs9h9KZ5F3tKvE
jd9wIWAX/HgsKiENXSkKG1RZtFmffMTp712WsFwQM7mTTP7sd3Zoz1NQLAJpuCS1oez6/sMlbFw3
PaTyOWM4uYXR8B9OMKelD5uUz6riT08VgDxVi+d9xJPhMJnoq3ZvoiMD30w1VerHKkR+qC8CK9C3
Z0y62Zpj/TlePo+jYIS+C25cSJ4JqM9TINPA202ocUt0u4EYJ2mZGAsqsQWnWOFS/LYQyogfuEjX
UgFeZnm1n71Q7mXIiM1ux3T23i/ZecPEjLO/x+4EVGKzbZTIirRjKVU2NqmOER62rdg+k5YskX7c
6IKCvVJz/LWpWkFkeyCb6Ttx7ZmPpWnuT1wQN6iIA18sKhG0sT8K+iSr8/CU3VhqegqKJvmvRjGn
NqGYIKC+vfjiSbpSU578+sutKm4OirD6yc+tEuH2p85ZNyreWQ4YqGIRl4z5cAquclFm7rZN9ueT
DKxkvm+kTkn+dw117vx77FWdzXj2m4lwry/KkMTFleA1kDbVi0MGOlM1XWp+ihxGKHMSybaDA782
EJjpdFz3jXOc+tBZLn++FZ+ClA8aGn2n+AVtYlYjkCRjmKNUnNIF1RMIfJP5Ia2kiBzDm5F2x1II
Vw9V1vRU6fBegaHOX+cYv++x56pIAH7B8Ola4m/c3zH1iSuG7kaua7fncNtBSEWPrAGj+gpfwEgU
+bLjgyGrtyLBXC/cBEa8XHIZ7Wyoi8IzmxipaHEywX1yXp+LS1yJKE7Wm8LOGsEEu5WumSuV5VST
3ejYHM/dssTf6hQA48OwsgNpyY3GWx4e1lYiyUGoy8kTGxBEc10tHYgrDVNRvq5m77b9o29Gg13x
zTbtbIJrp+TXPJjcKJ1qGU4eUXjNmrbKLCnT+jLLOrngt2lOAtjQevqMzSLnpC3n4bx/6wzB84TF
qQgtjk8YlJXIxvreprzfKqZOx9UfuS52pt/ZwlxioqnGF+GWyKDsBRAtoQe6P6mIqOapRd62Y7Pd
V3vfSXZlVTHbacuPQ81bsKXfekYhlqDdB0YLF7CPbBTN8oa4IIPgTb5uxTBnQyZCduSoUncE0oKh
9WpPfbfNmyxDGpaGYfwSnriA9k9p07euU7I4MxzRZr39NUpuA8yQDcNT07FEOXL01uw0XcGxcxw2
OG8o3luIogwBZe6AFGSBPnCtUyyoqANMmcMXREQPZ0lmOuejlxfQO9tUfAZBL7ACWPb/WBd6s3Gy
jdKN2Pzkuy9g99IsKZHm1pI1xSaxWqWSbcDqC8I5wV4NUSlDJURFkw2Ka2MEnR8SGIORLLJLUlfD
YJpoO9SWrDW8TojguWrdiTQCy0WvsAdDydZU37g3vDzlWiwRK0/t1J4hBnWrUTSYFv/jHzqluUUD
7b2K1svaPBpK4vvuTNy945lKZ/SkhLWFSYMT86+mhj8uiTQC8vepzjX8KeiBsFQ7kqH1osOa40/a
bChnOa3eQlnlOln/qIxo6fkWKFhYlFrt7lOfNMFCVVz6RO7+tx+d1a/TeygtiE6pttYZV9GQu656
EAwNkqzh8C4EqVhm0hB6SlD15/1JFG5N6hg75GiSE0k1gUrXQash+UABJAEjBaSpPLvGa1owPaKg
Ziq5iY7dk6w9ve8fv9vY7jXwepE2nMwMswSCWf/5htoXxjDnfbC3Nt4i/6T1JOhRwioprXs5Xy/4
tEnj+vmmfAPflhBaWkmKBs7qtXV3JWWD1H+FDl8edXXeYqPpdG7cS2VBA9yZ+/uRGV/BumZyDJMR
y0njzlqGj5qlsCQKzEljKezVhb9k2j88Z//NSho6Ec1veE3q0IQRPfsOLOLZmhGhJr4qubWtzgR8
lMXiAS+sgdp69dgJveMyMr6iiJyO9lgMZadwzmJ3W1EzbQ//z4I32birz3J5OtvcYC00E3q6B+8i
MvcfGOS6fIbjCSy5XHpeS236gBfLu2dgbmh6Ik1500wV3520+EllJ/TGxqR9YgxFYMQ6BBCjeeE3
/SDuGn9KjtfZ2E5ClcmT03gZE2WSsk2sQU0YtH0fGxKOBnYcmf7b+EKjKDtouqHSMYDKHhJXzmv2
hYNq9H9pOjbsgdRBkA0xsOPjlddqGE0A1BY2QCp7je8oDVenVkD6qoz93YGNANuwfu7Ca8oG930w
XmiokZCK5GbL250vjn95JXGIdROFPlNXTR8foJHmRXQ3Qi98HLEUKPi8qMaUVMjnG/mr1Cv2W4G6
FTey94zDttqqP5t0Dj8BZwmogSi/qfT8LA68V2b/NQyf+hCZUtiMrN6dBgNcwVJjqwT0WhhnWctX
zZit4dWEPiNQr7HdvF6qu29BO/67Cec71xZtzSIsGSD0mLMZOvCvbvWzI+zvFADd1E0GETjiKvq0
9lQgQrH8cmSF/KncWVod1HBgVG9ZKd4hiWvutnR2tzhcyPU24lTVb0OqsKpTG0yKHRGiGUwZdups
JN9Q1+sCADRLzH5AjVsTZGDE51Ce4F/yJpHunCc5+1rZYXmXkZWPYnvdnyYeldYLQjct0rtKh9B5
A5QEfMy8O34oOCJgzz9rFQ5WK0lkezf6S13o/se070fBvh78667iF+mxmAuWtF4k+vERZptW8kFJ
pIr+KbtFaEksOReHSXI9k2zpvyAfIitPrJUcKIK4Ul/XNZP4LdAgba05UJjPHzo9tL6HdgtG9MvC
qFSZQ7/guLFyjz/s6tafOdnGiNEtLlmow78aBsYPZAea/MxQOs/GVK7gfAZ7CK1c/hGec09BrUL4
x2Tpvmx382vykvIdg8VVQFf9GjgPtU4G0YmYHe8QnmY2FdJHzzrzV+eGwwTwQWbohI8EZI/9p1o/
FpZv/gCMu1NZ9Su+mflwy+3JgC3mIM7SYEE8fuQW0JVCIoJyqP1FWpAea7+xJo9O7tptVBj6uwYO
EUrP3UevDoC4XIrDdbA+zNhv1ViF3pGqLFtEHxJptKwLNEvzx3h4IhwvtnByZDgjB10WXZde+EGE
qHIWer4nj0NBs7976e7Wz0zH8oqEM/FzRqR22YrW7t3cFrfiKUSYFvCykhr0VIYzEi9IrcOety5A
VUWuku0m886ztDblzS8IjlvpQAU+Ovs2CkiOYBGT+SgR21FatZ/2Kd1TkWkvqUWPvF3XLAyxv3hE
/jVfiRO2ftTjKxa0FhKcm1Ae8iiMJJ/BCwlGBKOfBpoRAlH1b9JVnjpk+QTrqw/r6ZGNzVWQ+GIf
WOPu+yD0MCkElS0NubEnAxC6bvIiMBte5w2/CTbjGM3TfF8wycQj0wpCHpDjxCi6jW10rwZUvzep
sdsYLzIA8xfRcSeRfKhKB6nWXRA9nKLSfL17wlnUQLX4qPTCubtP5gO7VGhv5xyxLXnivYycfTUH
lHxrSwsdFiLQZwW9GBrmlC0K5lT9uHG21IQSGGPeEzXojIrZIkCJRQ6CO+AyBh4syLT+Ad8IcZrl
T75hubgxWBUrcShRFRhX9161T6V8Yv8tcMHtp2KcZ96D3+eofKKgVfq4YPg/Q8CLuNTTM1ScwxsV
FLFuKxA76gApCtwYOs77npUsAvCtyujTA326MQ3vE1wibIsoe+zfcHCGUo4D97OreQiuJBcce4bL
tFBbzvM7ej2EPUNhIpKmjS7hkjtAWjhIlR1S/MVSKKZ/sfj01H5ZPZZHAh/qTk4cIpynj+8prwuf
RgVQl8/x1ReEwkNPkvGo8rgKGmhJ6QGkrDjjZIJzDnA5L+eoUA3LsbyGVPpVDimZKA4K7u65SU2f
/LkOJlqIpHx5ONn2+EqN0iqwKbIlz3tXe+5PuhDnmwjPO9vDQvWkoNMdNK0B9yiA317wYLSQXSlC
D05nV2GZ2jTc/ahhF9tLjqdqaFufzW0LsrJeaYeHtXrv8QL6svN4eAGIY3SX3/yiK5EieQEV/c2T
JMRsVHlF4W9Mrds9zGSs+d+xiN6XTNKRG1EoDpmCi5B32kytnDDM/Mid9eV1fODjm2/3nszQlaOP
QqYWVLsKEiSGP9kej90ivf0t9wFgQiVheFHnwlUZgitB/oly7LkaIRacL1SxxuZVH0a2wXQaQMgo
cAdX6c3GrKhgey+Toa6fLsFrMkY0vVDJNfdnYHe8JLUBl5dh74UHWqV2n901mKztpEP7b+RXSpFU
PZj00q75jxZzRt0TCnHInPPKznUiZRpz5g4enn9ACRpJUh/xIHgGtBSjixasfJUrXlnX4ib4XdBE
qNWuPctozG6aYX9rX3rPBj5hqUiXPgq0UuQCEIjpaUY/mX1Wy9HS8g3P7Wc7oUprTtVwqukD+7Rc
PJh7t0VulYOP7fEmTz4x3rnrrbuS9PkzhWhRmPzbPos/vVAKbxH5ZJslX1oRXBAjzW5esXTwBOKi
+YoHzUhbI2WDfs+w7bKhsWwcJMa3dBv5Wur182wB4Z/uoKqr+wvmVib+kZcURldosgEeTPaS5n9U
nrL8dHIWsgaJ4YjPUztZh+LH0Izw7UvllAhjZGWQbtcz+bPBA/BuViiJk9dYJZgN/glBuLgziyp3
zDEb6T9GOSo8TCko9b5ErS10tIdlSKYOGy4xdrdEOgi/0LwXKvelKnJIau3jU3SJcOUuJSFpb0lD
j4oBi5DQ93v40/+46DPJJOOnC8cQ5O/30fp8VyxD+1TkKe9JUZSj4J/A2SJQOiV3BxQzLmHgEMV7
+etyHg6QUCx2E4nngfncxVmBf5p/fiAl6p1Cnr01pW8CiQ/phwX/idUxuOHHMTRYHj+3PMphiuQY
zoyJnAbkVqQ0qUKf2Sxya6f8pIWqAxMc1Djffm7pIVM+l8aA5dUodZeJacsiy74E1aQCJQcORFbK
hQIneqiuoxFkROkBHH2kXgDBZXyrOVP9YxlsfyMZFnC1qsPjqXFfleoMHPI8IEIonEyb+MFOyGfH
kGDQDLP7GuTViuFGqDgrsM88dnL2ZRi7Vsh7dHTX7oPJxEAcZOoXMQS82Vt/KHds+fVqAW+9UklG
aLoQ6xgtxLWTqPVuAUj3pjPJb9TKsJmStRTllKHTr0Hh2n1yFZe/OY7QmXeZmdHIuvJx1L+4ftdv
w+s10QEYvE0euJ7mVJLrsGRcrZr7tHyB7PpgpDapVRdkb+PjEzFwS9joBUcTmTm2+hcEyYXVKwHt
F3rpii6ScX3jnVqIeK2oa2ArbDZen5y7MxNrfZo33oWU+yrCLA2CnlD5E3xSsONINyx4zOXGS6FT
Z7+W5buMaHV3Klg8PrNuwwrizIGK6NnePaHyUNMfTeKZNgzLFhzh+PwM8INWeSX8HANbl0rNmbBn
swy0YU/W2koidQNwcvOqkIuWZlJHgQFJgFSgRFrSEN9rRutZPNjtvz5gFdf/WrTyciWcXSd5GcoJ
Czc7cyX4YtVhOJ+xdJdKhpgj8e85ly0t6ofa7V5AoLzllbrT33ye2g/16uCrVmurjDzmWA2d2Aab
A3oFtFhjQRQshPVv/tnloihaQIzJUP7M524M7m2Lh5e05FC7Izari72axYtAvIHrZtrV2GIvYHAt
IvDtdK3gvGMdCjA6+bF1Fy2X5rf13+1hj3b0n+VjhtxPeiWbYJpQxh3ULMnj8YeuRGIL8Ub/mnKk
0MQBDpWs29yzoQtTq+6D6KH68STpVeGycDoaiuKVDdSf/MvRUt6ilmZ0mA6bqfTFoTmZot58S4jm
4TG1M3+K1bZUfFuP+QDy4bhv/e2chvNVo0Gz5SI/NTSu/D862ZpgW94Kz+nUby4ce2IVVBfc0CXk
2xvQMG62C6NskaRnfHxoh98DoS4k+7i+E2CIzZlZ0R6WmwauwcXRGL+UVtc9BfkF2LCeRuw/cI5j
Q2qC5cOEMQ8MVKeim1bFSZBqHuaOtlNrRRqRrkl1OEkBsr1zIl3djre8zBDd+MH8Knjess/1+FBz
XE95ATwBii6edAd9ZXeeHR+8WCbRloUamjUDeeeqoVN9hOl3nzVzkbFs/9YXjWcR0xYrVlv+shdi
wagcI0fmGJPAKo7vlHvglL5mFFn5tQY3Ez9J0YymvGBZFVjSVuUI61Lek/hVkxJhT4/ZsEhh+wVh
Ift6YzWVLlv2D79TqbCjEMriWnR598mJ2krLSZESMWT/pFDE3K7+7X7gqWVNiANytjDB2sl4qraf
ZDDj+v1xElIEiIE2XJX/iIAqPXHVCv/SoL8zGY4D23np6XOtUCfPqcDILGJ0CVmsPywr/FFyp9GW
5SAmM/Bvp8PmUoOUPE4M+3Vcs9O2g+J3SdrBTPE/pw3b/0imisrv1SAheptPZlm0onaPEhokaQ4b
hh2q/lSdsJ9LtDpoCiqg1H3DWxP+Y3yP4M8d3Gro9Z58XzXPqlg6aGmaZkx/MXYic/duu1cVVTXX
QM8j3fECv0d46vcJ//i4cXxQoQzj3yG4X+l4ErHRGxBeDFaCeI6X75FI22VJ16ewe9cxl6Im3ire
xAUfGNdKSzTlfzdOPlZFAos2Fvhwv4+el2WR6a6QRxK5Qr1njysbnMeHN2E9vFeB2P0WGaOcZiAE
ZIimx0PX1BXlu/M0jTvji3A6fhaxrfUq1fZpPJWMWW4gnVFvOS2Nobx6ztuHDHogndTlI2DJgZaa
HF2WDFzysnAV4FbNIwD7bBeGCIWWB1jhPzeWeMkHM3zdv+55LOJ/yFsadS18yXrBFzGI7BEXCs9Z
8T+QJGgY0Rn4E9UxCnjMzJZy+BGHCU84UP2Cyf6blI00Dd9pzLmm1rE2wA1fkOOyFlkXaMLzTHDg
Vg/4CQlHUj8HNCVAAbq6pa0maMRRHqacFb5SabngWDDv6EBeMV/mOgsg0nj893CbET4rU/RpM30E
N6JdpULz7c9DOgADnzfFhJVe8Tf5LCUqIdIDZjOo9FaZcoj1Iw1zNXN2i2I2Yk+JTLaqs4auYl8M
0JiNaVS1htp6sBu9yHnQffCRZF1ik4cEs77ZQpCofwXmiOdoVnMEmRq0X+86WS0B9ecyWCZUXIhh
UbQVVDEBWXwXvCnDxFtMkPpas0lygTf/KyT+e0B4andGi1x6+42g/sf7dGYfTSg/qnze34rd0oGU
X+haZHbBPqVnYwiy7nzG8+uLIxiAQJ4JN7/D3hnJ2dudNe3EUSTInhWdOfwPmQJP/w6+77/2qVc6
2ioGYsa7pAsxeX1TxVl8Z07YAeQWzd7Vkk5B/EpWkmxzeUxDIKa0yjJromfjvwxr+p6zKOTX/fXF
/VmOvsTOfnDmVXJuLQyiIA2kHhnX2bA4l6HpG0ih4FtwmJoq6F44JICQsM41P//826B9IBQCZNwI
YfAhCX2ajvoRdkuI3VyoRDBapL6libeBQaYKNwxJ1gGskN08E+/htpjn1Mj6mR6UnGEttjejnzXI
NqtiHjBqt58x7+qDKlyWs634FEmRZooM+Vqa84Z0KwxVny9sGhar4KaLstTAXwU6IoxbYEL5h7Cc
QjX+FJ6lIDGXUibQu/QrVSTSWZVpmIlWlQO5rXsuoPNQiFSk/saN7EQlcVlhfwnOVJzoY+QAv7Br
2zuIcFi5R+eLHmTcp2KEpbGaWwj+detOOK5ZOEDxavDJMMiLCMVHiIitY3/m+PoG0Mo+D+3Y//q3
CqwHJ1ckj6ij+mv/gwozzMYpXiTPm/BnCi2HjLQ4oTrTEW3WMrVDJeVKHydsJCRj2DYFm7p0H6Jq
INhYPTA/kCyp8WTb3jMtvqo3MJBxg7L28sh4ynJB87ZrY2nxVFWY+LkMBlkFewHJCDXHdlPzF+n8
u73v3lfY7JPNxQuPM5LktRyzF0NDTZXK1n0Qtn8BtkYvAQYBafhhiyneDopXznVVI9383tRbrYOm
Sw7ySAJtA9ujTBArO4IcV4vpv6IaPtyH8uosPjOMxRicVqvrnAalpUHH6cU/JQVwbxoT5ycc82K/
baCpSLQcRJOk7YOJDrlv0cwTrAE0+bJaVuuUVWZzTvkiSm1pqOumcdrP50Gb1jiLkar+S2Tf00ga
bTdSyaSG1htEjj07Ws6tDJwTIIr7O7UHykmPb1f2D0VfB+eWc5RaSVTFzNyEmRNVDmBJ/cIRr98y
uiEENRlODTB/1GMMZlQGA1JZ+EOrSYc4IKZP7DkXK9VJ9Cxc86D61DXwib4ZdJFhnpiaj/N1cmqE
hAHz0rFcYJavxbC6NHDt0TOnqhlHdBRKpFQVZ8J7ii911j9FDEHpklssOc+gVAnqmTuiMm/EgaTh
IZbiRtJsj+gpvyM2G/SzjT0Q7AU5DA0nvu5wu0rUgceM40YBV/FMUx49iqdbrwXsD25ni+L3Q/Fj
OwKJSsvh8VyZnoi36me/4MXqjhm0t4UjqFczDUmgPidqxQDa+yUg7stACDFRtlAb7V4Tq8CZKa+y
l5BlBoAGhGVRpwNG7FArxv7VH3U9Je+pM0R1xN/VlrHHVMDpERevjVk7/PTn1in20Tg46se+99WF
9C++QaYqFX4MuE28xL+5TWnucLqU7/3Mx/TP174x7mQC38wQ0H1oCZLsDv+1zoH6Z1jldUbmpoYI
baU9b8T9RqS86Kz+wL3K2Jtj8knAdnELJI/FHRKlMT3cDrKRch8jtFRpAczs5yUx3T4daTRIq7BB
PBZ+/fAo4k3f5RtEVfiwhTpJw+ZrL/znovOlhkvp1pkGlwzpsSBPoA2jWW4SnuRlBiJ/SoSLkF3k
UVa4GNPw2naryfy2vug2H7Is73sxhJmVBdQomBFvF0OgOKhjAMApS8WFkQ1LBYxcU6oWE3KqeiAd
nFaDXg1H8UkOgmo9ipYe00eirqvYi4J3EtPG/pXdeG0Je1/sgnFERw0NK+00bDm7Tj79rc/gH9FD
jml3vepY1dqvPgZcTuoOPMPo7Ov7tovopSu8es3O7puKLN3ORgHPTdIXSSfiCGkNnbfVkvdwqgws
5XmeaH6t31UUB3mHWEJ8DvbBjgk+TBcKigBnR0QMFH9NBpBQUpIYlIxsd3/EwK0qHoRtpc3E+Fph
aspPnopbmn8NqwqjdCcDJEXzeJLzTQ055a1Vov8DMFjov4iVUelrHqHt3dd9zJpFK+rnsluMnREf
RXpyBtM85TaZlnX9RlJSOyDNgrORhGgrR85MjimnZliFGX/3mjaajwzVz7i5RomnnEToaQIrQ/D1
rx48C6xkcLjSoItkC2My5zpu08TpipGi1rJeYPesaXd4jqtL7YDb477awNuDoGq3LhSbzkRarIRP
pgeY6c2sNp99C0fs9tg2Q1/fzrOTJl77ng8bz1mRJZPZ0rJQRBIuxegfXYE0R9iv32yZ+lrZxYb5
oWZ7CEDyd49rxXS7tA4seFnrbrqDiRQfDbyyH9/Kg22TbuuHt3ipjizTazhSzihoV77Y+EnZocYn
HFvuAW3xQ+YOU2SFtcr5nPcrRmiRk6aeoo94feaA9vB3IlC0GRXeyc9mvSxyU/WCiteTAJRF+l5H
VrFAySQ3PLzek0RJfxdXEp9HzKLtM8NpgnG1qQQLwZfmPrSlTjw2szxidzN00Cno0EgaQBsXxu31
6/5o8HwNaT6AG1u6c6D7xKPP3LdHN1AOfpjZL1t5LVl9LZYQ2H8v3ndmBEcMdmyTfqAuqU0pXKO4
ov0OeeNuBalErWeKzgweJJSMHdjPD5eYkdaEDKAApRIGkFpq0XoWj8i7S8MYbnI1s0ZsNBMNuj3C
ykwx8w1lg9m59HDA1PkS3d4ITHLhliJ3XCxG+BP1VbbJ5anKOnGHKGxxONOvlGeC8b77udZgeZao
U1eSzPhAJx3XFtrj3GeQBrerzY6g3oij54gYA6bFFBDV9FZUFiT+95khsCqiZR8QTRKWZJxWQOw6
Aa+R5fgQTJvOmGTn7HOox21Ejk2IKriTIVcgcjqyPkEBPxgeNgHUQYYcy0Td8UUW/fauGb8S8PPz
b8Q7D6BwNyg0nmJ67ukDdUszNwX5XMvcxacprSZuqvpIStcFc+Q5vb14/IBfEfQhz03USgWKQg0B
1nPrnhXtyULc3fGVoORuGU01tkDuxDQyoH8L+MwU2q4HvnrbTp7iSUIgD2skAaCNIXQ0pBQWpuAr
okwDCCGVoSG0qp5zdKRgv2xIDC3f455yJGbS/ztEyxPvo7jezzGWRjmq8RBCbNVfV4PEb/0iiPb1
35pTM6WusMrYBWnksNZJ1RcsU+zYxmt9J8rNCykH7vWwG/xdNlM8Ki7XCT4ueAr5RJsKJ/iJUCqh
oboDZCzVrEkJ0ATQqNxHpqBD1nttFxAuPoRXUfEnBtMrNWF755dHtntPU+826h6z8dVTBGTPF+uN
Hlw1rlS8YXcjn2D/RttH2PlilEe48Gfqh0LUrs6AtZuLURPZRATG0JI0YH1wQJ54qlvwZwaFdVuX
Sc0my6+c5SoiKRyilHpYAwhAYNuf38JiYBxcNoUv0EGrA5Yz0d7FVyLAefI4WXepfC6q4zc3fsGo
ltdUSwwGUCUMlKF3ZoUlhcc7g3F3pKK7gtmm1DgVgbomnB7Bece2G/qpJfpLI1vousTcSf0jtKjU
uS+xWQhkc7k399+uihrJc+fq/V591e3jkHE3Putm7Neu8UVVa4SMmp6aE8bEURHs8CyqJ3yoA57g
bWF9eKRrwavdjYVRDakzRcJJ7L6GyCrgLHsP5frGn0b2/3j66AIBnz/9e/rkoPb2dVlthVYmcVYB
gPVoTgzp4zWa598d8DwF33msxpUjtuDLM5oVwv/0SHHCBp0udZcp3MV3xueRWUUMHTR+ANdTQk4P
wJVyLOX23t9x6arZbHtqxHNNNd1CUl1Kf8V24Fh3hwtg8M91BFucJIoYjY4P4kbh2FhhDuFJHlT+
1SuPKL56mNATl3XbpBZwi8Hwgr928TU/AuZ/0Laepgtq4Dc4xm3cegjsfyykPHgVx5526+V8gm2G
L2pZQ63koqkD7dzQKhwoMmLGtoQgR+gPbM9KO5aOqpYwJGOrvNZyqeHrj7EngGCnmNqe4O7kM7Eg
+MQMaIRBth/HAh2+03RE6exbAMrk5CUEsCZJs2a7mY9eiCyv0sGxUfG20ZJULMI8hBGfPY2+sNxU
nxblOmt3lpjecrv7VJTUpcxZOEvScV/7YzNKZMMWe8tg+LpCXsfDZ8tpqp+WkeYQC+sC3S4eyj9v
5O2DqQ60g/8QjIiKkC2bR1LzjvC/BKlMWA4WqOwzTHsRwhUWpuYuE2Jq6vgAHkpI4Qa/bKgg5arI
FLhbt4os8jJy2b6e1lmGU+187OTfzxRXAdRH6MPa4QtDwlKxua3C4sP2vD/yR3oEG7DzC2zZv+1D
8Lw3KFjWilzGTmTZymazfovsMSnU1RSk87QFq2RW3vcelNZBlXC2lMHfPWtqDfwDSAtXflbSorSK
fHjldqttZPS/rMZOyQ+KlQ/nbl0iU4JOccaUkA1TmmwEMtiPLczcc0XZOt7syjhmb04eSMoDm5sZ
ZECfW1ELAmye7Vq42pCu7N90LdFx7U+MHEO5ZR1fluBBgv0rXR6FLKHUDf4sfskEs4j2HP5NWTc/
HOK3ezI9DgQLl3XLDubdgwjlhxn9toDgETbFL7u7AnbicAKlWG3Fi4Po/nvD1y3kYKHFGJXKpXfw
h72zYoA40Wu+sUvHO6CUa33CHnE6ycjWAs96q1JXyzOzGXQ1FGDKDxSE5tKy+K5hdqQQbaBwIjVT
OBt1mD6kVrIthkGs6v/hRBxp8ui2ceEyJeB+IPv1/yj03014fW8xAeEtew+WXkgVabMQfHvTRL1h
vtDlar5Y5uZ8FqLNg+LbP62aXuYXVdF92gFV4Kfl4AEjKx49fAJ8f5tbYO5GkB3Rs/PoxQr+nyI3
HYcZoAniAAXw2sgT5j/IXhyNJ95a5YqOF8mpUCxwZYGH9No+LbiZ38ip1BMFQKfnQYt735Yri9Tq
f8Z29kRNeJCuMoSM6sz9hwqkk7to0wN36l5JPMqZbRPvoXh3XrNQN4DKwN2IqE9N3TiCtQvrVnwV
yNFIXFaOyFEeDOPkEbE1f0Yda3PVRROZoaDIHzjg7J4SDpnzeett/KIUQZEC00OHsBCKTZMB6NBC
XZkdgWpXQddBH2oglMy6NAc6rf686FKuHLPx+nGRqs3SbL1oqDfLyEyIxSpsO8IyVugW8/jIZ9ml
E75yMKK1QN5dtiqTrZfBS6BjyYVyhLnOgpcH1OCDU4Gmp//a1Zzhq6rvnhliQBU9GDYEgoWIb3kp
9nECUiwnIEv9VmcQ5VPqGj4L8yjw+gKEw0Dgnp0ksneOChWmFPawZ92Ma/jZrVUMLcggtK5X9ZxJ
szSX2bPowPuJnMwxOnwhqqqnyvingk+wgZdltpSBd+bniNVOkWV1wB7CsVgkOIDxmKgkt2rOhLP0
uSQfEGX3Qd66hinA/dslgDe1OioKWDM1AwOVm3Lx8pIxXyw4/DvjqWQ7lBiDOEjDJjddaLCu8/be
QU1k+wV6d8YLo+TJZD2a3YfZW3XcqOWxsG1MScG/W95PGmp151YXms4xIbtkh+36J4j++7Le2FL+
QPiz/h4roibiIREcXpA+gNINshoO9CCnLMM3yZljszBWxQaA4jf6oCTWq4j5rNm4dShuZw8rIZO9
m8kEydJwfs0AfGUflBJHcNzW4FKBjXNEIOOV3IGRZnK6sXldqAuvWTXrfEb6CUEtrhIaXrlrp7QD
1YidKSdORrn20NsczjSASzN0WjeELkznWJK+UEkDm9MZyElOpC4seuv88xWKbDQmAMF5zhqVw73R
iJry1O+PVCtnMemww4s1dim6+vr5zo2UvnQwDc0bGHo3z+hhu+F8cwZyZ0OtqhVniGjs+WUmbRue
YNdTgRqrsKXomAe5GS/l1ag7YUTKrv5cyhLo1vGZLrA0WqgmaPllKThPeRPCqU5Ew3IVKc07xz+B
qpR9PmKwHfgl+HJOwIRWom12+e+GGhlgnpRmmdkJaX/g2MV8LjMKzMr1vXcYygoiOrXxl63FjR5V
4WtICrqNePRZxjwHn4p/Bis+wRzcgdYhPAPmq+c8jGnVFpWxOTMpYCXSugIhd5TYnDV2ic86AgQY
I1B7m/W4Q0lNxjA4Lqw/zMPTcXjL/Zv85F5hHFzMMm3zGqebfZ402BPiatUNV+33NSoQMzFkyasX
WTmTME6PmIJrqnWOB9jkHsiv0V35ooEVUbz/g1oa60P80fcLsCt46wo5E6bfgpxRsm3yCilpaCoW
lPpL+38AZZwd5t63e4SV7pkscl1zkDC1ha2NKeZjfg2HRgGyvy0vxAYFGcsdLn2uJ0nCQPUXAFkF
bcHHckaD3PobM1kvDMvd1WllL2BW9G07MSIOUnmJB+1ECk1rasXweycAjnPoaI2A2Eo281ezcfJy
ww+52OEg7WEhUFrZVSX5Jo95IPxVPcIEfsfiM8iLcs3hfOjaZ240vaRnxakgJLGymnkdnXSIXtBh
+dTreka0Jwp/hkX68gLQg0tC8NRg/WX4Gu6Ohmmbr4+EkNOydli9mUx1WZdTIJEVEXKfACG6G1MH
jVXFwelu+gAS6CXPd4D9ZLLBlV5wUHlLkIOgQkBo+Pob22v93XTrdEV+LLv8LP1sA7yF7vXnquxj
ro9/WqvQ39nGGixYeXB4cWuY9eqXSLgtT2VxVN4MBmNfooizMfdFwX8Wy9ENMLkv83dDY9QvT6Q0
XCYjinD7UyQVDwOH0+Ij+W+T/AEDp8E/If6X7WwgY8n2EdIT7Kt7MxpwO86opbSzkTaaAH+lyVLx
txZWYQZiptP6WTUonzN7U/swcJa2Ds++q4zMO34hD0jzrc6puix6tWlCcvdmmGoy0Bf6XnZKk1p1
ImfDqPxLR2QsCBk4BVAORGo8WVItPOpN6IuxdFE7JqNZ8PLqMLS8RBKVEU4HZOjsKlNIDp9OUADJ
8iF+wSi52AWtS3RKO5O9CLDjIzOjQ4ocVgn94JJ/J2+JChYT7tHf4sPIH/j8e6ysrvZjXDivwDJH
A0f5TFrPrThGLpfbsjJHjpndN0CvniIXL08JO316bIAiLNE5TugFSTAtTaL5p0cRqBpD5GEXvfnx
5JMBoX5Fc5OwP/31YbM4GC3Br/C5iHSLqqN6rG7XvzDIpxyg01l6p5vlOxerFJ+zFC0aNqoIAf3k
IFwp7zm3QB0KC3kwEsbnDOBjqjsOQuZdE/kXNTxekx3bdoOoVajuGRqEvWhp7DfCacQ76zlF7mZ2
hYdiJN5MqO/QKDoXcFk+Fm8FfJhIguz0tTVsEnphhtZgxBatyM+13EaRw93cMSin8747xN2xDpYC
d8m5NqoH0c6+8StvDCQ+tOdJ/tfG06cXzRNaE6cgULZh1BZEqmbEzT6bEp9YiNk3W0210x/u7oQ4
9dddyYmF0j7YfoSbdesa1ORz44RlluIKzV1AMnSp1fb/NiIMdf0oLQZPuHH6eRb7JWc5adGS0tkD
qMAeHkhnb9+djJ4q+8eJtGxILjVvsW/gTR16Q76wbKm/eee3wFGmwZAYh0q/Ca/jRxX0Jb9bEAK/
kWI2VSYA/19ma48td5KUtR9gey57pkWD1EkRLGyBKxZxIowpGbA3NTF0/82fQ0gs9Yu1sjFWaHu4
TPbVbtEUa7CZxxl6/Rrv/P8BpEGnSWhLbjHnfXuyGDkaiNwix7AzYK+xfc2g9n1oT4W/IkFDRsxs
bm+4Etny6ZHa+4GmvLD/YvSEHm5CBv10tbBqIGn0EwwugMv99wZijoJ4TeHHzPhwy4dusG7lpR/r
mDUTC74S6OqqvSfaLZVWmemHVMzh3O1x/YfgZPZPV0jpKvmdF/bhiBEFdVjqjPNoX1/T03ynlgHe
FOksY4NYiML/u8H3BjRUZMynH4ohbIlyZBclty97Rq+L4hee43iCbko6uXs/nrzPukZz03Sm9wLd
L041epxT3F83X20uI1o+Am023rjjzqtrA4r/MiniNzgBNxis5bH85eAZ2SJ57r/RynNmfQxJo+1Y
uoYE+txbpiZzVGvGVLhIPeeku8yIL+ViB+YQSlw9TRoWFUJE30CKvLLB3cethKt3cuISQJRO2oCU
JwEj5yJSPlLhqzjW+pdbZBpf5SJOWnCbOKM5shp6q1mYyE+lcD47Q4McQMNlsja1Fml44LNLfMAG
X/slcEgJaZoYSNja+wbn+AfOKsfOU5TFt/g/Ub6TQQslf7r2dIs7rR95gOx3ykk1t8DTffvLpRFo
NAykXUHG/Jn/High32xqIVNq2U/7ktqrGhjJ+uEDCSrzxBZQu1WL5VBbIwyAJxbhOOBO6NGDkMJE
umAwPbSfZ1S2OwpJCiT+SqojML6Pv9mYXCpqqjIDF7tGMMUJbY7uvvTFEuz5BAwLZRJTexBMorFR
aXMFRIqMpSz64kI0nbOmjQ1G6EJo5pU1knPten5J0zwGWUYKaLKboBtJeqwCmBl2fvtwCLewMq3q
vGm7roaU/NcYLDgQNi8vGb+nsHhfVLc0WIHVrDuWdRzySw3JrTNRCka+6opa0bRbHDCG9gs/ZwdY
Mw+4mO1dGQUpygLb4QMt1z0nPdohPUjk4gJzmrdDLIIFdgX7It0AIrOTvwcgGHzOAnN7LW4Ljer7
io9+m2xda5lkcMohTrGfUDynuRsWWJUjetPuNtdQqfaFStW7UccQ4xCvfC9eeuy7pAUqpPRiH8jR
9T0wza/moCzOisvTy7xZON45iknRmzXP1syDVOeSHepgu0dLmtMTITGWxAwJFCJUNdFB1ix/v/b+
V0ENYDeYi9tST1W9rHDB2d2p6f4Xh16ZcNlFg2zGi0T8FIIDpvLAi4mrBrqU1HKIwHugaNq7ltFJ
qnQxzx6cs55h6BarFydsCSN+win/Rh/TIyhGSmjF4ervIJU+3ANBQeAclq6Kk/XurdRSdCEkslr+
YfxvPquwqJHbV4MSHdGuG48LcyGHimh2wr+yM0El1RngOraIPCyhPRkeof5VJPaIY3JiQBjm2BRH
3hy20UZk8CPLBY0utCM3MGsddImZ4tqlw/LIp/98sUJYn4OZYD55xh4FbJFT5vfMTwGParIhv/ks
wRV2H1OLrMrNv/XP6J+5Yd3QxVL7ipO0LydHh/eFELrVJ1vJ3xC5Rzy19Ss5DShf46OPU1r2rsWL
TdZKSqTHRyw4yUzpS5AgXc5XJkT2C2dHQE9sBF02AmX0B2Ry2XPFupgKtjpdKD+fTUDC7UnL68fT
Xo/M5nBJvVbIWxvyh1oDw81dfQN0C37/O/ZM4jxrEhOFKyiZ+3s6hOmSJJZacjniQ07ay4glLwwK
CqdXgEvPa7eJCwbZYr1gS4/1F7ejqs69h+MSEKPE0rx8zoECYxVKdetIhJwNGgxX1vQDXE+Qc5CJ
lChSzjWD46HJL+9KMfyeWbTfSQXKBtYzNTZ1oTRuWMLR4DNjAUpvudbXlrwEopLMXvHHQR7j8rea
l36fcwrfaZ+mVrW8vqPp37tXofEGJ4V8K+W/MwBt4RRkds4L3Jfcwdid4Fuso3P6x8Qmg6XbdOdM
2BWbaOGkWqw5bzMOZ9Q6iGqMGiRyn90YU7jwUcq+cEHntb2pbCFuvUKDe0VCm9DXf+Sj30XW/XD6
xUZkg4suC80iKobThqLrKe1gkil2NFCQmFB644WrRe5MKvcpP+akk1o0uNiN1quIblJFN30dmUEE
Hmplb6CQiiogaCV+X4E1LqrZ6AYDrVuQfiasVo/1vxCYU/L/RmGoZfQ5x3BBaiweL7bkLktyG/Ty
qGjHOgXuil3IYF+aDHVdlOFCygWRYhX4fYeTfZC09QIoKoARlbKDhjZoC7OYTmaAsuYSkLIIDTz8
sX4wajKCb4TD/iWBihr46Qa+CXYQk9e5QFuHzYEWTy4gnm8G+nMoaDCWBKM241esuY4tdl13fhm7
InOQMSPmJzBru3nbdJqvXpW7FLRKUygZqC5KzHzTMzyc8YK+0eVSUgEdvJ8+1ctwiiz3ruLj+SBu
dEJfFCCn03Rb97JuYJmyTW7mtujIAsx1XrMESHeZ1AyfwTpO4vbQ78vgC4roc1i6ssLLq51145uM
EnTzHVPpX14Jx30rdwM/W6RbNhsVRHAXE+1TPEjQ5r6VSnLDv89i3ia3bOfs3KrJsOO2Wf2rDWMM
ZP2HuFHKUBsy9yl9qqOAmCKFnEtAP922Kp5CiOn39A/Azyfn3zU8xCBNPaaovXL+W5eEdUAYNZWd
EmaqLcU29vBX3I0n01P7Fh7kiLTwWs9ip8gtPM6YqhLu9SJmj/Whwb+ZKWTLZHAICZEhV4cc3PKd
KaPu270xeK43dULqFsLxu5tttbLSXy/2hVHeUJBBy9iA3fuRVJX0vyowoUKYFb3MEma5/PbI5ZrA
PZS9jX56nMDjGBPARvlV62y2UXjk8PdfntuR+SwGrTjgl/LdifZ82LoFXu91OP+qq5Pg1bq01umu
VSQILZ60e/1hLbJ4WvwzpBvQl5v8SknA3PMbGy5/1BMyO4eiMCAXHR5xHJswCS+pxrK44jRN7IFJ
neWI6UYrBz9AQcJTByzR0QvyJnXNf0fZl2DiicCwEIIukvsbWARnP8dfWIbxLQlbZXsdiZx8u1NF
OkmPM/6dtVkm2m4oJPRKz2HzwzbmDncFDcq4DyH0Bme8FMFOoYngzEVrHhMpn75CJyxKTCVoqPOU
6HsTmwu6wdtaqqLh+7VhOkNpAbw72Y6x80K7A6uQKoB+8T2NVQnKh5/x+scjwI3N4qeU57fBq7Vo
L7fPO++evPB08xglDjF/9nY7QCj7Eo3XzWfP5mm1UkSU75M61pO1kb8wliAmPL3uE2x4ctd5uck3
b7jhJ/mVgCJdYHgf/OIl8jcKoo3Bw4y77gqnfMdT+dUGpvRAdiSw1J9DjFWsLt8aR/NXckEWTkHZ
8lr4u3mc6g5pQkJmk/umboUr6WnnB+eUEg1vtzfWDxuX3Vf93yPXEuSSvue9pQ7K0aDEgNS9lCQJ
BqyPGUTVz8Yo4SD1UtiXCm+0QCp/dpyDS/qofzKKEgeHN7molIDA9KYDtKfAUNwG3nBtb60mOckZ
trc0pJYgjiESgVqBnSEni7MTE9YXkt2C9n09c8xx0go4u5OP4aDvY7D3JCDRzJFsVM7lGlwJoMMv
WHQ8VTa9k0ICySCiHKiZaz+bjg7QyZpxsT8lqDlvTcMZ9vtnjllhECU6xgpNIuUDm4h8Z1HjUchr
wNNj9oCqlMjntGbh8U35uUob0DyV+symaIvt68GANdaxjDGHcYxK8YcL4MzT1fK2yD/3Gt1U/HLW
oXOsaauTUX5CF/6Ed9eRQaw1nUutsbksrS0u1oEbFuwn8fevQyY+iMnoE6zuKjneii+Ph2ZUvNmr
vgiThkLiRrYfIKXn1LOJv0VRsB0CmT1xInq9goyyhheRlFuMgEWQV3wZcHFu7+kblfB8NnGwWuqq
RFOrofok7LmCStTSawH9WVOmI3UiXNOjAesKGBD3PKHNPzfQZ43q7bUTOaAQFXZM2vWO+4aZ+yyi
eLhopn4sk/+OweDrbdv2caiahVDx50N3c+MCzfl8GUuv32/bykLnDfeORyHHU5HrrozAYwdrtvR9
EbvDyV2G7/HQBePuWnWVUXh2zuFeUOSZrN0xlKonUJKsMsoir3z30UnNy9f01YTfpy5ket1dipaW
7KdGe07ilZhmdsNPuh5EI4gPou3PCaAtcUSd5/O945AtmJ4qugjthXYyjZfn8bIvumJ7eogkSjfb
uu7m4X9yMpvUjY5VmHfBgzcmMznHuebtM2il/oVCOo3ztBy1vRZLb0d/Yb7duOIOV5I2gAUj9dxY
PPOTkO2Bcqq4uCG73Z0+4X3cYZVAXOL4l6/RVW3PNU0K60q882ZGhMVhu/BS4nCdE2z8/ZkpZvaP
OC3DscdqO6aW/K8OVjmLHFHz1u5SMrD1IoMzb2P1r9kx+W/SoMNKlxAhaiA3eUXiTXlwYjGeS+vT
9KeaMeREXi9DlU+QYI6nDu/KXOqgXQtSWA/Dr/4nTs64NvdagpuwI0EfiGVq6s5EzG9/byxEIzkA
Y0W3wB0hCeX54kvy7vF27vc9wFN6B7UH0mpnv5C4AQblNks8Fa+rHv2V+pwPmYcz34f2ONZzEcwL
Xf0NZr+XximLS86bCK+yZcQJZcXhSAv+2DltSyyAysRvDE90XeJ9vT1X1ZJnaShZEb6wj23WtK8e
WJs0A0S9gC1UkjxKr8ulgyx0UlJy/O/7UH33OCVYzH0Xiqn0Ljf8WJOG37fzCLXJtdRMwkVRh/5D
HYW8LHEFTyOLm+obewMeOxKHx7PmgWu3QwDOmG4Cf402NAsMirD7dKDeS0wpwExCT7AEeTL1qWhL
PipctMt6XX0sMf8jWbv0En/qhs8JJLJVOXQlxiBx8gZ3Gz68pc3fgu9U3OIUOJrglgh2r92GOqil
4KEIi4BKh8RcXMzV0deuyrNZ4XW2PaJ0HDd0swqStzJvQG4oPsybwarvOts2/+uaijaz3yX3d5Hd
hfuiAdIVbe9vFg8bEx0MbEDAVDwiKT8sNeFptuPPIyfNsRZek/wTyC3hr9MPWXyV2Q8Alalsh8lS
UjtvE5w/DwjNsiCtNhFtm/xKGZxfb0Fwd66Md308en5x0GxRJf3EVjixviQfhHnzlTlpQ0do7n1l
Egh5Sx1RXyDx+iWOxC2ab11DjLnOCgNd3ZGhkd4PHrGtMv/UZR7A8bU5kk34JwYPVTgRHCthVjBk
JdjYohC83FC1E8v+R9beCcbGiDDFrcAKS/7KjfTzMYCwqgL9255oFXZkfMJCNJ7b6d2Rd8SZdbdI
nfeKe1GvuC4JagJVKxX1TfUf19gGzyOTka3tM6kYmNsmzDpkCIag7Eb0gmeVTET2oQIKAscebVwl
xq9ek0ffFJiUCNFsTMQFEWwGLrHBGNFQq7CDIt0CegR5bg3vwuUzNqd5MM3ikePE0Fp6ogodZ6mk
TkRDgp54QcRuEoIx0bO3sG9BeFN5K8hlRaKp5sq0Gv79uAB0uUrEeY2TgGBtdAa7Pkezmjze8jtx
TJSmUEviCQQQ+sGzr1iXvC3gdM8V5v1/dVj0uJE/liUfey/aeUUEsYcZUr/dK6DsjkoejhIzDc+O
qM0Ri3vcpvukBeygN0sZPfO0EgIRdkqdr4jC3iSHvaACX1hnurpkpGnF/4t3Wn8fiszLec09ZU3b
smXUtTa58k2PtvH93L3Vu+5/S5zsDe7bQ1N+nZBx7GaIjnAH6hFY/41HTThfXuKbuhxEZUsWoIKX
PzvD1QoSkv0Lnheg3uBHlCLVbn8MrPFKnSRbHGJBaHR6QrggFBLyvMY4iaGi1JrnGxm3mOAGQ5Hj
syJjfoxeqXuU+e4wIdtPekNACtsgb/uIR+m7IRDob9pWOYnXs4hAE21bJIzb1rSEXqeder6Pqq8x
PedzK35W+3/OpeJz4U8VGRV4EB9lhd28pwnUR0l3jdmn6AYpkawuW0mHAY8aV53cF2hovCokGUts
U/6TT/78qxfReDC3WAK4ks0OZ5LCjNCyq/zSqYKVFMllAaV64I5AxR8fZrGiclTi2Xmp7KAxklSC
TenNzz08wHl3ocVrUozJMcGTzOWI9Co164pqTf5IgPfctTpFhDHOZn8XQ3oUfzFQyRcb8W8zgmAZ
5zFzfhZZWE8Tqa97B5e4VW3Ug6iY+QQJkj1YqjHTwsjZatjSR+FkmY1AoXRQ62XLGhoQdaQRubYG
VdQ6YOwd6ob3JW0MvXtMhAyUuSpdaDjkU6kfjsz05u1JgWtQzpZG7izR4yPfkfNaeNUj6i8o5rOV
mQP6GilgFAAl8wmHt3hq/u1pG5ORQ4ywdNWrbmJOmxY/c6rajttZ4X71GCfrrD+Lge6TPqePFGMO
OZOcv3VB81TVlQfpRPX09PErhul++1DqhWFWTAEIyhRQ78H4kD4/yvGRPQ/saurRsCVJ0uM+EhfX
DwnIISh0aXngX39iG83beHTNyCCVTMYOKuIQcJkyCwFnmD6YncdFD22RZaD8FbhSyOcHFuI/0uae
D9Soa6xXECQ2tZfMng6Xv7ra+6uz9nHvzu9wQfrLJ3YQmJU6UUC1xNk28tLhwxUZboA4pbZMDVX3
vL0fw+x+4/lvaMB2Yu08pH9YInPFHSXldIas0jLucEA01PgyGEpxLGbh79QHimRvUIq/7EiA3HwK
+IFXTXecf2YjoU7+sTzjviBTwRZxvzNLCummbyBEO6Fqs6JXZDUpTTvd1FTzUMtfPb7zZYOKLu8C
O1ihxDcZM/2A16dPjEGWZ/j/0ONbJcKZetHTWZVQ4JJvyJV7SJ8L7MiTft0OweRhMNojIKRknX+a
JJDnkXzS35cikEahnNv8d4b+DQHZTZp5JB0hSgWx78jycJTpylCXbGDzwASaKhRv+lK0IAIyqUuY
uOWJQndviFnU577YIAAYkPn2o7YCCteFNMvtTh54yt6COwsUxTWjjpT2cfUaQGtPWWJ0NE7hSMGr
TxcjNAlKb9rJ9048AMTV6bS1K+ZVr2+jYDGdBe2zcOGJg6YwW28V0jdvmiac3Oj9l9xMWYq5wFY0
8LYHcMM6sLo1MAniyvr5Xcr/hwJHcB3xDgXdNt3Sgf+ZbalJGIFtUCMPGlhgRwHOJtffYRZkixkV
RWpWfaebRHSVVMMpDHi0/YI6oaN64le+mP/444bV1Fu9EY0Iv2uoVFPLWgtV60G2LWl3njwoDeht
mP9WJ60GxsedmWylB4FWHdCkQZQsLCNQomGGe6R8IxEs77EaXovaaLdWpNMC5+A0q8yFfdltSVyS
bTyh8e1iduOoaMa9d/6M+JFVIZNzJQJTDohnBHuRl1JG/2oQvPY4vq7add/UBjDREC1Ng3xzi2Xg
mR1iSJikp8XjbD5PK6z4O+Nsi5ZGLSHAOXPWgUAJiC1s2EB3ghynwDpYqyxfjWqMx8qPuhIzesj+
RoUKo3iWrfcelarg6zVl5t4aLtk3GXJTZSmzebI/VV9vC+CKCjqSY7O3zMbuDbcLej0otWjUt/Eg
dbBFt7SUfxRrJanAftjnBUEyFkyejgMR6LLUXEZ0V73McrwrXYil7bLe+6i1e9Zk3iQEdMkYkVvd
SgQv1Bc2BIzBIfbCYFaW6Cq1y/UXwSqakrsJSDBsUSfmzfqAfGZNVXj+YoZxxg+r63kNFHYeWpMz
0vhXKE0D1Ax9Vv3AUj1pt3jpcScdAwlHB3uul91HCSDfmZBXFbMzamG5ZpHGVA4rAgtgMB/oilQh
7RF1Wyxu4r3PplnDzKHYm3Q1vKpLzM8YQSfL3vAhFCk1EBkKFcrcs7ARBjFhbeOVGk6+Sxjd3Uex
zIP1ORooNCRS7Voa/4nLHVUDJ+So6Kpo39qpd9zZ7ItkQWmThjQDjekII4Q0TQ/56rPRF51+QoLl
oirWie6VNTlIeuVl+7qOPNsXtFAR73CSIT/Q8fcqptt/02hauZSmmA4fi70VFz2Qyq8zLbNxlLNb
6jt9dwqNNnV06ZQP9viz6JihzJvhv/58blwFjL1/rQ4cwXHqDYG6zyhqR96qMW13JQiiccAN/4fZ
89BFgWzNjFzk+ev3Fp83ZZESjsEsP7QZruU/c3TI1YpPgggoVyPFVhvGo+YIv6WeS9IzSS0iVkOQ
zyA/l7YsOmWqRc/akjbeKH7Fqb1SGoNR2cM2hfQp3FMNni4MCNaDcAA9l4MEs80j2aolljPLyn7Q
2ohxk4I7yZk9yM6Qd6CmFlsHwvPGfV/pTAQAD9uRsVZdJdJh92OmL1oGMYTM0i/lZOO5/iCfx9W9
AaETNq+UIYiNw4QjSiRonTmHJPjdU+pLYqdxaHc3TrEVQlVzeqWKO/3VqL/1ErDlS35WQ6JWy3xU
IsvO7otIe4V57E119KFIHtAheFfpbQQb/SzWdKevWmLHJ/8rvxj3L++S+6RfaQLRJmM8dgSNkyWJ
ZnpBj0HP+wV+KYvQmvON4jx+oxe1SBOjSD+TdSCi97+0cBgYO7IbWW1svGAsIAc8jIOwILNS2Ydf
A9HSg2ElXAqwTK9UR/nCNIhKpl1DDVMiQZjZmUCjjuSI6QgzLVSyTKy4h3QymZp5ctbfpd15BnzR
aRkVCwoGmJndV0oCCaD6zVSU4BskslLu6hjn6CUzCF8pCKf61GAAxGN0ObwGxeM4CybFi9Rn2vuv
Pxw11iM/f3iivR5G9YcyIH0RsGPvvnavR5Bg8mUae1Ybp/G3+CfcEZ2Wgqw+B9vBK1A4BJJfmVLx
kaXib/DhrqNRt3k36ND4icxEzrU02roFZiA1s/50urV4JK+NumVc8iEc16FRpbHP1dOmdxQg2iLh
8d1RPr6TuI155cxUSGy6eUVImh5bHFo+oXNqKMNkxiaOXAGJE62GSA13a/FG8NvoYh2/Xqf/n8hY
J7xcGtdfQFNXXpmVFfnh7kIiKV70g7Wf9a5UGnU/J0J/wmddj6fVGtyzaQysoapkjPnAoNaKyCnT
D0OsvaU5tW49H7NIM9c6yH5MFueoVHDNxU0p8mRn2B1Yf+NJQLv+Lj9gEI1AzJMcyw6YRKPvVceW
rBUb61ebZeWWAMTDoEOOo5JTX38HB9ffhdENRNNUkzXMRZd4nmErqJH9Cxlz8jLqEftrnWrVCBfU
RqoOV0aIUUmKvXp3oX5ByDixskAdVSY3JB4Zy0QiHUKektVHPawAXtKnHJ1Cd9QFfLlEoOqTqis9
J23qWhc1jlhD0Q3qwKKGOb9pML6FoaXQfy4hoqhF5i9xzUQNRATfv0Q9hu1FLbt4I5ydRR9SqQ6h
KE0dvY3h+XNnrlKRfgCkXp3Vf9wEpYnJIc8Duaq4NLp6Roz5TKiNTANpxZxJ5CtJ/Dkk4+XGbVX2
3XuN6RClimGl2D75OgkBYE8Li8DhpQpsRyX3Evs7MedJCm/1f7dWJIxLJsuT56m75K2EMSoaxmCB
iO/Qp9FeQtJAkAImRNs8Q1tZ6onr/KhQ+aiQ7F1p3uIRjY4XdsHdONiTCQ4CBS1X2yekDVVXE8HI
ipBHX90LMfCAEiWXGTF+ECI1LnP/juxhcTmAS0WmoG6PmOQ1RTFvP5/YfS0DYrQhmZwP0miyLK2h
MR90SgybiJ1EtfzYYouAW0GV5gbRiP0b7eX4eZ2gpDnREcEQBDK7w/QeWsw0ci3KB+cYt436VgLs
xOQl0LHKkLbo48vel3i8KYkrt7ZLow+wxINRGIU2JGY/1MiRdFwbyc+R8kUXJdf7djul2/eCEhTZ
MJrdCtSlTaGZZ0oMSrqxhrc6tLna5RMF+6vF0GWoGo2WkEgz+ZYEEb4tn4aoaiSRgzUBKp5wZUFv
kvnJFNtMXrkvJDPEGfFu9niSYwqYdtO2l+5jKcndAXN+J4RppcQDZ5KacvrD+fj1oRGHvYF7R3DM
urSD8hJ0dVvV8/WVTM7aBEKSnxQmQKia1THgZGa5HnrrRCnUiEJTXNsfCEGkTIYY+7hQy0OSmV3Z
kD+jU+IOxuT4b2WqOA/6sCXrzQRKhcqLKYY0+5jgkoi32igsxRLjgVMfowSZAEIV9w2HXRSUE4fo
Y4fZCpWz380qqFmV0eZ/In2g/ynBPVXFuU2rd+dtMGhVohupvaFFv2C7BYAg1nziy07fyr+SETZ0
Fbv9Ug2LBvAlsthZKPM4H5xfh1Sc6S8vTkZ+qe6AbA7vX1Osjv4HpvLEvvTJtMK7LEeqiBPC+U+i
lFwgXLMyPxgBDjQiFcZxBQRr/rLKqVNr3zeGbCFUQzDDhd43eVGapfw40UxvbKUqD9SpYIUIp+cx
6VrEl9UCSF9GCNHbkl6bhcPRdTPyBO6Q8aw0G8IkoK3DJYmEzcGZhq8FlgaQAfAakyOofaUzJG1+
PoaH51IMMfMAmCn1kZfHw3Iuze8N0vQnF0Y6t6hgDvWJVF/fwV4YzL+qy1QDuBRa67JPid52NXlk
EPy1/WCdVYUl89Hd1d7mDrywivWoDoD3mAuXotivswsEcm2p+ubI74BrduO1SuUvq8ADm8yzAUb2
TkKzWKb3NcnohN26QBqzMKdxTje7vp8OdDWTwUJNfWQ+Cmgs0FcSSEV2OF0yxHB9XmeTHO+nXPAB
2hrAS8A9XUr4GvDjXaat0XIYSYzBojJaHlubOJFrau8q9+fNpYLO6OzywTZ5VtlIEW0WxNqPa/Ij
LqU8O0BZX6e34jsMdFmfVnW8k0myKgVMn2aAp3ocTC3TEBALk3AOob1pHF0qxkDHZqM7YN/RHo/d
d2B5q/T70z6CtDpzZSVyO60buD5352Wtys5K241Zexs2xFan2RGGkKW0PQs9b2NIkf9PiuV7ltfa
va4fF2NLjrCT4lioVZASeyodeGMyxKGwgFgdgGXnKwOHzPAeH2H9FlaQhHQ6S9fw+lugRPRT9IGN
aqPMaj+CG3yGqpzD4Vdiq0vi6ocmN+aY1JOqWIPXjchdtvAnyoReZrmOOUbwENPxUDqeaxymHAJV
xM8bWMKwn8J+UDPv7EcNgc87JkSTGhuGhPJHy6917yZOXkGAnnoMFWgcz2nU1s4Tqj1G8SzH7UsB
ED6+DUav8oqgn6nBYHuTLQdF8KxSgEEswkC8N+6Dr3asJuf10aoMTnax3HC7HwNkcMGdxOqkxBrW
Vy0X1nLodht+D7S2O9Vw3kzxkrqTyMjwHJyNucmAvNB3rYbjMx3HSQhkK1pv1xSMd5RUHNd9yCdc
TDaD/Z+T/YOG2/DMWEyF5HecnUXHZtiXbqubjXujmkjkRo0gGI4oWTeidhyEiWf5F26WmHmxQnyI
R5V6ZjQjYvkETFwYokxNweM0xh5xnrdFuu+p6bIVfiyFR0hBkb52Zkt6G43ueeMA10sDsLHTPuiB
q+Qe9kSIktf/Mx/FNrLHO7mr+9r/nuhButaz1BFaTnn+1LS0CwEgn0QLjUyh8Lac1NWY/YlGsnqw
DBgixUGh1/VrSG8lbzlwxlHCIV+8tCmNpcDePXwt54nJTe5Ry8iXU8VzYcXylF9Kg7QDQnO+Jled
xYTuBwfG4mV9y48f6M8SXZFOdyIJv+yKpgANWc+YSuQSaO3iXaWr7etM4SIc4vSI4c818L75XRkE
KrzmQ4S5kBXsfkIAX8YmwNPjexKbvOvQqWU41cy1xBYZ6fSiJpH7RTUgFwTQMVDB5Vyk2qv7uTBP
s/wV9vzQ7mhWpTjAZw4fyVtxmRAKZZpuS5Ah3oFo2Q2V0ZtbE0pBRCmWJLLIrRzmIbkLyrA6d25v
S32QfiXCDa87d0X1Sr0/IYb9S58CPrzN6sijA92LyGFoo2YvyQo61lXB1TpaLrpa38gFJzc7qzn9
cATI5s0a3qJhvv3WogpIcJ36j3CYrHXvOFWq6liiiL+2OCLEKfoTcfniVV/uRiv6MSOWVx0ILBv2
EF/Fi2vQIxRzUdmL7sZsIN4u9+i65pJ5vNNsLBhNHYw/Nq5czer/Ysbl5ro7BwONPDptSZmQF/9l
fn9h1kNAr8O/JK5fUp/G6j4wr/IxcOaG79EGC8+IgqU58BvWTsZcJ1+Ud6QZl2rW7rBbdcFw1R9T
w7yDrp8PbPRx1XecmF6zbV7cK0ibRY2pk9DY94FUZefCPu1F5IEzmdLX7Ob8JQAC4kSk1opeFt9Z
cAVcmOgA6xlx/4fgm7ncyo1cpCxmNT9ZoBPfaTB5IFgP/EIJUVY0csooQhkxAeTom9RxiNTw3u1A
sx8iDFkzov5A0zFGe/QLMPrdSOPo1jqgKvFMFwiwp74FnHGRUD2sGUNS6jRKbxRXkWBfbmdf+fjO
KnG1ooOuTC8JGuEQN40aHBh8o8hbMh7T5HvDs8udc+EqOt2egoEiA1JhW8bePrYld33ZC9J3DXgt
V+Jn2yD/fX0hMo/0NiyCk2QgXPHNhs807jtzsOZjbAYN8P3YGjC2SK9mJM3sPml9PPx6xnKIEQV5
P2zOlHIdl5nJLhorDvJHo3Grl6jVjPfjhoNBIuxNjAn3S8CMrGvxi//8AXrT10I0kH+44xU8jFIz
xzAfSgXlQZ6hsTY4zepEEkyzVu6uRE2pihQE52ZGcTYgJcPszFxxmzoCYbBk+F3mia/OwU4ICgT7
q+s1cA/qSAVTjwiN5gSC4zZBi2xdysRM2ldPSQQzMe2527792WllGpB0tjFp5ZXjnntYtE816fvY
dLCqEfeavqDFsTFeIBHXAOAFlcKyDx7UHWvzSnr01V6TbrisV4oVRqgHDWCoxhQ0iXy2aSommvy3
S04VXoUKlHWLYDzo+G1Ro/uBjnYPTwHrPB9myLhxWO3CRmrxdurfvyd449Q4Fw14KZoGEvyTOQ6/
LuRuwOXzruJK2KQ6Q2PAfjDbnjJJKFj1j/iyLwHZLvg/qvPdZQ/kqoCGXEatKYCT8ak3CDkTmeI3
1AMLr+3pR9C/IBNyuOcInySQiJSJuOwrQaCXRnQ+cjd8TbzSpNGIgVJ8ihTkSYKm8cz5qxiP2RCK
OkD6TIDW3APjornaHZ7CmwE09LD2xDe9+RTtQs3TbK2/pDYTQQ1AJq+ggGRnOScWpMjLky7bFUWi
sdI7eNGRD+lPzz3euNnznP3r7yRPoUjakhEprxLNvfFlXEgcz6re9b6IiXQV6T911dEgNx1I5SNf
SIWnpIS64Gp6odWh6jjVC01/LOHYhsXYhdtsbNrrayRbT7thYy9KAtOKdi7e28DYuvENW+xt1pnB
T0NFn7WLL1ifCQa+gR+OqloV1Z7fQSPgClX6JniQH9O0nRGJpJqs+I1H5K0elZfVW5tYomyAhCoP
VdMF59By/mAH6fDgxCi9X3tTY0TtUAaUzCiifNUFb7GmJPepfEtLvJgVyfoI3qpm1qYucV1ZvO3/
6bxVw0dE5aWJyntunr+6Jd4VMUEBjFfFz2Wu/B8paQZKX8VMJf5GNYIGB+fO2WFsycSM8/1lON4m
0WhnihZRhQPHYMOzmeazxbBwojXTbdx1Y3OHzA2s4DlPk44v8/K5Ikpf1Ua1kAoycB3vMLyUEwdF
NiUO5gZqwkuzumPy6eipsmCY3JtN9I949yeo2llPVcvIOioUt7Hu9Ge/tmwlQeN9WduGaa9PdRfN
Fe/b87dYmV2KM9Cdu1XboENKCI0E2tuCaC8F73fi6aue2FgdTXX8lZNW5Pu2DoeCODgHdvl9FKgP
OyqLPkCjcsdFn10QO954tvtZbsnLpWLO/Ed45ZneEQlT1pHCgt1bA76rrYtRyUB1atB9Y+2QzqwV
K66/2lNlw+NhR8jZ65mIDVDWzwTaRJNj9HDf8X0Hddwfkgc18UZbR4CFprOoRuoNbxXWDkKVihD4
aoeyA7/WWvubgL4ylAbSV/4ZewyL4JEsxuX3ocQ/7amB0Mox9QazxJx5HLF+I0hy9IpSS88Vjo1e
0pN64OjScd3iyg+aSXkjKRGIr3aY74toPbKtd6OwYZPSPHNZEQNATXFmImuf0cFBwdoAXpwlihts
uJ/JLu2v7a/oYfvFQ2L2f1TxDmcWe2luKCyotpWJgJ01gkagPDIMQVc1+vdVqjsLgF2eehkgYdEP
QIRsJ0HzV+a610608GpZCLSDwbiy5h+D2eT2zAv36U0X4dbzE1yf73rRzvW/Hke3wa0Rvvs2S7me
xKMzN6fdkOnORlpbdgukBu5AEFEhW1VDDzOsR6WW9K4RzLer65SQE8BkrwxGrBEobJrwzPFzaThT
raXvxLOvzioATaKdw1xWYwkgpn15V5rcp5/uCEA5cd5Q0TNhKK95INumwm1zpXR3idL+LLOJoHQ3
nzlrodhVBNI47+8KqD9R3MJfZspg45mTvhTVnLBw3MIeBXvIKFY3VLynCQXRTlll436kakgPv0dq
7CjnjSzYVDjR6Z4fcgn2gDVjjyvKXYDCplgYpZrtnWsFvvgz9zjKAq/gheYtUFSRFrEEIcjjPLmi
qV1U+3SoKHacEIcZ8r2oHipfRfiAl6x3RNi6a+8PiH3Z9RtwhAmzWsmcUBIe9PLaFSHY1G9h57+V
QKfKeOq43SzXzzri16KFJZ3gRnsTDfBDFEnP6FOheYF5HuKH4WLPShTndceX0HRFRXHaYH6sTgq1
cx3jYEorM+jbmFUsPlqapOuWfzpBA4k/v/z6vbchVL0/6rJeIaaK8sbvmll2UrjZJ6g+80n8C4lS
klVVJbkpVaE2WO/MdGzMyxRoeTMfsQtPqGJfx8GvuB/3tz97n7FhcS4JNNnDjMM5vjBhkeb9yxrj
ILSAs4x/4gevov2nLlVNYcOf9xlBp2stq3qELSuctYlrnN0H8SOU2YyOsnQv+Elg0DgI7UqL0ELG
O7/L+z3fIsnyBENZGZvV86rBmSby8yQCIvWBHhiMGlvsbWOeXX4LqcEE2cU+zzhGfcWgek9RqZTo
DDuAxSJK1Q4HD2c7g39qrRAnIMJ38j90hB2Oi502/hiD2jQC2Cu/6HJDXtf5iA6zEsKNyZ0992px
nYPmUTMXRpEa2S9hQ7LLRIREugKVggQcPgrvOwJ2cq+w5xBTQmZHb0K+tui8ME3lo0Lcsr6iXthM
S/BZ2JJ52QOUqtY3QdK0az13FWdEWoy+W61Q1imcmmz9zkgQwitXfoahlrf+1tGN+izZSDtPBGNH
67PD+Gs6O7RFVt1ap5FCrxHeyW6rPq5rLuC2nSQwuQ/bE8vqTsp2AipgY2bCSodRYObXd2NM0vxG
HLeLbjarE1+jgO0eQemfuRzbsQjCZxpH5jTicTTy0QyxneJYhlcIUY5fG6eEIgcYK3tjpt9NBrPY
APW18k0Rk5exdmrCB+JXEnXYIaRkeb7OHrUmLfUxjDlzgEBo7k+cm7D7a1BghdxK2P+xmDZp0UC+
OYbFiWTIMlqBgLrpgRyf+HBvpFNL8AfUQ14/0Orh/BMq9/lUxOmrt/XXxd2BHE054HpYwbWfA5LR
+Ocrp9jJKikPffq/uhy6pwpO2Tpyem2hxBI6UtJuQHR3LlVxbz47jupBnJHMPe3rITaoYnJJeX+C
8l+NL8iHSPtrJOnAhyOAA8ATAML0Hn8041pgKWEZZkd7vX6GhohrDPXqk5i3VHCGU9KOV+5DxPQg
8MwRMRM+zV/v5BX5JCrxGa9yNfrvSDyLeHM90sMnMr44I+hoYJD1Pl0BOSeHJ3Vk8MTS2HK1+i4U
6seSEe5PlAbTDoDaFbRQuvd8AAJlgaeSaUZsOqliNgCxzMt+o5/bAj/VnEClD579MO3zoyZcGCV0
ERdfhgtZ+1D368xTrz0gsOiges8bKE3DOec5SBI4mxWhU7CoFvxKDYV+i+LcFiFZoQSwb6QUsSfd
1CGI8bgcUCpJDbj3hwXDCi3b4d4FoLLGzQJAXSlyxRilWdMbrtbz/8Sft+zSZP3iuXmWJAmoHWKK
/VEm90eWEO1G/nbo+eHVcK7cMpCAz+AO7uTFoLV9GdDtiaANdxFvwwnBJ0U2qcAsP9YPvTBcewGP
R1XSb02UnbQoFmvvy+Q/GDpn78jzdQYWaAruEPdlkA4XAPkBfzg/w0DW8GUGK1dhzIoFQB6Bo7rL
DJFkEc9jylsVLZiT7To8+UFjK65CCXI7rcqQPQs0qPGTlfAxBHQQ/HlgXULwSaF2LVwppWUkeJjy
sPO1H4/mRRMU6CQUG5Qo530x5y3y0pCoB8zvb2j0f3lF6QX1MYEvZ66+W3NsVr3r2/gQWyfOkSRt
uLEnaTW+wb1wiSh4HsPEJt8TVzLcbYeKpmicqy9dNDGknP/P5YtW+QiQ5SS8VKi4BdKkZknhZz3q
pWbCcuI7g5w0xQX/7KpCaB44O4pG/535d6YVY3YlZf4udekTfzymI3s4SJLD+7rBmOytjsT3jFPY
xYwxDbYAgZyO/jqVjV014rpTx9t9wjQXjm9KrcrCM680gFNYIcfv+Gh1j/6jUMi5DiAgPN6fWd9P
3tO6oM/E0Y2dWzNNe7RgtfX+wHw3QaNaVIcEmcvSWYIUcefixNlz90ah7OT+g5rtDmOG7KSoPlv3
maNAMU2EAh9W2bSyLRvFW+CxLsNPQQJWSsrhBVW4sUKmMsVmEj0aHVDaxFAbudBohSGB9EbltMQm
OsUdpnlqWuXbvAdiK+3xk1Q1B0LinfePBXp3tdskEcd9J2M00pU2SiaZBa0PFNjVufqvd/IcWHfQ
1WZ2bvFiwKwDNb+h6Bqbj+RGkNWq97GjvOgS2OLX+01dX3qjP5Kg9VJwrIcawnaeT7Hodt6T43Ii
q6W57PgL5LsdOr1X85EhpcO1/spGRcNhlfHLnwuZVUChebHhpzUOD1u7Q43A+hIl7v3HIoDwIXru
CTeHqEaompNwskjCss+Hb5vu7YX/+VGK2qQczf/UGrpqpFFFhB0q68FQ1ROgvcgTIidbzd5KEl7q
S2C+gi1AydTMatu8pz0ZrVD0csgqNKg/LYZIzcUpAObhAibW5Qm6s8OUC+z0KWdi7gqED0ToSz9k
k2Nho/2WvxG4U5o2wAEgMyPDDwSsRdwuTqYhpisEtk5aCnlvt4b7bStFbrJKHywK/gmv7Cj2Llm7
O28tYLVmZ+VSzH9gN2MwaV6cXascftGy3/6wFvuVKACGKKuoUzSHfY5snLwnBfFS0R0iKVgc5W9G
HepxRauTfbF7A9+kwzgqb9CLFQoYkprArpZv3yhPdAuzA+N/BeUIJ1kFhCjaqKPW4vsgB3xpXYcL
+Qb4jyF5NdnY61cI/ScwlL6OtYFVDbZ7vGk5ZbuzYwbX6PdN0MMaqC1cGp3ZYlH91mH8XON8leQt
sVUR4/dMHE0MXDxnItbbFsSMJr/CMrUjWiY1DnO25hlV1Lj1tMQrRij4+9eXYtYcrkzXkXerA5l8
eCPSh7lUi/MudRzX8kUNmXUmhwUySo49K7F6cMWtChWnTjG46Qz/qaYoAae093f4Tg8qvXh+yKif
orQjHIdFhtpcbgwYKqF+jljWk6DRBFZ/J0Ls7qdOv4GW+s9N6o1W3RaIXv7Id2nnud9b5mhbUf1X
XXuFm+m2nKzBTmpjcKcWZyOX8Rkny3/Jsde6R1sQ5Uw9IL3EVwai5JPNJiMsbb4ecW40Dmy2FuBW
MAZLcmlNhtAWlDlMcacyhxwaOCKSg1gQwainvGMAVFMd6T0ESji6BdYGtFXDBs/8bF8T/pA3DcSv
iCeZowCzz/Fu/Brzdh8IXg1T6gsB+lmtlXwXVjouMK5ZzMA791CcfvHhJpPK6AcVdrXiGOkQ06Wj
UgBiR5MGBr7y26kavG00WsTtNjmE+pJKhkeomr5/bmfgu4q8X0qT2ny8J/xBy1p8mAk0V6vddotC
XprE0BD2zk7cErKtojPZqgHvLOIyiItZyLmLpovrGpqMdrGCOqKk4hRpLxne85tFF4GmMFGPd3HT
myZYeJr89LM96ThDcQuUiuxpLj0gxwyFVto8YwEpOvrrA/DC8lHPbwP1v1EzyD6/PbL/YyLT6vhA
ClbZHg3itkOzcr8TJ9hqBsqNR4NVPkEyzlYCwz/mjYqp3ULRP8+cDuw/Ka1yYJkmo1LC1O9jPPYw
R5umdq4446sMqPGj2Wjct4jig8DqSh3adnNAYKdcsCBkTU9+AqhOL3oL3FmX+ydD1IEhpsmpK2kh
yXs2xzS2HlLmx/Un//S6nLS5171zU+jGjTAitc9YkI5KxDcs8Aonb4SgMJWdGNMM58rUvskkNfNH
dqqWU81jg9qVenMXwUQnuJKEN50STQu8wnrH8CL8WbW2lR9aLEzyuDW8Uf7bnIuWP9UDtGCbG0wR
cgB9czck0RnQogDeYmZWPVT6h97SlznCXwdLPhuNmDJAhUEhXYIvLdYlgBlGicSvkUru9eVrpTog
sN4G75L8jFl3aIV/GfAgA9LXe4qJ4D7/ZLGttSGirct+2tGfDfRO6rT03QtfecEgPo4S41C9NK1s
UMsu0qptwkGLn2ngeaEAg32K40WBJo5WRAZuNoxgA4pRZXWGX5NDUE4y+qc10a9bqgL+7A6csNL8
JSeMcC+KtGysc1sRTvDt40r1mdpX9aYDvQ0pQpLwkO+nIT2RMzLJNyDiR8NtTybV4JeL0fHF2Rwf
A83/88y6DeTJ7EmrJene6dozNQ4TPvrxTGsspW4aFxrBcEXB4Mm7A5dQELVHqaTGB3bBJ2W8j2dY
i4T+c0OIPvgZCyboUu3pptE0AfnEGglm3KtZizH9cZVVj5i24Qy5xqAT3Gmd0dSE8e1e7b7tE7gz
O2CLOCF2g/x8lZI1+EtmBrDUoLdVCBBQJuulYbDn1PWSK9Jd0G1l0cuccvx4ype2xGTAx8XcvcSR
isr8pDLjFSF8h/PTrbE3EbLNKr38hieAEagMmWxwzT/vqzC64AV/xdAWsa40f0jJeTrp5xk10+Uy
kK9uQhYMhAZVqci2vYyG0+INwwoi9CBGRFXvw4SnNrod7PUJdtwcRzXTLjtITZA+h7FbVDn1d39T
qKL+t6fkCZCTTAPnNnOynCkMtZ7m96ZtyWzzbUxlud5ejRIaOMYAzL9fbu7iQfuI5WmgyFdsGWHS
LiUxCjSVhYT6SxTXw3TXqXOWK3PhaES5Z8XS/y0fNw/DRvM+3svwe+2hLn8cUmoBAOOtAwY1slnL
nkIpCWUvoqR/hpvAJTuVyj58Mu0czKKBILHf4/dcL3QrVfjOqz6IKO3F1s9yASlxSHU2mnrZMZxW
Ue/86U7QvBf73iTGQdB6HHP1WsUah2eDs3tT+D9CuteMehSFHzuL1usuRU07VY/AWkKDG67cENv5
SgJfHJSo1nBDcfv7ubQAuwVs2+B3qwaA0vgwL3W9fhDVmTeFe4fCqWIYdUfVLgK6HcyflUUMfcSJ
kbVi17eZfLlqWpJPl9Vpg0RWLM1xeiW8R6d7JD/hTkb+MbD95dTgbOWivZV5E1YqF5w30SEKb2HR
67wUc2Y9IjqoTdcXQZWEI7DbCOjvpznWKm6SmXQEc8IcJbycdDACtGd1ldJi2twqZg2z6VHUPUKn
RXY3nxnsshl7PmycZ0eds2BfjFUf7d22YlEKsaIxHmftLnp7DgudIBf/b42VlKVAJosCPK8Nwbax
VvaKluyc4JdN2lzmSE+I2VYI+pAFEKCJDT88cyEIPIDHWZSG7/ej85s3xXZ7auE21muAYoPrX11h
Fkoltnq6TJRi7Sgw391mdb4m2PL+Wd3APDtkvfP/PA2t7NAsqUYaOwOES0NEGaQJ432nkeINc6Zf
cEOWx8CY8BvMv14DuLh7O7g5+qd710tB3lSXZz0SyE1MFETL34yl0HFQW0xnse/FS3FU9iEwvlxv
1y1pm+qjl0SO5H/P5UALLQfVTBPWR2U6U1cnHfUwmD7Qu+6aUFui/dx8HWY/7UIJl2Kn/QZIa+24
20I6/RA+OUYzRspaWdDP+04IIHgaoAo+9HVB/CQq6ATGpY0WaGitXmyx8nCl1+5rEoebyHJG9hKA
TnRCOSSYcQpPuhLBNgNcmA2/bhA+5nw02e9Gmzz8OT4xrAuu7i8ZNfo9DOVuNyjtCXvaLcw9AUAB
HcG7y+xpfeAmfSrir8tZqTCP0VxFROsi4r9jZ2de08ovbf1pWXjo/6Dd1owzWB3svWUeQMy8JnW7
oLI1nweZKfl35PFVpbDL2vlB5MGfM60ZV5GVkBJZU20Jqcj6kaazShzyNuZ3DnEi3Fg5p91OVMWe
7Ulos9s4XKQV0EgVt1xy7qrZG3zXkgCVqxZJRs3QBR6BEHU0rk7oRfMHVkZoFSRexypWwIKqlmFp
/Nq+RQfPtr/IPEllyLUWCtOQx++AOW3x6Wf9+ZlyZnPqN4SWBy8cY+gQ/mDsgQAihXQ+CFyOhadk
jxoSHZ11Rl3t6MQ6g2Y1jENqq6aGaNWItcbNrkU8ko77KsfphavSLrhPxbdWAM6shhP79iKXwy0V
Eh0OWmZO7yZjHMA6HHrrbFjmFRwUGH1pytQl+G5HhkKvSpKMmYLkM2i/XM5/hH+1w9h6KB97ILh4
catqRrxi6Rg6Rb/8WRuuk2qJpiiTCE85edQ20i5PQvLCtcAjPafAQtwvVRvP8JtCuIGvSpfPu7Va
lxE5OgXJJxYrOWolkzRLzhZjTrjTZwLM/cUfQRASBUOtAe3aSP3yc3tfSrevw/qeN/i6VyyEx6Hm
cF5KAuEbGigImNETn2IMZy809Jg9UYi4iFKAcAnZAh3/Vq4TO1QkaHI74fL3tkF2TiAN9buZvBSw
QM+MsN+QzU7vgFW7XiJG8aH8ti8xYWTH6H1nJIvUExoaiWYlpT18AwjD39NEIYzXTBy2fKbaMMNl
jFC7BfqcZ4hm9Jky7iY+wcGsjpJ429q56znPhExUXJnqUYf2ctKviDdT8r8hMHwbN8Mo/NLaU/2X
m17dPrIbrj+cOcJz/bS1d10Qto0yegNe1WYJZCXcQqEvw+O0ZIWaeMgU+tZx7b2p2+Gjcc2CXyvR
Q5vJ3MyKGJrT2ATglK6BA27vrLbbXH/gqfKAHvGTJtvqYjI50RO3Foe35k/7rpUJU8/spndmNcDn
VvxKgzI+vp36DUVO53eOuooaYIhYPA8g/Roqdiom0wui/soSR5QA0avJ+Uh4Q9KqT9DvFzqHp7sI
vX85e6yRNhTo8aVlsGZ4BpSfLfwYJ3TntW+lE732KhU+R3+tvTOLWla6cX14CPQ/F7DvZvTLnpor
FyrfbqrfrgHryVCf0CyOFPGc27PnAtgRCJkQjvr4wImh1Nr6NoLpS3zFJxszmeuSYt/5rL4B5aeG
AqBQdN4mg3vshIv8mS3rSiP9OLiTkJDxhZx/tpgXcMOHRWoAaoAqFjs0qM3uVNRF3YgFOdH4jXRV
tgtX5e+Gg+nBOq24D/f7wtCglyWCYhX9nhE9xtC79S040BoFbAFEpUs5KIjFTfY5hNIC7j1W3Q9M
CLdJn6K9iZog4Rp4gqnpCfYHcImSgpzEihnu2XKfoaCnjUb7UXrQbb4FLbpXBZJ8ofBJfrpblcxM
MLaqzSSYTyverzabK0V3q6ZaziteCespoZHlcr3BMKJTtP+PW+XnFDOm+pBWsGNIbQGrpBJlT7IV
ZAOf3y8KoGm6csZJGbeeppJ5cIEREKIjuHI3BOgBNcRgsP1wf5CwSGoDdoSExdgY3Zrf1DogcQl8
YzyD2LuWndlxWmXIvto8gpESRTJpTAH2LuZhA5nPzQp0nYA238ks7IHIB35MX48KPuSJhLnX1oL0
bBrMjT0Hm0RADrYkYHfC4VYl0MQ8P1vOB+WVFpxmaOF2r+p6wn9K2EEh2jmEv6yPVTT6YGv1xZUY
9OxjMdt2gnv+nTUioRloiCtj/AnMV2MWRdH5Qrz5lyhOCsMNUdD+K6eC9BT+KHs4j28evQtuvGYl
ZgKqbgbAjFCYWj/47qZ8/TofGeWimOYP9Tp3eHI//QtaN5vMOQWdI/FnvahhTu1uPx4Mn0xR1Of8
ll9ghSs80RFiGprqqpWHjLUiPHpns8QJVm+kxlHrablAN5KbWmbiJPa9M/iNQ/8wdn9nlVIVjhmm
nG/nxqsrRhJbzIrOD9YtSGwtyywP4FQbfw80s4NvcyaMARMIgj/ZpP5V4AFRV4uljJa1dlS/ZjM4
Kw9uS3my5aiqnhwdL/kNt3yjhYi/Fu7Yuu4sQ2P8t9JDxAoW0oRrMWfDFkUxA+/rPJ0HZ5zZwjkv
0u1OqeWXKyN7f4pZ/x0giqgt3rkiFGUgGkbI8u2fOPuV7IVylfO1hWV1HWIEd+y+blPSRP6jd555
pwPaDZxR268t/idrifzTstww+NWU/Bof0O29QDVvfvse1JO7kkihDlorReuDjDnz0Qj/FN7gIEXX
vxKh56wBkn6hF3ZE8NUqn1s+qmQzGgM/PoVHvNnq5yNIvT+EcH//AMM6Hl+I7xvZMhjp1p/WLcjJ
/n2gRVo5ieT8L/U/cV+S1qW0XDLanmiR6sHFuFE6MfeaNy79IOYJNoeTdJmz1yDZI5L5mcDHwijI
4Gp1oP8omOjJNaW//7dRoigrNVCYLH44fMVDd07eU86ATzSMf4vXzMTx5uTRLHt/1TaxiAwSxNW9
T7GGLId5K9wzlpEUusEErphkX5GZJCOyrm2H5AdvstJs2/HhmP8HUepBglp8Vi5J1ZexGLuENpa/
szeyvpOYZQ3KuQUJZ9w8n7UYPKZieIkt293FGFTZF2pKil7OhfDAm8u5em3FTcZEouTagifgX5eG
kDh6lFzFedopaegUu3HmHtpojHh90NrQWaOyFxMKeLxqYxgE0NPJdNoFx9Dxx44Cc6kT7PzA7osZ
9VRhY7v3WcKo/Xeh/VmXHEa4Bg1P3BggXmEsXootVkLMrXkVuJvYGDdoY3X0vJ/LHy0NnxJew7Uy
HOpDAKbTdpEqAO4Bs1/PCaaLj1LviUs4ikASPyhKP3XvREqY/OBeigau9tRk4VaVLFe9xNDblXqD
ci0OuitXBe3x1UAOGdOXbOyEO/Rjv4TRSsYVC2y0N0cAod0n01pbchICw8sj6NSqAM2j06YO5gF9
gs4x0x9IsErL14gRwOQ9prJwqGSyGFta4Z/4aytaDJW1s3lwxeOgIFpTvyLum12XMhJZMhTqhAA/
3rUIl3WClABuwzW5a/gOspGl4y0cCgMcKaxsWixChcHLxQBkIiFeGg4w4qqVxGPOfDXWIfAyCRqV
psWZQJOEB8y5gMa7CfEgBnwRVE2gzhlnzR1M/Mw1hchIgfkSRgFjQk70AxWBHSDqpNIWh1k8CQ7Y
4uJvTbmo4+QBCPUqIsvM0bsM6dYu5RpyWu//vPkAUatvq64YDhGd8AiQ3iR9FhTTuJ44t7zDAKMz
RdESCoHnCvBHZ2bxO9V3Q/AY8uDLrqSty9fl8N9s44XnodPJimmf0atK4+BIjAaBcY1kYlX1bI6O
CEBBu/bgutpKTz6n7ppdEXVA27Sp86Y2vWr/MV4vQsaoSMepG9cKadEAfYQnXaY/jdPoQ2WZzMTr
enzDGplbUsVn3qx2Tr68qUCZ5ST4Adda1Rn5j/xEXa8IAh1NiVRcvXMNb3ftccCHdSu6eWbJd8mn
DwFVYH0ua907C9UGvRrQTRGrHD+TWpI0CMENh8kS1NGPnjGJyhF+iFu5FHCnpbW0Sl/CzAjzx4j2
XqCqJtug/HnWSon/YXru/e0Xv+dmAR78iRf+snFH68FLeYIy+P7eXxnjer90nSyagiPTtN4LuPUU
zT9/oK7ISFgcJngLNWqAc/KuUxJPkkNehXk6E6fpIqp1FbQ1fdpbEGL7Txm0TbrdlBDE50hgodec
ljTiP1nfkXu2NKpUrZ5iAwXe7EKEUiugfXk4gzwPE5XOsCgllDwwvDjtD5X78ldf9WFEU4QO89Zv
Gt5o3C24pTC9s+3AgodwPbtGhsVFsBxUbECQ9T9UjKGBdy6OPqb3rwQIimBoZ9C9ewuYk7YHAwc0
pVcL6X+fejrktlP1ApGS7RkwHPPCR97ep1veR4CdWoPeZDq91dBWPWPr+FBPlxAoeTH6jWJKTn98
GdyJY1Qu2GOA5vcpNlcym6gdfTg0zp3ooio8I2hNZD9MOoqlBcHgHXXZVipLQDKjkKdAkv6CFMLr
a0UV4nmORDATRYLXPMKoacc+zUEZw0uMP3sVvqi+Ni6OswDKu9euDY5qN5RE0iQVVXAtEcL+kSrG
uU/8VX+Z+nw7SVS72+kQUIIoNXfh53QeZm88USNXGuW8I/QaIu4j1e5axCmTi5xuokx9iT6Bn2Jf
UoTL0Qws6dHbYz5YbToy15aO0FlJgRakLWvQ/XqOzT0otdzwHWwffOrFkgFEshr9vPCxxFPrEBN7
Q3sDQcx8g++84Ewrpek/0w0azDe8q9m1Q2GjwVXEBF7KUqI3rsqhvgCtSaA80J+8O1fnVIgcBGd8
k8arZX6nUO3XxDKmtPjzJMK3l+NT4zzGtBWZcDBJceYbrwxx9VYZEWXmRSUoBjCCJTqT+X00kIM9
IkTVz6Secq/j9G+nS6sHU15tuSYbKiKj3b0kcF0iUx+5QLMlLkot26oME1z6ltRL6Dm0LX9MZQzY
wFSbTV5g5UfjUgVj3gIw9LrkgIbJScs7AH8lRXaY8LwC2D8tkKHQbSl/AfGCHZIYMr6fGVzjluh8
xyRzPZCMM8xNGM1NN14JrSqusT+zULsBFyz+g8FAfz7zmNN4MzxWWR6/sgYr1JMA05e4BhyezNuk
KLJpy9uuxaE1JmQLn95NoNDlBtCr5Z+Sori4PYWJqEkHOP7sQA92pEgEQHsW2lwB/aKlwV39Dula
LBqwBUVHr7k2w4UcJzr3k0RdwY4/nts+22o2+IUJQLEq1+IZ/k20bqLGMb5kbuo7imlyL1MJ235w
vMj8BoQaWw263H4nKzBpoJiMixS375O/hUOX5ZdRzfw32uwNg1evwZgsG9B3PlPNzcjiCzOpZrMG
lK9oyJE3U1Nn3eR+jqaQK/Gv+19oYj1w6Li92oThJ0UWq9YjnjQhn0bFSQ3nHdzyc3p158DpCQo2
thBcDRfDp63vGaqIJYj30fgThA6G+r6vZMn5zQTT9e0x88oCdKucxsrBLFWXwTZek8+Sf7GdM3Fe
gHEC51CU4CCZCCZBUM3zZxv1bgxdYPgHKblzrDZfC6fa5r0PHFhkFPQNGIYQqsLSkmEPHFKdub4U
DDOQCKxTWa2PWLdOTLkEvKg+jT9S1hwJHT9wkUkSvBJBBtBOkxhNLpOHB2gyw8joE8L+8Sif8jb4
qaJFZypIGcYWrEQBXVB6TZlJMgzGsRqFqtzJu2Ho8TMK55vO/345y1asefQrjZIi6pGOm3NWM6NF
EWiFCG+RIChE/EKxwzb4F6qYxnWzjy+JGzqzshWTMRJS5Oyg70jjJxv3+6XLbRFe01gaUBs7fcZL
lZiCJoMoQfkATs4NSftBxK6TKZTHfbtFpTm0VegWFMXgs5bQb2SRu5eoShas/3XM1Byd7pzlAmp5
e0e71koWX8Kd/3aArSX03V1RVNJ+MdOE8QgqWOzWwoZPoiRUGaHMohiozZHXlQfQRUlRpdBPLIRe
vZJbur6AQlZhYH2gMF8t9dzRz6B2UH6f3P3zgapz6p68oRYbA18LR4e7URWUongQWaOoMQUcZDfD
9Kd7FcCK47QFjsU5UwhqnrI8VTn963KDdDKQgJ6uTnJY3wXCLI3u+goY6H0IH6BjXPJNKfi2phFV
flSj8wdoitqCptsnXc0VOOcgzIwl1voC/bELRjtUhUTiY9vwWYtr+ACXX55kGfYoK3VZMY3Gue7v
9EdbunzCa8QQO7tFa7595JfBoGvW3j1bN4gPLvL+pNfB8ypM0uj+9E+vWHJdOg0thyN7G5r1wnMk
FBZs1dWGGtKBft+kPnq/g1cMI9ikBud00BHDbzsy7j7/b7bQyPBYEoSuXIjGyi8M01QbObwgryC6
LVUMOUPYLsGY5W2hDuL7abHsO9GsRDBMnj/cmILrQOnG2hjz+7T+KrJUo1nOi/YIpyjzEnkiNWG8
4ziBgrjup2GxGTmIUgWz2RaQGdRGa7t8ft5AP8gQfPhuU1eoAK199pUWspsBq3donH8IPtI4uql+
Dyq5Oic3g2VAbXN6ym2WU4tO97CKRXJWMaWG/Op3AhrQriNPcmVpAMHYowEJUDjD9wOVcsNLuU0+
nE4ta1pyA7nx8+Fwue9bmIbmtEJjoWz/ubajSW35QNPRv/H8WKS21UWXf0twCVCc0BdpwFhFSedN
4mPetqTQEjhClBAYHU2jO66aIRlrwJ0JMmQ74rpm6NF0HpRSVUhlGpIuh6CpvAh+1PpGqePFqrKM
DHmP43IgpsHh98ypx6UlRdxRAZc1vlXuABYIVrFoZmLDkWAQkcbWGNwQZ5Px4rv+GVrwVAZxZX9P
SsX+BEII48TNRPggpJc2KgPQZ33ZvxH7qxfGrHQ0nrs0rlJHd63v10wfemHYGuYcU0GNfx6B0Aar
/mLk6jHvcDE1ALyxy/6oYMf/aliAUOXR1zwYRLbNtwxiH6wyJUomUti0/xgSAgwInvu3jLr4aSdz
l2mpw/pllSn7MI9cVBEJc32TD2wlFVJd/8L+8pUilMzvDPNsmvJ4oVo1GT6xA4Lgc1lUo/IreIaA
MyUsZoK46vptSNNIKygFD81d9limrpAzoHtwhYky9zxjt8RgbTwzGWYJD8najyvV8vs0Mfam7JYi
66D9JDpebSYJuSJXiDzwya0pgqEK1O3eZyQGZOx4bwbKQnVqWB5NT9pSt8J8GMTjWLJway5QAtSO
WmKudJAiUkk104h5E0alt7PVRAt0aHUo2ie04U9VhHRMgoaADoj24Ct2yfaHZJvwE/f5NpQhmTda
hZqiuwD0BgsHBYgUNXRTvRJy+qFmi00uqR8bTFMNsM+TifjuhCafxplUxskF5EfjfptzxMiGas5y
cSHdbJkhKcvxYfyBEFx/rtf3B3gwDlIh3COz3e94R9LXt8sRpZTtGb9gtOd64MtYj/C35Pj7XVkJ
Igvq9Ej4GtkQqq9qD2cm7TndJPUBK6ae9pZNeEjMEnG3afa6Jq9lcMiC48edz36vtk42qkGG4F+9
u4LxZCc5fyJvLuNAdwCk9ua8IH7erP2ITFSiwGyBJnpVuD9beqRNyr6mSSxmVRA7TSnRv8ehV4X2
XX1Gtvtg3mTcym+uwqa8kupix8LJGpB1akwFR67ePm/4uIfxsndUxmRKpOd6Y5HeghP5Se6DLsvj
WLJfkIsvNjIzcKB4PKOeEgNxV58VwHJtCIv07U50XrnDQBU8irMaUreEsI+qhOCSXYyk044WOSxo
VNAkPZjvtpDnQxpbSJlfcGP6/IfZmeA1ZmXSBaq8rTuNV6NdwRsfSoCGJ17mp1XmfA+go3+uRIyH
u6+YXhrqX317OtjRzM0hBdPyC2uhjDA7QCQ28UFU4iTFDuC/vGGcVFnLsogyBQPvQYTK30xBTdsD
138cMjAHkQWQnDcHTs8F+KDviWFNBD17a7e2kTx8D5TYEe6vCoux1QOdtzrsHpcEDLY9rdZGsw8f
Xjvaz1qkEM0uFMRZse5MUJlv0zt+hfcbN+tmI5FiqBt/w31QgVLlBh5o/x3CFFkuxrf60n5cxEXr
POKFXHeiEhOXyXRy5nx+0EtLboBEmAd3OLH8+USx3nZj5PhAsqaqbefpFHghm70MoECJKDIyscwl
aaNa9O9FMgpTg+Q07ryrQadjC7SBoy8/vbMG8VNAyUlb2AmjOvLMRYF/JcOYWkq43ghLOe1KYKcM
0q8j1ez/WhNoMdlzEmErAouoMWkMUM/n6VIytPMEkwAYvaBw/YHchlj6Lah7lTxPVlMArPSt+z7o
Afq7hd4fPg5OlOZES3hz2LhhSfMillze5PTXJ1kA0gjNeTQIHPOkEaGVUhOGCXJlyzVcaL5ovule
Qm5SmZEHP2ODs5CzHSpEng3IS36klY0KkzIL7p2dkKs0K6yqmJrH33JqE0EhWtbljVnRqQI+Kp7e
eTT2cuMgPTIUABUwwEbEGToqG71RM6V85yrqxlCK66fzrRJGtl/mXcHVsp58FjRoTPQ/VqODHMpG
yn/zepbO6BNaI4POGFygPQflzCIeQEc2h4/WgS7c+Q6S3DBZQmRYgALLLZj0cCPysQwRFu2ZRifE
gRm3DAlC100Mk5EVxIXvTR8i5Qw9If4uSQVy7ywtmJ+p0nZv0Vi1wsw2HQqcDTDdr1A0+lzkRNa5
JAQg+GwnTs2uFft+PS6EBf21hw+RQ4EAnNa4Tl84idhjsDPBNrMCZIczKeBYStYnNFU5iyGkHtq0
cwZb3wiX2sOcTs2+bahrqJ7YJncEvwBwbw48VItV/zsRjliaSEM2K+McRaKvQKJJFACix+i70CHM
N5W5qXFu6/+LghSEvBinZ2oLvhNseWc36OBDwcJ5FdoIvLO6At+UE4qcpyvDeYeg+ewLq5rn0Qj3
sYvftpOT4R8jbxcPmaDzAHeP6cNtUmZJpP3kqGuUySwouJ14QmSvMX0tFoggRjf3kTKmstvAQAV1
+Ojt0+ubr67WzM0jQT1evNZZHk4qs8/427eUoCWmB6+arxoLtIs3BzJUb8dkaZWMl8Zj/avU6kID
jPIgiKnA4SByN+3L0CzCxyqB/N9yorpXs8H5BOO+wzkVd0AM9exvGVfpz5zVu+kWVVOR7gIxQ6qr
JP2sinWw8HoY6EthCPKRSOTpwc7hlMWyJdoOuWGv0l37DvPGp9dFB2J9EHLrFhbK5cpoGwZBtDUc
Bit3PLuF+79naYNRSg3JySE0Anr5CjeeKtLlRTOU1QspP7jeHN0XPfL9DG8DwRAJp4rv41QCGXeB
ynxe1Oy3hfsUTTZnWEFJOQJfZcCy9xtYueDmncr5tykp9o8RxWNNr+bOijMgqn8jZv6SCn4yFV0m
xQFhi+xNT+dh1u6RptVfcYZ/XlEeDb+h3xiODDTRH91cjnuZXC+vKmOPsdVjH5y471PWSNc5MpVa
C5QwBJrhQeItrWudAYVLtLGtuNxgfk0ZD2WcpKryMbzxdWKnaidgkJsVhhlWs9Y9hhlvm+s1Amjl
9oxfsIw2aw7gjr2yy/dGibLdDGwbdYEjHXwE/S7jjXPvIdDAmKRV95/9uU5obihGzKZOyn1GisT/
iGM8Wdamwbt24oohmcOPBn/zcFGIAkRm2XoZjf37jd9vFPUm/uSFfiLsc0yoDmDn7/G77TtMqxjL
oFQJUsmFS5bjvR0MXAU5LS/OZjpUdcUdZa6BxzoCftxSKaCMoDqEITGYVlfjzSPHr3GoZ6S4OXnx
TYxEVofLHKIPwYYCU99mpUr41hYwVVL6y6GKnxqrYhfcAn4b+bEOul66lBweyqCX5iv4AbNX+RFH
EgbwkryEjGM+YMNMWZ6RW4/5NcbU9xfAow8+Bh8Ahd2q7B9N8PLCZ+I9n64P1YolvH3uAMsJsaU7
jCD0lHD99S73VHsvSVWOB8iyjhvyz1azcSj88uKoqN/+PvtbI1sobKXtxPHv7CwGFozuI9KXCxey
VOjF692pJWzYjEacOEL7XVeRy9yV25iNaup/HgejDFphWnZPGs/TbNJ+yVBX2c8vMqZTVwBDmn/Q
X7Okr+zfc1coRqc65y6r1/0vJh8r/skxB/1gXR+XB6npwOi3YXlEALAKqHNu0mBrflCxVjIK2HyY
aSQpS/i0qnfqApIL4WqKxICovs5Tg1jjOczfyUKRWb1JG3xmr7KhrkX5c4AGccB9F3lq+JeIAwvY
VsxcmQNmmeUji7NrSr4gxw2qIvVUN5q/kSt5YgltewN1RyfMfJQ6j/SREilIfbQalM5llWrenrpu
UTrzB0l3w1LuxM1W9GIRh+qOt5SRsgn4eFangDIYohyPoSgQsr0ay53tqdvHBj7KXRLfGamV9NFx
VNZHg9O1Mrtt3DzEhi8YSo8ZqG8m9WJ2vbsTSBq2CooaZC384dXG9Zp6+QNq/SxDwQJ7gRu42ola
tG73RMsooOK8gTRY3tk9YKC7NTOq4rw17WwdDxbJYQtBWEJO4LHY7khgk7WAif+/7W38Wycg1TPk
AtYA/+Anlt3qstqx27A8bEwIz4Q475nuUOvA599DlwDOLixFJxKmAi07VajNllTL+v6N6eDrJEDN
aI/ym4Jw3XcV9ne6mkwFkZlKyMVwhNjSdw+37Y9Fyzw6zrnWuSZGrijLWjSGRmyPRiIo2rwMw5Yp
28l8hYP5p5nEurrp6zQlBgqloyEK5M4P0qRSOsLBPsIOYoM0D584cYp/j6e1W7B7xu21SaegY0KJ
li19YeDqwmdVYLCXjgf8VH8q/BB6Y6t14qouPJda/2oxsYk7r1BkSbVvvVkE+L0O7FDfyU8vIPpv
0t2uAsZEESjA5dDqqVHtATFVm04Y4RwFbtB4Yj7lWC4kW72ZMpaBMnMKfpElPt/6ndHTsSasuY06
WA4409nsjjVM1mHHwSitqOrdNy9R6gFcPjDujLlCqHne/psGHfOm8GIg1wPJHKDZ8/DIH08KVikb
ulSoO/C7sj7vDs/ejNqTm5crZQvlx6IKiAgKYYq+X2xV6WFz4+Z9pEUjqNERyax00ln+7ayrstgu
uqHwY5B/kSZvZYs/efulWY14K4Oxq+BTnRfccGrcwR1vdidkwRbrPr/uEMKPYyUYBb/gJ2ye5rZO
TIRTWc6FHBnQ86MIAr0i/Ggrkm4G73PgKJ2G2riE5BBkb69zJIZQ6ICG9fcNFtDlnlV4FLfCSAkH
atMsba2z8QUo2CYm6hztKgiedcB4wQrr5vMDuU9HzsQv04CxTBO1Ppq2Sio72XQy5z4dH5qGq4aM
Px1q9tLy920w7VC0RGUuXvr/gRFPQck8uFgPEiZrgbP7FqkLPcjOCtnMeEK87chcKQCH035ddTYR
VLKaMk8N2NhQc4b0GrcyNw2KWFztTTVpkH6qX8ikkvZr7YyLjJaVyLOv9c+Zs76GTJ7f1zVcQ61D
rexH81DEm+klbc0JppfoDsyuB6lqOCmNFAmgXsPMwzABO6Jp4BoPSbTfQmzbsggYm5pdBEY1wiJu
v/qC9z0v96pFg/pAs8qjyIPt+J+rUszyYARmrybDkwLmVfq7ZwxOXr/zbJBxbPh047Bu8RyJK/XV
8IXJzygjPfOu4HAiYwb0vIxLxzyud+LV8Ug0zeaov4ljJ+pYHIvDopFDo7fO++dH4j59YRF0XbPG
pIJZRQ/bGkdXQwcZyU6h2/6PueaBEaI7OZvJWvlKtPpUItasXWZd2A50ZUUfPNEyaUuIDs2v+GYa
BiFFBqMbdVYVIeozHecWofMPlk94UB1mjcgjPumcDAGAJZnby5YwKPbh3YWZ6YM81PvjKSbaSOdG
1db5qUiTIPXFj9NoBKGOoc/tbkucjSuK1rjV7b7aFNHzu09LCwhQMZ5zd8TRkOCYFS2AIKH0ENjb
k8jjQNq/XxFlsMOI75xnUerzUShunpCjjlSoBShMidayWaow42qxtDNjaxcFVVcOCUorS0etNKXh
YoJPK3phjKGlZGssD9QkMfaMxZSmgXXcR74IYv5XzTF2IB60dqf7fw+b/jv/AN2u/YVjkPeQc4zn
sMiS0Sp8m2JRnybTiCAYA5WlukU46rjqsJo3MkL7WesG0B1sqCV9UPIt68ue9wFbXqw/xoOlx+W7
eEkxhZH0f4TfQIQeenuVoPQGY5T0cEnVU+p3TJrL1yrT5Ll4tD+roOtcyUUEguzOlyrCe9eDqXAa
DLXH7O5vIABdAzffhOgFZ4cOPhERGiSw7nsJ2ITSKyTpa0FASJFK18lmvbJywENSvuPwOpTK9QFW
U9rSNY7mWSy2AghYqe2/RIrixeTxy263XBoWN0F1y00Vn6SokGoaKOKhwtYhMdjc43HdGHaX9y7n
dP1iSAzd9JQKYOIDXrhPRPfflE3Bb8r927v06xRuE3K4JNWM1OSX+p8LEc9rgi4k9O1TZxoPM+sd
BS2vlHfyLUGkmiWV6wLLS6jjxJxzB1f1equV8oQEz3Vhmyc6KUQ4sgiIwSYJTIFEmX87wF6wPx9x
2sVSDM+zz6vBess7GUsE4oD7n0qpNNo7RMxFZcOnCm7BK5PZlrSOun5/DY/cemDQwYlGd6HQBvrm
dJR4ppypMc+YBIPAQHPWS0vMak7rIVqZNiplq160iMnrSY6/5fSaDQQqWc8Bee9qgBh43FiM71d+
YqLPJkRVxgR7KhgSg/oiemnqLrD4Vf7JEvLA1ji4KsMRic8Sa4+8zjQo2THLfgP3VbsA7IwIBe10
uVJYylfWCXSnKVsclrKBPJAYaEhLafOXhPRk63F2HnTjkICnv5hnGqZLSOk8n4OXjKKrGmkNKtqb
+bDWVwTigNrmim/8/CPqPvOClz9UE+YY4i7AB2/ogS2kY2jlELvvSr5g7jovvkFQn2NZ6IADiV0A
BRjl/ubLDQbpb5hmq+CYl24s/sVn7l1mssfHcEG93yr9l/sAR82MV5mcvRvGP1io7QW77HWXq0ud
kE716oRAKDUbi8jj8wU4JU0jXJ9axdZoefX475jIXsJY5dvjwZOGSntcyQ01gtCEKTqWf5H3ukdw
NYEM1vtsdrF7X37Qk2b5jqRQnotOyH/MIOJj0qSlhpvZytnIr94HjxdH3ORXeLBkcOYKkQA8Rom+
2FlndprDzfHkiiSq5eVLsMTlCtlIkZca5kO6Tbt2lHNx4nSkw3+138OfW78DlSDFaJkOhTRBVfYz
d20AzT/HGcjgtpjnZzEnaLlV6upQlsWjT6g6vX5MYvr/GWOmsmJGeesslpOHjPRn+jmSlP0VZ4M4
fOw7XIL6OPmdqcwsbRMDrsIDlQJDhEKF7WiTQ5pzzkrNSVlXwrkibEVytZXuErfiwq7xQqZcH0vN
dE3meUK8l4yx8mCJrLRYsqdtgFs9tPNVOqp8JnN6DFJObnxzoTtemRdiRmwO7NQpJVJAtPPv85P2
9KLZB7AY9htieIHY9laIaMDaZK2A8C6xiy8g+iCyeB+6yYy/GGrtCMEwOT9meEJn+TA9ONJZlf71
yfFS782MoD6s0e9kclG24GZwG6RdRNKbXwZZwb+rg4WbfmIB9eqKPjAdYm9kIoBSx+cK4gp/DhDz
Zj3myYel2ddYOcO/Sn69DvIJAO2/fF3DgD2GBaNjlJ7SOxztDm6lOYTqU6S0xAqZrfYIrEQ63B7q
fP61PesfN/FoSXJYXLYAS50viyBzOpATY3IN0mU/ugOVOLoojT9EMOUjEmOdJPUdKYp4oKR9ER85
cHEp5SbwEhdRPfGRBo/v0cDLN7PFfXFE3mk/Fu5/ZWcJt36Lw36xPMcyQHlyh6Xs/dJBWKcnANSf
A/EypY2rOh+E3n3eeVdFbcgZEYGUkFjEMH8lR8WHRL/V3TPrXdtNquRk+cy/8uWhCSYjy97UlAxj
KkAO/LG5CjeurD58uezTkG218OHwVvQxhnrYanLUf1qGl3LrYgLfKH4ZTOG0hmNJO/4boKRwhgRx
DNMHraOsQ5261kcuZlrSPX26knZdZvKdh1cn83Yx64f+kIah+0HiR+5MGaqO+sHmANIKbuZIiaDm
s7Qtwx1pHlxrYRZjaHWhHyBbfVHfauNrxUalZSaK3OuP/txD/0vm9Srhl2fVFKQauPf2u3bBdobe
kAo+HXzoaeQYunzzIuT49xsOkK9UOkar2Uqjj30xfWeuDqI7U/TwZyH4RGzX2YBlBH8ZZYItnYaG
wta9ofQLnJ9Lbi+0Uv9cL7nZfNnNIgFzop6XQNtAqRTOhj5koyzdEFWGAent72aYaLFI0F2AXq0b
2Twl9SwEySdVB2mktkZSNSv13lrtoAGo5WrqFLSnlK3/Z174x77eRCB8oCYwk5c8FhgyKAPABTOw
AMQjkf+SBmhzIBJwXOJHEoDlRMmi52QABMZZ3F7ACr+wdCFKQ2CHk556Ipq7hbt6vCOVvZzwhGg/
GCdlgrEsGcwa1unNlCAaGuvgAVFfHL4NNdrB0e7iHRZHte6YTi8QSSTYFrGB2NOHx7b5hMYiPdxf
YDE9XNAHptYfAucWW86wzp/OYsUuSOzJmL6sohv23+3p7PEYU1qUgyriSUI664Cj1p6nazEveGco
+elF5kKgfpSK98Yij1DCJcMDWrr/dQi2GghpiR5R/vg9V3wAkWAKMmP3wLeqh5WbB47JVW/PWoa8
YLkEL9Yf4ho1Iy8LzDYNwS/Ymq0wzfl7cVRkruO3FrF00o4msfQGVkyop7s9fuc+Ux7hDEU5VTgL
RGGtxl92xOAWJ2B5W3wD/sCJ8J3wbm7LRngKlKKsGFf4KqSGPDT1oTuykf4JzoL1ih3wSrSUAztX
oYCiBeLXZNARnN/LYo1xwGtVSXCxv0gmfPBVmv7+hNhG5evLQoCcvR5aH17yuJ+IAff7er0u5EFj
B0ID6r7MQ7GAnyXosQzGpQZuaKvn8KMVBfgHJONI2AJzDQsb3tXXPfDqgth8wD0EVH/nXTYuP9H6
PFPdXBd/PJyMnwTKZRica2O9YKC1Ba2xcdG6CBqD2EoNLkGYD3o/YXJONNHoeK+FD9wuPx/PG6XH
CxPFPyaCRYe1px439RrrqOXnQlebuIR/G6m0FQbLDnjIkUb3HtdXeZDVLIa48cERqQQ/h9jtVd+w
7v/PY3MkoK6ZgDCynBy14BFkSRiWfp65y5YKX7MQOEA/8LN+ILZrrmxeNMbhtXpg9Vx80MtP1Ojy
S3qIE62Nb2PTAcRdaR0gfvhGloX3EZkaN837CnT0x7Ts0okoWKbZENn8JDXTdtp4P+0Lmfhzf/0k
Fot6dmqDOqxTkGKcfRtx43ICPBFimTnY3mp2FflHAw+WeRRPUF4gZxdkEn4f7M4h38xcQEOND+VC
2S81okV/7IQhYrgqYpt4MUxXTOJn9ys2DzJLypxwqpG5tLeLYUfLOdmOvwC6o2ZY9mInTh7A8Z6/
5X+wl5/ZVHq6kH/8fpCq9DcvFJqaVPEvu0e/ufb1rQWxApVTVJRk+Ld2OAf5qdSQ4lL61YAnWJLr
qTYpnMJnVXoR4i6CiqLXA36rZobmuLVLexm+FN9hFaQJhuCC44+PAQgsU0dXvcF3NCK6ogtoD6QK
e//dzBSWvaLDJ3kIFV77rj8gke+34Y+M6k5Xr7UWgLZ+fkZ0zdSZRKFcuIsotJnDnleXv6ArVxRm
M+kHg6W+5K8iMBLBiaJmYatp99d1d0UecJpl9c6X+2gi1G8kr2VjBiEYlmOU6BUjklAHem9tv1OG
j/jPTsXLQSqSKKzS/ZA7KcELcFtmWseHBNU2d8BsK2WHmkqKLhFT8fJ9IiucxaVa2l2ntfbkbBay
yLun9+U+aUN9W44oWhk1+LDx9xdrxaCiT0OQnYosuIp+kvm2EauWJs3/5MMJivViBi+ymGPcwib8
ltAsI2Of/rTLSXznymmQ3Us3kubzSLIOO9ybQokdRg49A5XqczbAt3bOMiVJOEE6iU8RLppQ1jem
tUDcrc00GK2OFPIb+Q7hCk3wPIT8lO4TDmfF/QlqVpIj6p/INqutG8qtSo4YOWQoLT+EVINMtGwR
JZNvyR/NZOinHTW4VeqdfzZlMHd6J0nvZuoBpFc4tTN1MpADlubvfiS5QmHuoMQU7sSVhlD14DM/
iIvWeRvIh8RxJKG+lkKD/UJ96TJyjw6U2j7BwbE4+0MQxlWmSg8ba8FVQF89pjoNsRsj/uJshVZT
76m/WY0jyObYRL9gbAeCWFOCoe6tJO3fGqxGKkIH3E3Dngrxtu5ikjZwjIFLm9FwBoVZagKpJkbN
JDWp2bznsBaCIJm1syJAOBINxZ/PCT3rWSmVTKSABilKrt+7x1RAWwdkZDsL0yKaNDMNxGrnJswR
Ort4s5/p9kBbnJ68MaSx4slog5Gk5aySw9EDTVkrPRnyQiuLwCQtgo01bv4eoDtyDt5pLqHimbdu
bPsNf3NV/1oGHz1GX2ALp0LDAE3bG6uTCaep+YVDyYT5RPO8NABjzufL/KnxfMWsgE7VB1fhloDJ
XFYOFYskCJ30ta3EurdyQyzo30ZsL4xYSzdpELhp5OtGUAfSWLmZv8/e52q/Yq6qB/DoBOgEdjFx
yghWpd/kzvLfkKjolSwM53TqcyzGdrPuVLIe0YEr7cdksBLw08Z6vi2TWwf4qsnaNrvKBbtFdA+s
6o5XJ9tVgCrAUQO4x+J+V29PeEftIakYgvRqgyjlSvRehJX41b4j9XyH+w0NmR1dMNeUYxa2kV27
eTFYRYHMe4nMrQOGGazoVWrCwZJVvlkFMWM5o0kLQl9RZw/zwgFUy0aOROxj0d+7z71npdl++p/F
TcUssvWy4Y9xdh4SuunjSLrlYyYNlDyYwLVEZTyeRA3HobU5XAVsvtWhm2yE03NmHnTwTc7lLWS8
aG0Zz0GzrMZDOJWcAIvEJxSQrcy1mkET7tXDbfn5Py5VOvofOJsjrLVYQbuJ0oYeXjUjKOYx3ZCr
JqQocFI5D6AmWyYbfyyam4EGihCpXrkMxjcfYpu3XAaedhpRr8OIYGhO+uCp8BmqXa9QrGvPoFZ1
EUymx8pfXZqe89ifCJnbX+SITBdC51ZTGJRmLaaG/EwtAkma+uFt8sJvleK6s8LhAtyLRqioarz7
xzWsErhvXIgqg2dQReO107G5IrUfymx60NnXMAvB8If+fNgCDz9lm5I03ABrh61cfBWumJ8HkbWB
UrGIvQmYj4Ma2H0PepXKmtnzcDxlTPE9gIYi/Zbzgom5nNUdcUvYAQgPN5Ln56FokYOPm/rBmPo9
7dO1oGjYNKEJ4Wyjtb+6lYj+MFr4dzYRHBDSZqoBFdWC26YyohqE4XzLmUKRgHMPZFW+CDyiNfyT
iFApOg/Xm1SNLhQ6Zt9p5Y3Lwgdv3eDAy1iMvK0mWSbRHJ1eQ5RdWoaepg2Uj3TRiGPtajDlwlAU
rbBWNwVpkJfEid1Eb7VMsM2T9JnmdJ3uuCZLrR1bTnNeObWw7VDNVjo1oC/38EYl2ixbYLtzWmoh
XOttv5Z1pr0dNedLcQXKByZZJabjMhIF6IYPYeKSY3IJ7UaG0ABexjnT+PV00YR7PyiRmUaJpUW2
uLuDEhC/j0ZdQmItMlx2F7H/Ds1BV5+zIWzHTPJaFpeSpp6rHny+Smfix1TGvdHRNGviTgsUsnUP
QCYeQoiXuXcxsQzgIjtmI/SeaxZ9kymTkjPoWCAspHkGdB/biP/EPBt4kEoBxS++mRYQU0q864VK
R/QdzAGBm9vBmVZPEmri56HS1uXWC6HPF+I4G8RwrYlUoaIwcJGhi5I3NQclc4toE5eiNLdBQIqP
cCuUmRhXfhcmtyKQk18fnAOTXjJ9WujCaiEH6BTTHHoZFAi/Bg4jRRMwjYejFptEg1CquILiDFbN
0MBjls5BepnZvaHOj3IER+DSZ94L3zGG3JO7b/udd3tRKTl5p2nLMizOsAZYybNj1Xxuw4VIulhB
/wZigPeX0K8pKuAbBI85QhT4nwUC6rWV14nfqwaq2BzkjBpv0E6e3uDM6RRSqCswHmkGEAkMQig+
fBOxL3CJkMBsGkbYRfd298p3IAwz1ok1SHLOZRRlAv8lfcKMEr4xc6JzU9K+kVVK3xwXCGKx4JL1
CyRgpJvteL6G/JZXPhzD4ZuCnRpjOBAyX7K6lZsMoc/jktj7CYLXyNvB4N4fKAiQXEiqKs3QwTRo
72muDGmgo5evLTqNHxHfphzXBDWWgbp2TZvoOxa7YRj1Zrwr4bXwlVW0i2H3jAAbofQ3uTjDh7Nf
cHc1ON0HARXXRiq7j8ozdvfZvtoIqvfP/LIWZO5014VJtGw8v5D1SNNFB6trQKnxsFQJMn8fvkki
Cyuk1R2qcJmiZcqZJgK779tctrzynX/XCxleMjXa6LqcUnSs/R8oPN1MptmsndTlvoZVSoZerFDT
42IgZu4rXlbogsCxKM87gyMzsuc90+E6EqYLhpbWzJ9QhcPAv6WAYCYThB2BCCjFa9wazCZEqo5h
XcC71nlSE6Nn2K+/wszVI9eeF08Iri8WEZ9qIcmvsLjWUdzQPAeLKYx48zrtIwbU1lnS4UHArJAL
wmWdt0rzOMal2ILvnzX7pPcrfYrQB/yHLFYf8XoeUNSRcjS0gV6CbzREfeA5RJXMaAsmqlzZor/x
dFlAeuEXr/xlPMkMOlUiljpEm374ijZsn1TdQtnH/68Swywj4tiYNp7r3njjWtq8Pr2qh7cGKHVD
b8DhA4WXDAR4+3ShQ8l2Ne2GZUIuCC/j5x0wBeePFDmFOQKaeLTv68eLeC9moUXdPMz0qMTDIeVM
4Jl/tmT6NoPiIUPcJK4874QPxAdwt07M+XlVL5b1Xmv3exI7HDUENg4mxHwxrJwq37gJ/mAQxGjn
ymjb6FfvbWig1vkkCoOYvyH5lMHgWWIRLbZyahKmeaO2z/tFn5Qlk2uvXIynkt0PUiGoLUJbhhXI
L18Kb1uYe6kK9PMIAVS5hl1mRqz9zPanCqnhqndzmXqkqK8u619yTWEf67vxY4VLRGk4wXw9pBGz
QiWSXuYlH+u2bKWZU3YmPvLGyU6kcmoajRGdHVgMQOO+DbWa5dSW86dnzdwffoi1t2uIAFc9dRh/
8H65FrfeBjGd4zrIVlAJg7gRvKsiDFd/u0yaF3oJjS5P0BjGRH6jF3m+HoLdl7qjKt98DwAVmTc0
51ozCvA2/ziYw7sz2C9F3Y8vfP88YAaO636LSR1iGeClLB6xQOQONx/eyhG66Q76MW/jGw+pKqVh
sknpSg4xVuBbB2W69CLFSWIQ+0rH9/zhmNo1efUff+zn/MbTV/p2SLZ/bN6K3g1BNTrPHpkdBRGV
cnkOU0FYiabcYeXzw4ZySgSl6C1OeQzVLeDghugB98lcdGfK3heWqUbGOKDFUviZBNi1pzWC2fo5
jCaS+zH+2orY8FZBJD2sed9LilIWfVN3FcLTtYsOp9HQ7ouGbkA0/A1qUXeh2QnpagXenlXcqP3X
zsRNj40MmfpSuxoHHLJ3K+CzuzFWzpFAoxonUzVssPTvb6vucbWrt0aYzVGlrrg33gOKxsZCQvSS
ijOnqdVnLNGlAxWNx2MDW+aUx6/f5r1jrPALg3SOGMAPlA6GlfalSCCI0mSFAgDFguP5SAXNd9nB
HwZTV6f0iaISdNMSfKgw/Z/WAJ1C1woeC2awttT8v1voRXwvAxY1bhMy8xabmjCNojVoyU7L5+DY
Ibh8G6gH09En7IV3nTR3q6Z0ZvvXytCTCby/LP+K+HqIGJ2jYEr1TViu7y5cXAHo1JWQ1W77OOmd
IXA6frrZqma+Yy9til2LKu79ks9xQ7agE0XDXQVNEmna8zhuX+KhBAzWKpdjkDGQj7CDJIdtfO45
2B/1BJE95HbUefGVL+VDDjS+rQxhRTF8HBOagVg47J+csJJ37XYlZnQUZIE4fwz3hA0upFPrj/ai
VgkSYa75KYG+1Y5Bk5ZlRuv9NoKybecBsTCRw0ndNY9wxs8v9UDZRbryKPwnZXCl2uH72UG2+Mvi
SqlaqM7Ci2HiOPYOcOeRE0CgW/rRlNLkPIZWsnsnyPz32GDjAvar05ES+ZZ0jcejlTmkbmQeD/Hz
gICq1eK/0uYUaAEMmn0jNJy85cCJ+5ioPitod8UeyhvVFm+Vy07XxhSuXeh4UhgYi9/tRDFL89XK
trcqzeLaAYjb2Nop7lSopSig4b4guZUom/wbBJrHhZscLrtU19KbnkaG4RmUXhg96axU9+8jvm9o
DoBxdfcPjJ5DqFn25wY+00dsgmvAZX4zfApg/0RZ5N2A3UFth4cqn7sIxmb2T9i1OXi+NzzK44oG
9pTt+mJZlACgJBS9cdikIgQT7yndbcOOC064uyRYDULIGTDG5Efxpiu2zd3S5tlJpotnNPYPEz3P
j+Ez1fIZOVQlrblo6wVc98WyZNnXhL1gJqzvKgKR82vCXQHw1Mlmc+8hkeSIgYCh/0QOO1wYTWlB
k+HAuok/sBUfVik3TUIrSMp9b1f10vPZQDbP111P2Bw56P/jFEF5nQaukxNhIndzBYh/+/NpliZd
S5kgzentrFhOym9XjM46M7OBfxHspVtH8iwkASRt+ds8Apnkk2fMMztHWRwc5lVQoXyA6KB+28Hg
9R6dFo/vCV5NYziAnun+Y3fyEyUgpoh7FAwjMv4q4jyJcX2T6mbT/DGlua+fkBFlprEiRaw23z3S
71X95BG4L5YoXAYAzJ80YH7HiPWcXHYTfBe1a82f4yngyUGvDllF+Lk0Q8NsLsLVrX9n5ijlQalC
hz/m9g6th+wxVvtcjAiLPpRE5rSa3yRAhDR01soQtD5o1iSi0QeS1GTuQmsiYy3aKLXS4dXrcqHN
0p1uHldxxVHg5p+ux2ShUs04A7RxMMTc8QcNT6X4lJZ8Ik4pj7vT5biKFQ9Lf9063YbFmgFtdWM/
yOD/LGM/GKtQaKpx61k3V7SIjp8pcaq+AVmGeJUWZHj78VDqTgVkdxCfnJXdP0qRDHOOSwrWwUFH
Xc9522/7x9dYzL7k4oR+qbNz5N+0PVQerT1A09Y6YduQHJ4HFyCO1+WGsqEDGP0g11j5mweXmmoq
LeljmaroszKTKFx8R60m+wDToVvWxZwtucVDTCg6okMC5jAQGhxy9ytiUltGyxwl0JGCbPhfEHng
hjgn586o7+jj2q4NR+1+0qxC0/zkKlmaGEuNQwTjXMIykWoDJK5GgpZxMzcQ44dFQZsu0pRekwQQ
6aqMTr3WounRFmGlbhZwF5M9lvuf6n34hDnalsXhX4OnLApTZ0Uds7P0Vguk69gZeo8NAyyiV4Vm
KXuqrv7JHrVOB3N+WMtRs02kWFjMZ4Otw0Q2XufZIoHS2Ein839iU7auQl8LbZ6OKxpG7wTUVvYJ
arG3cC/SwdVY756fbKtMlrg/L+nQ+TjWc8aICyHm5Hdc1hS7JYo9wUwFFKQqksvfi10n1T8HUNmw
jNVhN+AUKzezgz7LdTJPTGlzfZlONpUCDqA5z27OGGLyjO4WtEA0xzFB0yHI52w/erg9Y/DZA9jb
PpX6HioK7qvNelixWY/oDkPaZ+RHsWYXWGHh/zAKqrBR/1NyqYssD7cLAEz759pB80u1M5umeILW
9tx44fvy3ZFWFiGctnt/HelRaE9N0JC753/QQB6gWxT5Ud55JxnZBN5Pq7m+lzkW7E9zQ31hpAP0
5/kqVKPumu7iQsINJm/S1lTo4OFouT88z65/9+6SJ8fz0MD97PK1lnKXfTfBmVu0ue6lzG1V9lYb
1QLxEWercVNj5qHOGwW4sel58QJXqKKnw/ruxJPBuPiluUfAyHbMIbzNhgk5Vo4uwD9mu6TKABRt
7AyH5rQzspA3UKVO3Sgk0Sn+ivPnMZLEJ0SgxTlYf1Bekt+E916zUUs1vxryo0cKrclIlA4lMsSR
PF5ruysP5ogf9ZD/eWqGxbTeAGDiMOEQx+c68cfj5SLC85UevcwLaWtgURvmcSp4RbM0zPL2KpMW
PSV7cg5FeyxFl/RrSepaBQwMfx68BfGufPIfuS53vcrMxDPoehddIVGlhVeHHzgGSKTt3uj1GmfR
lKPhCwYz6ogTNq0IThe5pZUUGgAflaMekXhMDSl6Pwm+RQm2HH/MYI1IjE54UJ6l/56aDKX4nyAE
cwhdsWnIapdwqmVq14lOTocsCS3eXtn9R36yKTaWlBCEfpugtLIJVw5udJG/9Hr+Ujwt9pKtYLHt
lPsYS444FzZO+RU2zl9O/OwmDlDdFejhdzJ1bMtTnifwM2k6t1HgMO90PYfTg8uyolW2PUgW+IQ4
2a9pO0fm4j3V3i1PHvB39v8nIclfGNQUz0chVASzZjp3x7jFF54HPeWMuUW+QYpvIXascg+9/kZw
KeGnEzg7yN336nzh9rPiTctNAzsGvpPHwmDTlcUu4DGfFloIuBLO2/a3WpZNuaU70IHjPdgrfAwI
5WgjS9VRTy1rKZCjKlWE+npOrlFKgcCBOoCcq2Xe42Hsy8QaCaTlfNRNgcOkScBaTRLp42bzmHf+
vwUxpK2vPUiT1MNEWkauis/8iklXIhCWmXcCVoV4qLclt4XfCZ0xWopGXljekBubLozBT+b+HzpU
/IIf0hZY0dnqsbYj53l9+E6rnxJqBBNeKgCDT9/2I/Vn8s7ykyLKgy7fq9xZWuI82v4CT70DY0lh
5jj94OFHW+YcdofVSCgSefKLBQBMUOJdvYOhmvjxfaYUsBpYHinsmoPL8LUhGwd6tDKv3VSBx1S9
97ADzEBmZgsxxqrKOvRa7Dn3uSx8XFMteU947kpPCMLR7z4TPeoEKaEryvIPzAtEHVhCPYgZDMYO
ZCvC/PNCGRwe0N/um10JJDNSUGpI8tHLs5Ijet3RzyliW5luTi7X2tso8vlW5cxPe4/6zaJXCgEN
cdiWCMvJHoBEqe5dPy1lAE22cyGCjgvSIwtGoZUcSi/4B9jSkLXZk0vTsuxRfApqDtuZRkWcbxTx
a89QRTIY3+udL8w04cScf0Q1iHqr/jXYcIw4SHEhZ/DyanpDfSLJYs71B1VRErnJQmRsbNP9oqVJ
r/1OPcW6fshs+CmVC7YkV5N4OlDGO6tennrbuRESwgqC4Ijh+FbkEHe42g+hABAaTShpUwMr/Jsw
m0ufmhnl/IfBXqjn5RuiY03qf3LNTxFHnTqjW8s4Y6x0vVgX2UYUiIFrE1FkFms+yWbD66JjkbGO
XEIZsRljAWu4aXOG27s/HaAvrHnfsTQfOFr3KQSxHo2NKTh1bYQ7GJtn9QGHXU+wbsFvQi0xK8b6
3g2WeKg33BVfyPLwFw7t7vPgf9ZxGKi1+ZEGmRTfnKrdKj08LeLrpA8BoYsrzFXMs3Q8LNpC7BV3
mSM4ko12svPALJMbjedfK5rvzDerpol8C0xYw6JY8g4gEtGxa6Stzrb4ZbVwuqIN9NYGuTnAGaWQ
Ry3Kq5X8weaTElAzZ1TSTh1Wy3qvxBvti9vFTRl73/jmPh4oP5lWPdJFT8p4tZbkOlXux1KZiLGf
2y6hikq/m17imzo6wumaMv9GumI8PpLPsn02STWYQjbmDORlNLYe1HfmAadfLaU8i5/TuMJ3XtA7
DZu8uUKuuIX/mEZmcfe7gkDl35MhWFWXwaoKOfSiAt6J1Nyi+wd614vKJLrAAgmavNNP2HOqF3At
TVy0b6JuqNiRvGvLeYZB5Hgs97AoCq+o0AeEdv2k7qfS5auTJPD28ahbofe4YFKwJiGtiv/bXiS6
W1q/POg2WJidcpFqn23nlJjkgC7SIkIcd2dPNPNWsDcyx3bH3N2EB35fYu6yA9/zY4IJERCHf3wp
oGjabTzXbGrSB+SGXGopmXiGxr6+zFPUEUTNu5k8uDyt5Eao0vkoRK+ccgcFT3dbNFcs0RY+8n/a
A5JS49S4dqB3edMvDU6r2QuK3EZZdEEayOpg6YQZMF04oPnATEtUqjTBikg8R3lx+OcQZS5IefkH
q+atyThNruQ6gz21d3wzqWq3t6hubnZxLSwP41D45gWCe4I99WuLefsyItalH7BG4B4Hp+1OEf0K
r1HDFFd9/SuUPNAD355g1Jh/OTh2BH8mMzluMoF8ceQhBd8CdmoiZG2spqsKHsq9tlNx0/TxlqNw
mCdxo4i0Kbr3bxTeJDv73qBz7e7aH7CzBrbXLaE391ymrRkPM6QzTLOKys7T2pnTRU278eZiBEXR
0u3MMbVC6r24dHzmGp624YSRDBSdKxPtuIJ1yJjglNYzYMGcJX41sFEi/CqP+C6SvBRJxZYW5Pkk
IW3KN9Bbfsjj17tuzliDQZVOWsQI3y/Ai7GtAxpcQegc6d8Z9jCtXB83RGkInfZf3B+WDMY+FIXR
lvtt35WMM9DQK1xm0oQK8ziXq2FqKrXxRXZC1vjZCLLNbGcq6meC9ZBc+sjuNj34pSNYkO/hXB6G
fXPQNHTeTEl+OjIYTTV69doT7jt4TNaj33cHzJ0zll6U2aATrDkNqTAINYalyvHViUEN5sGf5vHQ
u2yKcGUKrsW0YDcjQy6g9XaUata85MB//nWVhekkuEiVFME/dL6WItw/XO0JAOgTrkpb1VlofERg
egNQXtfXkudONZUCLatTiLbM11X0FbCkIr4R33v9vSRPfhpI2P4h36HjRdEboKNX9mbNqOrVGd89
w+W/aBuoRfo+TfuT1pe9ogBx6T2iOlOpkXwZv24BQghZMBwQCwB3CE1ZYVkwID8pIJkQqURK+0eH
0z7yzubCHrBDOmex85cQuCGx/daWgu3kadjr2gpIJiUVGyTYwntn1fSPv2JzZ2ehfhYeBtYHW+Qs
2RcQfZsT+0ITJPiTipnAhXSkRM0jHVxX5MigBBM9jWve21RTcsocFCR3Csm9fYxCTKvjLBQ/dL69
YBMTkT5p4TV9tH2w3AhUp6gsHeKYUbZ9/0SRxBFDMz1oABKy5YYdi8nxw2+hb6iJlYzVMaOOgQo2
FS8Qp4qFeEQuDZZdPIlqmqpj6FHiKeug9xza6GxVnrqelyyvDaaFSRJIXgiAcDi3Psc9p7kW3LVs
dgOY3ECGowgodVpJTQVtNWS95rqmzYPU0vA9fT/rCfzIB1ASR/cgxpIQ0O1fl+Gc2l+DwPfPtnuR
oZACSF+HEoE8TfTlIQ5Uuqa9SZTn3Ywr4ZGkzGVS2HL/dWEIrDKUNpX8Hr+1idGY+ULj8eS399oZ
YWI5D7Fs43MHUgurXzJ/aCyrRuNVl8IovHyCeSevzR9XBv1cScVKixO8+XiPpf+wI3at8h/Se8sa
l6IfCyeYDTefyNxWKqnppX/21pE1w1TzXzZaImBBs985vMywFwhrlJJZ5QblsPcPFOeoZM6n5rut
+C3PYL3I88NA1sqXkbrNoyG40NeDKZl7WBJbcJ1nXRVC+2yGQ8Rswr9tACXufc/4PHVeO8BwLeOU
YD7GDFZBfYeWKka9YhdbQMpdvQsXioqPKtGoanu81OrpRvHkKSpsmjxAd6t36vX+m1CmanNR3/PV
OsnFi32FUfdF3OXCsXSSp9YfXLaZYGZ/EslD59+fCYEGgTXk7nPImc70+kUe0Cd56mgOB62iqH+v
rKfVhRfaK+EdFpguhenU54//oJDggvb2ZemsXnuSgso6MuOmf6vm90BsR98ShoHKF6jgu76rAm3l
KMljo0hBmY97dnFfE2e2YRSQfa12TYdYfDt5OhBLk2pcWc7ioRthGQVogAY/K9lbh1ppZd/cQQmo
5KV/BuNjyt6kDrYA4RTBK+YsDAu87+F8MZMOYiZyL1Ugvg7H7Nhxh15s26YLJw6gDRURH00Qq2w4
fnFTPZnB1iKHLtJN7j4eIKZxxTm4UPEW6SQZkN4P1eHVQaAB2tUGhfP/Eez7thrwiAC1cWhwvJTg
OQVr9FB2C2c5XuQ6PWTCZSuzmMP2JjzmW/aBi7G7hTZaWjkRUqIMk6ZW1CgtOfK6E5i224+Ymv1i
/0kCjd6ILf/7sC+B1u4AdFCbvFl8t7KkES6SEuPeZ6SDgx6zlXBC+cFvoW0fTq+3ifPKMnkwqNe0
H7R20twtewAqxgt80EEQg4s8SeMo8rUDAXlyqQ+ZqCaClQGKlH63Az7UdjbYISUEXh8vhE7XAWhJ
4t2N9dMsEaM+CWljs72jjUKpBrVicYwvDrkSzXWiX7rZbfrUy8vhysarOcLnRpZuIvhowxWiwwkZ
cZBMnkNRTh3cyKCvto8t/1rI8pTyDnl4mToWoJGawYJz9oKWWu/mmP1LTAILVL5t5JrU306zX7FU
fhDI1+itekbjdQ4EwV+zEsmhUn9gipqPX9woLOUnew3T6f8RbDCkxBtQR7qVeHPGWPe8LpBc1YYO
U7ol6KavYdNUVIj/NBa8p+hsCq5ynqurYfyZdGBzSKwhDio8oLTAj48hFiRjPHxuMIrmvwLL+Qhq
TPu14GyYpez45Ku5lO7GW4SSAqBjsb3w+cd7SZqK/Xu6I2si4Shcokm49FkrQjtmT7WygIGmpqIN
2kM0iKE+wEPQ1bcHZwScQnfVXheN7oZS4PLEX08cFxIdICYXf59NOsooBOZbs3GrXZYWbM8+vdb5
EA30eVZc8NbgfG5b5YQjxliT0TmU3lRA9seces8S5l+M2GeB+gDP7Se8Fn618dSpdh8iw9XCwcJ/
ib5zvx9bR92B47sP9rtyJ4NCxBTYuNfhH72tS/+rj+4u/LXSxxB4U3QgUoJNLHHustF1vKkWzeGS
CRhd75xobf0dTxNHz0RcwhGi4j9ROEkZHuMO6lb3Df8lR1zPYwQS8ySUxhC291LLqAqty6n0JmXH
qt+rt1O1qg7/xPsNBJ73J9jR+wIrWqRpQx0XameElPPWmDrVBOWcT6iUTYL3CFHGdTud5sHZencS
bzwycE6OjpkcAegbHZDCqbvf2ByvWfpyakOKU0GrB6ctWhU/hIYNjHSscIeYbnyvV+vrN9XEmokP
iFUWEYX6xu/nqU7pY5+LE66POwnJTTQIpDEmwD3Ra+bnAN0feOYAsG4gxpemC+WwYpDfIJwPiU5/
NxxeeOLCFxvD9Hon3ArqZBdWbgKwvUccfgp/6HDvkayYqF6JZ8bB4Wuqwm0qGH2YS0n/P5I4vYA6
4Hk4TLJUVkyjf8sSNGDZ+xHzVTdFkbGw06hZ6dTnkLUImBs8QmZbZ2IPtagX+nBK6FcjvdjyGHAv
q2/tvqsbC3UhtIjyywHCvDb0vy3xeRzkJqXnM9K0Tjji+cSyYUawo9TW+IN2zoQjoMe6xvUPf8ky
hSncL+lwkXLEMYGraTvw5rRuwM5N3Uha6vUIr0S1eqGh6yyDopXdtxsUvLLxjyfB23Bsmv1knw8+
BA9ExCBlXXQFkW9XSdqKwJiRWN0aMycK9IseRXqH/yj+12u+PiQkGHSTRVhKLSoUfR2JNrAZzPzA
zyuzgGtsP4SuDur08j0Dfp5jIIR6hyexRLvEiPaIpYer7ISHNkodH8r0Wqm7H7chX0tEfZZE02je
UWbqZwBOkkuFjxFDSDPr9HuO15VpBAUKU5aoQWkV0ZPsiNJU9c9FGSJXUZMDK7nONAnJt0EuVEIY
88EvxQdZIbjgR1mdCqmgPCdEaxG7Xb/hwK5UO1juEUhVKxBMltQW9dJSTCnNH6QPHcdQGwoBrl7U
6gG36zGRPqEliy0Cy3BM7HgUQ3KQM8zxdqV1FkZXRhdRVyAuCYTtba4DfryF7d2W2tgjiTHYWKhn
rG+GOb7HdFT1Ob8avYA6wI5gDOOh2yaNuf34wQ09YNmiXYx5YGafBUjpHIqW0EtyUTaz0UjHLs+n
le+iri5d/stQZIFGdsU3j3GEIPDyQo0FBzj3QRKp4VENcFvCuOdWz+Ij4Hhh2dWXamY1ahlQSFIM
youB3GN2IltiICjDVCRhOf10nDizhLdfh4edkDLmTWsvo+CECNLAKKgSSvTIgQtBPTo/tKsKxN0Y
lv/yQGpPGi8nmTaolfm8/gjzb+nhkOyd7KBjUQQTYp5YaarP+e6yvgOd/qPhttgJzngezDpo7ZQ+
Wewr7evcZQ87eippLE6c6MFzqiNaKQ12JorOySehVC66DbY6NJYRJlzgBDXBb3Zetghn/H5C3bQ/
7NucosC+XTZbhqT4RJvIziZNI0qD1AG+IdNpKmQVX+u5HuN7c/6q9RCUpwknXaEPsiQPKf3Vxu9N
AKK4ak05PVeyrzS+11UY+wlxOOK5Up67lhyCBKe2nfoJMGUvFmTQPIjYsMii3+oYkoHcrtyOHhJh
CJPzm3orRWvZ/WI3V7w1JcXo9MY/F+b+2bVlB0RwMvPXfmrXtWLfm4Y30/gBF0pzvtJGL+MaV2B8
vjOl6MVAGcWIJKnrqzTrjubgl2lnq4bIhQNggks0+BFubXrzpO+AN/AQla3rd01GyadG/sG8ifPE
5PvMfP276ayuF3IRAeWjxlMreLhFpCEDhwLQL0Uwar3Ajx4Y94imayIQ6qqmef38Pjgk26jnG3OM
T7CGLvQ22q1hu2VJPQZkAbR5FEcmBGUuuI+y4SXpi2KVVDYHL/xFlptPKyoPUf7QfYIP8PpF+H6a
441Jtb/NpmVwOc2baK5oj4STT0rAYc+0bWFKSfLCzqJWqyOgdQITfJii+DaHtmMBZTOjjSKU723R
Ze2ZIBUhT9YIBeCefZVDBdp73P5tCOPAylcSlEgsTl3GzTXS0j6Lb3GqIwb6hDjp57aAcEHrz+fS
mtvy851Iyjf5dtd3+Q6aAFO8Ggx8Cw5DExy2ltJRlWw74GOngjwAUrsdCaXUQFMEGOKon6Q1rJMm
eMdS8mEjP87dG1KIn5zclXcqDZ4RXAUuyx8+rE0bY8PNGbN5kPgcQTz1LaR1AHGjZ/v+OIKUrrsH
1HUCWdYvr3xWKXg1+jrSzJibpbT7Y3zNJvYbl01CvJG+7ltU1WqFA9qdSaeGu4xisJVe7pufYhI3
b9Qcemybv/b93tCUG6eQg4nN1PjZw1aOcsBjb0Pm/1T7hLKFG68T2HbcSAmXsuv+9vo7zDyYgclV
CQwGnVKg/xKc7V1sb6Op2L5HFywSwmUcqxSKy/ougz67/lG84K7/1CzI2H3xlP/wLSFTrK31GyEN
uTWIJjHSPLinQsxQKfAatC3L5gxVjUBlAJQIrdor/SuIVXL4C1VDVNFQbtaHhOEI+I+gW+TZ9a4K
/wNJRDTEwZ57FswgAylbWZhSwfx58hIwekg46YPUhNmjzKna6hfwC2dYyyfHYcw/KniRUlb1H2VW
vY0MWRXugOdZNqy8RIJEMFQfWXV3wBgRJTkDGj54hdnKTLSmGHkzneCXMscg5JzfHdamKGErEB3j
lqFUY/W26OFV5uDl5JrHQ1eZwMpXPNClwUeU89Npk+ivf9WTFRanV187u+xOqfmS5u+s+xZCFHXA
sCBWTgMJ6HyViXNXLY/121AUvrYjheHu33O4gb3IWZR6sgD8EV07zh/nxz8uNhmNzuh/oMHKhwyv
s44ND1OirW00DaLLusqlgqUVX9UR34g7io/PMBToe4PP2S7JE99okbNwalZwDcZ4A0vDX4kK/S8W
ZpwEbSB8SN9k9Wg/T9elN+ml1x5JZ8nKR673CLTn8OGfy2Yd3OLTrvYXVdeIsmL7PrTieYUzxcdy
L+c6QP4N9OzA1XePIDl5RonIiweiLUwVolw4o9rg1M/z+4SRrwl3arzXpIX2WvYTBgI6WemMqW0P
rov/GVS3ZPBjRcx7TMn7Sj80txOX3Jo/IXqw/1OcgDRn0MTtxjbA7+HIxuqjc8p8mNt2fChRvkTw
z9EeP2ILTNFfhf/KJQzfqyriGDgjDG6eJmGneUpXrEMD6Xmb5dH2D3HExNqT2CYi6fy/VkHY97sn
9z5GhZqU67sGmM2D+XcBH9ykIvnlTtiSErG+iDfDFQYkEnhP+Pw39l1YmJn0mtw4hIJiTOWu+8yW
CUbVoKJaDIbfV7k4j6fyfgFpTKge/9eD7tYoJlQ84UqnSLH4cqbQe2kYaBbkmv9i1wbfBKemxvR2
uPQZGIHXpd7F3jhOB3/NcTMIBSOIlX2d8KvZR6mxp7QfTFsiqOGxDsEt+5vkxUpDFifRXiLryBkf
h8PWSpNiI+P6ZWh+0byeimg6RfADb0QMvThyOhGD9BLwDfBvZWd7PZMPvtgXrnW2svhsfWDnxTrX
D/PTcP7iaUIAYkAYhmuAkmFEwP6pNND49SqAouhZu3snuzMhDSvQAkyhtStK8BwPBYq9cYkN7yQN
3m24LKjlGxyLrI0ZFOUG8nFqkdz6HGZhxyWJT0J9efro4LmN3bk/uRdeTY43eOxZKecdp6ObLPwS
QGR2v3FgihvI4u3uDEx3Uz+H4Pa8A1M2jyABZirHp65XPLlvKC05/rvDCXCefFkMmaU/PMroL5ES
enfnZ6l9s3Gmg/C2KlbcHQDTJ894LLEYjQG++/GMz84/QR5jC6mkyEDw3uVVS4d949/W6QoPR7IW
ZGJLXSZlX96FFM07WuFmQ8mcMftTqE1kSsEH5bPEHmpCvsT/Z8BXjaU9Ke96nsUAfaBVGfhJu9K5
cke+fDxfVmdCpntEschGg4GwiiQPNygYhJAh0XZa6+snVtZLjotzmqtAbmF1sxK5fwUgJks1R7Uf
CGqCJUOiigfsXfDrYvdiid5Yy7p3SRQEVhS7sraJT57jwJbjWPL9/W6P111gcgiTXqLNZ06hkltr
7JhiVlIwkmv08zys+SDOVTAtGVXxSeoK3RlDzju3QM19JKFxSD7dArDShpEngAkjZCOz4T0niLWn
vbyzJU8ufv0NMKBCZeDQojiOgj1Lyg+B9U441hxwl7AFNBu6l4uXUu+yQ8JCXsdxc3rIjOo+ksJn
VEwNS+ulcmIbOFlEAZoOYGC4RUex7gMYKWY8i2fpbZ8c2b3/tAJSVDHb/kEVsZjVUPlev6OtSyX5
EPz7/zzS2Cl2677qddYs4Q7YjmR5JG4E8UYZLXKr9BgB8STbhY+VdBRJ/BqY0ULNDx5bDhg+qlUI
n05b9pk5oVVkbZPDAdxiLLriErxgw29P5wNzpP07uyYzbYYOdwGNLj2N4Xrm6jxCv0qBD5aJ4HW7
x91mvcFgX2jSpxdkXfNYc6Rqhv859jAQJYU+6bl+lB8docIsi1ZeN+yKZjeq95nC7DH3oQ7tBJQh
X3ZILQz8fxI2OIU8zespATYOON4tIwoJBg7Sa8+YKE2L3XoM7fnedNXnv7M+qLz/o//VJ3K7frdg
Oc+rFsLb1fUW7NtBn4ET6TZWpcf0Vfgtc5hkZ8NT+blDwkQ6Qo1QzYKWXbjYyi3Pp904G+AQYW2O
KdYyeuE+6LrquaOPOqHsfQrsg1NJiAXuZP3ZcvdvpMf8wVMiQmohrIg0XJS/tsqTXPcjz3ZyUXlf
N7WN0ibaNCMDse6+VA1Lsv1zzevbQYE9CwMTZtFzI09RIoh5uGrd7pqAGnQ9X5DcX2CKAsb1w4PB
My/b7y9qLm36UIOWn4wTicI23aRABd+R72zIpnZbqDiSt3BD+S69PiNqWiG8ly4dyxs2nrOE/Yqn
h3Ic7J8wmFcor8wHwLAd7Sdoqq/06jppqKq5kCrVxs2JjY9mwpFOYQQLUMmpHVs2qIZlK1hLYuGe
LqnqMnTYr4ufopTJv+SnrTmBbfrlHRwwreIfHueXD8MyOxgjg+Y5ZrTh55zA+o2gKgNDfXaZCg6M
b/nHpe0sgBILcISLRjO3vwxzB86kM02JgKNiWyvFONZbPRf72j8wz2aWvmveUm59CVs95bAjDTuj
EKbtiCyXVLw6Me5ocsdgYOej6IAKnB27voqj6QHkzp0/WGODpcRjG8/O7nWFeIOW8DjPf4UWAn7P
+k82FsoMOVUBaHCGHeuPCuSe97B7uVIjT2nlHGEd893J5GBFaJV9ojYNPPVJo8uVvZkutPsPGYkO
+EKs0nADbw+4IaMRCINFYhgq7G7b1Hc3FW2peS2q2gZb6nMSQpznSwt0F+eX9x9KOlIsrQHxNfy2
yXM2Zlxa+rRtLLhMcnrhXw/r+LBJwD7dOwwiStTOOf98h1UqrYFtAHDZ8h/NrXcqbyJQwtqEUfYo
nUm23LCA/er2Fh7hvwBr4fK5x5/yOf2bLewJgiyVDFibQNnDExxPylqVHYbW4STllgLx/PaedJBG
tFQDBIOruiHEnI+o34WRz6Ah2Q9eW/kCQeBSMSxhmJiEKxvYhg0wvVi9yGF6iAJLnz+resknvfRr
rSFLEFVZ+KGjPavtf2DkOS22GRQ23jWdbQZ3TMRczPBmQNtKXQPjAzmlHdjOXVbP51AjCDJt0FIn
0p0FsEhN6aTP9Lut+scISieT90bb8IEZM/D8ovFa7PdpWlkqU9HcDDHY9bsqIcFbfAbyDRiNLDrG
Ws/QZQBXRpXm0NK/2nzT4M7EiZs9xOxTzkgXIh1njFBWcq+UsVmvOLgJ4ej+PdK8t9lXq2nZwq13
qh/T+N1o848hG+0qHqdhQIbF/gwyE06qRo6qzEG3OlR9Y3nLrCHeGZt71WXhje2GQaZsHBlTXFo8
ofpLH9KBsq+xGXOaJ/UFba7zWxbaZ3QKxGJj1XopfadNv6QY/dh3fmxcfl5uwRQ+aMWDnxkOkvPg
kibVwzt2lqqHqJPp6BlFnaMbiGAKfyQxA1Bd2M/beHvxPgPFJV1JaXuz7eLRvz8jcquZ1VROUZL9
u4NlpTX/8U2jRFqCjAdjO+lrI9+XkPK3CCIYzBVd/miOCs8Q0bOqTKjBW1/XbWwIrs0ehdMXCFNl
hhv7gvl00WKcM1cBvh+pvqzCkAT8nznVyLFQOjbFL37jq0rjdgEEI9cEvEO7ak/RsX0AGID7a2Wv
HR5aJO1Ijqgu3WQudMDbHBRwb0P/DSHHoHUzSfILjkX5JP0FasK3KuLN8+JRBRyxZS3FarIeRgMp
etnpDsgtQwtq+B5l3oRVolC0PyCbkaNg8Fis41DSIBncu3LHlNnpX6k425WWmHT4uiDDy1OhMUyY
t9w8+knqRimmDHi3mFnJC93EhZn//XtynAinvGYXR390yccDeIbdIsTONz79yLA2AwLKwDgwEG8H
sdq6OGgS907NiPFULZBxpVWrkfJ2z5ZFa12tc1FZyriw9WNuDsXH4QwKL+NlzeyaJVOZ3v0xofSN
DsdSAoqjfjW77y6XLeQZMlFB5h7su9fyWxR/tLubkrkoP8NF97hKJW4LDOE03Ac8Eu8uLWaLhk7l
PLCI9QCYR2aiDKSZolKJqG/+aiJ1djZdlGS9gQkz0wlKi8BZu0IGseRMbJAaI9eivKX6JKY0TRI3
C++S2h7XrCFd1qbuPgbJh40b5Y7Oo/tu6x3fyvk7p0HnEUFC3twh+xyPTI+/TlrNmaFSOe/0gehL
pz6kHN+B5fAS4zfQxh8wW0yUSPJiN253NVEZNJECpnC5xz4NV0aP/bfyrM08pkpcWRBFuRDwIezn
tMgulO1bNONAIQEU7RU+LtQN6kRIyPNIp5axWaOWMAJO6DMgG5aZskINNHrL9OAFOemE6qIkxJ0K
iWwtpP2jUrqL5C00RsQrgeoxt7TN5+vV7VcoInA2fB84SE6txBtMYRuQ+1J0aM5K28grfmX06RDC
CfEjczWZxk7MMhbCYLgOZGlKo70Xi2w+Er1/VYVDjKc1n65EZ4yB7ZYkXtGXMGIqDd9m/DQpcZ7r
MqDJweGjD299iiM5TXCaZO8mqXNkYt2+Sqw2jIk25/9fcHMzxYdkAkUnTkeXmAujgGoMTzMbN4eK
edWmXEOiCGEZx0Np11Vx4TjNRu10wztkQPJEXHRqu0tnQhgc0CcITjab3OgRyVZTD7d1fKN5PVTy
V10Mi2QxRhTN15iLZIK6IyJ/hf1rOxYDcYIyP6nNOXR3djXIo2PPGfStLL/A7WIqZW7AhE31MlvO
xXuSDncPvFprTEJVfjFLZ6e5rrHlTu5udcCU18ZHp2Voj3rJIbgJLouMpkhHTHNTYocPQLuLmwZq
kYKu6sHv8I67dxDRrcIcNcCeiQSQB+2OMxO/ZEjs3PjZwPLSxShc9b+Z2a1VOutYY39PPaxVL08l
IFG1+vGLh9AIwQDoKq1QY/xIIWXvJ7vDO2bdgkdkhAMw6RfABjZhQ3qtrVMvqtNqDymkGy4G/2OA
1D9XfSLkrDyQU8mXi/yxZaWm5LpKYj9mg4xnShHgYeVbxcfCwShWcJcnhgwYayVORqmB1de39+I0
SvEpaqHF4wamJArm5NebXHgJUvRU5smX5/ELI3R0HuzdifxGnm1a6heOXs+xPv4bNUnmY8tWyTf/
tJ9p3C0zSMZUYYM0f6M3Qng6U5vZv1bubQp+M8ntrdliujsVehN6azFlnTFBQS7vBa8WYa3mlshm
WmlsaQ29R+uPqKSbDoKGB8OzCR6y6QNbZkcJ2yitpHwWxU51w564aiEUx3cVidl7tUYOE5UtaJ0P
DiBhiv/BiKe/fCs3OxNDjOjCdbVH6mSjYGqP9r/rxpgx7jAsCGtjP3aYjwyfs/1y7BhXB4AU9GK1
G+kpTXY9U5/+Odjamtyuw6a4TLw1OrORu8lyKT6yzeppctlC1EIo3GIQQuMaIZxS/3zp5v5s9nAM
aiMJW4MC5h5wDUb8VjAJbwdBglfH15xkiRBaUdOlxhh9iN0OIJ96ICcVvaRL3TA0gduz/R8KJPW2
01iHed3OWFWIGGdskWxO5zfdI7zhoA1i0Ox4hSLw3Us/tG8pNvzjnt6fOpwD9FQMZYi8tw4m0bMs
WMCHQPTQj/PaRiaFXNHUisqMD0+KpYc44kCS8ijBsZ8iLpwrXCEyzlqJRp61J0/ufZx/pHOmY7f5
RW7oHxfCvtzzjSlQIyavhlbKZke1p7CBWcxPXEBwGIv4+q4HkSRVOWBat7CYJjJhXH1+fZEEBmlu
s9iIX8cj+uwvlk00UHCmQpw7DCGw+0CNksizIpR6TUNteGpUGnb7RYGalPcQSdwDToUfQCgVIiff
VxXlkIX4Tiexf0J4ilYdZ9KbNMRbcnYJPcq6/LQGptHwUVrT8qkQjDB8H2pubGtRoRqGReINlSYu
UJpzojk0qmwLkY0L4FMfFkkxkZ+eZGuxpub9saYROvoLKC2wD+H+Ji07GtssktL/l9NKrW1x5PEK
OZQPmKKdqvU6Knwg/UdWcBEDyynh0mfBSthwb3mTTj0lnvpBL1VKc7x2Rvq0zKljbhs/shXVTe/n
JHEAN7G+Qsr65E8tvC4y3Gtqwu0/CnOYZgaOIFBdhqGI7sYzUV9NCpJ+Bx7Wl8gD4xUXmaSEk3+v
FO9KO1X8/Pn+B3czLb9i+Pxvq0gBXNKaNEJv/CvnbG8rIDchz0D72HdpDpP0M7n1R/ZS7TkGNaEo
sOiylYJq0ahtTttUyL/ari3phl7SkAJbvsVimeAyAJ4aJ9WVjnD7K+oRODE5gCrTcoRc6AjTX2Dj
YhzN9Yg73yBhSz+m0kn39ImQ92XEhpRViuXPKmqluWCFgYtleezOxY1v5zPFiGarSbpq1ZYaw1fA
LkccUR8PXEEv4advwz63QAcAon8e3VSqFS3RNnyt4Cj4lFQ7htF+OlGO1jDJYNK5GJK7KpspxVYQ
goWPQC8DA79pzUtLo98az3PUPnNhrR/o5bFn0mdzEKNKwf1nqqhAyxZfC4JDmcM/1OSVYMLJV1eu
u3AhJPlGAO24MqGbQ8f2GjNBKSzp9mrYwQ5EoWpEz4KAIT+bYLMi+ICRmDQmg1A44k+ejwBGApJG
XNhTKteHq6jxU8kZ2MrLRBRdy55ejLD+Js/a8eerCQkYp4MVMh0pkYCpIt27tLce5JrchxPI1iX0
YNd+xWNI7vFn3IEUpgKnzT7ZMndXX2Zc2KAYBWfXymWkeJ9glsjVtlYr3tJP47ond+vIcna1l4eo
VOavq5dgWulHnpvYMnhuQulCOSiAOuR2hjtnJidAEljaSlQkoCU9Za656GUWd7QW8RlDqce2FlZy
hW7ah2ushFSxpe7ZNYb7fTIdpebxyZJACd/ZntDft8gN8m7BEbVwnkyA6eNUbgGcAnbVWjmbndda
mySTx2hoH9H9KCX1215Ta1p5sE6S0oXaYihERiskeiZU6kKzXtVpUGawcOJdg4R61n9nMCiIHAPj
AQgl1LsavBOrxTaxwmaq921ufeeyH4DrDhkV4J8GZjClU7R77o+U4Wu3BSAdL3bIi/qdw2QQBabY
kn669k5AFqz+GP0AaJaJEH9SJEnHqavrDvm3yktarTuvn4n8p6JB4BFB6OdLKV8yxCmyQmiUvets
xIXxJxVmnizJN7u5yOHsExDCNc+FgwcgNT/X2ZOsQz5DwZqZqcftbhiTiQ62yRO3c02Zu9+2D1Vl
ZgNcKEVBzWkTcYlCu5VOsFda7I8X4ZotOiU1FG0ND3BayX/EdxAYMUI5XMkzPvKHHvtZU9M/PVHx
HyWE3O3AoaxdjpZxgITzeSPNaaeMyVbLy6FvyTyXD3fftwOLiCPurrrtI0XN/lmhYoZT6peViy+D
E1vp48GWttcrRcYBNvVihGqyUoJ7D9vbaRboiea73eQF93r/6zPkEx9jMNON+6jN7z7/If9+T+1Y
hGf6/3QrGBzjhzE0xAFrSIF3TgQljNNolKdDi3sG1LOVuIph0WalYDL+FrBCn8QWDcpsAaVrJ+ai
Pi49PxLokHMUUwNfynp409hAE5M01KwcoZ6KhmfLRxw5gEKAtVb3zQyCD1GHLTS5KRoDJz7qqxt/
DOW5UhktsLsodlc3YKxBmNfwcqTV/ECXQME+3uzYZS5FVPQ2f59xyTpULl30DyQQrFDrACyTTvgQ
hQuqEk5m+WKBZJbdTP9JA6Xv0r8rNAkYDxQ/eoQtVweK7opZL1rBN8u9sMxKAxo8MNMSc0JWD2lQ
auOUv/+5Om5o5CxHgEX8pbrpogeHBmLZRqemzk46QXVliYAmdnaUuClna6BHeNokhU/KeapTLA0H
kg5T41dYZ5f4JfAVDf6u8eT2m2bVbmef6l4Y7cFt70+N/SCMKWswILxLzVEflETZ5/JGixP8odkE
I+/1RWaJTN2PlAO6PHR1+Tk33nozPokP3kd2Zex353RszPXe+djP84gM2wq+gymyMJVLLUC6XRiT
Om2vGnVKEsQLyanr8EDauEmuyuskgMDmeXY0xCGKX4qJMvno1wuYbeJ0ZeFUWaqCkSgMWFCcKzX3
A9JaCIXRAHmgKPjDFCn7JLcNj/cJw0fJ21cc3cGcoaIUNOD9enIo7qnIxf5VMymXypWLHnlp385G
BImQiwNuJwelRePFDkLQ8QntKNZjWPXpvt//ZaG4076HqiLOZUYZADdez5+muc/vqlQnT7UFi+HJ
EMTsv2i35ajGB6ekDQ8l8CPfaQw75b9L7ReJ3qLXgmmOzjAXfIyUCW/MbI9ntfyeqvIAfteuYqDs
t3DwhVL9Vkw4qdHnHHzyX+o7MDyw8wvoPPmT6fvvdVwq9x94CLnwjdNgir8sSf6C5Pi+cUjIaLe3
TW6Aw4AEGi5Cp+Gi1KydxQvEfW6DcmNlkOweAxy77R7+6mtKl/b4WeIcPXTRUnGNJobL7pd4mhbi
ReF5AMZknqzx4GOFYvrN4FRytWrpZnY3m8H8QAhprc6HEbYwz92cDM8NzDS7m3jMvQn7spVeFbWv
q6lUH1D/sVHJ5/RypPY7dkn7PbdQ4hitqCMusWH8BjN6+T6RMmebp0NGCQeq0S2nYWu+U4jgQ1XE
BnYLwNwWZLzOEUo7UbjJKEvjcLzbf/zPeIPBsmsBdbcVEZCjXaUfoQw8htR04TpQAURwHWRUvmrP
rFuThZ+t72kJHYuLq0/2slDoNWdi0B3PXGVPzgJ0NKCDG1gFLhpJ/8uouv3TMTLyErr2nGK7n9I7
JkmBxvnOdJdEOMj1qh+jIDk3UPIy2PDGTIW7VZo8099/Yb/qfn+OdfNrcQvpZhcpNSubaNV11WtT
ph7C8ReDhVrtWPeri4WwsJfeh/4v2exhSB9lDZkFtmNCBF1JHVnGocUZJ1aMyHahARiCaEa6EB60
myepZ9mP5YtWPr9hir1HMc6u40O0Y03AB2W/os/xt7ngHb/YRchLDWQGVPz2FFszIrDRLU4PKXNu
0IlDnBBzlhMyf3PI5F/S15Rxf+Bz/biUdW3w6BpWRLbWtGNxiYaLDbjg9c0AljYmHqTIgrsR/jkk
tQzkgkTxVNm8PIyvZaCuAnLucwm8HwOI7Qk9jug4uujbwzXVRLrOcfwGe06wAGcrECmyPFJvvcI1
U+dS/RvYJ77nUpMGmZvraNq1QgS3LaZ46GrpUJN2CNUxHYqkazqMEYtSDXiUke/EYRQZu+RWsaZL
ljwrEr06JDMR0q28W65Hsu8H895R+H3lfWvn4bYjQc9GkJxKsKiLpuqphJ0ZNUsCIvABrS9iSmSF
uv7It6PNBZKpE6wtrNTdmu7/zAt/L4Fnr1fyC3VLjAVAEJ7rYFLFU0qnFQ+66bPP2i8MHI4tZiK1
t4t3rF/kVLoRqJQv6Yg8PVbp1OnUMse8bziM5MhVhAAwEDYf6MJWwURmfzgmlm0NGJZcpABRp3nz
j/UP80A49fFKzSBuHYU4TEL5v1RM7HBTKAfiratMBlWKJCaOQypJ2mRNjYlpHjoq/MoGRR/Gi91x
SJ2y4F41nVViZUDmg0jayb2gCSBw1ZAE+SVZWZ223/MdoIDW88hnuQIE9ta8bw9DJElmWLb/UPep
6n4CH+dNVZOPHm5NgITFdv4uka3D0QD98xpo45v3JEHaVAzfHVgDE7orM78EV3X2x3eZ9GJ5VzFz
xjJ38w67PV9qUDOQTBjvQmjp40fyC5+XopLj8bR06gEp0/pM1PuniJZCwJ0+BZXuUHxahjxBoxdp
R9+7/yu1gPyL1sJgFPsupECypj/Vef0qPs7qfbA6JWRR8oQD2ksAN0ezjtB2j6h+O8FqE/J9aqco
0q226NyBkqTGx166ZfS/UjgDKTYah3J/FA/JC0FqMy0sk8SqMKZqvrWpaPhYv2PFiS8iIXEpIdyP
xwD3tiAgUkZdiUvuLROcrZXX2S/kqxdC9Vvo0RlVXQVuBJIRvTlwIwwzAN/aE6y/IeoMM1GODovm
ODmF/D8kBkVmjbi+v65R6WOJuQE2aGCJ6DNdWABZZa1p7qWU9eeOwRzq3NGd9uZURSjAVxFDOYJv
XKRjHztHkOSzPZV43keTA0y0noaxf5olyoFXOBy8BObN33mj9lMqMNBwb8Q+V/ZZdi6twjEgIQ3r
4nV551KlQG+G/86V9L1Tq+xQI6TvgRlGAxznL+8gX1OI/8+x1IiyItnlUX+//4m+1PzpufjdIvOe
9poZCA+YCqocFRxxii+IGYFVAMdkDNHcYqvHbri3EiMN8wyU2LawG+tLaWYGSmneMEOAxmxXKkiZ
MfROI1QYMR8d+Hdj5bchmluYkVhlyn8kPpYgMD0yclsfmwTX9N6cYbGjgZVpX65VJZIebbDA3Jtq
bBJReDmNk85T3JDt2KIQn7ZAyF1t04YSGSiGibxIeyLpbkdhA7SK35404EPhfj1tKPpy8tw+oYlr
80roc60kdPcklgOpJ1r0GamUnO4sZyzocP5CxwPEcxrZMTuI8wIbY/fKSs0Gk7Kp1uUPp3Dn19gn
yH9fO4A49ZJLV6tTPqjaLsFuxGNgMjVZV+zjg8a3wQj36/LghwvCDCK39WPnjWT7BZgY2yI2pMlz
URu4cK/H1na1NCqgQN46X6phMMv78IE44WU052ecF/K70gM0S0Njxzj+Om2a7kKFP37fPxthqIAf
PuCEY0M4YDZy84kVmnxzhODbYSyeGjMLMzZCzzLcJn4BIgJurY+KmGTRDdsIa3G2eXnAfJgdc/8e
EzHnRloDzdjavhurN+2FhG+bYgW04SjU0yhUs48T1BgLkNtMXV1lQ8xe9Nici0mjI03fRThV3yw7
6xfFJ5qUiQ2qUpPjfmb04RWK8vfMSP+J+VpAvaVbsGEhrb5WJTesgwKS5rKaJkn1NShrwBzQ0jK4
xtCuZTDJwr8AWedYoVTNTV/Zs6kDNFExuJgWPnZs6J8DVHmdETmpcQH0iA8Dcm+83xv3MM7t43F8
TZSQidklP+3iSLEtPhcmb7jKOgF2ni9zfsBIOneg4Op6GVObzF0vQOtnNSg6w3a+mkKU0JBwTF7W
G7Jk9rAmPQeZ3MVa/HBt+nCuZ93FhtOhs+e4ciGuDzuOldUPlWQj6Vn9hQnISGF5H/u6TaJPFjjx
4F+GIFijgAEHw1SREGFHi0o9nmKiS5zVZdl4IE+OBeq2Bbo/M5j4m39Fl/asS7logClaEcfiTR+7
AhFyVJCOzK2EEgbiq7tQUKDkHc6bvDpZwprBBSrP8DJhLUruyzQ1MQKgDWS79F0gpS0nI1Ym/U/L
n3XmH6w3h/A+0hwgJw9ZMvboQg6h6581sRj5+TEQjKNfaXJP3X7ErbyBT4TZuQ3QTlxu47bNktgT
itomFYag6lS4XZIvAZt3QJDMHOJ88NIL+Lev1xiV9lRsJCZXXliVtBMmWTh9fzMnbpGIyzPUEFK7
4MsiFYtrCf2AC3Wt75dT6VIkJe8ZudjNvgEaZ5B/FwVL8+atAboAtuMVMHJAEvO5bvuA/y1erLtr
U3Qhv3iOdow48Ck4hFV1+g13Y2fQAXTACdmdOaPQCHMmqU5nhBWMJfxsv45B0hhRXLYmZORUasaL
kDIKGoFQ3fmnloJgRBN0QBK3gMl/+mkhaCz8ZEFl4sOZYpOR0BFtQSzJ6r5BecJSL4buhEWcu+LL
3ba6isKt6RayrisN/x0Pd3s8AFaoYA4VnP3iLVCI4f7WVwz2Nupd8tKMYlwpEdCx3f3Mk/dQAHrD
RzmdSxHJ1q7vlgft42ai8xigDVAqBRlIhTaxqp1RXDRYkMbXLmsO18jjwORzg41XyrSMXikivB4z
xZs2osXU+WUtefVU11zI/TKdkUPb+1LtcV3qdDd3GWBqDkcPc5dENSRtdKuAKg4cjCnHHCpKosnz
jEiYXsQdQtgDT6tHG5FlFKqdCmKk2uqvnR+EMIvEK6IjOpTu5tbsUproype2JQpvg9Xv24ATmWDd
uHUJvbvdNoZyj1l0zbwf9EsluSyzxcER1849YX6O0nGCBAJDCt/FMsgw5/RLCVgh2Itnr8FN+yWW
3V4ZVarPWlmY7gD7SCHrJ9FwBlxoiwmO/LGOm3jvbaae8UT6KqYE6IlLv7gns7+6cHer9RM2cJQs
tXOGMD+c9aYOb8wK+DFqxl/kNgmhj/It3/yOMaUXc3dH0JNZT+IVMk0erH2MpsSF/9xkYjln0AXw
0TncO+5f/xjmfsS21C4ZAVB+qjP7fqab+Q+e6OboPyZ+90kdbmr3ZiW44iJILeSnO0kHxRlyxSy8
giCZlaMbsZZFHRpntPOyqagbxz64i9Nz1Rf/coP4Lp2U5eTVwnukcIN1BrdYupqVaIXDYdmWj7uz
xYyTy4M1FlR1ua++S/r0B5Hw9jr3HTUgrarnOC6jw1EfR7cymE4JL55zCyS5WRtPBFKgyIEQhtch
KUvZHSKhJ6KHMdyYxYao/uppnnLat86Flcvbtcyi1342uRHUrzo5QGbyXhqElJdPg9/mx/iKuzV6
uRr/s8+3KFD7/Tvl1uaWxK3AStqfXyuTdrHldpu1ZbvmeTyp/jKm87tkcfIB7SgAd2D54G0sul0h
xS1jyi9GTwuWTyrhlthjkBTgacwbMwv4N4GyWFdA6ly2HCPTQn5fUp3cReniWQTfCmZ4NJOk3kdo
ddYNry9lkHmaoaCT/LdB5k1EPWgQPP4tMa+28UOYrHbibXnYekT8zrhGuh40tEiJey1TDwRuPeQb
BGliTnar7sj69Y5MFoHQ+mOfYP1Jbf9og1VFTRb7fveC4OnZ4cpKwlM/BYfHWrhal3/KUsU11uY+
kXQyhObPz2wJ//Hex2ACttDRNxYigylf4czttSVo2fz3zOBadI+zoakBfl1dKuwK6H8LTvTjbEMD
8/NyquoLG8T+9lFhLKhO+upS6CVwygqtDbeilPWgPf5O3PtdNiwnwTWfoI83yB8LMVr2cMNPNA5Z
pUHGCh2ZNFl7KuiqrIZQzNfCmWo7gNLn78PisWIOgs08wzuUSFatTMZ4gbyRwCzbNPvqlP6NPyjx
PPAkNsAXkwjOAIJhfk/GjnoIa/QfIriydsQ88NZ9Mm0fI2ea6Pp8zwGWk3jqiI6lXpMK8OOBj++I
JRFvo8SRhQp7Ov1h1mEyc5xxJvM67W/fRNVsUYH6CI9gJP1WFTWBymWVgHYjgGCyFJC0mtg4yFVM
i2cFiisNcp1+5bcW8eO0H3M2ZjllZ26j4eK/Y4yXoKQ/TYrNkIcch96TYNybS+WphsB6G40sRhwe
za5Qm+M7wf+pB137dPQLiencvfPir+uQAMY8wf7CStrhC1bTOxgQch0FpkgcP2qaqnRSXVQxWi25
MjyCcUY00fGc7jMSm8l9s2mjNEXJThjqkTRK4ET+ilXy3eknAWDSQnoFSi7E/8xArhyMq2Ugx1dv
cIm7Zg9xlMm94Y5GN5LHs70wnn2Bc3RBZFxPj9ugzNjPoJrgY/JRonB8QAL81imESgPVVKqJTcCR
XSZxafFQIIsLP11rS8bvV2GS4kT2CeIkBoAqlchXXN1of3LbctX9Bz10S1nNJMF6oMgpSCrBJgNe
ZHTfbw2GTm2re0JWmrksT0XGkYF5drIoGU7SOrCto3VRtv/GHZlh5jmbWC1zMcmwUAaRA/dv0nI2
XtDeCpC3XLOd0wVkmNOJUdzr86tLrjz7SU996jh1+y6lj+NVRfhd99vThGQDFl2OwlSErjR7X/oi
3rocxdBULuDN8qKHbWxZ0dlJOuvvO2pmlQZZdwkfhh3nozPF6NFPYnU0FAF3n5lSgRJkooC1+BrL
06wdO0cRLctOpwtgAev9UQH1W9Iw7iZ0b8YboBI0OBQI1StMsAYu+Z2BBHzw9Vgv8VjmncFteJvt
4U1pHsqp9+vU1FjXleA8XtcATJ7AsJSvTO1i2rhx6JhV/CAx5RNF9V39oFzBhWesEiZDzGPpp7Y4
kKWeEw6CcVaZ0pxikv8AmkcmGGFwubAAQ8hpvqTuUfdqIszNgt9kDHlAbc7LFCn/Z0/JCi54BWtq
7knmZl2hP54qm2MAmPxfeVGpO0JPTkTPQryZEyjkkmOL8LHDyXhlmlhePTbilrlyJ4WCwN6lTX3c
M1FI3dW2tBg2VgugtIckKRAnK/LLlHHpoG35suBVQLGA38EtUZB064EC5zY2CvGYeaFZtEpNgJJs
ASKsBWJtT2fdsDh3p9w++1/D4K4WhWYNYN9yJDG6aRMfkNzXMeyCVWwHeb89wJGpnLiNZ/eMTzIZ
uvcyoJHA1nEBE6gUV10siq3Hqz3n6k6iyRVo1X58Ze+dDeN3OYwssTuX9SbMQj+YhllRpi1L4vIM
8lqVbegyyylWo4p2U+/Vbi8pnPwvWSqvhg0QleydyxDPHtzsRhUOFmjH9lCHQ45G4GndghsDIFd7
bu85nYcf+bSij/7z9qN0YKJN+fqFZtV7W1nq1R8Y6q58Hdnv6KCiCCSGNNXUD6L8gT4AK4sqLWwd
rFoasFCwYd2Ek6QjhQsB7ZqvomKSiIn/54PfGHNyo3DfH92p8Xa5g+4E+vAde7BBwJySzN6yjx0N
bUWcuOYlkBmVm3dLMnbHYP5FOqIpjwU3b6+ZqgSXDCgxVMbl8rlExOHmhWEqRCkOc/LPxJEsEDEp
SGsflntLTEs8eoth4hd67sWJ2h+Fu25tnhPIJfEHMAFoTuHVXvnpYm8CmTpoK8uXyZ9IbTR7ADxq
nE3K1rR9XoLLCM9mAEi4jZ/9Q75SVLRYoUWwid/O4be6jBp82GiQh/d60S0CP63fu3BhykL5Ar9A
CsDNglml1ZvFM+qzGUYiWye8cB214+d2IKsUqwRXx70YU2M4bRMHvhC1zIx8DlOM/LiH/mymxNeK
K0QZalLMcPq/i4O5XvxFGxrLWbawOywq1fZGEW9mWSel9Xlpxf5aoprJHgxqkk+hjoGHUMLQikwA
cJ1pbdYm9If9fSS1wuB6BMZzO9DPxx3Xm+U3KrrnKKGeJOnua6EraPAOvJ2FFFda+T1uf8k/hyRj
smtGcbaeBkJQhmznJPTWzeOAfU9SRSUz2s9QUD2cfntOSuoim75XuT0p06Q94IKWmFPM1mCdlQtn
YF9nrswMCa3eQF8FI028qwhOqOEDgCNWgDkux0pGet6Mr3dcSg2Ufvvm3/RWCJxtCehZYnPxBKiY
H3jYwoYCshPZcg5wQylhp0Jwm+iEPnVNGbvwtYvkoS9lC9P1w6KR62+c/h/k5Z0JdTFBIE3TLvMS
PJWfneM2kyYrF+ImYWLZYjcKbGIwgrAJpEamawZC/Ked+VUE8eH+yOp+mOTH3iI4vydkPP3HAD6T
j2aDN9BnvIpGFuRI2zES5JTil7aWEEq54EbtafPcLewr6uVZot8rJkW0oCts+ReWsvn22/tNOnG5
YGQJjOMjco5osZJEX1TqL6Q0n4jiK7KZE+gz6SgOhKQQPA+tckAbjfgSwc/CyciyAWLd4uGxHYrE
pmujBiuwnS/ZSHEvcq5h6dbfjqDjFL9DLxlw+OUKSwU3FGTLkHC1Xmw3mLxOYZO0OR/PhacdJBJ0
DSdNuqcTWqb4bFfdFw3UeQwuCoHkdlG0A5v2jSTL6LSv7zsdcaNLGTqsNJgkwrQ9kqcuytTw2qwh
5EQ0cqAU58sOgaOCCFOWMij3IlZZY5CM54Qm8uFQtEigDJkUJ3cfztcL5EUhJfeY6aJ/fGkhiA/b
UzXLpkWuhy+pxVw64sCgXU2B/fit86ovm9Q8g9V7gYqKwkr6bSdvfnv1EilSJ30817ib/Hf6radt
mSP6DDNG2+y4gZUrLZDu9/78OMvieBsg1AeM5fNASJRgYtqG3/C4Qko3xIEPW/Pm6spso9f9rj/u
d20/AhGim//MzuykKKNnO0mAOQWfLg6LpqcE8jP9/sHx4oVl4CU9EFQWepfJkaUWTiM7nDyAdLwh
hCFYM7Ua64mVQ+z7IDPbuGmvSLYDIFJODSmoupPP4WxCuru4YocPp8vfKJOLuoZ99YrzePB1qe9y
JwG085okzQg3SdRZzuHCtwHzpZlGB/eO0P+4gqfVaBNqLVYvThs8THUQ4be72kvRydhf7UdilAXF
SSK3MPCVOvJzO5Cvrj9Y2KB5bcs0mGYkqOGGifXNlN6M9ejELrdvLbqemV7xqbLeZLsc4gkQ5aqe
JDYozPEPn+lKrEIiFu3PZbuURdZ+7e3i+NxgytID+33oE6jXIxiGFkovibYVZ48wEqaiyj/ZIasK
FZD5ShYvR564QzgIvy6Df784d6dcT0pncFb3ZmIiZ8FySz33L5ZsY0RTrdRCtGPfzUmJZNnLX1is
n/fBVRFpynpGD15HFmXK8xU9CO+euuNHu8Ohmp1Cx/eOygrIX0+yIEKNc2Kojl3KNzyzIoj763j3
at7/37deRMLFnNsaDXUDsMbssHKQ4ZrFsyu5Sc5O+Rw7Qugxx2af6au5n7HzPkheKLDatREjLsPb
pbgDHtXX8sI8+tryQ+bb0BYBJT63VQi3IHBU46RJqycHrtQOArVKvswKWgLbfN16dmKCNtbmfOHT
93YRYiG9LFNTxFputpyxxxWmK3nL/J48FkZYwuobGZznKcEBw3bcIS/lAIrZbCMO9DIp5GTOoZda
QJ4Z0L6QV1J/oW+fRdomvzOuQho/t5jbfH+RZGphCiJR5n76RYWiKf5uGv77PbCBroWw77Vwjpwu
llYCEW4iJG3PcaOtie0R9deL04nb9+LzAPTRnxSD6Ne0rgtopAW+lwrRGFqLURHsTcGa9HSmkILi
fG+HOY2YLQtzy6ujE7KtjTN1UCRegKXTrT68gCyF88HzIAaFczKolly46OfJoenHbNQ5oLkYfz0o
vJZ6o+TojZRCbvfx6oyIv0LhYlu6xhg3IsjiW7di65BOd3KU0yOogbcMcbgOgf5BmmrFB896MrBW
q6ODRI2sJLWpjqGprDYYMLZd/2Aw+FwK0GNNTSYVRTRZDPytvJURhc5P/eer7u/2HJG3Sih/l9mH
BENWoMzIVresTD5xzOmsn4ly2z4rZR7tXpEzsJawqAELAAzIfjY4woJSRNEE4LEe5TzKtHRJNfXK
upTTCHxJvvOaV+x2/O65krymFbT4LphqruVhlacjN77fFfZX5YhdfHiky3kwTg2qb8kz/Q0d0MPR
P6P9LRVrlTGjXiBGaj0hIVfnphGYrISSJiJvVWKBnJuZVzxSgR+9QQYnbPY6NnUTk/RRBdMH8Bjb
WWxTmRCQxScDplUxW3X2MRgINoHa+etqdZBF73SkJaOtNB9N5WspBCapknA7oRq6dny4LNzCs4nX
61dkDtF/8qIYjGEcv/DQEyb/VZ1dEDHoonAx8l+TFnYAyc7mqScN2yd9ATCB2BzMZ4eRLiu8xWMO
S4t7IiAi/HaegfvPLEjnOhL90CpZEn7qRvA+G6PgSDkJRJgTJPzxHO6X3eqmEYVPWs3J7YgzQGSQ
ZiqPES+jSiBrVi/qGVYHGX2xjngFi1GT2wZckCqyyNOd6RySCVcluMY+b0DVfCkkis7em7KC7mO6
lmpNskg5Pi773HhURVvj81rCaCf2A4gpET5JMLMFZ0x/pN2thlS5knuzDS7+I2jPPECtz3whUepN
cPjccpAEmtewLGJtMQoUG6pNYH/7GfexQbESuK8eNQnD8Dg+GQrmViIfVwvOB+V8syMvwBPGtiWI
2p2km+t5KYPp7kF96v0ZIn+w29k9drBRoy2EHnVEavrJgg19eV39YLU4jN1be5DBk+N4zHPni2kt
0l1nexMv2RR7KqCTY2udtxHK/+0t/Gc7IGJL2CaF1BZ4JTaf3oTHTOnqsSP9FBLZAQgnKpUGw6jZ
CAqk2G8tjfi+9ss4O1B5N26XYBsB0UqoAiMa55qucmGJaNmjSDBUeqKEEH1AOctPD/ZYBIiYliZ+
jbcKJiPiwUBpzZBesOdf/GghvB3mkqg/8ssACEJ2RsZZG9Ire5qmA/zXGdqwJvabAscxxxH9g0Uc
wDklfyFKbba/CgHxnYK62an5KMLRCbiPPsNlmDxOPlLYzXL42FaQOi1/Uf6SXhCwgrCfCp7jbKn2
IMYIGLpUuKJjUiYDg4ZzPFbHqhDehLp2WOrAUqvt+HvB6hA7aP5/S0iDFdoVEYIb6xYxkqKua7xZ
yzQsk+M8o4GzE7aTKFrNG/kdq9OizdIYNd7PaQ+VAbTGOIZSwVrLiAF1+Xpziz6FJHF+FoYyiQ1k
RKowy4nPMJnD+yacEbTsVxq+zFKfQHunAB4hrFVil0udUDMPvSWgqXrbaJWHvVsoLENe2Btm84pJ
HggH8ekxT8zwKcHYiHunvOaRBXt8OfuSHpOXsorVFvJELPP2MPXtT8/y6p6Q0vzNdLlq2KYgi4C0
Viv9MgHW8Uk2/Xb34jNoK8SjVRa4nkiKxQxKBZinEzwySMvDiGqX2KLR8EWwurGnRbljK3ha6ElS
ev1euGN0NU3sNcl2LjntF37+TcNQZBJhIVjmcf10qminXgzn59GaoSx8Eb0flogGBJaGVWh0I/+G
VgcYKF41+sl7Age/WN/2s/mvPfqHGlo22vvdcByQ0rppI55A8bm2C3PdmJ6eh2Hu7yxxpia1ngUv
Sijefhc497/SXhQYQOL6lUYozCtsw4aLdrGhRhtXENuOIbrl8iXkdFudH/chV8OZCFkdQzV1MG59
NBUGexLlNpUSBH7UPxnH0PLVzA8O5nbhD0prObcJ1YTXflrfl0pIrKzjXzsyyoncFiTJ/R/Lc1IF
YZr7EXRnTDDJ8akWC5JQw4F3ZirOqFK6CJ/qjYrE5+q0NwUy7+KIbT6/yXFYV76oiqNpV3JzQ6Ds
rIHZWWNafmdrDNxrjryVXyJB7yCmcfoR5juoeTjeG1ZE9XL4ylh5LMEWVmePgv0YZuI9G+lDMVgC
cndVCds90bvakS+2hQxZldYdT3axGrmXAtecd7af2WEEgeMAu2Hlx1g1FOYrWhKKswaNSViGODfx
iNmDsTdp7mkvKf78kYuN2xybXx+GCJ9jtI+cXlskmNgNw5BeHjprZX4dzr6nOJCa0pGT3+uEyAPu
f+TWS7iMphzo73JMkKjfi3IQwy10mo0XyuXDQsyS6NbPxrBPLnXHChbc9nX++YDjyBU0TwrTAihC
5V0v5UCyAOCgbqu5AGhahB/mBI/+ayZrbxcIvh3E1Bp4C3otONdjN70DoSq6ey/TWcdl5cdCEnJJ
oIMwT398XQNkcnTOywHmCWsW7cQCGFHwedlneQd6vbDRM/BfRLeSb2QrqA01Mo1BH8/7wDn6PI+R
t9UhByWiT9bOuLLeJ6JYWYAHjd1/70ZPMsicauPhnH6F4OqYAmGLUVPDXvQrPqA730QqZmN9tJ7e
f3Qp76YWHWvr+4w80QO+S0ytZKsYhJATHo16dIfUbJccuJ96JSkWWYJIhjLp7dGhRfipT/TP6RQd
UEcQhJNw1xa9IIdmy9i4VLgKGiSBpxa8dm9rbdxLqdz9lD6LdbdkPkkksBPkV05X50GGTnUUUcxJ
dyAQgGg+uk4w0ORmBtE9hYuLXy57FbVWGy7p+9VYACX2lX6UTZs2ngWKQLvQHNrdWK1F6tO5e6Si
I4O1WSlBOTbgFWHnQuntQq/TwXF3pIKrWkwtO0Aqoqe070X0ZeHibIMP8hnVtDLP67eQPdVkoN7U
wY9dLq7xWRJ0pduQ6WA76gEb5BEG1c7TaSEkhbR/OIN1wGpKBUhV9o9qFsauMIGKTzYJkL+R3TEH
+fezZcJB1GIT7h0wO5KLiRlc41NL1LJ1nEUgxYssMcs0/o7cXH+4WfV4hFQq6XX1WzGOqZ3ZTNmG
LXWOg5L/O2bd8tjz/BEH8rIfDh1D99fEKptrxdX75zGGfrh3UhG30t1hXCGPdUcW7LARRxEERdk4
7x18ygQZWVP38uqKb+KIY0vh3VDWsM4TDLH99AICEKhJ5MiMlfyh3CYw9d+hwXpVn3bm5hMXrxek
7AEUa4bmIxzIcU++VhghHHv7m82/PsM32fjJcmGKu1EoIDrnE9VLHUmQJcNGMa+SZ02YClzcnYdW
T5cHSV6gGbqUzDI62KH7ZpvfhrOKMutp/A9VRwWzWo3SS+uSMEFEZAhMnb13W17pI5O4UOXsKQ9o
0S0Z5UY8TqOSx3MNGIV/HHBKG7XUv7P+XKCQPDwgt8nucrm11sY+kewhhAKTNuvkWmg0CTYIzFeX
qc3HdbO9JyghnRw7qYLfprhq5JznsUEr+2eSwgLacsQpcBUFjbC8Oa+7Ts9o6scxDR2mfPXjpLHl
iPdcVSnv6X6mo070Xb0z5tXFxrqLJlFr6o3gBIHwrjCTlIjJ6XaQb+CwI6jTjt+sTHs5xRerelga
TNYLWHNM5AMynUld9QX32v6rvQMdzlQ19p+S3JK6LLc3LoyKInVLGmt4uXntJ0YjKvSVa9I2NYKe
2FbjL4Y1fTOfQN/LCThGIIMXC+STpTCnlnppgbuQ2kjykiFqPt1vT70GWGBYiX/i2qSoPtFeoRp8
5UwOuqdLpiUG/VNwG6kxdWZkKHEOf81ggLtNxGHlyBSlh7q5+6OF9WK0+RwHIS9a9ujfUT0zhuOJ
bCZ55wnzXVAm5bmjvkJbKnVeFpYAOFgzRMX+ajMKrEfbQzEkfGNIi6yOjLo7o7OXOHIIc7KnU2mL
PBB1phP0O0XCsmth5G5idhP6i2lMRdJmVpji8WmOffBBW6vmbPf4UpnbjiBecPWZ7cWJ/Po/WeOv
wS65s8gGqxjEyK6t59n6ROcf/TISbictosOWesouGRb3yFmVmCW0u2ygmUIbbGQ4IBLfsOxElM7l
4+rPvSeSHsRDp/sP1KCGi0U499Va9EToE3c2F4fuAqT7ONZGMN+v/rIH5puHTuySBDZw5IH2HAOY
piUVOcUzht74OTy/6M7xiRV/8Fz0HSOl6npDzE0A3/UQJ3DL7amP8fa3Q5uXboIrycoLlDJrZZ8m
hWHmO2tuY9UVtON+FODaszw91yMQ/WpINMuKCl0uw7XIdeYeuKS+KspO6uhDMU1hlfijWOdghyY/
qf8g6SQLwrULfpgCditDw43TSGIETkjGLBbLtdcz9Xe/YJABJJScH22bMJFLc83Zkify17/gHRY/
kFUelBZ6zEhwTfvKyDmQfiXCgLOkhnMpXS+/zdwnuOLSYUj2gs9+MnEwAHpiIqD5NWDaDcIVWmue
/Qj+fhvVPtn8M5mGNpStTXlFMtnXESjUSPHvNg5iaGFg8oPs0Tkqvs0zJLbkoIFKS7ELbFpv/E27
OmBvI6UOL1sFONZXxYkyg3EbUm35dO71KqbLgNilPlB2Q+ZgQUJL9Hn3B80kzY7X5kHRwo8MBxu+
dwxNGCrquKDrzqVMOCmPOzEMQSSIKG978NpVnwlAFydKZYEUJWRmfCt+igtjuufJE3NJWt52vKSM
ZqHCqmu2sc4LijfQjSQSUv2Aak3zlEqgE0vR/o07mX+rC3QeIBrSRJiOOkr6c1a0zgWy+NioKIBv
FK4UYTDRxDIuJs1zFTpc4NISJtjqqh3RxXD28hyEVrf32MMv7dCOHcLKkVyIDEuqXYtZTYwTExdo
34Rfc7FkiS/YJXUcEr5xCdequs7pp5dew1PFOP/PX3Sl+R9Up8AWHUpmE1TBl3BezNrqNwLsctc3
PZNJu2GXsKe8QRZq98la7Glx2a8BdCZT39ILTWJRNhh+AJrVR2kHET45D3sZL6rNQdKoE91HI/Ip
QduYiIscWnkPrJDRPxTLaieOVFTYHixliILpx8kk3IqI952u5FeW6Ae0ptk6gfw0Fi+c3T6aDxtE
2eWInr84Rj6zyVfyXE3q6qTVOVXj+7CXZmdE1wokhu0FklC1ZjlPJN8qDtDdrTowzko2Rb/8lRcK
ezRixCY+heoci7UCiuAFHpTvyfNOND9IE+Hivsv5Wg1FzUqReZyz/pSqZuYgVjXiLHS5iA5kN6kB
rPw4Q0oSXl8vZINzqsGNjMdJsNSFCIO+PO/9zqPCxKN/7776s8eIgbRV9IaNPm9Q4/582V2+zqDN
nTrwNw5ge0WT9UF/U0mBjORlVa1AMMsocILQryFFPvGbDWDk+ULiSHq4Wn/8djvfRDOxEQCR6/8h
nVtsX7LftmUyK/r8/Hv1YpaD1D+vvrcR+gtWXoLu46jjuArYR9UUm/UHjvq4S/OZosVBgW22cSW2
LYN7LgeVW3OQrmSjLk/635Tn283m/bIKFBPBMlVN79e8EMhpB3ACMenRyoQEVfGO1t6NPSAe0Mcq
sOhdX9ThtdRBLYnpwdNpmJrN/yj/QA8zI7hvilIztw3FVCHE+xDb6lNVCuuw1oA/5HaZRQ6Jz66y
qoJiON+nPeVyYSEfTiiZfRiQuIkj3r9oU8opkaDCq50BEIKbFETXP+MZJZRMeOr26Iti/fDvluOF
5Gt/nzKZ0OhHs+M9uHUvX7EgvTp1uRiKLsvJCtsw2RJZbqBwkY4A51MdSG1yYHmO7Y2ZaON4NUw7
IVpSgld845egPI462fp5nO7DsB0mK/B7yqg2cOp3EDhGVLmhFhlYlS/5cKL3v9JA9SG7wvPFR1E+
0naWxn1F5R2Jo+mTuk4s82EMSfFQl9rzSk2Y4DfmNfY/8bHrgD9kjOkdnVurgnGTsVSnMWPQWmSF
7O6E7/Rv2lAiWyynJOYWTeU8ZDQl8F2Px2t2vRe/kBUb0OrOz1TK+XbZNui5BjEUIs0HhA3Nycym
9XBrLm/km98v0vMqd9xFEI3Pr1e90kWyl6gFIrM5c3fcfle5EhvI1ci0M4XF4i1x4IN0YAD/L1cM
H9TEjIt7XBTBzjkFmgfZZ8BAXxHY+6soZquZCy+e5pCToDZVgd5KxmyIWPqNk7v2z6zSLw/CLiSJ
qFFSl17iwHXjAvUAY79sEhHvEdTRzzjW0lJpjwoOMFSPWv24vaphGOJZ3guPax+aGJRchVJysICK
bo5hYwlNv65Fw+nja/ho221X2jRqL8TO5Fun4heSyLYZyd5dvnNIpIvXdB+C6bmamA1cYO1doMot
ydbSLa8Tob3W92fyWWNDRNJ0JkhLwwwZS0T4kPl6IM/azudKx05mhby1wcHjvI9HOnDXsSXjU0w9
jgOdWxtMa92uZpT4CkqAx0+aC2oX8MuoGyKQbvUQNsuzwnHYOc5hXGHCC/MLZEnkcB8vROBeixj6
X901YWgi9abkFDU+ZLUTruDlkM41jgvkDY3Md9q5cRhCcjp2uwrs0qN11GORbzHjLqMmxFqdy5gB
aQItAFo97R37NCe0g8b5zJykS0HgnhS21j2gqYg9hOmHSS1zFDn3J+BNoIDyFwNtPJg8FyXbvGfo
Ieqs6Trj8olQwkS/6XuPucK9cSu6XEyVDSMeSV6y9zPUXCj0C6+9RVu2+YV/zTsgD2mAEPCR+Qok
YA4meyXI8AhCDVv/SmpUDolPBx8EDNmreBDqzI7x5/lECWG5pX3G6hfYYb6+D/E53HdUH71U0Lix
hiCTcSKPT/syipXfOXXqjhlbd4uSdo0E4bpzdeA0P2lgt6rEYiJwNcIHb6cqiLRhh5XvOuegks0B
Lv0btVhjipOm+gKqGCPI+AF9pyT5dmndvt9ywpe/Cq8cuCw5GkQOLX+GC5V6qBE3Zwp/EnwQ3k3m
OpW6zfk8+DVpst0qZEoXcvKepE/wH/cZvaTsd89mBfuOyWddRx8Eg10cJFbK/yB3IeVhP7V6PLpX
phTExIoMkepFJmPXyWVMkj6xO1ngRvjXjYjxs86bh+ADGNAwKSml78Rk6zpT63LszSJBrccMEYtU
6QqQ/3UxTeKr5N+1zIDpxz4XcDINfu5BoB6Ri4NmJtLU4IWLM5YJHVhtweyqb6YUQAErng4aUTcn
/9xq0ZL5DhaRuIFqZvjU/8gppISDN7JaaOL3+5SDN2gEOLsa7lG/YCTz78NSFynB1jySLoCoI5JL
HYqoK7+uKrGaxuQ+e2bKxvGTIhf/4SpMv936VVTQ6jwwwFN/5lov+A7K/7nO8kT3pbuWFbKnEpok
t1GepKM7SQKGBscJVBgwjR4K21ERXg7SDtDGFL1wZ+p4I9OeTfFpo8IhdctWA7ffjxyP1OBHDzRk
nWH/NCZkEHKXo2CbYtUTJjXGyY9AyYXiN0P7rilhYQfBYQzClFTdTyTLTwnb1NHrQOJNTcEjS3r0
hm44Sgu0vOKGzqx/HiJnE0PWEYUgq2imgY5Mj/SFmUSd0dbf67hnHts59aepk3cB8lqzAW9dsHLG
R+JtBCV/KzbZ/ri2ZJ1aEAGwJriJY1KE+g7iiX986Zkd2Qk4go29APXxTqP7NJGjVp8/xqD+Tl0r
EJc/t3NlPDIiNSlJBB15+YoGQpT/BODjwgaUcKtwtFB0PMx4wxxLjjMHtmqkDa+hUBU3VmSDyDt6
J0mJUBeONO5nklWW5Ss2YsSWHf44fxb198RdXavlDpqKK/jquLM6S8TUWVl7sqQBb9g373XqKDUR
YRgD86YHHve42/XR8p+aW+as9de3jC6ZuQbExB16wShHfADm5xwUxPjPkAE0+2Jgc0GoOYtAWmA/
GvloYaViipRRQENPNR/UPtf8hlSZIihWGk7hP46tgGYQCZjQXrWJU4mm+Ulheir6rIrr9JfEIs/O
jyLqQjpOusCyNHrpKCqGckbMM4ArY2egRwv3eP7zV/v+TwfFz7/Dl52b7o7G3YqnK3c8ziaXJBjj
tL1HCUa5qIMdCpQXKy/cPFHQU3LRgvcJIhSiypAWUSHjelA+ThHajMi4tAvdVG66MLqaLUziXS4Q
hETVwJ5JjUCSL3iangXNu5HHVk+SQsLqqODBKTnOZ/yeIlgDY83/6vJP334AoFaJ1ak+mFS5ZkUR
D0J7R2u8lq8GPhK+C4p0s5HDpj97YKNhQhHlGGgkiVcbz6puumYq1t/YlVOsPAG+cy4QP5JB4hOS
mQhI2RINakKrv0YHrWKWgLul4k4lUtk4Xg75NPeuzLC+LHfGoEm/0rVTR0KKKqSrPt4Cjfo6T1pW
Vm/46of9gVhCc/kijXoFX2o6cGf7OvcL1IB+nyJ9C3czFejfKDNlkRo89FKkoI1BkVoG+KGHC2sN
lGj9S4aUNDhxqGLTd5MK3tvfWDRr9Bx3jUKGKMvKFXsZgXsSPDIx1BdZc0qRdsA5o0Dvt/ME5r4u
H0S6Rd6nerMgsqqZ/pkAW7FPobJD0vA4nJEt5K5a9TI5a2SPJojG5hEhzufLBX1ytTJ9j2sUmjSL
mZ4PHDuYDMjFevvQretGH1m8D8OeVKimoXH3vKDUHZq/CUfa8lLtK78cpweU+iJH2Giwre7y/Edj
k0Ls6TwHS+scfU6wZaxshkP/y6jdfmBX5QpYd98SO/hkZXIsaUR7GHJEbK7htkYwprR7YicgRCD+
6O+Zu8f0fHXllUcNqpyAkeByhoRGpdBXN7Q/5Xzq5wbJNkinLeBPSoEQ+iDDSd+a+BzAWNu2NlTY
Oy9QkvAUMRZJL6le4IasAFD7kE/yIJHq1qDzsVP/NvblAFtkvUWv4q0ffOLM4rDByRUNxDF5E81N
wg7AfX8yLVVPdAeWhpXzZldBwh/fdxcRKX97CxOUkAg/zdno/eG1kBJ27zmSckr9UvvZLuSM1UOX
rl9d/8F8BDLAJNTeVKwzrvChZhyw3S7BJA2OZ6aTs7hnkYg24Qv2Jrx3m7upC3oQnlhxR0ga48Ax
JCzCM7D5J/VndpLaJN4kIKdDUB7zlPu+yGRTeeFEP6WKvdlJvjVtY1zmDnBNADWMmZbgA1K8hEr7
SnvJ29PwSPMfLVo6V30mROk576nATwftgxk9Ef7xsZd8GzNSjKXbclm98t1jrZ9fUrch0d7aViSA
VVfJYXURdB6deJmIaVvjCOULlkXmE0akrKT0/zgkG6n2XWmX7RFNTbbX6KGiVJSQFpbSlOBHhusf
rvb0L3HktCSyKSolB6Ck9ZvyXWGjeqnyKVQvR+OZDdjjXEHGsD1vWaMPjTadKrz/LhOxiMkwiFIb
QrhePe2KFyMtOOZhhqj9CSvGbnKq8YDnskQYYiQLdbA0Hv+bf6/xnqKugEqoQ6RqZ72H5NS39Cne
W0hyMouO295B5fqUr6aAmE2FzB4Sg7ywayN24www1ZvpzjKa7V5IhD57fgm0wn+AZsTT1leozGmh
ccq17e4rW9haFE4MYTqiazebWANyyOLgUXZ0cx5svNREc+hx4m4bK675oAIRt5YFpl7kSduymN/a
MHZzNRyqHvQicp4DRB6EcEyPcXUPYOgs4T1HI5ECStIKy5OaIURxfxGf1Mrno40VBB8kg/+nqc53
B5+Ib+onjglnDIXAcdsnOJp9+R8wYl0DYYw08ZTsKfmCrYWTr6RCstWzLM0Hn+Hy1W3uZkrDgjO/
JBVJIX2bXMY/uCjZNTqBNSk6ErBmHYSxKf7x9GxT7v3Z8h78t/sfwDWQSvXyDEQVOTDudYzveUkk
Dq9ssA0azHqDFDRzTiZhFzwcbT4naL687QaLG1ZbDF97k8fC/EjhuqUFgqtFnmTHCRpneo3ZHc1f
QQPoNoAAWJbqZWpLKe71Zlu8495wIT2s1eZUCV2ZIU9PAizMjDVmC2ko3k0ReyqCDggM/7Db2Pp8
H82K/xp0EtfRsRFN9y4QlHQ3WYGOzQ8nLtQuT6LvpXCVJlf01bm0QOTjbCR05mxUugMzv30b0ynm
9d9zDANFKBskIoiZ/WP1c9ChDUUbXAndmkziI/e8Q5dCiqe9tVsRGaOo8Pzrmcd2rmb9ZD4tguaY
vt9LPEkV54lTAdVxMPCAv30Fo4E4uQzI24focfHrdmULVLktEiizYYnDEwEPZ8kxcri7YDmFuLuR
Fo0gBTJtcRGRI6+C96FLI/PrYl67MhqdIhWnmlonQ0FRGhHj9QPApa95/edhtb+DzkkSv7zPyt+Q
4jcUC5FmhvAVqoA8ZhHIM7GT/AaN/HsxCmloTlkJjhHsk9VdmKwoKbDtOmMnZfAdPqVPu/BJ3NOI
1FBb1pXK37IAm3W6kiuCYrZv9z1T3t/oUlMxBg7OYrVMJQqhiZEC764um1IX4nwbVhjLuqSYu8Nb
6QIw4jvcMvrUFWhSi5n+LmWUc6zbTyD654Di5CAtUHfqmZ0ail4PZ6t4GE69Z3MvcCmySboXeuHC
mb94WLoS8RnIeENqURLVEGryY3nzrkYKDAp6EIY4LnbTL2zvoPB1dVR9kImbiUNkDNcVvL6UMJ6U
Vru3gCYqXGxLQWzMr7AP2C2t/be0yzb9gQF2KKnLN+U55vRttdh1dnn76m4fPdzuC4A48Y8bvEY2
/kNo90qItK6k+nVnV7w9I7VNEwDPs42N9tEVdXH39NZCQLoWTW5GY2m9QN7fXkhWu2tq6vfmMFhQ
gb5Ns/fBmakahELMyHTm/K0dQuquYsOFE8LU/Lls1F0mhYKOeBVV9MmPsDJWtwREkYQdOiFMqVX5
mSoBo8lHSmND/m3EYIRYWTsiNu4eQzPGTRODndVnZg11DljY+4vsKsT8CzuqVzkrfdRFwCKMr6If
/LmJ/k7rDVFuczNxynWd59ALdMdPuMoVNMAsaKTtua/NvSV2GAUP7b6fWyOVS4gZ+eMbKMX/ySGo
28nfAZQeQLOm1JdS+Iby7l4z7qm52cA0C2vDitUmAiSmWQx6rCsY4p7+tkySe0geJUiOS9VIPHNF
qBftKgPdmWup6hWVTbZNV8Z1R5bNxPN2iANT9Lr6kPJjMEkb1ocpYvC/kNBpy0Gdj+cXerB+3Z2K
SK3vHsYfWmin4VdfrOKDepvYBQgtFbTGkZSX+b5rTivY4a6yMLZoDCkcrpWn5EwvMQ8KK/J3OPSz
KKe95hovlJX32511q8s5ANa4NcFS9kqVnaXT5vHpfwXUEuwvJXPyqsl/9s/AId3hOySMO0J6ItQv
048UtNBKUtDlw6DEc2NF/dFNjaNcX6FDJZvOHqCR4PJ3nVEqB2ZPHxTUe4tAZPvzNRys2umGqMJ0
HBUrxBTmt506UQhPbMTjP4We3+HG49Pw9WGGG2S/wfd9WEYftkHlgeTMCjh5oxgzIUGNncr8i56j
tvKUcTCOlKsWpeXyQstLD37jd9qaE9QNJ/rRfLb1Y+2BZ+7ZPeAlD4wfgOObIJH8vAKswo+xEY/X
PeWvwV97clqgjZbELrSdPrOzENoRj55s1htYTbq8SKt2gsv/sxT2YjPBUYhnCnlv6d43CkO0AtYb
H9wQfyKovG5ezHWHwrNZOo/nLGBtHsl2GU09u9CPpZ+4HG+aQojl+OtWY6e2XjF/H6xJMUsS7B3z
i1sBv3Mv7/T3Ojdl+d6+whb4dinJgzaAPz8+ZaWbuXRjoRGNNxVEBy+kgGU34pGpICkq9/5oppQt
AbYUS/Z20Fr38fUd6fea/Gc5n/HAa5AjcWEnxbgBiutkSIzGUoEjjt79vmNdycxvpbbtlUor9PaG
XvCiwZUP5m5lTMFJF8nK492BFyt8zZJzGETU6W0ka11TnAU3fxP+YmAUEXebopLXFb8pVKS1GkUQ
zJK5BzzmZcD3Ke1DMp876x3+ZcDXzIZFm2UMR73/i80j+VKPETM+BsQpd/tL7Qf6viVFhPNHt1gK
uBb5u/dz+c/yKUKT7sI+Lbw1JBLoY2jzygLa22B1IbT7/Yffi8PMeXPhyXkAwcGcDLmdSKjd5Q5q
qo0Y5Qnf5bVcqlRRTVuL4DFdMhrdcCVJhwk3hL7l5ZotPfIs2Lkmgw9uKwtF5z2HHErE6NiwGpgI
a7p1+TZ8/DZjIsYGqGWFKcvDMStYgqY6N7Yul9Srk7a0foC87BEqe+sOMhckCmyTR6+ZVuYKQKoR
R1NTNDXijywolRaKjWCSF3OauXXIlchEHg15g/6Ve3z08gvIScRLDHN7J5zggBW4Yyj4zcdH6/5F
1bY5T45J8IfFjsmrojQsoQ6fho3AMhc/shB0YVC+iOikq9WzEmAUlngwwLctqeiALkChFhgQiHJz
6nTfluWMJh+cvrL0YF9GypQmKGtfmV66GE7m4xBGGY+MdS2iI4WG8py08yvfmp3uhrMIIwsVsLMM
cTL9CI1wwxlGpJJr3fE0srOa3ZQ9hQDqZbx3W4RFtcndyiPRWO5AI8aGUWQQOw04dBICunHoQj5B
KctEnLsDvBmkqFcJPc2omMDcIO7RjSXJogqwm2PdJ55rU8ICdRxvnnkzBkMsXF9ORYuFiZf8v12F
2QWyhSWut17iH4f/PqYst4ys/iWflOQrDJrfwGa3ckwlz+0ffXcmmYgT0fEC8ik/hd04QlyooXEv
KGRCqT2coAerIJHBagRQPzpuu2/Pyw5Qa92F6P36bwDDuB/UBlynASCAFEQd0qRqJQcU731dKuGn
x8WPJQjofVJlVrXWZ/SrKjlebbjk/bTApnYmxGIUGHiYm4TLQ/cwtq9McB3fOR1+bOxO6FSAzW3D
Eg1U3VBlAS40VggrZ90AUoLEGJbz1fuXt45qh9Tw7+7xrZPQzKnQP1YH5YcJmHzTI42Giu9WXKPm
JWi4XaYZer+Rm1/bRiVN7Ct1cCxpUPvBduKCS+T6PCKJk1REYgfDsnsUktKitPNgttE/W756s41u
heNi8HMMIztiVvlhJ0xreV/LRyYM3HUlODdCqieK021ZFz1nxZAKqlo1KRAJ91MdccasTFvg2OIG
zdT7IzliSMoAdpHgpFktDgY1c6zz5XEGnka/UFXYwtsG5li0MyBVvAQRiWJ7HGXE4F8SSw1QiaA6
Yv89ZC/M60XCb/uHtHtiJ6c6fjhGolTEOn/qNvmenvbwW/WGUoTsp59NK/GbNmOa8xa6ovKhM9IK
phnHIC9rGw/sfFbGCddFNZEBY2UQnc+IC520qJ15upn4qffOUORPtkussBx5wR7+tLtHMFN+T3N2
k6mNJkZOOVVlzFHdBuuX9hU5oNaK2WusHCRtKiOPvy5P+Hb/VaXY61nRh6c3RR9ucsf63/W+cd5s
nqkcE7L87yGV+s0e6U0nYILmrHPm6cE/ghS81W5dyyejJt8kjMe3fhwc9dWb6Z8Z1pmjC2i5divI
NaGRqSDGcWI0eCNNQOUHioSMNgKCXTzjN46jCbY4IFPd4gCMARSsZel8yF3d8StEothqURpWj6Zg
HPR7GueXUvFc2p5MhbsAcRiJYb2beSqMTJjTDwEtJWOqEQt6TqsycffMohSwlYisaf1Y+cP5M4uo
8ajaZbCFhcBkMQtEitwibdW4hN2lCCertnTmxTS+EzKHbGBL5iRD8r8+KWDPV3WeOZQiYweId3Ge
FgV845ldvjm+8cpYkQOgeZioxx2dWTO96Lr7gebaNU3ccSK7WnRzvWV3A4Ko+8v8yQo5JPYgVw4m
AUpFQz3HuUn8Sc5IhfXUA83mdCQXOyvAinPS96RqmOIx0fglUXh1YGOZVbpbGWkMGmhgAWxfwa1x
JZCnsq4B5aESzHzYoiidV3MA46qTO8TvXcHlQChlPQCzEpy3YZoqL0vIhwJlHZOlPcjdMVeg0ZCx
AAkTzRD3lqjEcXRoNNQwfLbfG74IsBL+0C8XGVqxvYbmubZ0YduXmYkPJjws3lGbkSImTffFlk7n
Pi3+fmoSL5wkFyJYcgot/Ypl/pMiqsJ0xJ8rWKp49DbNm+v+S/OcI+JxspKGDXtDg82Y8jSet6m/
yy1tjNBSbdiDqBWNir//KkeEIKsy7N3cVLpTKq3etubk2YfHhLwSt7Go3Ln7BNm80wStcsIRr5fH
4pP1SDT1jsoEWv1KO/0L8IQjEvMIxTVCq2rrT7dti5y6E5Gyl2wQ3AKhubxINT3yI8owCj111PTE
9no1DY3vbmFX7kj9+UwBlAf7xKcr12hwUJ5d0SV0Z2eAZTuIrwgM3CTdexh4uWH8xfEihJAzbJeZ
jGcRQvMnPygALU1T1tCc2KuVf+8wF2tMRwK+6a7f1/RwZt3KTZRpPzQxCBJmW2HCo9pPDgOwSx8Z
kmVp1mA3VsGo6OQuu8TlrfRnXaMmeJMKG2D5oMC4qSPWfMP4+3Qf/AxIRX8sPrIyh99Ya/MW47XC
GyGDsseBRCxrGJOK2f7IlqFHIdgzpe2smQ779pHWg7u2ZYOjby8W0AT1K4BwVA8z5bfN07SAMObd
ySgi6lojvtXAAYtRx6bv5svypUY+hc08z/R4ctqQ8zQncg7OMK+DitdVA56oiJGRrPkXtMtXNSdT
WEf/Q9wzkkvoQrZSulZ1j4U1SCsLNfKs4oJflDziA5/0/p3fX/xxDNVH75JiL1E8mpY4GY4k7I8u
GOKfGXWwB/9G6LFH/Cv/pKOeILRR3Hd7XN7c+UaVbttj3tx9Kl7bcA/borV1idUbAXfG1D+XL0gI
cgPM9kWJwHh3HEq8Afu3A2VjjyTSACZzT2WiVSiqv6YnhjVWfO4t9+9xrCWg5Bn5lC7p0iuZ9QiY
JFDH2MT5fGKVrHgTt3KVbaoyaH8+kMJjCXXmvrYyNBMEBGtiGICPQsv/JWHxU+oerdqI9kRAH14j
z/ffoWNnNrNENuqhAFjNI08Rt7p7ORiRb8kS82HDDMXXhbxJ8qBITgMOkdL+YtzMSyBYUrIrdBvr
HHAhsJ3l4v5Ju8CJqx3sLkbSNSkFiTkAZsNYpFlSWe+RiDRswhHW//D/RHH1seVb+WYRI/FYPRgV
KlOULvS7JrhF6gsW997FWa8ZY3GOnBX5kNhu+71j4LxbpvF+8I6UwFZuVNe1+ox8w55XHc7Xjlmn
0UziZXBJfk+1UDIwBb4q0Z9mhyzfXEgplIh/nUiF7zb9PLjfk+kSj3p72S8+e2nLzzemXK1ASXmn
jUU/YLM8ee/nUS+wDx9nDX6inY+E3WJp7lr62ok6I7maGBMPmJyz63eL7aMBivY9UFQY15sjgjq8
n7EJb6CLpLTghQHGNe0D5G+73145VlpRKVK/GM1LWOf7pY4rzsWRXiToWsqgbGf/C+sWWUCzoqzq
Fncn3qH+ogVGltU49zOy0060AaGoAYtMZsj514W7IITmfdqL60i0vJAZHiBk+FkTJ5wmXh8Gj7LD
bQOZ5xGPc3hEHkF5PVnjf5GWnKykqxlZt9MHPlm4aAdR7di+ZTQjrYAuhiaVBPi/VXnfmet78Onm
u5MDMqmb/YrCroJJdEyTycJM+Eb5CMU6hPUkWf5fytoXj0Djk5eCA2zDg+4oFxY98yOpSF6d50EX
76rdLa1ZhOwxEwrVyO/UhIqVEGxr7agJsT/q4nbxChZIZHEQ1W9AxgkrhZi0sizr1AHUtuj7fuYb
4JD48pkjRTcDPxXdjQ2aE3lgckr2Iep+TsgeXgbmJyPDZbgISyy0h1fXds9y/QUS0oRrsG0/F5X+
0BLTFRqz1ockxqFPZeOZJVtNhdBn1qNRF5mwhxBh6xonsdnUdHRQzEjtQQ4YuhjQ8wTs0u5U4v8h
knMb+5pG0u5J4Qoz4PI2s3hdTDC/0KC0ZFUf242ifXWE/KPlaCMzcQySTYOyrJ9KSUaQAk7+9ECE
sl09DtqaJsgwZN6Jedf/dfM+aBwo4EsWhxiA/3JXcUgD7Wd4xQOF+rvXqEzxtqidzN8X26nldLJM
WKPvhhi2s5ysNWfNmzU2LbQ7Wyld6v7+yJeUhVrBcaxPZDz2K67DfyvNd8XUcq7IvrEmZoWNtACY
Zdvj1RY5nZfObl6FpQCUI8aXBLFzJp3ZQaL3uzRWoblf1AwzbIH8abWYpJJH9WaY50fvyqjRLoxp
nUlBM+SZSpKYvFyE0d6Wn1XKvgVaZesPTqfo7ULl+zVIix5HK0CYy631qEUayR2J+jycMTHmWLUC
pEDMzn+eBoHjoqLqq9ZUU1craPlbXvP8QOWtKN6zAxNm7rl9r5DX+KcP5tRMIldVdudzXUUPJ/Zt
LiGsU7LEnub9zScO6BGmyuGrUuEzw+NuxC26OMzyBuhc8/YNfumJOh16B+NFBAGEJArgygwuQNLQ
eCpVkREPO+YlgRCBro8UUthNlMR27WKgXyLwDOhJEb2kOqGnrnHZiBbhfgZKtq1mul7ZUo2TYMyd
z/tysBlclDr6aO5pOV16okns7cK9ychC23w5gXKQ8tbgia4Ne/2TjHpky5VzfYi07V1ntI19bFn4
g9MAbN96PEsjeHQJ2b5W++ODBARQN0Ywyc39G+tWDoonjIFzcrmgk/Gk7b8c4T8fDrFClFqUO9Hj
OwbbcETQNZEZEPnHKb3gsx+U+5lZ4m2Vz5ib3JKMsq6vQnIKG7Xw6erlIRbfd+sdLAh2Cz7x711v
6P2dCzUynGC+K/fN6cXcP70CBVI8xgHPGf5UPMpzSIgf3p+fg14TMcYjKQbpyq2s637U9UlMci+g
Z7zS/xrQ7IILj7F7vJmuWpeNzmHUyOzRlwjt1MQVNjQwGBoyDrDo6V3klIY/P8z4jDgoSTQIgO//
+hEiN6E6t/aX0PjnKKYkZx4jjeqTrTzbcwLOyAskN77o9u5UPw1/MEoNm8bCsxycyXYb/TefL/39
jHA6jFoYUlDbhahnRGulnm3a7NWML/BTgkHN/oK4fWxalaXD5ccwG38K6LaREC5Bcvx1dUQtx7Ef
84WDr35Ph+Chejsj3Vbd0gU7Q0X8gmFzon5Zrdbrq0C2Ky2iOOy29Ka/FNsU8MrQphk0zrD//jWS
X6JDjFGN+R6Vca/Cuwg8BJMuJ/YWUxSnHuI4Avgvoo7FvXGRF+LRl+pk9uPBcUODjDz7h/f6tvk1
FMo/B+HM8cXWN+UT01a0jLIrzyOerX7pj2vN7Im7QXJQnDPx/1gwSWXeZc3u3l9FniGOUka0CDbb
DsZMCJawAgwrWpNOwXD4IiY7B0Rr4aTCdvoHxAplHhczvVP5L6zhSV5lUFvSoLVNzQ/ARnTq8QOt
rp/Wi+B/IFpMxdzZQBxwV7VPAz6mlXY6y/e7Vr03r6RhUmDSUSau9mU0x52sAw1z/PrBSm//XetQ
ZMIt8FMOPPOBpS2+CuL6j/u3KRNMn8hikOcK+sx/5A0ypmma6E7B11kXhbW8UEYPMPfOyKfavZ9K
nvHZPbhgxIiyFToif1uYksdzO6jXmtSFgSTwbDvrlW0z6Ln8EmcSmgaWVMfFysUDSZ4D4A9x4tIV
fIfq/E43OOgUP3R1JO0TeuqxAJMFnXqegIlmex+k746SRJclCavEpbqhnncq+CKU5XGzAlwejWlN
vXKrd8JGdadnFpy+TTjGltg0k2mcQu8ZTwqWnZ3Rb0O2nNPTbcCpX/XG/mHxl5U0Dkcc1DbqmYis
bDuwxCAJkFkLLaiwOj7cBsjeg37v/0Df8aMRb/c2fLDTGTaNwPbCgiJFaUglu4mZBb0QPot2eBrS
EXdBs0Z/qju3eElOC/AbKOyyMBB/STIbuzFA8ZQt23jue9GhTzPWbD3cKgML+xGKweRj82GMRJ+q
qs49m4LDue4yDeaKzTGQm6SAba9KgTHpTOhRI8+n6SIVGBFHWv2imhJ/xJJM9e++Z9umndjHPBDE
Es6ne3KbHzpMuLZN42cBOratBpEv01XCelN+SXaCLd4qXD9kXg9l8/FQODIbNO+Fh+wFrkQ20Vm5
v0USDVTdss7O7UGGbfa26FOSgFK4Zy+lntqbxU88BsRL8OlpuOXD5TeKPNQ6rQxdMCKBOLIP3bCq
F+vGef9dcUGYP3roOFKGRNapnKGnwiMyo/ge9oBwiHIKun6wuIkXgB65c0lQ7G7X0kOMebNy09J4
XUjPYXogr3LRjgXr3Zd2NyMxrtO+g28Huw0IYUFX1EX/Q0/ZL/MgI/ZS9oadl80vOseNnXRZptcK
FgnCK5ciODUMR2O3dFs4P/9JrzYxDK6Jh5vE1EoCMG3maN50gWySXKZPQFCYc83WVz6qKp0v034M
eZkjdevFQz9tQQeHthQWuJnxfKFuEkn0E8SqbQ1wNuH2r4w4lyQX4UMqshu2LvM6fdertr/Yy+Xk
kmTqrB+CoAYdok15mDjJgfznIXOnbbBD8hX3LmX5ZVPsgTwD65HjjoeyfKaxkPjcurHkXJwtJuQS
f3+Cgh9HFPcvROQ4KIDt1NpxGjSHl+cGBqeicvOSI966BhHovsqiXaR0P8cDe/xLe1qgs+aNcuf3
Fwhp4sL7t1ozahufNJX1+C37wHTpF4fx1+v6nbZbv0uaSZF82nwaH4Yxj5v5r8AdTAYef3M4/OyW
Idqj6wyUhmKPU43LUOxbVhG25Lj1/SYqTanVc8jDUU0Nc7XZ+1v/XTVfSlzQXM5KQoyl4430VeDB
sh2jfQYfJnrlp2265aNFqqzY5H9rjpTlPUiCnfI5/bgGoawRjmeZdHBDfsli/DB1JhTUZN/sqwDx
fE/eRGm90aohVOSjoT/pUmleFeEsKffslVMMqZfr4L6udcisUE80CCoEsdCeU61PeoByfd3gG6aT
As+HAhbpsXzYTgQ4BL1sYT7z+JJl0N8xXcZD8+5taglOos0qEaEokLhhAneZ4lizOtV2OoTQpl8D
E+bsY1X8B22a5KrfcSC2hATDh1dTq6d34fTJ5U/+zSxBH1/90bpKWOuGpb6ERSnQPxcIwXtdIoY8
MgFk6AJjDoPebfiuTREuQx9O4adHjsVuOlMAKPWjF7wSJoFVNQ0Tj8ffUhFyq2MQmBVuXW49LSq8
LtKun62PP576XWJoDpERvvbhO+Yo+LXoAzaNZWmmYzG/HIRKS/YeNoMwBbMWlu4yjavZoswqsVj/
/zyhSzW64Hgx7ai5SnEcONONdE1bJxp3YAUjIk7Qu/kFUI2i04mnFxbBUAqgAfbdiHJ+2uP7mhJX
gkHslcvgdp5vvC1/GvdNNIQipdFnh9NNT8CQCGhS9GxeAHA/nNr39SBI8CmHfXeYH8jWvx/eC/6j
INbTCSjQ9AwB/UiMKO87kzmkb4mlx4B3Jqk9D1CYYiZUzMq6vj/7LMqfPCkJV1++NjJAmLNqeYhk
4Pg59ho44WA2+2j5WL3MWmZXmXFBVk0febNbXtYwDA7KL5voAc6Q0Ti+HXHmsY7b3wjfwrlUDMxj
W4O9mBt53+HK2eJX8XRDGJPJd2ovstZPahKXc+tLwS1aEQEj8hGj7Ywhlp6h3F1DSdUvF8vRbtPU
IFF+YujJWYtmf/5DyVZK5+s8w/uvhKko9Hkxm+opXUe02ApHEcsOzg7Tn4v/QEtviprhxLKYhJ+h
ELYvgGdJkTCHav7YM+51EF5Ukmd9FSWqagCWSlN8r6ZiBBStD7lVw9F0D4a4x336Vmjkm8lYu5Te
8Y8M9DML3aES4ing46v2yN3MyJTfk3A6iT1pjhCr2cPfW4FFpZMCvIs9JwEjre6KVZFn3MiZsoU6
qcoSjDtkmDbnHZfEusrUw+eGaeFJb+FEsuLh13AtPuXyPpWZux4UUwVFvSMj+MtaunH8wCRkDniM
mJHydXGQsUwnfcF/DC9N7xS4de8TxeMuRV5vv1s2kwTANcl6IxryFeUyZntWKcFyKgME+iA5QT1K
rmRbPi4pEU3Qz4WNhi/AED04cKXZOjA24vRD6tkFSzOWYRzoW+priVRIDekD3mCdi1hzMtxnnUjo
purmIvDbcVrLjpEqdtLT5qMInGjVZwi8en6kqBAXgtl1dkAobZG6k6vUFcBJjUuvLOhZ6BAKpxAg
YT0L+gW+ruAGOQNNxtv8HqKFLEeBRa2ONxo++fX8wTyUERrk9YUs+764Y08ot00Cd7uIk5OFmQxF
jg45VVj/xLMQc3EqHE5XTYXHe3k5177cD+n7xM+6oEBKSBWfPzaci8+646PzFmWfn9R1bJkiKK6t
3o+jEhk0qFeuXK8t0HJRimeV9j/g31ajlIriUU8rGp43NXknjpq4VhpXdMQ19WVji7ZF2D0XsOl0
0wPX6ssb4ZC6APvbNA86qXZkTQLI4II8IPtkzyXS2H/Onz8ahZq0l6akRLQXCnWpUK2aXpyXYsvs
e7khQyi89W66LMM/U+Y0PrmIa720R/AKJJomavDnJS430ATpdWJPIaLR1X9xU7Y9O3RcHHtioOjr
GEkdeM8b4ndCCLnV1fGc11pFwcYrHcUtNjC5FRX5ZHqIO9ogoKh9MJ6Tu0aKe1zxWLPmpveHmT2X
gwvm6OaRMKdZb0vS9pijCrJ/Zb9NUtB+c8fqesalgR5aYDR34y9cSp0y0nzxgjdqT0zEH88kA8cc
N5/LQtL5ewe01laRD2R9wlq+F1W7qoWFEn6998KdIBZ+baW3+wPsMuUwgUO5+hmsCr7nkuTSMMVW
k4re9i1QzLdRH2oD1CqQjwcGdESnqtHZcFiaW1eaAdS6ceQh2pfa/Wt1cLqYfE3J4ugiGNR67HdK
jT63WPwJ5zSgRh6FF523r1Y27PsyXqsT1WZjvrTO8qwQBsPNjftbUiUCL5OkGON7v4g6kfI06uK1
T8drxm9PpcVpaR5bJ6jwIhh+6gBlPvpicE8U5qB5MHv8yQ2fWBpL37403VZkhyXya5S8qQR6hHTg
qGK8HFkIOxX3N1QIuo7CAPsJijwsD7jqBpMWMveVXuV97oqvTwCLWHyqTHJVICJL2OmcQsEiqI6o
9Zieojxi5t58gBg1oHJ9razH+aXLo0dd2g3hbzWae4k1LP0VMDoZdv/p8qt0MOBJYu4ypQUmYm/c
QTG6PjZQ/ghTA231aARgSdZhnOjVCpocNHFzLe4QouNI0trYjq8qseEKEBiYnl2x5HYX6nJ9EJzp
U8hTFUwyqHXpZDIPv1zeyLb33KhNEZ6x/vdFKmQawfK5TSi3i+KUAW1pRmi0KFLYd7jIzftJ2Yjn
FWFYM1214taokJbdLIeEdOy035xYtP7jQKgm8ljRFlK9/NhrEdW9kM+BgcEvkWYDl06Q1u0787Bg
KsNr+es7Zx+3lNGMyysphpiDLTDAFIx0OtIVj1WKQZZGO+U2AEkR5rfnZ24CLR/r1B3+7YxLpocn
5zSalIVY2RNTsphHmmrgNXqVNH4FUxTK0tcQflBpC3Bum6/F/pgBrmOmG9lTHY+dNTc96hl3yec/
dKyEqn+m8ArOUbuJwamR7ZldV2mXqOKX+6s4ICu9DbnTglUJzqQosBP3GSQG1TwIMjeEClrhIoHA
7DstqCxqFJ6NNj/OqQLQHPSPSWNIj5X/XEZxs9nVa+pqCd8QJVpwB5Z1hGOnbNc1+QZplPK09x8h
9nzfzHwZCLX5QVi53dhh8lfx56wlvBQWmw/q+GJwfHDg44Zwd3sl2KkIvsqoiOci/CMg7Dq9fICO
uZyIBSAFuAL/hyI0bmqsWFKR2buIphvqXnAJNERRfXlmHZhRS39PpBPdAhGjnJwYAOKo/+buCUEI
QB62LP3eRW8H8gPJZcbDG8/s0P7Hu0P7LhMfjZA6vyDdD+7qleIyfw3Kv+GENeKmg5ZZFUyPjioW
o1m+jxz33aGsZjQrGYls1izXxsnz1Jp9RLHyQg78cZY05NAotvxaEq3+anpJOH+l5KoGgkRoZLiJ
ofwCrp1awQXmqDUGAjKk2peVvlcK5DVJRVKeIRc+31HOI+tUppXRN8PEans6gUEoPLIAp0oSlMjS
PMkZ/CunH3BHmR7a9DxXpUFmSzTjM2ikdDtEYpseVO+pmhMyPz2TzRscnRCJllv9S/KEZ/AEMr73
M3tcFjFot3+2/b7UOwodcqD1n3AxVpUnmr+latusAg/ejiYEQ7b+cpmt9mfiWIn0BRXz+m1/E7/W
Ip2jrEKokMWbx98v/97r8AucvorBpSfb1PasWaDK0RssWii7NLmO67ck4sEhGmsCCLdgmx+KYJuR
WWBB6isVigte6kyV/20n/g5npBHVDW7b/IrcTQoS0ZdOlMGOEsmb9XkgoYqNwZUZWaaiMaS0OF5z
LDbKNrw1I2eo3g/d8ZMllO48lwZF1sw3fszZwYi1SwaipcyOOM6dT7N2zZ/SliAXZwYKQwJvDx35
90LA4sv2yKftg8trM3/eEZYEgoLhjAt0odl00Xc9uSlcZRSM7kItY9X6fX4l5rS7+KkvLvr8mo6e
STOfpHJdeO3TbCNho7Q/YxX6Zfmtdg+RmrF4sb2KekvAZW3MiZdHvi6SfgSDh8UoTlkeTR1mcQDk
Rkpw7U+NznbRwysuqq3aert2n8ZHducxKdXQiW47nBTE+Qpn88mJZ5DwE1r9RbRKQeqrqRW5a1xr
h6KFcUWvlNXIGQEzWLHOh07hHJX58Ixq0XoKmAnRUFO/8G3c2ITptbMMtZI1uEK4Oe2wdDqEuxOg
z5lS0V4LG8ZDTxOt7qhvuKbzC7myY4h5rvbfuTHECmovqZvq9UdXbkt7Ymn3QjSIVSIDKHQys5vy
mCctViES8kQMbkIGnAU3N/3q2Ks+ivA4tjWx3pkFAWgBzQoBIzSDLTeJGj3H6fN9lv799YtUq522
QoDQhbIQcDflGOvLUAKFv/m6SJWRi6dDTtAE7HZkEoyZqceL0tfbc0kjYjdnfvkx4YvJUuiOublz
ERUwYdwluWF/2QxQu6r/Ql7fMTJRXD9NL2TLPc+v+NEZJDqaV3fb+w3+b05OGtbuuk8Z5owLbFyY
j8FN9q9kAiyCCsueMY+kR+wY9gQ6QqzvQdZgZB2FVhYM7X0gmejm1l4CmsnOQGXiQKdGTQast34O
emNcq2qHHWEni6eLYnZmvKgCKnR/jsbAsa+H+/ZrJcu4HB2HaOUbscZmLTs+3iZyqlbieIz9+zw9
OFV/5kIrweqZ2T1nB+pky+mBRRfmlFfJMTQ2wWS4ylnqmsRsZs78VoB4s1qbeBfnmg5RG7bLzo/G
wOXu+7bVqH4i5/dFgeo1o3ggtKxYVZYUZAD+bZdy2sEJcGQ/AUTkJWf/qUtZ8qYp7AqfRqNr3G4Q
X4kK/hhhY9H8z4T4JL681yp6P09DZ7lUCpkNXzUVrry7zBPuEpLPRI3Kt5tGi4RRpAsmrwogkGS4
+YNKgPG8KlksmRamBnFAnIXEDJvmLdLD2+6jSHz97sN5jq89NSPOPBO/Hyz4w7bx69bmNOZnCJfG
yRjE2y9JXwa1Mt1RGzgW3xN78EnShNhSX9VWAs1YU5lRPSMqPnaC5k3Eu+UL19DYszPicvS35ZLC
gOt1W9KJnG3yBACmUJynU6Lf7ZDUrZAe5r6ALy3IKIzKuViUCyIKZzjEFqfsvBeplAA3h3GQJ1PQ
OGVYD7DHpGUBxbsegDNPA6p9XJooWRZDKLFP2NVlIJkb0a5pIj3mRqLPXI5V9/TGnxW7UF80B6OP
nEt1iHpGlC2Q+HkRgsU+iB+PodAFk0ydqfdb6lkZ8l/u0fKxf2mW7/NDNq6pfYUrB4YeKZ8EwSTw
DNKc/zXKJdz3iTZ8Z++lzXw2q4NskVqdg8UKwT6o6atF3LbicXQIwe5JPe/JzwPgGkTq7u2vBYw9
4ET8ExB5JedI3aiOu0EatYKsOObCbNNEqzz6TbEJ0G4JhqYt8wJvKhDQBZsP4K4U7xKpxmt56RNR
Gq2b9CJDpm3VH9JPhjnFkOtvtGSog6O3kZ0Dzv/3s5Y3q2ZhQADDMVzenhg414ZO8JiPwXwVy6Nd
sP9a7iGPAk6uCl6ZZj8xtqoDWuvZje5Z/UJf1AC2ZYTnJHZC5MCOZCDmG88VwCPpC2q6ytipuGS3
SJCScJ6/JVLa+zzvmCxNUCey0o63Z3gOEvbdRwzzll95XE5IljaW9iuJmJJIpXeVSrRNYg5IiRKf
Xsgoe7LVtPQf5EzDQBhnfJDvkRpDeoTYue88qaC8X2EGCVzCrKGjcPOYWwn0jDhc5rOtqDisbf0/
MS6zCCoybkNXYjovmTqHkySheGj1z9OIEAAfPOovEfkF7ez6GRvU4C1T6jSpeHqE05pcvzWxmf21
mnxV4mxuimEHnwVk9wy0jjRaxykNxHc/ERmvdsuDsE6vVttRNp6ISapdwsKyEMSkAoANVzdxH3HO
TzdhK5p3eU5OdUdN1zv+xLmgtI4fLNWlmyA61EjdUx1klyDVpD1018siE0YljYdWqWkx2ecd+9nX
1pWmlNFtEPZwnH1Oq4CLYwQSkz6NIYXqmVaeX9ppSUJ9MH5/WefKzA+t3YJSqY66OAVEsEHntzrG
5nUgyP47kz6zVF3slu5RLzcsQYUhHui51u+GQ8i5BOipQfgTKlJc/UDjKj8/RowA8EVjdFTADgqQ
W9hjnqvMqNTKVwW0j2HSHTe25Ja9wkxsDAl7B3WQ+/vfzgwO2ApdxsECIrM9fBVdD6ceuXewUTF8
Lj+ROKLsKhLKm5VhJpeN7EveuqsM26KWu0SYGMNuSgjBX8pzCEVhgM7Ww7sSS7bQQd/CExZaTJ0j
5Bqf0+npEadkFu6nMOJSQMKBBIVKnJkdnIpk6uBVZxesVyxnaXycLErs51zsh5X5Y4mkHot7gJ0T
bxYQdPS1S7PmSNcSRskygcmTyO9Sof/S9I93tvSbqcQNxr0NvDQBJtm/8s9DHMyc4Hl2MRJAaPXI
OmYw1Q1hq2iTi4ibSH+txgFEuBaRlj8WgBJskA68C7hdO3pzWSMW/3SbkOFXC+PBIcSwpFm2m1Ef
um/EAEgM49Opfiqr5SsK1ntim+RHwrpHtT0+1oP+dYkWIj17YPU1QV9xPvi+f//Avc2dyMF0AbXQ
FWCAHqqCbhl5yi7/RFgzhA5XPvX3TLb9liSsmrYhhUO5IzVHxjfLMrfzRehbGwcND8ZoFQB7INQC
njqVrPEa+xOGhpW/jwKvgFxS4btrtWRY9DjlqLnUiQ4Ffmv/D4QAq6wpvFlEqGUoyt/5fwv7xowP
5WxFzxP17LE7c72rsJtdLbox0Rf9Pj8Fry1MCfuHdNKsm2n7d9ta14dzbW0kNWy16ERoPCn0B0Gi
XmKLM64lc87902XTbffxwt3mFguhnyzDBUI3HmqEiOr6b1e1NcncBxUmLuoA0GC4Ja7rjiXXWTZb
5Z9f+o1OsBGECFMFmxML2648cXCvGj/E1oFVreXrsFKWPJWdQR3+6ytwk+yX1/8r2bLCJuQY6HDD
ZcAizDH/fLB+WMx/WM9+Z5kcslMhGxB7LCmJX2mWVig58ugiQBbKh1XRqp221ldLqbNGlgW76JSF
VPxcZxhircl0rtom0wJfE4c0CM7P2Bo0IZABfsnpgIu0I04+OlCF7kQQj+09qtpa/JzELkI+5Ca1
kmcLm5WDMC1AK3/nHGDMiVHugsHF6aR29FnhabneUWrrh8ZAHo71Y15utt8IooZGl3nuoHfKTLL9
MSDa8B9rH1jOFKPe/1rJd+mlSfvH70GCBn2lCNnf/63Sl9RTHRzWZqV92iAWbwbgK+VwmN6qFp2b
90Ut/lhSvyWWud8Qu2uW9di0fZkMrJ5cdZzYOe1jZ+ELBAyY4TQzhYJsKp01LZGPiGf6B5xgmo+S
0aNsJuszJjr/AdwWRcIr0SUBWTPfo7Df0p0hOCVfIb+uB+Zm0674vykk/bqZmvr5EkrFrBI94fRG
u/Eixs67QGaoZJV9gVbYyTF11/R8+rA/OyMUFQfk490tcLuZO3FtEiN7gRlyFPPJP9V09iGnf9fb
bDRO4lxTAJOLifdxx5lAiDjJWEM59FuAzeDYDDWV1phUujJaGhlV9BtyqTj1SxTmZyKpJ176rqSS
oiXJRWrFx7mlLTAlwHrQoZcPtvkNarC66fnrknZNSzy99mhVbLFv0OjxRP5KfVUkuKu6I6FiWIFv
s/BKNsRZVLJq9Dvi8BxeKzdoWSaBLc6WJf2bAD+2duKXGrGzvrjtmP/njk1wPusMqIRYDOXB0CWm
DsKvEd7clWgjq4rq8miw4b2IfueETtOB8B98a/xCpWlIX2m6Tc+WLW3ukxaS+teEgFh/0jo+3u2D
8hI+r6gmsRRdyHQ1ew44WuuDgUd5YSsTZ9GWBiJY3NwehiczvchtZ7hfjtPpQGNFe83yMpAjqPZL
Z8y/5z+9w9U8PjZEQjzDlHd8mWhXszqePD+JL/uLqClUrMVWvF3zze9SfmjJUOhVqiIB9PYZzg8L
upnNansXWu7eOHMxfk3EMirAL9Bv/1zxfEGO8ckp8ASLSBYFoKk3QhEwjyQpTncqST1JHrVcC28i
nzYZmasBkWCTZR54pZ98fRnz0UMT1yg8O2GpHmJffB53+HnZrmRrreeOEdnq8u7GdRDSzuZ2fT5J
hQUbLHEJ61wnBUDfaVqKD0IKjL9qXk+XL9dnS1Kz5MK4P5IRWDEQqNYWZDdSnG4YjUGByJ4XW0OQ
A85jTZE+mB1IAqwBkFkUCZ+CCyR+WIjf/Kk0dLrbGQVpP1Kl6n9LUUD98hrlt+0fXD9uILjWnd9z
eMxyKRWbqp6qg0yTaS0zn1LNz8biGon++6isBlXFbbFFDo6yGjLr7+kKSA/zmWAJ0WhczUlyPs6J
eNs5vl0vHQdA7G5J2bVqeMzhHEbD1yaVXjLkGkU3LboLBDzKIsBd8DsA/t30/9ceWRP4PqjAso4p
BVqVbA5xFlmNf2YALPZDI0hVS+oxISuq3pkNXoN96lS9zO1lvL/G83yz2E+jDmn99ksxx5rR6wkR
urgRtnSEX2CSUci/3OUx8lEaEc34VKZAVLTbcCdl2iJuw775EF/1wu0+3neaB3rPnyXo6b6Jjlk8
Xl5BctNbuMVg3CfSyqahDqKR5ydQPSRDmKC/E641kLpbdvZ5x9Qnedwyx9EIa4Brn5E5hGsHZUSD
nf42C5JhYxVP33qJgcAYQaS5saYhmIiJoz8Nnv8AlUzohCrlq7lyLH40xqp7M0+uIc5bJYH9J7TM
41TC4n6MLKwXUj/TSFc6N9um10lwL8Wc5oQHOd0ErPJfdKG5uAnfBX+SHeRQbAfvGJ3tDyOTda7K
n8cXzq2rCGxIS+h5hj2pLY/xB4pvrEdIU33Sv4ZBfC2iU2es/cRlWlHK7UdZfArozeS2J9Et16Vq
LjcXSZlB9j9J/v2JGTt1b+GYkharoXomjVIRn5NV2F52RkNXxiqYeLor7Ur9vl3DwN8tTxp/tOLB
NBt23mDwPwr/B4wskSWcTDdqDeHvMHYfKvtLHQo5kocoIVsjDmX9VZno8RGyvccH0WyBmUe3ZpCO
0vlwcf/DPHdoa54x/oiRMhTi44vFnNi8H9RgAa+acreqbp90mLYtZ06KR9ZcLz5ad9WpHSKjl+Yo
tV4y0eP0bBLFr9KRXKnBwE8WzoT+0Vthr0z4YSamjmMQKipDyM+623vu3+LCs32CXKSBvYGU//Xl
TWKHzDBssrvhLSh6AzSSjenxpPZ6CRPlAW2GHgXWdLCE6ZcBeZ7qkQcSn4wIsTeeS8qRa0C8zDZW
ouqHsda2mYi0JHZkuzWj2Z10lAfrzUEAD3a8kaLAc0qEoodu0Zx1UEaK4gAdKhfVsHhS5WpjtfNK
T89pqvWEB+8SRxqVr4cOlScXN9tcEZPEamm0+8qM88kGJ6HPi2uVW2ILatojYKHBvfKXproF5C/n
q8rK4sIYdEfnAKHevqGP88gn0UPsewTNYyl4vL3sGPeLoTXHAQnSK3rthhACrnn87qj0uNhVUyab
wALmFYb28jqJXY4vB1dyaFP60DCgxYbjkQRMMMU0TDPKZ1dIIVqLQJDylQUGhOhPNOhtjKEhs6TE
E3YmxWps6TFc2BXLLl5P3fvqKRaJMXc8WPeFFGu9VTm76k8kCs5fs/V3gtIcjcLZul4gE5W/ZEa7
KxWmZGr1/xP0KhGCXk4p59rs1osnKKJY54OBzTFA9z9Tcs2+iu07LwLbQE63Akm7WCo2rjEB3h1Q
4ZRrrISrL4qLUqS04BSbX6awl/2252zEoCxtjo5OBsC8js5xEtaiQe3Az22sdF6mpdwDV3fMFnRU
kVoRSLMR4QlZQkxRmqClynnYaEwT19+mjdM4iWhYF9cPoDelAur1ZLIwvRDZXBZ3TZ34zPhwXsXC
gMgiVAhnq41Nhfes9MNgp4qj4dM+D3LHRYF86d/D87Db/xhTPLbX/LqSpaDNgFvKKX7NXRBPrkFb
I0UUSLj0SheIxUiBpn5pjc5qFLHBbEZTIlz8KMQ8tAouZJF3+gX/95XvzEj9H1lhEs9njH2bAQsq
RiY5M9I0WStgjNu+xPYoD7TQ4FwHPc3H9az/fX6GOh8Juws1NOqNITclhb1FLbTBpLNMQyi1mtHz
U0WN7uBTLNFC21Eps1X+V5SjV9qnM2DxO0lleMsc7PjJt/PYwtB7I0dPOTJgN6o9+7inFuIbR+wG
jBOyf3uM2OAIFGflAT/eYCoK9k8Lh89Oze1P0mSLIj52Qj8ayIdTx1R5NQfp4PdKboKKdx+G5NrN
t4bV+gQCUGWBD+d8SsQWkke4yDdAMSC5Pdv0XJE1hAFC6KHDMa93QRlzHvQv2nX3WGRPMNElwt3f
EjpGlPxhfMFk+qycma1VJQrbSYwEGhv5RdBnk2Xw37fTTZeMAKEHbwMDqKV66wqNyX1W/mXF62Aq
lywoLoTSb9CHNz447QlBNVg3WTKRMRUHCwwiaCQrq0I/mP9Z1LfD5kMSymNdasfklx3HXHOM0NVH
Yo+1U75dtDG8Y9zPCYV/by1rTb14a+fEm0xvF8l6oIUPP/rrMfYtp/RbWOpP2fbqy+yTGBs3PXSv
QMLaoDKBYHWDdBb52JXiUqe2Gng5gn9tgAyrKEw5hrFhhG6Xgbb66KT9r13b9mctqlDD1ph706sT
+ydX/Eivkps+hYiXJ3b4S0YsbwOpSxGmU+v/KaSt8ZV/CtYuXZyystGzcWVaOCI9/PnVZQ/3svru
ghCCF471B5NERdl4u4ljWOzD+PKbBWGSGspfjDcH+eqjP75spPEt/F4GqRVWYhkIcvIkyEa3D6PD
nV9jky+hltnWpXZQRR7PemfpjCwAyIdeKWGrisDODySqcCZB5IWahNAiU/ca2/W8H8wqtMT44mW4
SXzbOVdhPrR6eH1T9HrFbrO5EpS1n7u/GMbJ6raNLVSYZRIjCdufuN0gARHu4ok6uDLDyXdbRk0K
BzLTgbKlIrIrBOs39cdMbBqt1B1RbMQKHbUVSJ5RKjWvV4CKxtHyTqKC8vV4WxHQHWyF5TXxGCLV
+I6qct9c5Zq7NOENIywlq3psqrZ05lnPIYTDeOw9f175XQROmQFwckf75Vdh6t1ir1HEzUZEkq1G
eqvu+8sKonIK6ca0cNbeZTEWb+dBl5Y0A8tgdQgjN/l7OKafBIArW6ALkQbdgmdX5By65ioWqPRM
FY1hFwXTf6LISN6x0jhxAn9PjZgXPsIZ9Pt2nqai7hbO7/g2Fg00GzI9pSm6uqifx6bHaryA1t8C
hpa21LIaDU8E8xwAEAhszO/sjJIL/X30MiJIC2ZvrIS4hWczqNNSQvPoE8mRV3DVGDLdP4FO414y
Vy0e72a1BDnxubdKaD4Wer2js/H980fQlktc002uXbpZhJcrvgmv2F/+oW9iFPdf9WZo9XxZtdgP
JkGsgaAFupXeMgtoIzkSiPzpmtP/x/n3w27Q3rrhtbfos8FI515HDgJcxgZDFL64cozHrfHrbE3A
s8l+K5Iikp3oxbGEwNdOluf4vdreMJCJEKmtvsAMvQ73ITiHQCKLr+Krhf++VopdJD868OUL1Npm
REZs+aZ9/0TlQ7qxCS6t4VhjYsOt4ZjvGJJv69kZwANI1jL62+BO0gTLIX8rdTmmD2OE3SSY8unl
i9R83KGyWutw6i6Gr1rQFvJwqYkGO9c1UajWooSSbNHQi2QzU1e/6c3sqWIynfb6sxomIhevoNLE
VJ0QV8PtZ4Se3YYsCRIRiChzUS3iECzRyEh69XSTDAKemtQt3giKJEyg18NDsfxTBAAOsG4wBEDA
9/54PK2uTqsZP58b+1YYUjWAnE8+w7bc8vx7Nzkvdu0uHPVXLiQnp+zj6hostACqDkF2Dyk+DDYO
Rhk6ktefNuKW1sWz1lUZDx/F7bPSI+Bl/z3MeHhP6g7humMueI0t5RcN3Hak/raVmDkX7P7VnTTH
lv2DXUdDrzveRlCFiITSiW8t0ZTuYpe0gUMSo1EsXTUGlaEzgAInnmvRpUMwa/YV8vFLU4qI2jVt
5X0H4uBXeHmMskR40tVayoSZeT297haVCSVcI/9dwzCr4Flzy3BVMDDNP4LIXdx1diQwfcve3Hi5
EmOTlaWWNL++6KhhvDezaf3BGu/Dj7dCKDThHxSqBBRAdJ2+o5/9UiKo+sKStUASJeS32jY/v3cp
9Lq4X47kWMDkeANgwd16jTzhQuNKj+I8CvibdP7hjZxoDjm0WHNShMOwmT1CwaH2rNmBCpc6GfIV
tjC5qoq2tB0HDiFuxdDhvzJFbCJ1xFhj3gs76RpqXpRUwKI2+O186KHj+FnX4VqWpvDemAAVSzpV
TOZCXPWpqAUpzxdi+xMO/axRKrqGeT1f67oCemKba/RxYWC25dTGKd272557QHHuB45fOQ2otAsj
pDuffASs5/wx27gQko1KLEdf4rVIhSu/qyNOdjndkzyc3VZl6fazuDSwXagbBKAjYgNyZEfX98b4
vinqgy5mf6l34Vhp20F0HWqGLkKGitYFMzz4NgcJJuvBVdSLFzdIHYdEQZrNiPlrxZXuHW/1tp3h
ZcXmCK4fdMPZ7jYSK5jKjHL/5kaEldnB7U6TgIobNN/FqC37aq4TKCH30dbZ1IudEZOXqp2UXM25
HHQ8eRtbG7vLVDjULobMsDkBTYwSU6pOe/BhjSPlepQNMyXWvQGuSVvj9H5vUEHs1qA1goQq6rvf
yWDlya+prv6wEqEdhZeULvjZ7mqmGW1sH+98XM0zwGIiIyCYYynwaKcVE3LYEaHB/qSfj4E243ZV
nNPFQYZfBSy6IzFn3KZFKcTio567IpjNcGfUFP2b3L/THmwaxZCT8cCjn73DNOEs1J8XuKGZHgQu
bZ9KARyhehE+GlQ1CezJgQElGA4mWEVDZ6/EJmMTauBt2OEpJ37VSdwVbKWlP4CVQ0i56WE0To3l
rm+38dPeg8Ro0cdZoQKonIHM30EOPsohTCIEPJDdBrRFfF7Loh0uqZd0HbUZMBWCYd75f1xI7nhy
LAQhJ2AcyRLUzgyJTELeh17EKTm9dRKCFHoCi0ltlCvGugZNS0RX7202cVSZNVTeAwtb/DMWx7lS
VpCUO9O1T5nXPga81jFtFvYTILzdOIha445p7D8HYptGg9JveCvAGefO/19m+e4p9tf3cxI7hKd/
a7Iav+dLJqC4MoGWN0VCupDdwsT93req41ZpZbPAZhVXMmjVsdtoJQuG5I1GW6nKK9S1ZLggDPt0
p1VpX3gFuDKZmqn44/caApYhqDr/NX/WutMXAXH7cD4Gwdh56Y25gnRFG/vln8V4b72xu2eGcYro
CVWTxA65BUjEUPkYHtp7j7r+IRL36tylyhhnntg20DevVdxOqgAwdhBXgfc4TGM5UfrcayrjMkw4
IN7piV/l8hYBYugG/pCmoiRh9jSBBWQ8pRYAy8jeKpOaI8iF8nqjT8mZWmr4bd6EqhDhpKvf8/AV
FCFeaF7YX+90+nqI7AVP9NOkhyLASLxT/y1aVe5qGSxCSJ6Y/QIxq/kxYQj0yqZOdqMvXEnwXjCC
DNPT5iXU+G4bOZucHCnj3k0iubvNue7TlgDLiz8T8RZ3Lj1EIdd4Ke1zaNapm6EuDPD8NpOPcmiR
QM5ZokdtrsKPBkcj5DZ4rFGvca80+PCo5J9Iu5HXI5SIm3/fmBjpdKN1M6G0AkgCGuBTTnN55bA5
khgbge2QqvDgmKmSmsRe8UC8OHIuKJGBl/JYvGPQikCmPaRTa9wzGFLq+1KDw1FeRAFtkRY6Q6bm
vIHsZD7wqImK29/VxKmTTI9KqHefOc7Kjz5wDXvNXydj1LQD3w33ogaPb2r5epwVB+1P03jd7eY7
zaCOUBRJytMUYPb+u2u+H5UbS7spR9XaCXWCVDJtXwk5j/Op2W5eyvwu4JhnrUYrZPlLNSW86JW4
F/oH+gTF7zzDA5xC8TYjqXIEnyJhE9UcGgChprF+tX8qcAts/ZpoUvuwZjetLdm4gWXZLbbwUZ9a
UcKnTaB4DzHtdCFsPMMI0MMEKlwMgom6X20/Nx2Yhx4sPaaZIY9/yDm78WXddVbZdi3KEG+1xNr1
0Q4lNJAu86CKXVg/aDFp+YsIIp5zcuSO5XTGiVEgTmURU+JMaoOzxqPno3a6qxN/iQkix3Rc4pAL
csZnhBdxRoTXgAxXgKF+kfiMfEPLpsFE0g5VTH3sIODp0UfMs34tJyPHXsTBHnDagRoCWHvWO+73
QpLuBr8KFITNZNIOjrOHVTqUvH2wPKRSUoBRTxRb8myqlICsTGndYyw/8ogIxIhmWjNxg7h8XZIP
A+b7yTac/XDf5g1wzjFRRPVAexZYoLqGKeYI6rSdqWqydU8ZIIqQgKC9hf9Iz50fpDFrk7S0oML/
gwrCJ9rZrazj5StF0EL7btkX/V5zoxa4u4mVAdPpNB9wlqy5CbrhbxIrVvDKo+nJGpcIpK26MeUg
WXGP/KvTE2oG/mcShLZqPwtZ0zclMqGB+CtUycFjF2OJNY1xUoACgFVBfDy015uT4OFlT2//dXHB
yQVSv1MYYLUHffGrB3HibvewdI6/pfhdP8kMVerDJKVXTG8zwctoDJiZWBDGB5cb6JPY+Of+YYoh
cbJ3bQl0/wpHp/TBBCR+XBYjNDAVCV6fOVOSYMpkh92Smomd088ch1kuX9pLWzNpkNlswlRAj862
2nFzJLl05t+4uBIGjqyf9VoljEWxZpHsUTXAHv3Hr3Pqwes/8RX9UTWQd7E6qjiajq3kXJbht0Re
hKcVRVr80tZtzf7WOyCh+L97UC9Ey4yLcGkGlnuHQjebVqz5tKi+sMhiwcPLvjfr+QPns1mq0H7G
tri7etDYyAd1DGfr45o1hGyPw5Vc/isM+yj8AeVp6QTeYjL5QIRchTe6dWhT9Y41pnzi95LTWB7/
Fv6of9t5Fz5Q9C4hdYpZ+7yX67zPP7Zuz+0FPA7Z2TZ6leeF6as/ywa6Ay1azk9+O4Fk9wuREJ7s
RcejKs6Min5OhM/2cSXumxdecTOVnxOYfevdDBhDDnGYrJ6PgRX2bwny7be0YHFhNhnqz7hqCjMe
Oqo0+QmBetBBj0bKWrqE4WBkvKl/Zcp0uxASiXTbzZIBi+KpQYDLwVtsbSMYF3IhvQc2xxMLs+Zo
9LD1a+I8DXnrLs1MJLjYTFo1ilXziFkLT4iKus2pTfELNoeYYr5lVraXyieDhvj/zfTbWGX4FmwS
iklR7l1jQHz3XpXp28HjCWefdSjX884IajBCBcLgopXC6iews6OLfrXPNiaDCo6ZOFbFv/gdVzg2
jVRLVOTpvYNor/4HzMdzF7R32fdIQXKtY/wFmOjKZUKXgMD2/+yzL5711xk4i3pCOJpC5p0XKEzq
ufC54dhKMVaHajbp41WxRQy8Q5i4BxghSQQD2+N1sca2iNX6mmufpHmrMF/MsR79IHgG+ZCeVivk
8cc/uBSGPMKF7t8Tl7B3diTUrC2dgQw/X53yT0HU1jRmyx/qdvInb1GNILdWHLv/p/5u7YzsXJXn
xDuL55RvfmeEGtDWbml+w7B9JUh+4CPOKyQ0ErN9EXmHUfB/KaCs8wMjgq4fhRNNyz+B14hLZjYQ
nMIzVf1H6nR4vOURpPGOl/95m6mj6vPOnl4Ouwsl2UhDjw10HWq1ukWOg8uYVP76uxw7LuZ7VD79
/3tWRnm8fkEWBuTj3crfpK287hZ+QmiXXxBoiEO7hkgXs2g3cF6GdI1sHNjnj9+cNlUoK3buhzmD
YM9TWuebZyTUvEB13MYvv7DlN0Z5S1hUAs1jD7zrq45pt/68m/ewIRkb4oTRRJKmlJc72+QVkRgL
/8DsaoIsyldF9lrIIRptR9qHfKG1iHyuQQEVuPqCBmEuxqfMyB4NjKTt5NLmS8hkLHt5t2wEb4bP
K1P+L8Num97GG5Dzi4Ngdhjetfi2c5f+YrgZ+bpijauZ5wBxeK1OKcWb0QjgfHTvvy/hmzGu/V8n
jvQztvX1Y0C8xBdg0GC1meKFATiTySdG22L+AH/Ocf/dFGrif8XnycJjuB7u5sYDJgLnPgrsghob
rs6ZwPhngQqtn4Wh8XEhSpr9UZRmWPsYYYcjK9Wvu32KfYUpJjfUCH0yf/mf2gg6WUBbRepSIteI
rhmPMucFz+r+dVFZwUbo8XBqMv1x8L2kkR/cS1kxsNLdEwz2uj8+q7nKeaLIHA/ihU8bQdUqTqZG
Er7RO/aYZYlp9UuFfILJ2EnxqwxDGGLWOZdQfzNuulHlIl8vmCYapeehgzZoPFZI3rZHkQEIQAai
Fhj+NUuJjmXBRc7ROYdN7cq7iYmCMrp76fTqemG66ylMJvvnT5pPdxTwoeHwsNo7zkoPnn97Si3L
UN7M8d7SFbvaj0/Mx2HABHo9Vcyh6NisqNlviMwSZLH1In91O68SqkjiCHtx+nWNuZwNzqsfFWC4
7YKAqkAc+8H+mOnRZguGEC1LUsUHiOyRi/oZmvZEwhJGDu3LuZecMRKkmA2sNDkeKif2yuEJqU9C
E2yGQI2ZDiGqRRB6oe88cw9lGz+MmbHEWtInqJdnSL0CvDvUyzVg6tR4YyqeBGzbKfXVnM5TU6QX
us7ERW6aC0I1zG0nH/7pn+omYKM/bOHVKGCUrXtZjKZoT2Q6GtVepVmpctXDs3l0oTXEVodCRBCj
rXh9n8DYYMHrHunanlNLpYiEUezCL8vWaqqlnq7PifRT/DYrzXs3+pI244g2arPl0elnPPoZ606s
sFdRaTyPEgDuSYTz3EEOTjKRxwvEt7/qY4bShfDSPL+icRyMpRqcOk8W+sPva63UOGSyCh+o77Ti
ZkN5NUpDJLzjzcc/EytRnRyGG27a2RtWUQLZZ8WoezxJCefMXbt1QG6UA3gDuzUywuUJ0hKTzMCy
HC2TxtNYY5jBgYx1Z8KHhqILx9HFx0SQkjx5Rg4rSxwSFzT8mZTGMZa3ZI04xZJ8psjkEbjdMhz2
6ZP7FPpfeBrvHgVzoTDpsqy6PTR66KqgHsgj3tj4zomnhDYHDxU6voZM/m2PygUxtc94VhpIsSBE
XjIE6SVFYa/xdN4AnQR7rEXIHQbcKlPdrFJyQhYM63vY868+Fuwpz9Bn/xnq99nKAZ9Ef9RvhPJB
sJ2Q7Gt3ci2A0v3yT2smJ3YY1sJcaXjLEty90BdmyK0IJqU9OG2gV7Z0uXnyomyzICvDHNBz+kfa
N4Vq3zeW+kDqKW4oaa+tAJw882yvYMczVxz6gJ9LjCWS3V6BcyFv0YNQldUOhwO2v8EMmE2Pujqr
RFu+lK9QZBRaeJ/0dr/htHJ9QxSO3SRHoMwoLDoOu7Lentdm7gLkV8M0cswX6QWlIzQ+Gvozpexp
qrYol/PCtZ86Wl5YsKYSnxvWe99lIoxtJGsnvpRInkAM/6z79n97usa6m0aXq7ox8qeAFiL9OlhH
1rW9Dw62WRy9+BPiNJdwQ7nXu/y46sUnzCZokbuwe8oq4ufj6oX+0kRzyzZ4Bk2Uv85jEl/vP+QD
IC2MZKB7/WHiJRweHP383lojl73MgEOGiO/534eDS06+zkkvzIoI0EoXLbjt2Ne9lgBsYYks2C0c
k9oQcc38H5z0Nb1wJqsNUNQ76Y6PFHB0WQ8lLMkVxFsnBXVxXxYRKblU8lRyw+OO+vz1EbAod5VD
kRqnS6x6ykgFAguH6pRsgq2RKpokJMo91LKL2jxbG1AsdL8rKASMwzfhkGuBpCJqMb7fVHrh53XB
e2nYbiOzo5SUUQV0G0nvfrx0WAX3ELxAM3nC1pR5IAeZCkq68+76NufmlPTwv295J/jEpqOvKd7Z
ZGAmCIVepGfs+TC0Es4/Cf/utGWQ5Ee5y+UGXhqFUVvLnXSQQWxAithnT6LyU2EG0n44NtvDnTXC
180sKGmtF8Y5raC/RzfFD29YTmTNhO+qP2q/D143Lnht4K8+098B924WVOsa675RVDxrHlDrpKyp
AUOcNQQSRxERPneV5bEykU+Eu8Z0jlUqYZ8lMF58rXrxofeaVkcMw3ZL8r5286V4/arpq7/ir/lV
4kK0MSYy8YscDy9EjFqKu2Hi/QOA8Xe5WfXLOQVa7o9p3etr1hGgJRUsDlVfKf0kVzwGG3sh0tao
Zavc7JkjS5DJzK3P0aFLhU8++LShOhTSzYWL6J7y0eswu4zGAqnjGNTE7A2Tdb1CZtslM4N1NRv3
4ZrXJUpAQNOQ4iauj5IW05oL67HNuPeWtlapo0JWa27/8af4bnUZHT/JqBJfJh1Ncpd+8W4+nvV9
WjgldJHZ0gKrKD1ETxekGGkZC7qEsHjBSErEDCnmtpFzvSH1uyN3J2vIA15soRjr6ph8lRqVfYVL
bLHiKqs62OB4Q7TP2vzmFONJuaHA2ao0/z25kGFzgqNC4+IjIXIe2UnBgv/+UOvz7jGC+/FQduNg
64Yj7BDjddTbamSAm1LhKF0rQ4ib7WIAMebxQGWryf/2DbJRYo3QZ4k7vBRV7ymylVGfOvpOwHHL
zhdXVvlPXL7L05qnA8k9i2yuXhnyhZ2XVuAL59ld5gxGERb+e87HcT12F0Ex2U29BAfjPKz8q5iK
Ol9serr0fiR0/frkmxiAAQTjjxntcOLEpZtvB0RDU4ggkbWBICT33VMklvrNFQ4Y3rzTymLrxXTL
8+LEFIPZFcbnXqAzzd5TIXUrAQbZzsqL6NEsTQSFI7/S+LPqH3K6ymKSOSRBtcL/SX6GvuF4yS+W
6LOq9WGCEfpGhm/t5r6eWWvRa9TbkPd/77Trvjyy7iDKRS9T/DOR+0kP87bl02k+Layx7DqkPE4U
O6oXUgxWB8hYn1mEYjnAUWjXgxUVqj0T1eC2pRf4yuLHeaaL3p2GwLNIKK2QsK0Sq4mlBoZIMf3x
bKJPamtD2k5TaEkcWSujJr/klqKOP8fnh5zFKRDgocalaGEmfIDfhD5Ek+7uCtBFGnBH/Rp6rx8M
fC+6SfrQsuNZ83ZpK18DbBxdityPdAH0Wa8H4R7kgwaZ7vv3AIps7xgrQSKBUsTH2qbNEQwjb93o
70whRilZGF8Yt6T0AkK8ajum/0TWdJ5pO0god3CV2m7+IYW2Xc2kai/OQr3A4L/lZ/4oFm+f4d0w
FUKcUPaFroTGhyNzv3SqecOpsvf9TOIFyU1/8aSqUylDszTIBwH+4r/tPtjC5ElWuQ7PHpo4fpwE
y4e4DrSrp20UpQW10CkuwsEE5A+GUsu8c+FLjvWwEwa+LI2l8+o9AtBwzTheSpoVnsMI8MIKqLJi
gItdVJnUqQBJDpsEjrQGFJuumEhXZC9yte4l5nc4thqZ8MCZYZARBPhYrknpqBPktB/LKW0zUWDW
okPe5BAHJkvKvWn8Ff8t02aTbr/4LRFD62+Z4cFACuPWBoEyYAxDEUcLMVrd/Fhe+xmlpAC3aO49
qRIeCGmeoxmVhOpxHtN8Irco4xFkhdT7f/NCx8YnpNJP6rhxETrQVv4U8qEcnBfKJBHlrIwoOYqH
0UnhsEefBMLHjZ8VY8NxcDJ1x6YfweC3Xm+l2+xtRE/7PMsc4g53jYiphkXi9iUV/BWAnharWRq0
A1kzXdICP5eHsa0gq1SnDI1hdVTjFojaYxtL+VggKPJXYOQXSfq8KxJX3KrE1Q83rHkxD+KIOXBC
x7kIiMxA8u04ib3ILwGwg5/3Ck2Bx2XdCICOrplIbY1KmTeTv3rRRk0TIBBChgTubxfirM+DoBaQ
kdooNbFG4TkwHNIMuoEyBFe2yqZFcrsmYX1K06ekmjv8wxsm1BrhnS222AUsVMRuAOGXkAsb/hsD
tqYZBeuOz6oMq4sIHGvsJchL3EbDFbJyzE0BK6u863MMET2QBnMj6StP6qPzOYATMkv2nWXe8nU8
+A5SabUoiXXPhuo4fgsLHrzkM/o6SAHOCpEMylwEZWkwM/n86z0GxzcuIVA/V23QBb0PxbQ8Zd0I
cIzTsDDI7gi03RHEqn2JWPwX3ZtBj3i0lWTHsEZrFHc4kLy+MYyqcF+yQY9FGSPe1jZkNYg9hGqL
66punDWJvyTdkl7fcmJYf6YU1Yjm6B2ZXARqbJaPurklINP+SDk+d45gJ2NgftEKr1JuPAY63i3K
NdlsxPGN48rmJCROV2KNnkyFk4JGiidSfq4GNoSAfXbfl7jR36czYo3mwDB3N7zZjE+OkSHP8b5h
ChuLNYL5/HKoX5kycp1PEHjGOYwkoNFE4mcVxMhMEgrrPoYjouOzEDUd4MSyArKyu0CCiHGvADqa
e5grvHDjPHV45NMT51li8UH2JioZzn8/evGYeXOpPDL88oEqP1bASXpY0z+ZewIb7TCJuSuQGQIp
stlrRuc+S3rPorxuqwC47WqnuGiJN7prn0tVkdiX+5JRoJ7ziQmeoOLs4Z0QdcJdAVwbC/SMtvLx
cSsGDZKtOR3B0e3bgV3Uste4h+rDjpXDrMc9cTWMG1+F7Bi12p7vGiyC2yN1+viwP5sklq+uJ+v1
ZwXd3QlSrKYRXt3TStageDfzvYL58rrqe4BSWuoQFlT+laaO5JfzklfaVsIEKBFnS0a0TMbiAvVU
i0dlQryc3E8b65Xfq20LBNKrTNlqibcf92lkyKi5Hi6W/bDUq54hiNlHJ/abYEWxHfAsSK90kWHk
uONEWqJYpqywY/ovya6ZS2lDfDaMGQuLDjAvKlUIekBVWceIZLORhwmyTNcoP4Z/AG0bZaaYC62W
BqVJIOwVCeSymcaf+Rpjt5s6Vz37suRbdd3ua96dk3+kFuquVvqh/LtSRkviRxR8R0UYkLEeDQ5n
7euGk8gVF8GC3LLH4F847o8Uay1Sbrb2HZRLLL3S86R7J/f+OoWk56EXTwlOSZ5JyvX+KR3NMPfr
yv8Hh2zggCDJY6RHcOo4Et4dW8/bXmDcZe4fexosLLutyyN5vQMYGm0cPkkrVJdPqzx0nfMevNBs
ifVemspovYgVSloP+YbEVbqPeKWqzThxHHzahew5rqo58a8vchvS7r19wMqKET+7WgRaSoRzbY6n
KNQmnrJZZUb1mDCG8Jtma25Tn+PXlZR0nyv8jgKciC3Zl4Euul5adbQEoKKy3FdcEQs1VYCRXj2o
P4tz7iDaVj/lEwez6mR4X0802GLm8C5TV0SpMSXw5gRnItmHc1PPmiEcq4xelMhYnBee6koplKlP
Hp/CeuGqtHn/uf7EfJCL7Yyqes+8bf1OMhOzWyMYIQDn2fldABPq2nn1FEuwqLdoHcDVLHWDQRJp
JvIFlV8bwCiRolfp4FG6eRnc9zNiL3zzw2lPYFE6KQIUN5wbBpSoJJ+p7XVvEZZUZBQPEO44W6eJ
JlcPpOhLPZz2soBTfuN/wB9mLgfQazuM6BhL189oULPchej+t+C0kTFmXx+UrrLnc8+eCYgRQOSF
5RK+/RH52XQiEc2yEhdtNFiG7GjCBPhSDOqWsWBwVUcR0Af40bxx+4ZifPPcY2MNsRBqWbapLO3t
wzaI5VCcSoAvkXbIiLZzhLVgldv7rZ0oCduUhs8kANjBEgAXBygPhS2ljjAHLH9nsh+39GT7hTe6
te1pPIiCrmEAm/o4lqQyyxJAAHYEVL1wCZw9sYmXj+EwQ+jd7l2/AgZ+SmAal2rWmaS76xs0AxK2
Zzaet5deOhqrsacIzIuPmXnWm/NvNxQILEJ2pok7BkIn+OvloYMfn9J7Q4V6tNggxa6LA3V7lqiw
qQodriBEWWdoGULWpaDXT+ferWQeMO5XxzR9uelrzj96OaACs6CG/F4pIs5EcfHtuVKYljJwnGc2
DZbPOnX2xeAB+5ui9hs2g4vJ5viuToWUwiyYHO/3AkyTemhR1chStMmq3pOpkBhEXTkrW2Gc11tY
sUh8u116zEmmaNGvv7EdjmUb2OAm1CwOiHRVLurxPwpPITQaCj3K+0zyFEep4bAxLvquMfHlMBS9
8IuhLnGYfZayt3FKFb82fzCNc9Izjd7n3wZzsJf6y1H3TvN+IEiNK/E0TKhZRwds0ltz08Kv17uN
FKEX2vR7tQWqzjw/nZEP85a3PwFqtqBIz8392SNPnsy5fRJEvh8PVtAI/QSZciOe41gadnAqwGlF
PslpQZZj5w3MOj+0vzN3Azl5daix90825z/2C3SOWdbxrpMPGY25HCCDKK4G5GmWeALARvTbwL+E
pk/Wh8c2gPVsP+kA2Eg+mJweYdtnXMROF2nKf+zJb2x2JG9DF7E5Wel9EnGS4a/ZwM4OTKDdUvjh
xF52X6eXhYpsNIh2emYuGCxba97e9W+md2502WRTNWTH5wuVIPTrjKLlZ4Fb4StXhvT1rpMUryti
vHgaJ7/SD7MYsHB7T4dsE4kkUn6PWKu/oXrMSquj0Hz4D/ZptKO26KdgXol4bOODhCMbxbMPMSrt
3OuQjwILGV9CtV2p9rw74j1s/QO3Qv8XZ/TwaA+1Q0eiD4rESlUSyXV+73J7YFWo+3tdLmrSSTnW
S2k2+8fyOxWk4b9+6im1Vjv5x+gDsU2wBkynaQUDoiC75ASv0pDluHC6U5w8LfcYhiI5DR26JXMh
UDLjSFByhLSfzI8TgNln082i3kGW7xiF22SBskYvXQ1fvytgQWGNckcXpuYHZaTKzBfp8Lr9GJgI
spJKhcMmstnghZiGuZl9t/fGQfONnfuhzF0lR5c8Y7/YGK3MeY64p7cpIw+sG2rhZtoOCVQA+tFj
3Uz9XX1vu0xXWz2zSx4CaVvp7fyZdECfSy7EBYq3ITZvd1KkS/+aupyZqXU9gNjnbp8rUKsiSvph
Zog8BrI+f4OzWw4FkoH9oxJpg/Ou9CNHDAewcG9l+fdiOCxFLU5/Hdw6LzTMdfgxOBrVbXF7QsZR
qIg2D6je6b12050BqVr7iunthWJom3QOVBayzsdHWBZ8GKLNIqzM2ipScDWqA4VUcdVXeK106wIy
D0966HGhXdi8VRLs0lr/dETiC56lCNIDcpRnBBViFlfkPhCIMcxlpgic3XoHWcKDb+IASwWXadtN
m7WAvEDoc1mRB0uhJHEX6trlPYxU3IcEgYK+3z4BNu/TYCrDrpPpW6ZaonxW6ZYqmrmmkJM0Bs+3
NPx5lGp/JQOdREJhLok4GZO3g4YGCBOmpavNteNaP38P7Vg//tKR12Tbs0g1yjUq3GyF8Eq5+wM6
G+px4pwoDeNpHuWXlwuF6XviStvWhLz/yuFoXRh0suDn1LeBVqkSK8XzdDp7JS+rE+O9ZopN41xJ
lpGr0vMRMqhqY+8LV1leE/EiNtoStVv1QwkygquOjF0NpsBXKCk5ayRKNrYs1H8ZNt8iH7DHLgLn
fHYLitCBzxwGU7O/E8tK6hEXqc56077Jd1TqqAd2YrbO4OWeqE2AiVyse+r+tcVRwzOIJrIERj69
20X4IjPUooib8Vb8pa3cOGcVERqrG6L77kxjzhZCQrO57xoONqhhWG2IzibPGGder6Vh/rgvjJ6J
oY5k60vb5Y9BOMgyg5LjSprCWDsk/ZPhdQEAqjVZD5CKULX/1FhMkScRQ9UJLopB6RcuBEi2P8Un
Ns7OdgNqo++YPJzQf/K4FFxQLexzFgn6R8/rlBmdh2bLC37b0Iq5gAGi27Uz4qnah5OETFt8I+BW
AaRcuohJzPHT59kO/JJ2O8LY9bz3DhMdY+kpjxI1x0oKBVVVvW6v+0PGEzx/LJu9l4QPRu5IJ5PQ
XMaqUkMEwSK1idtrn5G/SQGGuZ+8kc2d94cvu9elrTe2HowxGLEQJcgwRoA7l8OmMTqx4U91bVIv
oc9rOLEsqmMzZfj2JS/2FAcAsQfOAU4w7Apr2yKqMMd838pgU4g2/w1Mld1bUrcU0uk9e/jW8WY7
bDBCUA/L2ccIA0NpuPsDTZjDQOX+/pDl1WRmAUnsc/IDSk5MS6txaCLNNtV3iM82e+Y6DCNiyogY
p9xE6qaG1cxV3OKFHLFOYlUC3COaPfbhUYwLqL3qOnD3QIhQeXK6JCGNZEnKHrcTZHWeBe0IRQbN
Zv5DKLL07XhgUT/8A90lMpTyERoyHLEeu2CnP1+5ldF13FxXU/ADjCwYAlxJevYHRznrDEFpxT82
JNxgveryCz8sHnL3ScIgM7WTHzFP4M2KeHfsThTbpqT8P3w/13734A/MG/IXHcw1BtpX8cOTATCa
ycexSRg7zl/HQLWEOixP8ZfUiVR3mB2Ign1u8sD4OU3+43PPF5DKcSgY+wyNWQLngM6ysVzx75m8
gh02EW4aJyFH2f8wq4BSMaFrkD03p2xUnrDGy24FRqaUA2DV9GuyiDSg22ZHhiYVYuuSvUn+Lwdk
Uf/er89f4ybrEswqkpwqRGBApF50B3AzsOPYRE8hGiUYqHRAQ+JWFS/C/iBgYhRDoOrjfKEDZBfI
aRZUTuroczIr212tsQfCpsD/+khkwSL4aFCzZJXapHFWMfa+eZgA9yjJrT4p+qogX4YESFq5vTlk
AQOhevbMlnT4KU9HmXMjVFJZuvRLASrgYJLjUPF4PXashNRU7cLPfjv1y9CEKYNEOARv8UUK7Ztf
LvtwOF1fhJ3XAy5G+6Wf0TBazz1xgkp44lPLqtDYGvp+oAcGoewG2/d0WmuAGS1XBQwH9B5/4Ru8
LKuJxaHUXpHkxY98RxAIcZPi2DKx3+8gxNhCc52PFV64Tg+i/8JLSLnNc8ubkiVmO+vaAoC8mH+T
gRCLHKs3etHkVNi5XwORHuwPyykBtxH3KRE+D/0EgOMN6oIxaxDp9LR2lMpoP5ixarwcwsCA90Ri
TkaTesu1UvNIYI5132LhnLcaj6ZdCZg4XXYlkdXabz6LoI719eUgO9nijqVjIf2D4r2w62gkkREZ
FE61lhcdFriVO4aJmVSbtW5VYFVhTr7QP6Nq1boJMjzBYetdkBbTpPEgkyNrxiqe29/4hysKtlTM
lm0RHmqxZJWk2kTz1FsJ9wGhYwxrr6GXYjalr/Mr9UVsM1orVsBnJXV9zwvsJw9cWv5iTQuBwyaZ
BLDJ3OCR8k6umbU6RD5LZVVc1vb9EWIKI32jiocWbWXcndIndyPG34udkKyJLNGPPkQC4B0yIRQC
o4kIjatO+YCZBMrJpNprebg+CHd9LVnMr8AWVdHMEVO6dumW+FRbQBGyaOCZuG5S7czUkdg5Vnz9
TxDPPjZyczeiw5hpJORgqSXrURFy15F8GYcCrfmL4gv2t4KscGC65TBgmQvnFo2zlgwgGRJWnSoQ
Uhh2PMXhpM4r4v4kkaHevmoucheJWsO79PQHsQ71STAAS0+6JnI6RAVwstUChpn6fd/ltYRDJK/H
TvehmiZ6I4KD4uhUrZhOkxpr0vjY8vxa/RIJjrHvP81dTcBLR+hEcsh18qYZ/56dGSaJbuIqmjUK
VfQXjJzCCmuReuuKIQcLEzxiPLgAxQ1SocrZR5nMvWMATjbJ3HLzxl+y7+lz1iB47um4pCLXEyuI
zsRSStVoUJ1Nqngh7V57nHCUTCRx441xEAXAlmnZkInXYh8fVdw9vGGnoABtXXZUVClhL8AxrpNH
IQKRfl58KDtFd0okilnQ1gunosIaw/JIlQQ4U6+a8Ib9uxiOftWxW0RCnPTC77Kb4dejcrkVQpd6
bPANHJyD4LXc5HJ/IuXd3lcGR5AJEiXZjUsL3DTr8PaFUin3LmNtV50NVBwh4CXnt7oasJ8l8UsX
2gAVIZ8D/mQNo8P3WQjMQsKw8s3aWtUTnJiVhbmv+aaLgqfTNCqh9aE65Xvrrjw1cvI5bPDE1kxr
YOce5m/l+Un9Ywv4vZosJ0kb1XFIieEV2jX4ynGGvZ/2rEkiuDIlnq95ic535tv0DnJoU2Ktb+LB
9oGANiLSnJIAaZ1uSDbsLMnDlzz8FUC57Qt7le3yconqSFcHyh3Bjo9ViothUU1uU4l/S7D7GSQ3
NV59r4rkOzTq8nghtMKCMz/+05H51/LlPXfPmwpdG1lzFlsKLimeV2e89ZDt/o6Dgq8yC9cRrY6k
Iy4OWK/a2hvPqbBN1yT7hMoOGysx59jrcATD55WtK0CRHUbBvSyznlLxxX1/EZW4Jtpp3Okg1tJG
X9M93/cf+2UUpr9ChP+YHnIAZGB8Rhk2Je7rN91EWnd0PaxxX0UTc6x99uOnjlbbahq0mmsWj1U8
0ezcJxiiAaaQdNXefbPHMv+Si0AqucUub3eUKlvLl4ggpOGTeUsITBH00CLGWwUMCRjI/Yi+2WQ4
B9RwkdX5evJMYVjsuZK1J8AOnd9Cv+m12Yd4auSDC4cPULvj6qS3M8YG9P9v+q78uB0D5+ZKK+FL
MMERT33xlyFBLtmiimi5EDDvmUOePTBPThPPy3qoLxzCJN7E8mkG2uxqWysizG4pO+hpcHiWWq2k
Gsx6x029lXKOJq6//zOpIRZZ1a5/qmtTbPz4vVdIdsbg4+NpIN2FeNOwK845NR5mQ/IFz3F/YDfE
4K4NnJQcLdbw2YzACvRG5afNigNp8Gnwflbhqwer5I3mACVkQKX3s3XeUk4/cWkg89evc6dmUIUZ
ILBtCVaCnf0SU6ou5nd/oEhirNv6MBRbSlx66zwF295bs1EbkvNw2xlz3vroT8CsLR05PhaCAUk7
Zjn9XwuKRmSxKP1htegQueHuNN29i76ecHBXTSX2Nf3xfwzv3PFtJq2NYxbj6JNwSEN3SGdIqscF
YjZwzKJsAjTdaymUICF3NTUICgD6NL4EGuT+BkJuO1e7rUVLSV3ACS2Clxz2I5n8CZLr02ibzppT
jBB8h42MycpKh3KxWaMi50cL4jlYKFR9fu+/QeT+iAuZhhXMPtZ/bfMhkCuM4DSMPvNFCPX57IJB
cXPBp5C81oerM8A/iL4vI2d42zNAWuVowU2w/tUhLFMFxRSiSiEz9PoC1xE9MU1//Op67EH4f1v3
rH8A06srohGoiVcCwQ9cF5V19fPjaCIkvpoCpsmZRzwW4W9TGNVCPtMSbBMAtnXWIVPOUprpSt3n
3hFbE+KLmp3mL3bEV/G32Ib8KxuS+cuHWmT/KN7vvNznSUDGU0ak//zaHvsR7H0a4on/Bs4MB2Xg
7WYrsTTibypOlcjLY0lcaCm77iz/CsjfII9bkOTA9Oon9RKEUJra2pnovyboLSa2ZYX/z+DLoDXM
QJYb/eupB/4nP+ZbbfYjypNUuiUF2y5J5opy0pnXIUfJO+mG/Z7gbg1pMb20Oq5OHjYY8jnVxsiz
N6D9n2X8JtJcs0Z3B69AVgpH8zxiysnLb8hueztMqtbryb+AWBt1o0JYCcPAFHqsfbw8vRZcxz1e
Jlj4G+5c4VsajP1zawoalF94UMn+u72gyTpy0TGmDHjBKLJCT8BEo8c464cAecE13ayN/K4e7xZq
w488Lak332jDQHHwg0X3ilANdSZakCEiH7OqpqX08HYcvpzJNAr6Z7ldBPqDIaIp/csSBUD7jB89
G7QSXjVZZp5+gP/ilfWZwiwHKb/hu4pzzWBFy4CA1SNefv6+5Hkhjs9dL/i2IedhHZ19gdTH6zn9
TssLytRrdXbNLLNlvRma4NRkDnD7StZEqz7TxSEelsAZkNOlVZgOEYSe7Uij5s1J0dyIa1zU33bH
fgvqe9rb6FwSeFkiI32KM+hYXOe6FgTohS4HWED8YU+EXCZoCygROaqTIqUoqsyW3pjnQVASrmTh
XRd3kWovcymash3Kmp61U2chrnv06f1icLwYj8zTg01EGDJmQgiD6FLsfV2qL0CsxPjvaT3LQT7D
dJZGRBl1oMB7BR3t21mOtPUkxYjL/FwowVgEfvVB28VOlso/xf00e5CU93SqN4UbI+PHrt+IaIw4
G1RKDRRMA9IlnoxIbXVKvAJLO8KrU11f44Ov+ko4lN0/qCnCUrAGxcei3XQf7KjX+STRDolN2yjT
8VJLGdDfsUbKCAaVStcD+c6FkhcHre4m/muB05+Jd4DlpEdLjE6ii4tvGUrSp4TjU/zeMsPNVhpB
iFbLFNbpoBjxnfFyzOyhQSIatqKPzhHy/ogsIy6wwerjrZ/9SrcILFWXv7XzZEHzoVJ1Ma17wzH0
E1TUSCix4ldOJ/v4Ok8mco99doLikalRsaRGX4bjLEU0rRlRbq//G9to6vbt5cYEjfB7BYm6+8ad
gYOYfYNqXys2maeGjOVYIJwyief3hx6GsCLgPI0Tp2MwH6kg8jDKVzT0sUWFOKvgNWje0unO1h2a
5VAf/mqycvHil4CWOoPm5DmtC7HTqEVDbuRn2/TVNaTu8B0LEYmpJj55F6s9zx685kgZJYh+I9p5
S4QxEJs4PLEE4x4mirz0KwKhQdtguMs1vRCm9PqWgthQoflhPFq4x05CtD7N8Yr5/D36GQ8jLzRH
Ubr8FjiI3RrUZrdwCNBaxw7ZXHoq1ks4qtC8MbJ7cZwAx1yWLy2Ljlewh3k+a1wVbSJsngP13VxZ
c+aBAqtuR9HjPKTZ9GglRN+6vPOax+VOCjOURLoWN5J8W558nJQsmDXmex56vyekT1RuBHfRXsHZ
Bu5KoUckYbKaBVMsXGbgzni6Px1KXDltaeOsSYLDaGS2g0BnNIK0YqwNZc67Y3zicAK0W9ZB8m7E
oT5BfvG/gezOxNL/DwuKHWj56KSiILu2lFpNGTHBhnt4s+Dt2z+vhFrKzi0EzDqxahS2yK/j9QRW
FFNfRXt0snhsdoRx9T+mqvDxdaQXatquIY5fmSMCw7Adn7BVVPbWY4b2oc00Ok/zrg0m9qOGw8wF
19il97l/Hvx4zNMWzp8vqiqxbO+3IQyh2L61PvesrEs3d5b36Vl5V/NSwnRh4O+8gYaGIph3E0aV
4Xrv3fMGA7xbreBnmMmtfT3BOlGZALL3NQZvsT/dK5DETXMcNQp5oe5dcReBhkFgYNAMZK8YcH2f
lNs5yeXfRIAjJijag/Qf/Md+U5jp27txvl6XORBVfuI30Em+L/Vz8VK56TVQnVUIpVlI4jbzWIye
/LVlyfxMjfqieNqfELMSp6BR/DRBY4jfD2tN2RVwNMDxj2dSpdM+/so7994TYhyByWlT4YnbTcFn
jCODxUNUxZ0Od8+bL+3SLAwkR+JxKb4q4aBVUOpJpSejnLGy50qWaSwg7ZjkguNUHDCS5zjTrv93
LsnlzF8MSxJZTMg/jSIl8o7+cSD9xs2+emVVIs0BBQ+hmhM8dHetyPcd1QqyKliUIVhmuONGkUuN
/HByZYJisbRP8OIXO4G2TquqIAIgo+nmleqSQ8Lzr09gu6hnyUpjbxikrXfOStk1FETxbvDN+fw/
yAaKX1drWru4mrs4GGyXj4qGWoA4iqhIMjxtyW/LfKAs+3zck8qGjQaoNoizuZaZmhwXqnhgP7XQ
uauPDl+4H1HGQ5Lflcd+U7Hh+9u7M/2BBiX/vjiHL+Fi8aHiO278UKL+ditxUqi21y+7QV39F5pM
lyQ3gm3BozvUcCz7UB0qqqRoc3aH1CRqsVpHBRzXFixu/YkEEb27QR40qvLr7R0vXQw2kCv3pei6
WyIRtxIWxLdhgjuXW6dZtLh1XSwRpx+4/WKPacYUvyM2VUTrfAOyqtQgOSTHF0yPq6K4tcwQz1Kn
p0VR0Yp9uCcI+hrDumHE6AcSVuXBfHiN3HLTyVRAOw2SaWnjZdptK0gC4ZqUcuHZSG49LMHYqkp/
7W6q/t/DrpVwxfoKnsQzmL+GO6rl45/C8YxV/+GflTRGBmvb5EXY6YMm3rbIJ+uEddED8o+4fEel
m2vs8hQfDoFsMphMurewzEnLLT8UkDKuUTk4auXpvRJag2+wJaF0/3cIhlvfiryoPACtEcbn+BrJ
NFL0cPelk6b0tHC4ls8BRgaWqWBM+XjVhv2uQOPPlWkfHeCDBwxplViyXfCJRLeuVOq4+dka8x9D
fNk0gKS92bbfWaCoq1l7yY1VM8rHU3fRr+6M6slODCCHXYTXg8ZSn1ql4wspFGbrsrNzYvduEr9c
Sx4XklI9SUc0uLg7WUoHAMKTjRCcVQ+cPi2XFp4826qwr+ucOzwTJQkYRLeZDYg7gBVjAlhtHYzB
EdDg9TKgkBUSnBzdly0zTDzAz5u1M7T37AMHnHgFYMlODZmAoHwHRDamW2LezFDkPWl1M/Lx5ZjQ
0Q7cV6wgsNo63hASZi/BjiI6BHzHssjev0dH7e0+ERqL5lCL9eMC2mXRG0ds3mSBfC5VYCFLtekl
0ZAkxyc9JF8WuTpBlwmfCsDZFP4cKeZUSBmVwqKt4q27ufKsPELZPBwvoLZZ/CWT/tL0YvRI+vgH
8GBSYIbRLL8SFTLs8hr9k0kOv4Lw+sMg9w+3XHcDs4KlYjN6CrEIKgrR31DA8O7Y59tNqxW+k1Wi
0fjHWRb/6i4odsnsZuNwuKxcpI7a8/qG8eq9/rI60BjAV5PfzBznVGwcAaAha293Y0VIP//Esz4x
uLPvOgkgV+YY8NAAMREljhvcQMHo8yj+cS3nbgfSL4XThqI6LTA5qNzNDbZEYVszyE0ZRI9dl9l0
HpxD+3BW2OUBK+N7nKapLgGyhVys+c+WuszQLecek4mPKUrMKSBeoNiOwqmo+qlrVvtEdnUKN9y5
SdCL6EEOZubZFIevXQ2RCy9kdKfjVXFl+0GA1Lgbo+dR41Nb5NgG5ZGR2BqJBLjmcC17nJVO0CUs
V7DCFlDZWy3cFvjNaLg7O/cBDRk2i+1ZkC4gN1OqgSGj9HHuruvIIBsaXr2PPeMQUGsHtkjsSVsi
vQGTPdlEHJa94YH6DVGYnqZuCnqsFtdJRbRzULbhX298eTB3f0SF1nNUY4oVtlJKc6JRqXdH93/c
iZZT+/JfwUXTD6oxb9s4p+b0efa2sEviRmjySnuXaqP6EmeoW2+wIqmXzgQrqGhRatfBMtmDiQu3
Jy8fA7B4ATNYxfNXzDaIqxWRF2KuLsIfgjPYoDiEB5z2g1tz03KWopFn0iAGxwryExIbtYjszkbM
Ncqdb9Ey5dBGBkgRJJI3Gzt8KEBcnR8sT+jX2bRuQYKMP/S4aYaF1QLhmcEtN2GQfVi5azzii65q
nKcAIr/Hjhj6x3BLFjZRoz5WdX1ZfMHaEl45jL4aSK1k5NPAjH9oYB5/tXlsPL5V3RDcPKPItqgJ
Dc3Nh9m3F6h64x9WU1CxEzUftkHJRWL2n2Q6Z4z06FWVyAhOtZifI2MJ0HCPb/CUCcMrQPjpCsCl
aEP8w+a/Vd/4/kmwo1YxvgdWDfcpoAApLQ2acoyYc63SRkt0yY9wVQLkwQS6/BY+PjbRBnVWqtF9
RVHudSrOVP7aD8lPMYWH3os+9J3YC0GbK4EohxkuqeJnZQwYMTGpluA2E+GR/s7Pzdm9XUJrdO6T
U7lbh/Z1+3SHMP9vUq1xtzJU3QPnA7I7Ky2tmILnYZbVql1VgLKHjVitJn9o09sbnoJiSVhyYnfm
FQUGC3xQJcmgcgRqtIg8RORJanD3cqbs8xPe2j8y5pgbmJzcejmnhf+Cyrg1cmDUpKnWLsmf0quM
1YzmmLoeSHfLNtQauyuaX/dC16klcfiLV7YwtTyhexqiqLzRVfdqNE7RpnNvOpu5XuHV9Z25RIJA
jRW4GhBHfxVhi6VrwBJ5z7oPQHwls3jktf2KR1lQldy8bnalaZOH1QrcEvyipPT6X920q0GPyMyM
t4H489/W/TbpuzTMoaLG6EPoICAhh8/Cm3bxaayA+BvUmBkxXQkzPrwgKMTDKb1/lgFpHQqhnXtP
xvFGKolbXwmwz8ImHiEcNkQxkm00FN7YKAT4lBVqxXivUIfETekKznOG46bi1OXkndAdIJEjUyUG
8mCSblASXGnH6qW5Nyn9yav4+z2w0Saq99oxv2qwnil5os3U5w7xJO090SNCtUHVobLrKrwt0s9u
KkZHZEu6G7VenB5BecH+nvQ8YukB6HaPB5QevBeWh/oPQ05Goeb8yPJQBuk0tXcKoec046kEv1ra
BIQqyo5J07t7EoU+5b/2q+ecYSWZdrpmtc5ENCsTPuNvWpXGJPaUg7SkaRc60NGrpDmiMq6xfEJv
UOBzzJyKpuVrgnd//QhuFkD5Ik6rVpZcs3UytMCmInH6UFTwc1/JxI+c8280aDObThZExzKGJyFf
bOKM3At12hlepaZQAFsUUGZh31/Wa2YAlu6HnwBqGJ+5tdHX3ylgSvNBU31gXwioLB/XzI9no+ch
MItQfOTJT2ED2f/O6TrW9dF9WpxiFkQHYKPEaBGlfB6ej/z27goDdYffI3SW31iuu1Qti//z+mxp
iEoEE7PJVL3/G9PhluOo8mxN98Rsr/sdrSwjA1AZNjyU5JUMjS3w8W/KNXc6vr76eJwO8oLoAQi3
0kLRy+XnjbtAAeqCNEaWOBBV8dz1AmA3ELbft/kDtDqnnzeWym7my2JUFJwoXro9yUo1bF+aDtqo
kqUe64E92t4+/6yggVEnCOykR9GAw1oeouO8u04o/VQY71BdmMm+HIeHRv67hOwLAj/3ddUPidA3
0sNBmIVr5aVp/KTHxwv1FuEP1K1R0tf/1SDmt9D/mFNzM47wW1jDMiWnjNH8OdHsEGKBrXIUj3dU
4opleXaxBSxppQUrKr5UZCQOi7bmmT4ZjYO4QBx2MVNgwzt7jvTee9zPOp1W+TNTywzuHIGhzxhD
hO2AHCDaEEGhKR7g07vdoFa50Kwf27cnWPH1JyeedktJiV35pY81QKQMlV7WPBXw/zkJ1cP3FAHY
0c6oUvfXcHAirEMyMZBTCG0gNILY8Af+l3TTuOvBC9Pq4HXaCfDA8O27wVNjFEwbOlI/Onv+07oB
mBUCVeYAHpa8zlSuHGIhNupYa47jxDJSCMnb86wU1d+zCccImVWkf/5D8BnFPLFm8uN0bVytTuKq
mVKNBP06EpFZsp5qZpueJ6fkiHBqxeb84nIiR6TOc4+grndgvL+oxGIaaAltv0dQF3Jjka6Ie31Z
kvkonigN91eIM/Nqa2pGrwQc30KDnSutQzkj56LggjguAWXHdMeX4P9ePmGXqN/Nlf6peyVaqYc1
PlKwf1etZ2uI/dIGDLdEZCxWLT4IPRh4KYRLVKwA3+pKB675zEovJxy1BGRxe+Zc6uslM2waX8G8
i4KVpGrubgxLozinXZcGFkQpxTYyILTu21VcFBqptKcG1GfyiTcR5QzJA8HiJ+T5OjRfAtPB6lQI
pxXcB/6fMgA7mLFLZVNOinbHOechLbX/rRxYBscoCg+VqWLG8IDIHnfbjGYFgNKUIcES9JKefhey
ch8kSG6RU1tsXZ1WZ9gDYSdT9L/wX0FS9tvYxtNqUKuMdunFeb1UQrZ34eE027ptdJXcnnGCTp7z
sgCSRGHY1olVRKtUIfQ/8o8gKi38dbiTCFAHGJZcTM0wL5pAZlDf0qNfRfF+c+bUuLQ92wK9XqEQ
gqeRDn54BEI4JiMv2jOlP7Kba8F3wY9oQJeO/V8AWBkOklhqzq8RSC8A6pfFgX6jcduwfu8iY1SJ
cR0e9v1EhN9TNgvi9b9h2dOAybOJ/Llz1QSPNz2GtVU1h5e2MPpFj3O+JpXis9kIf5q7eKN2gPu+
28bt61snjSZvTDmSjujn6wVzthetmu4qw/VUVNqy4j2bmmYpqlKHjdqDGZxxHBWVUQOFydO3DnKs
b0BIRsIcWMOn295kQmjeblj9fpo0OHOiL6D3h4/Q5l6JQwkzmv5OAaQCM1pG88K72dcbzddR+Qi6
Ya+Q41Hg/RXS7VhQ3YWtm2HmpZkh7Vk41YOZ/TDgAgfr52SJ00zf1syLEwjeBDYSBz1J/RhNWwkf
WLhe909YtvWJHcXDevnmSl7IZLi7tYx2TNwaQ9gDcxn5O4c+2Pz9QOY//HFWG70zE29zfbOxPklV
hy+XE7XudbtCnrvHlmYbKEIwNJGTXzsuiEadGxHSquYzKtee4s2hZTzajPUQC5idEzpWxU93VAU1
ozKM9S+LHNF0UiRJOH4XWRA8K1eg+dy5zAj0BPuF82fmSl5E/uFM3jJ7VToY7a06AUkazsFf7n7j
m59+raI6h7eSCJFp/k6MUPVnqt8rG9RsnC/YEEF9YAVINIyhH/0eoxQ2rL27OnaWjJgo3k7sbOpm
SLZsnj9ZIGvPcTt6Yh0ww1R/6rTabY78ThbpcEKvjzEn2tm1S8+UlGAPNAov7G1K67h2yhTzb8RD
6ZeR/oNCI/sQxcCBcfRuMM62B8WIuPk1xulpdvqhxDSf8Lj5q+8/6IQn87820UPP7xiUBkdg6rcd
TDtnO2kZ1DCGiNWrzM7C3l6Jxz+wo/UHT/HZWnVk4GFWv+mFM3jB08MV4owTBIwb/OWiZTMmNh2b
CpzLcCqKeySPsIIRF9lJyW+vpaC5Sb0guJ+1faV1fVKnnBsTAHs842AWmRHvSF0KaSrNEKH3BQCf
mIKCYPwdE+SlbakeTRSHYsFwpcATrauEd2CaqabMJhLQFZTIyLZlAVztX1Pot2USfjaHB75v4EYP
xtEddo4NYAXUknepYy7GzZW8KUnv8OH2/B8w6yDUioMjE4pIkSysfyZgCx5LhrucLB6NtJWaA7gM
ufJbvRKOJpPtkt0tEHFGyx44ome6DyRnCR0rzjj0ejMpBOr+Vd5trEOgZ74v01cWPwLoZpJAxcKz
1xyuIhGghdiGFU+5ulQEf5eezt8wdNt8ore1eOj1bpaMgDnIFdfa2kxePMu9JEsSjUnw30/gAAtR
cnRUmGiEi/NdLcPekpKoI3QT2APkuhiEKzDL0gNeYRw31y+gfc1bkCADN78kYdqTqSUIckl0IPmR
emJOSpgIIYSvhN57135VLVjyVHnGmG3RbQmUnjxHHNbAdsG7KvAY8VtJLgMpuXzDuHlXTCfD1C6A
t5nuQLeSoNFKATlHOvrBb7tMJBlo0fJ8wXmbGVZdwhZ06tAK5gWH3Sax49hd63iLte9utsqAmvrc
zw2mkyIySUPl8yEuR7vDAcdAfgYyiG60vNEhelo3jlJ55T2xPrA6vc53Ym6nAzlIvHoY8IUJHSfJ
5O25MGBeRXRBTzHt6CiFEoM4CWqNFZzkow4ibj8THvCPRvHgaanL3aimy3XfmGcfX989QBVaEz7l
aZVO21d8tTyq85Rxdoc7lqPeM/0PsdMLNPpQqyRNdkeWHiKS8FVCkVM7y4zJHAsDaatwaITA16tK
Ps/KWhS70+vmQvD1tODjYZywcwN+NAE/9FndhAPQgPpCYBZV8ntIOxo0VWy/RHzuqMyycdc2H3qG
7iRSPrAuykVWCjDBXUbGS6xRR7zBuIVFjqG2cQ+WBVx7VvYccB67X9e+86zLtT49s5TqDs3rYMeb
pKdk8xtP1YJFYkhUeY/UGcSV//bvtigP2Re+kwNGpF+5Hnb32A+mxwA4tNjQutWq5EK2D2F9Rd/C
Kd/374u4Uc4g5NLWRcwDnBXFHaVQSc/a/IWq4JoOyCqwyAyoycqwWU9WxqxRFN0Mv1fPVMg1rn2t
Q2uawFxKGZqTrRBiyBXp0GDcICaZXzq8+pw8/tHKGiCE7aRGSZG22fPiZtMiIkJjp7OfYJeyVD6L
dzZi4XKGUqCsdPG094dH5rUPrmj80vRpBv533z3B5m7bYmN/PDRfSQKUnMC+4oOzLcH2xIQe4THR
mStR/kMfCU1DNF+1vbPw4wZQh0PC5dRuu6Ng1F7T86ICLlLDejfsk4BRveMxLC/1WVewXZaC0bl+
drQqXSf7MwgNsZzrhMjX42R+ICvl69l32MEeMxGpYbnOULE+DNe33cdtUB1sCm5mgseElCjLXOU3
6sXnqYKoMB6oo2G6NxW3g9Gq6BuPTCpJFhvdm534ntOeKASs0gKcfcjPtyUjHh/KcbJFmdI4E1bx
E6jjtleA0EpoSS7Sb0SKa8TcB1slpsxbKWPY+UaUdx+E4pJX+LBSqslWZfwI9sGs/eEaUyISL9dg
QfdEFVjUNEjYX/tWTguUqiXs4DmFSgyDCR6LhULW96cGK/O7nT7FF5jiTHc+wrM8GKEWvAPJgiXQ
ZXqrv/LlnBBfLmkKGgCAD9csqOCBGJYrHA/ty6jYPgw9066J7xQ6pJyqvbNM8b1yUYeM2uVbKIax
pjdIIsYP+836xafDC/g66FtmR0TrpRQzC0DJOdYb6kmlBATZGj4rqjCsboHFT2o8GMfJna7OJma0
/+ArqNYeOUpe8QdpdJEVNfCW9fEEdDorGTzr2AflWD2GzKAIdirrOylesSDGwmGPwP8Y4OHj38T0
zXIZMbNBAAZ30soRE2VgeGcqgoaRoNR2Eg/N+gMmpxMpesPUTtItgpjSk3svI4QaBbKXUHywJEN8
ubvngAoFTS31iPqG9JRpec8AFUS/f0ckhrAKgU6/LVKJfux+8hOKo1CVFt7Q/y+xqHPCpbuka/Cs
WZKD9PkGOiyGINL/jXQNPSshanVr1atjjfPgxdIQLaUqKi8w5UK8oakB6w94qlnlpfJRlcoqzgYN
hmjDZNCR7qvX6qhrKfIO70xpXiukHtOubHah7AHsBMKvmJVMyKKU61XtuuT2wpcbEepQAJAvHMpe
iwZNumwUNCUGy33OYGdc+NlRWmvxBmB0uOdSpp65HBnZ9F+oGXaJ49A+APkeGayMpBwBUs1qKTU8
dvdHP22I3K4nxuN4b6tAkmZaB9dKOvOTekP3ZKSkR4JJZ/0PrfKCS7PNUhus8x7kljOqvJRlTVQ/
VUCHOOrYtdxb2pQe8vdGI+JAnkrfqYZ1sxFWARHXjd8CawZqkivulmp3U9yrZFuvmF5xoE379QqD
yGzYJZHieixSeQXqOLW2gPnkzu0ndzeZ8LRSQcf5jDS63JwVuUYtoicsG92IR97Z/9AZq0giGzNe
kjjD9zpZDEOKnD9y30XEmo/LT4i9x8yGRBFGDudJbdSMENKt6u+rkvEaLFBr5IWezo1SSl/PEQQv
ZxfJ5I+VX2vVhwM+k234D6IPoJvhjHhe3YHnWUzfPpQFt5gS7SPmrquy/Xfpw8RQP+K+q0E9rZeB
BltIhbKGMdLIQuyPxCx835yQ+N2G2O+0dcfET1wKKtHj42BpQNaBTM/jgoC93txfoM2l5f0kRUpM
6cOdbD+5FJ2S8zY6jTbN9B4/JDALFinzvzDA4u9Kt5i0wJpk5tEb/elIpEXiJuc7y/3RH2RikFxt
BJG3rArtgjKUnzdeLKmGv85moXwbENyo3X7O6lxTSUYvLdHiOO3ymCv9QrNPxu9XDAYRwJFBAGv0
8q5Ip3WKlJsjjGysQ8OPO7ydvc1jAPzLTslb8macwGwOqWG//3SEU2cPPFwamJ8Zwp9mV5Xq9IFN
o22KtHNILH1gNWwedi4EUEetnwUQngXO4otP57gzaDhW4c7SQ4lgBxCjGuxcgn2/4qC72xfpAfaO
GGt0XK5ZDDVrG2WzmNbumsj+KQubZdAXRmCcs1QCwoxeCOI9HEW36BuZwAaxJM5jpWNeNXYIaTUb
xPaqXAQmok5oJo8H0f0tGpfJDiw/6tkwPA0RXsgBQMu3HeLm/I//qrYuIpQenPxzHT4T6lm076Wc
L9MLo6cbwxEv/Rp80NsMGicR2qxhgyxc/L58EpvhwgEBQf3sZ0s9dmVnziBPSIm/B5w/Tw8fg/qN
c93++NuxFuIgCvYKEcZZe2w+YVsVHxUzUEAgro9ufM9n0pjyveW0IZzwShn1w1l0IM1vITSZFZaA
t5juAk2IDCnOy9f8eR9j2Nt3qEPOInXs0fIZa9m2wVaW3PouFX0nQrlHikvpPV1lvoTB34z+gKnk
EZx1AT9+47b3rO/TcLbhvxiBH8EeWk/6BowG06a4ZTmgiYPHhI+ky+gOc6+eazLYNcJapifB2HUq
0w/bVCXaSPE7F2D7CGSvKVlIuIHzIIT7U7ckhS323oHRs76q9mT8wBCUorDmQQn8Lq9t1dSk57hA
Exsa2g/VXBS+r+AwIkY6nYUGju9n9Ic+OxPD4aRqv5wj5oG1mYmHdPTgaXEtKVc8fHiTy/fE/pTz
T3sU++GoaPq7RyH4ffq/krkcH7UX4gXb/KsABMinCc69jKxHDhVtlybN6XYk6WgkSL5+UbwSwJaX
tmidoRRMaqTNjPbyM/CzO+GatHZjZ/kB3urkKk2dz8G+ajH2KF/QdSVBa4eP99a/mH6/U1iPlJ/s
9zjebSpj3p2ApYDztsgCD18Bu0hYKzuSRZCbGvXT6Vi4vxb4ca/Up3hhEQYCchPCUTvU591OlBEA
YJW+FTx1NUqKZ6++NmvUeeodDFc8eRujRZM3Ycjjv4Y9vH9DyEkesielvYzBg2/weyoZzb2RfgdD
iGaRs1+5f7fQiq0dcA5nDmwBMq5fJ/ooO4YIRZSE/Zr3UI9Ya19I8/celM8KUSFUWQi7uAtCriHB
gBELQgrXqVk9rigpH0VKJyi0ZINrvQ1ggCrfu+kVwJP3tcEUx7idqZEri9+thrjKS34+hUKlvUv1
9ZLHr2n3qX05OdXcDdCkqfGXyqzWpDEWbzEmUY1nQBeR/zzjm6E3LpxkZKaYf3sqMUq/Xm8L/sqz
MftAbIbFdTO9gk2+UtVFULGDx+aw5IeXLBkux8yloQ/8xbO7HHig1xiNgNUFhK6ZGV5pEElKN8pw
a8lTFVKtSndVhpStRa1W2d9QYNbScb+UyGETtjRH9uQ1q3x2HoDqJ3jwW/LqmkFOKr7j4lOj5m4e
WO6qln4WvkQl/jC9hkadF7gGJBev6DuPs5dCjUNj0HcOtUOb0M/C25qode6YasJ9ySoeurw3SIzT
7X5OrSpGZ611R54j5z67x0sN5oHWdllvp0PSOefq/p+n4R4JbDzp/AHDtElDOJ7wtEKmQihVkc2e
mDQHs0QLTNQ4L3KGW1EpdmRqrVflLXAJVQMaLLbplawCrb294gcK9TFBNozTFHZGitEkAAfT+KGj
+cSGqW6oPVQ+MaE3pkBXmXzzl3EB+zMPxhsdeWCf5kVUfimtliyxg55X6Z3DPS6LGCknASD0QyEn
lxAn3on71C5KQszQ65c/pYjVlTIPQLrccbnFP+0ffK+i8uu4k9Q3RrWnsDk4CTfeNKhu99fyvpIb
vLpksSLfAMmKZ6oaoeMlzFVhIHM9VJt6RbyBjoOA4bhnWw9Gw0cN5DMSAnu9BLWm6cRksZqiqDmP
FkLhQBLf0K/SAyg9PqYiifOMulNdk7M1f6JaJwK7eWRBXqTdoz/9a377h4yqFGqQ7EK5uBfRljSW
TwMhyqDkVVXwJz0u2M2rBqmBN+2iQAAGfrTXj3ORxwrAP/i7VpIMiYvzJPZjqCjubJcQKrFgKryC
H4Xe75t3oI2GN2eDqTmFkyrG6BhuNAOkzhhCFHR6QbH+wOVAxFiEUjfRpP8h6PgJW/LtRUQVT1oF
HfeX9n04tqSzt0DOf9LxvrxoJVkweV4hXaG0UXjau08JXU75i06eQSJuezu7a/gGqey8zx/myfRV
1zM90n6kvpkK4YIWFNLDJRW8AAWcZUZgPOyte1tdb/bZ9lk1cLd/GwaLuIiMs7h+UOxAYxo0vhzl
oNz+pgKIJIX+8EHbaXzUR18gPalTdnm7EufPljmANFASu9R9SQdrYP48YSQBOlnF8EkS7is63i6s
hbS+buM/18899iPpUO1xQpXCNuQGi7v3uriGeKxyGOf1NIy7BSVU0oyV2cDyB5Yy40G+m7jQkh2D
XO0apKwzpbzL8JCteWviEtAMGjx1f6eiSmTc4ZNQCl49wCyVyeXzTzZA2vdityHv5ZGKXmWcZ2Ac
QZxCHlwFDarObE/3/twz6MCdU5ie/WY/1fS3qupPhCpF8ppUysXDA3jH3sVV/zgSZYkg8aMDiokr
IS5pKwdRnkSW2qfLmrXyEbaStnJYXP3V538/b35f0GOnxiV1uWdZVT2j0WyUFVk5QujfHBQ9yHTh
v7GtkwmGom4YpEbeYg1wbIg9AMyfo+abObPRvCsWB7TmfE4szo9t+jo7qbzITrQDPCCZp3l1L+Z2
XPsIWeu2YfOe4lPuPtn8K8JJsJofIesQ9Z1RRUPlxMw4un1btkcawJ/0IkEU9xHT7IvXT46w94WE
fhPKP7HZAK2FjFxLYsxp2EGRjd0IN+MMMYLhs17x76yf5xUPpj5u4IYCImftW/wZQVwXOobNz/ke
Z9UAlIsGhsCcqeTYlrQp2DiUFrPiLfMLSscXF09JxpX6F023G9tfGGfvbRceqR5erWMGwqSYG7FW
blFgYVDNDIJtk38Zb8nq+IOeU4MU+RbOhq9ZbTdOJrWQRcVYigUdr7chL15e/n7l1EhGrXaiUxKf
M8KWxaLldPaaAMFUqI3lJbDWl8830IFJglkVqbtrUrNJ3KlL+TJzI62Inn/8FDMPYdC3d7tPu+2x
RrLhLL8wVFeBnQNglwK1dk5by0x8nRezN1x2Qj4DVmPdac2u1q4ewTOehwab02UUZdV6AYTpJlyk
GkrhMsL5to4f/nhh9u3K056M3cKM2Aw6FpGd+TvfSbJ6ZmMIUIHrdmeNBYNRFbOKMwHmzL2jP640
ciNQ1Gk0KIR04EiE43FiLgcp4MGcGjxAqRGOLd4ZbQg95NbzNnlGDlLJSk8Qlpi0jnO0J/xkJcPt
k+ncbleNi6kk8g+LGZnCXnDxtyypZQwl5+Rufvqwa3tA7TweyiZ+3h6k5l90N/hIxeIfI6REaMYk
4sWWmR7JEaezRhKkvwViZNgzdfc04mDmZyZSOfFYV1yKFOIh5YrIfMypmNpWputJNSdlWrCRetmh
92eiRB7f6sbFvLjOxihKF2vvoq5pVYku0yoFpaRbS/MYp/i3Aodm0M5Exis6ilu/eCgi9WD96WGE
ThUzCIUgHrOwfBD7UUdRsvKFIwulygZMP48BvVDS1icKJ2zyESzwn3Rl0lPyr1RGFikutuqnXTFK
oX7LUCvVpR5P6BlswmwrwdYArTrhdTr+tNrmRLi/MIuMI8EAKxaoo6cmrnalxsEP6ECzXJIl1fnx
9+OXZ/H9owuVXIBsQVGL+YM0ZiC8FgrGQgoxG+shhKwQAs35lTlnDbfsqgJsPm7VzYgB365RfILE
PrGziIXB1ydxFcg/ic3J+jpj2ob7LUde/8iTvZ/WZbRH0eamqUK+CaCJ+WriN1VPqj+/d0xeynif
j4fqfdH0EVjW8g6bNnsDqVuMIHOfzRYaHkUghKGRmsMBVZiD6BQ9HXgVoPgKHX9Q2pyo53QN7RGo
6Mg7NMEUT2Hrpllv6nQYgECXViVkjWimW4N7Y80U1I/5fwIRw5PviYQtLomUzJpsC2nNm7AJ0v3W
RkZJVpxB03VskvrSESWEM9MLY8TXw04Tw20cPFoORWGP1ZBfnNlTVmY2NiVTpSbQbA8lnNNte0wL
bo1uCB4O8RyjUFzzoFrHahyIihQVodkzTU1LaHNpEpXI3AFIv4IDmWa/yi9SFvLpWd05EEuN8Yao
5qH7Ut3sg61dYjm72iIWn4yaHYj71lg8bXj9ecs5wBihRWHuxvCEQUCMMke0b7cXj9aTXpat/UMV
FKxW3jNFIFLIuFWiHdG6l9LTWWM2AAMRXzHKnnLq1R2XNg9uY9XMyCmfYKW0r4P/QFo5n+Jo8UXV
j4t+DH/OQjDf7keEJVYhBDPEDw3ktMS6PweIxC4Hw1NyVrJyOyqj3ukq2xwRk0Jjlq1yKeCIJSQe
ei51V3SazM9ny11OpKbboX76N92XZvrGY5nXeDlYmsBsDhPimAGW4gtUJ85prxUj30sr3R9NBKpF
1oKTue0k1+zdc+wUOlq1DrRkCdVu3m+XW7Chqdr/FibbUlBj4n6PbxzJoGku3QkRcpXtKNbjEvH/
n1+TtkITUgtkAslGbX43zBVHWnUolRa4K+oeIM/IML0OUMfACGJBoU/wcFvlasNEexxPoCVlMo+p
BZt+REHsimRrgsIq1pseSf+M8IyYgESlzfFjcPeMi87GgeDGDHGHvyFrfYnpxxGdN64fgNdx60zx
YiV9uM0ezIgKCb0qtKaWK7SF9pHLBBhY34HGdClKWBm2vjUYzHLzf2ku+m+izzwn63xj0VIVHbq0
tgzt28D1ZawxhmpEGDylBDSUVz1qn37S2F3zrysp/ISAfm/mrRNxPB+9axbP+aHWXX87omaKM0xS
FJi93fKUbI7xGwTgsubBgNTn8GHijM3YNg/EheyPQ7PzQOugsPmnGHbSXEUOBQWguU1t7GX/SSxu
B6/arlgcLFja9IUv8raSRj58sS2EhLq/NrbNaviLiMeD968s1b0R841Bv9HoC6gDmhVc1MI906Jb
p06/WEFiRIXiNcp4X/XSI6yTYAoUd/Cn2P+efC+AZ1ZXNT+sxftHj8fpjWisGR0Wjry33PTdnGua
sDHmCbGx66zv3WYyy9iBedMD77oLZPVUKEjCdQVtDwfrPyFDjFTSzBtCbHmGaymw8bQ34hRrDRp+
b0vDYg0gd9QEkqf4wubxhhU+2aYPt0ddGPW7rnuPEq1ZYr9MceW1tARCd7IOxeP+0jSTSYe7reuL
aVbJTTLkWpjzVmXDLxi11rEx47Vv5yYYnC/gRYWzPvdgDG85f3FNdxE0riP1HXML7m4/EgBgcDao
q96WCN6viMNEPqqX2ie8wsxmRBwTaWomUpR7vaSHhtows3YV7IHYOTMMqQ9NMdN4mCoYZkeUgZ/k
8yWCfyDamxZOayKIW6v+l1VoWtJXRTQ5vhmI3EFOgG4U7QV/62nXifH/9mzhfp/LNEir2SF8GDc3
DtWRSEdvGCBQxgrap2lgPEZmzOBh2091yeBDhBUJxfs1EokuqKii7avtxjJGGmWzGyl/pYxk5aEf
JCsB+h8/XF9fiR3EVAp+YUAUTFukG/tm2k/Rf2kgJaEaa8Vs9cPQy7cvMMRzub2pDc0nnnb0k0z6
ZLt/MPomc1WLuTXJ0cdF0eQ5QBKUfZ+HcSbpevoPmonZu9dDoG22jqFFflRKPR0hq5vJIvs/Q9Ky
KVs9XcpjsLzxNaZhD0JNUSJMRyUhhdjUITqEkVQNeIXO+lswGYyOZT64zKEmvgZj9H0vIcTyObte
EgfSW7p1V5AW66pvAMjebEPsRHO8E6cBitmVXzFsEXfNhAYs7JtZUksBt6yG/OqPxeBkwB9qE4C0
JgnvsUUP0UvfTThqxrvs9kxDQR+14VCEUsHhN5cHL0jfUn/bEwLx+wnUvvyTSQmZV8RVl1b+lggj
bV5j/hq0FoI57SD3VZL4ldNe6t187yqqXZLbX/UnouIRHjPcT4eO5AXBkOnqz8NwwcFC2TNhYvPp
tBJvid0w3AnJmRpPmYbs6f0SZI47Nai6bWwAXfHYw59WQfVO4Y9ar8HGcRrtgA7hCVXF2mcSakhK
AxYE6pdBhiQ/4S/EdJMW99hLQGN6AKqQt57leSp3GOqlATmdj/eVW2UE+lS+x+B050IS19k3Jn46
6ezRnovOX65lnXf5mvXimC4hsJyhlg6V55KBzaA+jLEfeDmBp7M6Bld7PHL5sHaq5LtXNSXK3LhI
W3KX4t0pvOLwKLqItlvq++lpYqRL4EdUXp7COfeSGQ7Ie5EGg1dvKHXUMJ4+1B5U/oczCtvUyj4X
tvS+ELGF7rRCeGbyonEirrd3oRP5nEETUc5bNwUcbbRarM5Rfr56tAVAYxFlMren8pIHhfybSrjK
XzSlHiHJ66CulH6Eacoo9yBgoCtGWkItbHXyB0dgvIo5ANW6ydrNY9BUNnj9EcoWhY54ybqZhu2w
v+97qBzNPF0sN5b2a1raaLP7R3FZMv91816qspN84Qx7aPIt2HMYanyew4z480+CoHo0GLaGnUVS
eu7ushrF3FLvksk8JLsGwcPQLn/1m0NogCE+iWi4tGqZ6H6zjgfSEkTYu/WBT0pI3IkqDymtXVcB
TcepIKK6RKLhvuBbGo+rn3muE1Ovnran0zEzorkZCrai6La9oqo6Wkx2qfw7WrEh9RsJX5nBOCdC
QhuJjtjY15x0oqyEkROQ5M5ywJ1+QunW8RV9FV3HkL3RGdepEB+v8DGyMB8oqMrMpv+pMJNPcthD
yIqrJp/176UtjrZdrRWKA7f7K1hnMdsWVFIoD8pkPnr/hDE5rWmjq5hX1vgwgZBHcSgRMK/ybG8Z
Jx6JAe6gQ6FGE2Lmk1p8rmF233IkUX8jHW/VKcG9ex/2hNOluFQe/5tMxSnsSOearzAOO0Ud2b98
56hr8rQ4dQG4n1zzXqzy66os2BGLEnT13e/3HSWVU8iSsOlnvwyP5fq6HmUtMG7xMoz2LHLBPI6e
GSP0FvFRBz5rPppPL8UGWkm4lYQNg2dJS5jnigfVV3w0oXhnKC/5G7l9CnPI4hchhvUmzqVO0WOp
tEsndUs4i+eXC6l9eshpAkF8lbSo1IDteCstfnxo7xHSA0rJaoV8VE6E8CwrYPQlekeWkkdRGaTR
3kkf7vrLG6lpglff7oGgbhGS+bNueDWbWJaHYSe4oN2wKxCk1NcTsxWFFqRt5J7tgQflYqvz/tHb
KDgM++C4o4nBKw1VGxWH5TMI21KLeqZ47ULS4M7vo2gsiqFapisngTzDFwhjkuIRZoI89f0OgPRu
xmi3/hUQ7+c1bFskwYnOxo+/S6uX+KV/AzwITK2vZTBWv0B3teoYn8cxQsKcJt+xqaq83DOA/8dO
h4txGHFj1vXpI5rjVk/o403r9rSpgwwhNYkv9fao81w8CqEvEekvWT/xR7XaoIvek24gvSPUsSNz
Oq80vIdi+RFiCm2CA7YdbE++oYSBBGNpLU+nMwDj5LaBCuu53Ilc1d8aXx8xSByhC3P9ttRUh5LW
rDFzh9OTl2bOoMHfE8StIj9kO8n2Tr0rTWrzb+ILeJGD5gFqyiei+/ijvvvuFvc9FzVPZjDlN6av
sFQesnw+a/jzXvTZQxHcqrTSTSc95brbjwoDyBZkNkAAUgHhfz0M8trvbDClG+ocYhToCgc9+Mz/
ZAeX8OK/mxQ4B17XQjhHkffLPmZ5KwmQDaGxJjjtQ50e02eakDbVnyLLnBjEIxAYY1+giKq/ioTm
cL4SgHZczpSaCga5ubjfNPzKI6KaSXy80SEdKALxxs9KA7FLEP99TePS1wq+JCpGx4iuhwdlnBQ4
11zMhn9nkRpZxc3GmDf2LPfPzb9B+LQSpdZ99V+XbCjdOB8i/aik33nRWteARxCOpKB3n9FqEovq
cXO06J81a19D/YjL2q/muiyVNDtVQjPsS8DMoo5L0Y7dFEtmXD8/J8z4LHQdP6bg581RXW56rrmG
KWb7f25zMQ6VsaLfC2Hp7aDXZswa2ym6lxw3ANYckE8xUN7lloh+82jrlptgOUXTL98Ym3ekEFRr
zLnd+pZNEnSpxUm1vpGrgEd40PMoGSTT/4gq9RPP7xoMhdJwpXve2ratZe2zIkVImjSreSgaOyFw
uIVGdS3NdLmeptLMLvXuZ3aUm5FCNd71akiAXe7s+SH0mxMsnIk2GAcCgg1MgEmPtGxfAs37A706
RgssA8RL8viN+m4LHmTeS22cK9hUuvAUsFV+/krqHYq7EtR7oRazy3uapC9cSsJ1ZWZiCOSEszdZ
64Q0oWLmthr1OAeuetvPhjo77Zcy8SkqAlg8sT89MvPrecO8y1I+PMQ/7WGFEhpNUisS7zcLuBDd
Jz+NXHhGPyN1Z8tpt66NO32SyNRIAzNSUetg0NFEYwAwFCUhD/eAkkQU53StBMD+VpEbJ+4aoG6Y
p5RQBwj+P6tiCo9OuDytte+Mys/cmohHoJi8VyDKnqSTEs34KfJ0l40Q2ssQ96649uInGmhzavdk
k5isp2WVCp58REMFW0RyTjFb6/1dhQ98t9X1oAChulye0cWzM5o6zNUtzLqKTGCZLf/bhQw2+n4a
qx0jxoPymYLk5N1EILhccy1cDW1qrjtrJ7/9kgnpvMGTXrWNKwyUMm7nGM+F5XDAppcNh2rFR3LY
q5POfj9gnQX3XtJNLZIu+HRpOIZ12mcE8T33HLGMvWZTHvrQ7vcugarQTfxa+x31owe2T6W7vBnn
BxZ4C4OY+N2YrHtzybwP2hxk3hsyFIsOaGY3lOlcf5OkRogp1zJFNMVmj2JotOnQTrbmQIT0h/DR
LaCcZOlCvgMWseHIFuVryb2HzEIIXIFxglIj1mUfLI9++DHG6pKL8PhKumjQlEmHQV0ktIidrbsq
wcJ0x9+oSEVL4FK7WQAhH6sqxgUn9jZXCMFiKk/e8qLYsWwWZktfm3QcNeWDw7DZAi+P2wA/rDfo
gCL/0fN0WV/lQ/GmV6d9KAluTNB+20qgzFZ6W4e8eTNCpX8vdeXf/8txGY8wElQJnwjgs/pIX0sE
WKdLuZsKzQ0GneHRJAnA0Izk71STGbg7NCPieMyRX2V0g9AsQ5vpCZ//LfrbwSlDCL7JlTU+Q3+k
zmic5/cmW4xHl6FeLVvi0khwuXo7J40T/argm4RWvDl3QE9KGF/34mRLAKarr0izSpIwk3DOVrjY
hhsyV5jTT1MP27rMgNUCVSegbevVk5L0ySsfKlEBL4ISer7fHNUCmfxumV10sYhxlVCQombCWihi
rhqifQxjzKAb014kPBjrhEVW0V92k+qc+yD2QeOHAKgIzTyUPbOeC4Z/VqzlLQPnzs/pOP1Q8JlO
IBJh1iHsZXkAmkQH0DbN3bZ1d3p6mcwA/Fe6fjaTBJ65EnOPFbjY1/4T3GCzj7Sm4RXY8d/t0njI
PP2s+6un34HHncUy6PS8EmllY3yN1DBApBc+CDE8MZ5lETYGrGwyr2sIVTzBb5PQlUy2hHlPbNyL
lyhSRct4PnjTO9y4sN3IRelnp2Rc26/j7vTaKokqw847LqXmzadEK21D1fpD54HOBY5EAbjwmcfD
pEcuL7/JhpIcOk1Kzk/C/9/Hffuiq0U6i7mO0yzljabS4iTLZG0K60J0cprDZesP7L7KmRDGQwxA
lmpZlzSGlQufRjVU2U19a3WMG6Fb7A1fH82O85GjYhxolaD3RinWuf926B6dqYH32BzVYYGKCQwT
lJ6xn7UvINYd+SmRdwSkgkl6eI8sqGfsWtgwWP3XRPvQobTeX17lB2pLw1Ud/Wt+SRmJ9xY0Lg3V
S1eqxJ8fx/VHtdm3XAMCXifGRr/wAy5mN3VWcZLOxowFSI2mZ+/WcBbAP+2QeSPesFLiXZ5txijv
EtbVLQ1nvzDBIINI1dXY7ZjQ533sjJaSJ3t3k5LSsYuLefm2tM2wpKL9Ax4cWISYCtfIq9ia5g2v
LnyC1ovJfakckIkztgIwUIWDJVXzBaM6xgsdS6QpFR4zNChEiHVmW3IbBtfj9siNeod//nOoUqcy
opoAO3g5XuSan8/0vuf4+3CR/g/dlSHkOfb6HLdtQORb/4C2l9BkfSDYZxvlyyN8mLkBlCtwP3iw
OQI23vBZhioacSUqKqznUDFsuN+qeTev8EnBK/Bfe6oZOy8IOq9HH74HiVUGz0PODmgcfpDhkiM2
vj6Iu/sO+lD0i35zBbnFoSMJH+DyI5D77c3L3Omcl1JdZufl3VHAytJtM3u7zmtYLpEtwDSih9wq
SnCt6wcTf0CllTZulmePv1lzRZcHaCBtIBxlbvwJJ3QEN65vHo9tPd+lsu6Bl6G+oMlFnkoqkmtZ
Ep983g30gckrsyEzPF0uNjm5/QmrUaklNJ8+1u5BsSIM3shQhaoeUJ5qQtMgxdbk8+0pIjfM+bO0
PkfqXGojVHW+WGLaDbYykLZdlXnBtBntQst+x8A2VoekMmHDnnaQVi2mEWk15lJ1afuowIkEyVzb
KMs1RpKHKrSDXMRzN4ZwKftYsVoXkZ9j3uXGJCx7KGtM2+/GbjZWLjISJXPYR3R6JKXvPPHaDpdN
dIATedB4mXNzO511d/llEot349WkZ8mV6aikknoDYMMe3WbUZWjacAiimmqzlvLu9K39EGXzCKli
Yw4dTDsnyTQrgdlk4wCHm/EkyMOlyMR+Z2B+q2ZAWY21sAARj5WbmXZcUGu5ZDZurBgNTyDBt51u
8GNwC6lCZ+Lh3GxTmCCUBIQbx/pUtsCz+9NFJRhT1N1YfuiPsm8sfQnLJ9F7TB2SK0o5xCaBdODl
OPNJIjRdGP451xSi2aj9R9seNjANxMr5LBwlAjD5pJbsJV9cVBPB64kDSWG58M83CwOPr+BblMIP
fcYAvo5dKePJmj/wq+BQKkzGSUerHI/VoI7hZVYlZrHEJtPDdkcrkmXvdVcZEEPi+Tcn5cmv+0a3
mH7JPtMXBLdGR5le7Ln53pOfbKbA4VEwEUphGn80cqpHfxzZEeA2Oxlj6GqHMvnXCo93b41e3Jky
WBcAhdIzCa9W7t7Ebc23nUzRc2Z7q/Te3A44bIi0DwsA2ZsXEI/0skiI1mnQMA7mUqgJFEG0/8tm
fgPzDYL6MogXc0XOc/OfnWiS0O+zoLa5ba6Ev+qiqRPaAqsjs6AuTNCFR4T/567WL2dsl+6T27Pd
lcDV3HN2xIVvUfPHb6wcBReavlmhSh5QGMiEVfwzDRIDqmTsQpU63fLpK+QfaBp4rA6FKT27/mCt
VgCYOyeUcGajGY6ZDN69VFAR3V1B99Ak76o3AY/h8aYNXtBtIZqz8AA1n6M/ed0GMTdB+8h6s+/E
vjj+5mTGuFL973AVqmIi97WyiNsyGgd/cm6kFqDJpDIfE71Bi+S7SLJcv1sE3P88eQf75YZdZ0hb
uoORmQ9RVuB58YI9ax99QRrSBvQ247Mp2pQP8i0jNnT+XZGrrVQAVHMo/sxCjGrZAC4z9KHfPssv
kivGLp+jdwEF9rlP4G23Td9oXnDhyqk6EKcy0kM+v5BPOsTXOSV3H1tTuraLKiDD/CYmGed0mW8K
09WtGZdZSS0feSwCihuaM27CtT0tkB2jorPE0aZfVO/DiV/qC6sT6R+vNylRKtE3yn80zbu3Zkar
H2jSSCpwR/lFF1ILQ3e3YO84Ds5RIbBYtCWfygv2sfdlyA6SbHyitKJSF/pEqMC/1NjPXn4cGO0j
8lQmmdO3BcuaxF0pFOAH7CIaJY7PGjnIXtU1RBrAhNrDQCQZ9Fe21OExRwbuQkjp+tRZ3LEGTNYk
ilNVqcBbhwpmcBVEUm0Hn+2+QKp3TA+m3hoovghSAC0d7O+rqa9N1WzP9tMMpTRA/mquTv7rcpAz
/6asuqrsO0q8Uu8ADyIqxlHgchj6yYAN+ED0Kzcg2xMyP8ejYJxsNHGkaxiecP0nc/5Qqlu0tlI8
orgnn1twGzP2fCx+9dc/vo3xxUL5EGQ0xPyCM8gOYSbFE85OlU3VpTqcO9JMbFcvE/ngkr0gMot6
wKjpQFEmfVThc+0pFmrVpJoQZGJrB7CAzPslAp2Y5HnuRCT0pp04x4XBsQzehIekvWfgK4GwfHET
UCR8ACBrsx6ZBfRM501A2bLeDorgdfoUtymoxyD1VXz1Z1eW6fnSWKDbetkLFDKRbsgTxNSjbII6
ZDzgbjjS111hgwg4TrttPcN43e92sygNG1VrapH0vlyum6kwu5+0N1PHXWWScZhQ0ApUAAsSOcBj
tz3jJsr5jCDaSCYd6ACLmorfG+uyrBVY9dQOv8x7KJ1jjKOz5biMoxLyXDbrIeMxDPj97M0zVtN3
w05AXnDcjJ0mndXuLvJVmlPzmDI0POq4ktE3TX/ezt/TfaXwX8GGIHpH/mXDmia1WQ2F/EIqXIRy
wewIb+1KOg//PG3/j6yN/Lzyohd9y7ZPDK8cpmeryUn4WGz9CxE6KTrpqfIZqd8NlLFdMNjov/nM
VLiMEYm293xeMzWBBGk6fh+NoqCRHD9uLJrAdxnZgta6+4tqkd/r0Tmzwtl4yCP0evPeukJaIYQU
TkN8JrRLeK5FcFRB/zW1il56f2p8m7tI7iL3Vz+E01CnZRIXOXSy9RgFkSamE1VxMfhnhPZbIglk
/a/TUPBOVgou3jcW4wvpBZyT1ODrVp9XpuBXgjKgoMXDNxOAKmUpYvanwKF/Dgr54VhnOh0k0EaH
239od0OvEgH1vhVEGVDsiFKPmeW0C7+v4ZLWFLe0kxWOd7avvEjMAX2nggc7sEC6t7zHFgtz98VF
41r7AjdBk3YSslL6b9dTZ3CC8v7RL3CWx4jHoOxDHnZRtWgqMcPv3FW1elYtd/MZBguj1oWb6rfd
KE0AZoYeiwYmA5tjXAihomw1/+W+S31nMSpAqMEw48Oybn/k/bLBdUbB1JgedOc2iXenyRFOacxM
91HgjYzLpBAD34x3TZwxJ8n4aXzBtBTxQ4e8xqWaR+lk20KTt+KatfJwR/9SNb3Yn4KMIEgET4bi
Mwr9iaPKFwEPH3JLGRoimldwP/vYUeMZV/FCAoEAFx9OHlTcHMTLzuUM0n1kYcngtN0A44jdlT0M
7QojktV/kbkvGUVJEVSmX2usuqKXYQv8oSfUIHaDKZe8xaZJIKQ8Rh32j8bdyXsvK5mTvDWvpesR
JzBxKgWKhTqH74AfkGiaKpt5GSfv7t46zrlqz08uOtjo3J78Lmj1LzkO+S3gCfqUU3t+gAe/Qn6C
R3c6TKGI4jxMAQqn9Wn6Lkode+OOOQqfORusbbCV/I5gsApYV/k+qjc8iq8QnNbp2eF2VIpR2zUt
4k+caN3BY9yJZ0n98KeHVhdi8q6EtQQvrloaPn/aT58fLgTtAUUbGWeeg0EKc+BT7CNHaIiNBVG/
d+xqLexW0tJo9zQioxY5eUMo8FjStLSObqqON+1kGqLWjDT1Ov/344WS7lSVimN6RS5PbRiK7UFq
lWEsPLMs/1emuFKJueu9vXgNhDcbNhZNR6sbdn5w6/Li+Ye66dExxbManf2X4g/yC9sS9N+Xr77e
i1VpdJSf+fftnRVpNyBOWL8uYhAkWPzcuRiHNKyWOhpXGVDOQ+9ADAZ2L/J9LsNvCk4Qb2TevdEs
3Jo33BgwVhnPDmBo2amuhesit6iuOc5MW8ZSGvJLx1XkOm4esAJuALu6K3lJerLS403hzskjGof/
q1IIvKKOXrryzaX8VTcP5z2T55Z9WH2oLPUdd2E4Cu+/KCaX9qSX+LDxyURtwhncWjGYBkDoeU1c
QOmekGbZxOlCifUquFNAntCSsZw2XM8Jl1bcuPIv3oh+b3sl2AHcQyUU5IcTOqYoVD8y68F8DNTq
8VgjBsWlFmrQ5CAZzxHRMgIGHqYhTgI8n329/6AzUhgVBJ4K43RAIWNr4y11xyfAQzSu7QNQn0VS
uXaN81UMZa8XDrkBbsDdxwlNJKHe1oXVh/zpLJMX6MsBggJydUazZJ6O6S/udqZRbCMudfaZze2T
DiCYQEZebDxwQQunAqxyBQHdusRfJLsunecC2czN7iLtdjHmh8of+fNZ8Pic0PoWKa6Re0dEaMn4
7/vgctGeQfH5z4K8bBZtMyNMSjGmqgJzn+ltxKOS24h6UyU+xKx9JbxhinwRZxDmmpeKRrOqZwqv
AF6QCenizrtUvp2Uh5VbBkD5cLl9mLNPsThCaqdo+WtLW2f44NJbrQ6pfSqu4CkErwp4dMaZ+Bah
ypKKjS8KYQUuN1KLVqkMmnCagXV6BvMtIdVZ3qwiY88qsbGlQ6KR8BDOBX0epcvidrfnTV4+P8uo
nJ1Txa3pN0SWi22NROStnZtZWjs2qnD+kQ3S+69+2CH5wvqfUNgvHciLyCd5x5CLKmX9Sn6tdK0N
wjR+r55lafSIFtha/ISkBUFw614EqwE1qEu8DPt0PZU0F/wEU+QLp/iqsepLAlolNGoy7/BFiyYh
dWiCv3QGH4XHRtdU6T2EN175I55BcieOl5AIh4ovyXADcDW2yjkFPd1x7PZVuXfYaWlbsUUP0oLC
eMq11ZU6mVvzu9OrPF0R5lESYQqEBNJV80/CiawlJAgj1vlivfojBdih3ouSN4/xWDctoUAPXze4
Z0e6PyBex+7xUoYQT0mmgUtrbA+fjqXTdQIxw7iBP2QjrbdWPiU3lXfOOBJnxfTvYCFG3gwfExvi
+72MXPqI0XjGwCrSZHupzk/spgqqbS3jURRdzK4awpOZVVwE6xIgpE9V8cXDVYCRn/jSjiNKK/Wc
ixcmgtLtsA3mjJXZ5L7CyTwFREi1ff8wVLzvXuorufDJueihRYUUBd+ksnHl9pG4gzeRtKTZvZpm
WCMtbR3e5x6a3slIugbCl0ph14tSVe/IG0Dln+HAmfRCLrWWvFjy4KRbdDdkDxFwlS9yhAFvEOV1
PkGBDQ3rzxNtwZiuv0Rm2/FuWU9T9jyZ6HvsHJ5BolprdC6UXlnUgHL4lEZBpqNca64pNMsknYw7
7U8aWKBMCuKcWIGNfLxyCXtpL4ViLny9w4kavX+1Lwb56rwJ+wDCddwFqEuc4wcUQVhehAvhFY+O
8HvJlhCF6OD59OruAw0F8I7YGBjM98UEvp5V9vC9L3P8u+BRey16a32/DFQb70BPUaKvFcfHiWKW
ikaRY/TezLTGPZpEI9DobUyrKa+jpw4FWy5B+aiQDuZnPRnSLqyc5h0sBduzsZGb5CYfXpztyxuF
yhykaCFppfhm3GhUbier15HH76Jsao420hwfJHPln98gE5kehnZETuZDIBumG8X41eYKug8rWh2D
SUTTSfF5QI5LdlGaYT5koTBGrO9gGyZ/p33p4evAGqwcoRoJCXUFkRJgdn+dHawyCiwQ0+im/ila
bnnFNNrBMxLAZIQUGtmr4JRluO/l26YUoc2eZK8n/O10IZZOeKRXfd3Y059dakZKT1Hvt2RqqklX
1vxRrvawAAG7/U4OWlcTQ6o95Dl8ECnLtnIjbGw6tLbNzAxcptoQdn3ErfVp9wFesP5I7L8aVA1o
SoUUYZ2s89KaGWXDlgha4YiM3xuJiAq3y8ov+dgXDD64hPK9YA8GiMwB+OF/S5pKw3nc0ixI3bnm
CUACp/DrGbZxfAIApCPEOWuLN5f18O3p4xf8O9pliyQr9OFmpO8a2n6vu2t9m7RVlykpc9xKCCSu
5q4ZRhr/jjFj3N9nzLnWaAhMVlVCDtjg7AlqWcWXfzfY7hosbfkcCDi1CKMb56ln0l0ttZbM6Qiz
JWFYlIDlAA8cfcWEz3rDi3sInLWKJjuzoM1F5UqPRhJyCIWMQZ5iWcP7Vg4oX3VQ4pdaB5p3QxGm
bbs018wWMj+3YlPS7xbCuq+9kMwHzDouqxl5EabXtIk08UikiDtMcXJKqmt4Xnlc2GNCwbo7G1o1
wiDusFV0kn1UmVoboozfVtc9MeMz9kJNnTD76bDKXYiigGlqNcLWlkiJ36FVMNsglvW8gFmkHJ+r
0FKOlzXFcHB7WxtY8/i/99KqwkHXqjfO3SymhNNgBdfh0OAECh4bLz9RWdBG/aUZzjriiqd5/jha
83ruFb2gBFAI6rbXsbtaroQl+ldk0rj+Z2inQUAFRT1c6/kWyYnRjCm6866uDMSforj3r9esfGZq
vHVAuwUoGfVhXgBwM2bSuXtoEuIaxV+nO28wuen9s9x1iVNPgeEK3Ir6BFrcBvxL92u/A2EeiSeR
Ixa5I8bGqF4llOH+04LKL+Fl1NYkcP00TaVDbBJa1ZE3LsKAsML0P2Wul2rFq8jyDNh6Db26uZAA
ffpbP7KHtPDtiwAEQqoJE8/WIK3FIr6rbqXXnt5qPfig/+6rjLB52tsm3y14rdmGWN7bNPm2S2vM
N0KVJoZ95IzgjwOI4yzY0j5QVuDfQ8WLh8OmFI8hYs7ZitUG/1dt/WUD6e+Oq7ZqV+iJ8ljQHBU/
aKAJXMdcSL9u8JKUYdJsdl5piH8j6/VDYMYNILgiU43KfJB9LOEgIRwkcdSu4XBg16Pfpb+jBwxp
sKvfNMhnW84JvwKHaEp1N/3YHsuzhsCDQeHFoUvJNizxPwjthaU6zyRIAobiDTgfcTvER0UPO9mg
GZ46MFvbH7ZS4i9yQ0TdaiRY5ug2JJ17ZZYqBQnnTWEnzncq8ruiafYecgXrKJiuP+aNbgpgiUT/
sAoz7aB8PxLNnNqNkDuUzHSknr63AbcFrGXIZLjvDtui8q/+PjmwHRVWQOLefn44dW1aj1x4/YQx
3Yz522dnu3hM0Aap0FQwRlUsKNKYQIxVHxoH2KGq7m8plnZn/+emuA19eXdjDbW5+awxgKBwlFYD
FdB51FPs5g/Ov2nNLuMWWgSTKtigaT6wE/QkCkffR9VAIW6dzRzcgOT9fubU5FQGXAtx6LlL/7bc
bj8mTRU9k5lKgCI2uJAFhtOyF70MB0pzfM7l+O3s+3qinRj6rsDLwTLBhzQCwzmnAyqpabMSN4BG
o//f/qCCGJGgy904whPJdpVKHAhjYq7OWTEO9X9xu6UIoijjRlEYWE31T0FO8WSOt5+tEsE93mH8
PMyxzzd4XiisWnrLmPKUoZubeY/9Z265oa0RZTR3uaTA+hu9BnsBL8zM58ugV+whMcpqPkTYXGgb
vx5rZVfYeBUSMDcJI2PgXdWtpP0hwyLNoQDUGBdtnd2LV+fP+PjNj8AKYrZ52H1wBmnurOtBLn+6
N2fSCrdqC38TnjymGOmeBrLlVW/DI917cteRiwmQufd5ccLUN94pNAtORWsK/USiRt0KqXsXHa2V
5MPPLcaXgRRGpHUzE9n2FYsH6FaZSS2R8PMDxIMj5QLsz1nhKEOMja2swxP+J6fKlBK3YEGsu0ut
5RP1XW1V1st7KdlVPMl3tceeBk1rSjbBAMcHV9LJt4LOKEvw1JgNQg/HolHEzrV1bcyZVZ7VRpSM
4FQUsVauWCS1FrCaPH+ucq6m2ZJkj45WzlN6rIYFyWKSgAMuFdvbJQPNWz+pi4lCHbYn2Mpq9tkr
tkT07mIN1LTzzZ9VetyRouHN1n71x6raVjddtWYkWBctNU+mZsbyLrurd6QKhDv9cLMfVTLFfWFX
PdVHUESZSEOGBJpye8cwvo/r3FJ/NgsTiMGfVEit7CToFDGpP0uQe66eVElMuIidUDEOzVpJ1p73
AnAcmopZoKE8fPRRhyWLDgsD4iprWS2NgbD+gLZd9mSBch/Ua3uRMCUxIFZvu2eXcEgfu6vW6Vg4
n4ClRjLT13sf1EjQZ89g+iBEYpVNHZpFkztPE8TJTmm3x7OL4IZxFsIbLJVhV5tuFHJJ5qohCKfQ
EZiiBFvGKcDgHM5BCcR6SyNIzvbsnXDnTp+1PTPlckQWXIjDdnUBu0NdXXnlVMT3esiXJ0Ejr0Gw
Flz4s3ZP7yEJpWQq32Ftw8/ZoqSpkiiVOwKdbq5NmkpSaUpWBsf5L3Gvvtar1gt8BU8kjMkUiY3t
QFqF/S0eHVXMot/wyw47S8K1SsXXeG3Umzzk/alIMDXpYWwCjkXTnMNH5StHP/YCKZOkkTq14m8L
UbFczJvUmBK5IP43aNRocJqZH1u46brhOjJ1puCHiZwFKjkDeFDBbXFEYKq2VI791tGxCHLml60a
w51qWlh4YxA7913LW+E0VzTUtpj8enSh1WAQnY7Ffc5oiUorEk0E7gPhYx8wneLyDRu7yoH6PHss
oSlIw7ycsAZs4d6SFZm8Hz3nVDG+z0Li3e3pyjPiYmmAY8EL+XVch5o0ohXWoqCFntqKAopeT7HP
RcVYUPPo+M8KoorN4yeY/t9TbJrp4XwA0OXgM2/4Pwaw/nYWvwm7fQFWzdR+VyjpvLudUBzYqD9e
k8/GsAVBOxKkkY7v7kjlLwuJ+8yFxoD7FsNiss+JeuAs+aff0AxDof4GMA0ClcTYh/zGw57N22hE
qPg6h55WsYL2NdGM5oGhcJSUgNWKNIzOU7nh1exCv1rJCUbvSeMzphOozcPxw+mnQIAVL8ekQ0r5
u/4wkZb/P8aSdkIQ+f3XDcBOHP7lI/cpmEBQmw+/7Zp+kXmq7ct9coCtMinWOZo5SDCO2ykSqXIS
VdC2Qnl7OyltXEjRazT5+6zRqrhBDnSo4hiMn+cVAUmZ/wNYNr23e329P85gBLdRrtgBnlo+CG63
s7liLRerdX49ooGeOM/hw/gINP0tQRih163XiGXq4m7XhJm/HTnpsc24YXnbxh4uRatdCgSiiRJJ
x2B+yqhdh6kheBH5M5I/FTO0CRW8Q/iYP2TZfruSIcZFYEW+oPVjjORDvY5Uu9qHBEGpiH71XGC4
8J2YQqYLKn1DHCg1QbSmc5yoyDM9B70rxFqBfG46FOUb7m74qzlw16+9fE02AhsJlSVwHTdtFTdK
haui81pfFMMjzQ+F7CYw9XUjcAatL9Sa5I5IxLdxuhBcOqgX0n3a+cASxa6W5DH5wtn5KFyGwy4o
7yRT7TtbPC2q6Xz0xmBeDfX2rLEsBBozdTER/B6d0ndyoikEzXHJ9ykxnFyrVQV3oK48MW8EPQ/8
+HGQsso++DXT9Xgn0FItI1r1tViHV21NdtgwxsmoTAl4GzIkylPhFhQCpwEXaOjmwUKYgumOHvzs
SfmOJ/xPz1SfpGf9xtgTjNCGPasMlpNAsTch1UQXTRJfSOINkWFTd1mr9S8r4U4DNiYUOlrOEfwp
nJHEObdfDG8i7vTNxnwTUD2jS5MEVtYboDHT9lbsAv0LkRXfd+zQBaa7GMTHYHp5TDwzfdDbGBfH
UVAL0ZlfBKfd7bQsp2E6OoJO0n9o8zZiIbHIu6Ni0nlKbzgG1X0bQiWfve4/moR9smoRlUP7b7Lk
TlzwPmMHPC1qIQ3qxuumZjMY1WFEfGQyh5PtbTI/c/JCKqKy5Y0ZGju5nU5LacSdpIjkdfR7SyUW
ZZawQ169pgG0y2d6drQsfZ2v5cC8MkSkmGLGsI3V0GCqGJOyQEQJNalnBJauIW3eMDpoNf5tj9Lh
gTtWrGXqCnelgF3wuegi4DSZ6NS1INIc5zaA4axqROoISX7NLgtKxaHSX+5hFa7GmE5gmSIiVTPW
+FtXbU9cef6iULYkgVOgZpD9Q7G9eIRfgd6lXJaIq+y4GkckfhfUl+3qgMoZNv8kOc/76XkPjP89
YJhDru7zr4T7pzogAftYo+Z9X0poGGxd1aVaANioylSwUZqfTNYgO+9qTGHbAOeaTJVMegtA6XzK
0g4iqKYQ1bz++Ni4/6ISNdOfAV51cuQ9ba93ZtFg+9qjA99yhR3ZSuSpqT1YzJ1bOmCeNaybDHix
mh+tMbKEPdGHGybB8Os/nJXAZ8R21AFODbP8rsEF7Bj11kMdZLBu3wWBdKuycHnDNXMXfjfTgg7V
Jbldv4NoB2pIb3ZcFzNo2bL0rPrp9XysGhIuQXRzqSGutu5ZtMqAFGI2LloB9+QedzHyv1CfaUg1
DHkJo2EeJBxAymI67SXognkYUoc94n4g2FyB9TdBSY6HPW1gpIspamMgt4/u2rCVPephaJOyVe8S
+ws4HZu3vclMXH+e/td5owaid31r5Sa/NQB0hdhgxjZabQ5TI57JJ26vx/iemDygsKjHREMzwtkC
nbgHii4mnjtXdPr5BTr8PInakcog+UPOQAW5bJAc3COMroT2QcCbfSYvXoF/4ejwB7MsjysrTxLa
wAWWwsAgNpWP23+wlmQG3GVMvHZzYVrrr9lKCvDwMowwGWkAQFnccNH8zB59+dZ4JrTtfwtahZg8
LL5QQCF5AbeyxNigfsSXGk9+QrzLqKBxgR8UbgY6AGN+wNEXCJrihVEyJ8WhpRyagLTEpw9M9pIb
CeMvnylmWJRH3kZRNZR64jpliDCI2BTmqiyZou0xI9eZIkEZrFzztfZ8rumLa20z0WGc466/9ngq
4CXzlUIZh4OckdF7xGd6OgD0DdRYHraw0bShxgcKM4n0zOQ0sBVfrkren9KAHmexi+gq9EBTQ+W6
hNOIyKR4YQmpcs0ffJWIiEn20p4ysLHJGWsH8qptH0gaCtSWCEqm07SjX5Aelisd4JFXWH32oa48
3s7AiMZ5oQhbpLSjuuFgqXbRYjFQxrGC1vVVyyHSA2xh9mbe6aV2/Zlk5ZFJ88gcL5CyhnMuN3+H
mDp8f+4xsU1X7CYmAL8B75qIAHXU/TVhkTaBUF3F79XmsUHPpl4W54xihnrY9umca4Qf59YdXiG4
ZgZ9BKSepj7pyk+iqW6F9vprMavvK4H8pp5aC7r59wZBUt6UYcEVnBzp0xDUSA5Ns+2pAWMBIyNj
pymejP9jJMCLYNEIjlAA7pJjv8CBxlSFA8xftjRiZrPCO9OtRwPF3JHAne7MUaatXy9hUIE18K37
tKY6AjnzxxQjE5QSPvX/m6hrjPwmyzxcrPA30SxSlFIsGDIetJ6NwwOe+EEud2THntHrUAH0f+9Q
TF0hZ12Yw6dPnQhekbfmVrRR8tn0S4xinBJsuTRfzWe1o8Ads94PvMXbbo0Qf3KH2vpvt3s7y242
klAX/s2qz4YNhhbrfyT4wM/M5DsYYFA1hEIb4Li9j9K8I92YvD8+rKDAfZnAlx1rvpWqPdFBn1t/
JjUB6e/8ExcrMVdM3A5I06jkcBqmE6Su8riZlAjqGx7U3CyKlhNxlF2fMT6Uogk0CHOK4OYYa84z
FZJAOFcO6Ff0bjrb35bbrdFupOZNzr/93W1X0veesHlBDte7YjXUHzWQeePuOvnk4kfM2eTOM1KD
C0/gEFKAzSnqmj+cOKCobLkRCbaSZuhM2WewH2A3QLc4POmP1YYq84QUugzjIX0GPPsT5EatnOqE
RqXcoDhNaABLUBQck8PIPQJRo55uEW6jmSnQsgb7D+HLyoZVnabZbFCsxYRyZbneVSRrWGt0wkCs
h4SUEF82FskVRI1rhWhxxCAaF98qF/zVp9u5mvIeJ+HCRuveVy9/i8i83rEiIioR/3ZZKCr+su+J
uT6BFyMlgLyi1KBFEjn2HOd9LZfLtkOKxdwCSrJ/it4P+p/4LfV2jzS7omUrDF1Km651UGtTZTaZ
hOmtQj8FEyWJAimXnlAthGFgmqw2034d4H64edS4ibuGh3VuFZPoFiOLbv/Iwllwp6CDcRER8DUe
YfJ0WpcsfEWP1P7LrpzORIHjahmhjnJFqe0oIj01gNK8RolHuEpsjiLGHJ5U+Vp3nxKRkQDmpzqV
S5Ch5LxP7nPBXACC1TAN/izozsnfQ8Ah4TUqsLtSioVoxED1Vz0cm2HplZuXpj+hYUqmVg46WHb7
DJfcnnUnqMsAIE6IdPVg7bpeQFG2zjXSr8oDYVqLLWmDfEJhTV7mjaYZ7zgOGBPYW/BrMxJ7fxoI
iidezjTk2L4TTKwB1B8MAvuKf6xOuJGhHqkT3U+LS0I/Yo/3zTdPeafvsDOmGcH77DrBHGSegb8J
eoPdfGuaxSnTZKYLr+errULdLtSDmbHi0j88CAg4VzlKK7lin9nOJGQaC/uhDu9pbyYJ+Q5OwpQ9
RbduesHReopvyyn2Eugm0jjB4l3RDgN5jT75erWJJpy6OgKVz1/gBvtVhBY+RGd6WcLGXDD7f3o/
CH8WMfodWtV+4Ma2X9bbQltflBKd/BX7YpwPrRj0hzS9D7i5hYuHq7X0fkzsiWUG1RzYzwh+EEE3
JWviEF62G2m7j3NeBttKn7na1czSXhJt+ZDDDVKO54+EyEbMLiYScQ1f+m3cjum/B5HLhuOBBAd9
Bs3vqhB6cGGX35G3EptERCZDjFM2n5Vejrgtfvp7K8i/ANHQfkdgVpjBWv8gpKAPSHIjkP/O98UX
dLtktGlmnzRfno6VRXsCNBJ2BoIttTw33m3TPoKrwPzjCw5RUCOP0omAcF2M3bfEEWNd+b/78uKQ
c1DDNrw61/XJA52YCS71X6yeV0fLq2uEHbBfBKOcKyyQTIPTmCdcq1fEKUIFLp5xONhtGK+sATHf
/zWb2nLRsz1+qcpOmIfRU+eO5wOAA69A2V8yJwrctJUA9rSUHzKBos1vSXUNc1VU26Nhssrva9QO
R+JmcO5QjbhGhMuLZ3zeGmYDhCqubhRweBL1UZrt7D90CKCqwbFKfooPJ/ru1Mh7fpdVEdibxZ0V
2cbNW58a0V7vetmeXBI3jbgeYkeSFUrljIMtDTwwpDAyCFSgnY2NU/tmZcMK1UyiLR96e+Pzk1Vt
iEYzgzMdgciXqqEPP/V1JgPA9zq1muw6kfG8IdC3dbHBUcGa9Kq5lJRyyt5leKt1USBAMAS+A7Og
oe5NOtJdc+3fiGhW8UzJ7IfmB33a5pftbO93/Y59IMwlnyop3CwLWA+r8zOW30+sbsNzE2nuF1JT
DaBI+h8Zb7MexTZquTGdQnHnMYR56GrlnnxnG6obfRPWBFYmlVH6dur5fTpwdIxX3IHdyO8DXgz1
LHZab2RLhqaprpvKLzyiWVYWRWcyNNtK7Axj3b1o2Qu7b7T5xd3/mdw1Ju+Urpd72jHWUkfBaKBs
AaBZut9M5Bp4Ef/wZ6862bYenVzqdcr7cC0u4N+NZb8LqQkz5uJ6lcO98SuEjJ7+7Sp3TBO6Uch3
5j8n9zMH0DuZmLGuj5j0jVBb3S+8ka4E7E12TY+MWCh0zjVAGZpQtJW/5qKm6BvrlM6HlOskiwBB
e1AaKpFEhz78G+/kt4DcY00uHmUFBTP0x61PZwZ++ShGov8FZ/MQyrAjR0Kq3VuLwBqG0zTvdVKj
/G13hN7vk51P+Mf9V1krxpDNJZFguDik0DA6qdzJZIT62aB5TCUHbar2t+WKnaYKQkLk1Vyuksrs
UpnhgKLx6uzmuZq/FKAUCL//non2lmeR+J1D36kG7w5HtW5arfaCQ9K+wwMc9sgAdQwqcANg3ge3
U14hkY/5EGj6WldWDdMVUR5V1nlRdyZdqvkxsGgwU5UXQVwg5eBdlI9WcVgukZq70/1/SsQWg0P+
153OJU6ORs1zcWRp3ATvJfn8xzENFFeWUCU0TQgRzK+ZGRZodkKH7B+S6NAbCQWV4Jeb8Wedwiy4
TRdmYvcVm4g6ZHhjt9nIE71DwaZUMQqGfsKhXgWfsQAwFzgmVoZXk1QiFEH5epYdV/sBijZAN4Rn
Dj9TdDjF981JtaIjIv6Q3leNe4dcL8iPxvnOa8dmPG4lEQ06ZB0HOYtvarXszwwbn7TeD6dF+hHP
l9kyNoiGghMdWLubJhqcoH7s+xQWMnXYYOM/IxM671KzDD/netcrCTkmz0epwj5e0wrCvmLNEwtm
mShhEE1beCPCOS29Gukn9XPh49A+bx6Rczmo0nwB7E9duqAOhzhzc0eeDDNUjrotQRFpLJwC0PJQ
Ou7wQfwztDPDPgdIktyPiZvkk3/Hjr6CLNLPE15mKe7qYZE+2CMrXdl6+H2wR+jtgIonjSV6PPwn
nKbhja24pAti8QVOywC2ruPWNFuikhoj5EuO3RB2Bg1z/LLsSe1ohXSx48SBW0O1/t467xW7f2uB
1XmVmvJ+xKNQwsmNwg7sNufJHL6ALy1Sy016k1kY9JuN2Hd8anqcp37psb4X0QHpKdbshMAA4vq1
mxxohB3uNj5nhW9TddPSOkE3eSXoXu8NmQclHMm6wjDcp8A4whz9CO+AC+u4qggRiXY9K5eZHDCg
cwsEweCvfCWeKiRc8uHwm5oqNgDGxWCwrj+0ImccuL1sPwOQPPXdRjasR+U/GlvpZK/kwk/ls9FP
xVrgxpibqrUmycCn4BalCMGZFVPFP/2wRHy2yH2t0jcaFoKIZ7Xk5jfggoFaDLYAf0cuVuZZKOY+
0GWt7isM6TgkdQKXZErVEwP7VSSyLAFPALgBmDXpGJdYQ1XQ+bLvffIoht1iuTpFSgRnrPGTdSzB
a8Bna41YnPRzg2JbvXrXVRuMq8IVbDsgfh2UN4kYW4eqyRdAat+IVLAIveEf9NO2dsDbkKeyzI+0
uPyXjJHk1OVAuqWrQbUJgXiWNEs7zrNw2812o6GviOsNv8CE+VAHYjgB6hqnNMJlenEQ9iOv1LD7
pdxJnpL/82M6/cMLXmNdY9vPKQhLP6a5l3c8qTQ3jBJfHP+jw1CiordanWYZjyM6RaBMRYKWdYJs
so/3TjOp56R2euczyyPhf+kMElb98M7O4am3qEhe40IsxPW0JtL+EgGU88ZGJxLhDJXNndncTqsy
fkHY5S00otAhroAd/MFfhRUT90DqJ6zC5z3417VphARHw4UY0iXROEOMiqS/uQ2/PDbxvaor3oKy
DS8yknD1h/KDGvJzfVQUIH/5UvVxi6e5135ker5rvQzvxF7ww3lFZKmhN+TJ7xg/Axh0OzOoBaf9
syiI7eXg/6Ab3xQtQApyXzff3INHD6ftSLmQfpu+l4aR4mKW18ZPWLhQ9nyTSJ7J/M7paVIXOIta
6/O4hSRsrVLr9p6R311CYkTDkM7s02e9ZpXBm31o6702Ehsfi9sOjmJxs+pVNxfxWH/94ELmGKqd
oWVbUZtBUCx5aEW5tMrY0Ly7YnZir9JAoQ3IdOJPQBnV6LpDcDP5qhbVyDkKJLq7oWiOvjRsN42p
wRqtmsVVJKyMYM3qvOOrmIphxH8AnzUFosJxwAJ57fp37Y3ctatkMR4paF6GWeNbHu6J7NeWZk5k
CqqIdz/PbPUcyf6flYH72oclxRJllcbcekLTlA31nALzCliFxQeBcGOnGUwcGT98DaXiQV+XXD9K
/+LQlpOzBDUtuHmRPdnD6IOkKIpxLBF0bCEySbPnLJOZ3MvsJ1FibXWGh3BbgTYfmL/4bmsrcPhq
6mtl4jwZVrZ5m7JyJE22DIGMsTd/PH/+76pVSpQk8OTe576IdgUOS5OCh0z9smzh6JgCXjaKBR+s
IxFyWJ5zvYw3GQlMvpoRjFNiasvVNxN8JV/tYEUyEdJG8StlWe4W+ZHrF3QVjyxOt5xOwe62gbEj
O4xyzcGPTc5c7fyn5c31V+0Fa2RqVHxUYaRl+mzCKa9QCu0bHTSJudD3qx/TDe7vLCVQkyzuC8Hy
CUMrd5onzoCeoAydJ3v5njN/ZtgSu1Rabck38cWoZUVSc21C05rlkc8SjNjsWoM7iI3NxXz50opu
+IaLhyWadxABuxKFOP3nCq5MR90WXKydcnMR2djSj8RzYAP60sABafn6M15hBDkjKaUbm00t2BFs
eFwv3V6kG8GBnQWBo7GgEKiOjyEM0auEdPde2CD+fMs0YgVPYiVQ+ioaXNc7Ng8inhUjxN44UFmu
WHb8sxbvG9LqphvYrIiher3MUII3GECjocray6fjAQ3F6zgZnTW6jiIj62mQM3kjHWOAG6N+jATK
eXmr7g49y/hJpcmuJ8MFnyktexok4h0xpobz7w8t1CYIOgqoUUTz3Xq5ROE0MbKLLmz2TXYGSj6P
aPNyHTKePJ13tDoqrAiBXnzJAa9xrPWbGM2BFLn2Gtdxoabd2Eb+lridvWhI+zzK0EofzITA1N2l
ah8dAR3kqrk5LT//Fceo/6lFBEQIW9qKH1JXOYytm6Y60h4oo52bu20aj8AeMet28pwgDHeh2LIL
0fPj8yOhaZhHjv+sBHwZjYgTWifbEOcjW8ELfaR2i8dbG+FJZHCoiIx6K7tcaGSYwNH9u6sx2A8p
DP9WJHdnJBzitTUtoDZRgXdGQ+59gXOUCv4nK06VPlIC5RSfzm7HfVQ3c50n17+CfTYaits/RCks
0EI3tV8kIxYmF4MPECLgrhsfc0yVX8gbjTBJRYEgql00NQuWvtX5sKl0B4kRwBIzDAMExNfovdOK
JVVSD6Ll2mz7XpFN+6LqqDUFTg4wYAc0KbRcTDpiL/Zy5ISd+1HQ5g1ZV2/csTeqpH0Nnb0wYECq
3aE3qWNVyLegzWrKFeZegiV0c9V9nnbvOKrktvg9UjZV6Xe311YoHhJrvl4oiiiCU9ycCdbZAlUm
2V2N9iOs7vPgu8Nlt0ypsz8DMg4no7FI1KYzQsw4BhIXsnQ1dIWqM8NfSv9jHLb34yU81OTiIHNm
UEOXj9ISfGinUCElrNAnwaep7DpwpFPYCjoh3rpDHfOUXbcq4uT2yMTO0UtkWcxzkW49iUkI0t4L
seHNz/nm3vLWgosgtDQm/GkXDZzDqJHnvDBQ6hiMNUKebrhySXd6RxRnJ6WOfQVOJY5iV/YFNyA9
katA54Qd6+i3Vf39L+58vVAcJZ6qiASlZ9zr1q8xcv64Nhs8F0gSwot8yfE2lbKEwiEzVXlyx6bH
WzfuQ5dfNbDT1B/nlWevGgt0lHWKQAzSdiOeLwOXpZ0ttbbdqRlpu2nVRmaVdLcrpUABgBPczUEj
ILuYZK6iNCt1uNsgoexSM/nqGkTjqYZQwJhIPMPlgZ6KAx1rB//w7jYHUzIyqQtKVTQUoOkE16+z
kBIkyG8OWZt8RfLu7T28U/KbmnAp9PiXTuO0qFwwtZihwsf+/R22L+r/+KiBCbaUtSnRGIlM58PX
uOudTZ23vb8ZdTxTnUzx491n73gHLKcyRNqtXsETylmA1WbG+8P4qC5H/cJdH2g2G/p/2ngOqE92
oM5w8Epc+fviKsDg9IFglkGnLROEMmSOloPMsuYJAps4/bzdbszd/Ycq9KZgTV/apRlSc9Nl10F9
MmlEN3+uk7yFLhz9XpXBn+F8WPmBOZ69WUS04qoTsiXkUWbvSiCZKeU46omp5Nc6m9M3QBwmGm3a
Z6caukGFRlUftknASbWush7hkjph1rja3Vk0noUt9mQAxjapkzzC9BhwvxqOeIA9KXXf7j2lAZQr
CCGoFC1P/yXj1fTRnU0T6JCV9byHVyxhf8BLVN2bUhu61u3DjGbzwM5JMvikCBQgMY9g6i86P4ql
Y6V+cGB4yNS0HtJGyk0d10nSdnC1fuXnrLINDbX3b2IAEy+ewsoDDflFn365lpz2LYH8CancPtvm
UQ/D0TCLd6KCJCNJWHFYvSJcK8BmoXsUi0+UjUp3TXpsRFXaWmoNpGTTdp2Dx341PpEY/3ykso6W
YLVuXQVIYjBvbnFahEjsAI7tKFSuO0yEXhh1fBckuExz30vrYqLVRz/KI0zgytzGRAjfB77Um0jJ
lN6CU+i2wvJxnsT3E9vwutL+M6sht/cqFVs12m4d0LqlqH/5unwYLTo71mL8od6rdZQ55i3nXAK6
G7vhboqt06yq9kuQbTIOfvddmB52mVLlu7z7NWlNwICI6IauWZsp+E1O1ol62VbqLcPX8+/11sO+
G4pMfue6Tn2CFgtgQsZITmqhq6Ge+rcnLgLuLz3+sa+fauKPxPZRsksDv8uQFn1+gvfX2JID3/v/
fyOM4y4f9lbCvBVhEylTpT5kbAK5sBR/ob2VZkTuZPNTMasbM25m+fjc8x0NJqB3TkoVelyg5Xsv
nviQabxPx/0vhS09uaVpQL+G34m2kW1Mv5vvOqTPLfDd9NZoIHFYq3yXTR8DetxGgPO8tiHF+tKK
D8y6ttGE6eVuq9CHG1Zcr/nKXwNR2jSo3k40Y/kr0s7SIRTAi+AOCYdjSIwMQ/98so/5vbb+IfeZ
gR02x8SGTh6E3cXCAMEKZhKAvp7jI3E2+dTXFJ69hh9KWvKfPAo5hOeW8JuSEQFlxV9ilMYJN+uD
vDYhCM+zTzu9KaTxRABu82va6zwi1874WRpf88l+Y5fKYlPO5JZu132SpfJIMqzUTMGz1YDBUGRS
WdAiRxgSlgYfpwlFOhCQElFXcAn4sal19XpuQD4ZW1yCfpjl8HtIidrhgfXAxnXRrtx6tkq/goNp
pJbSP3yermp8vkQorUTpC/JnWd3ebO+DMY73Duok8PXZ6j4VOrV0ePvLVVTLandrNyKjEs6O6NDQ
OWAyXVYG9YAJdGuPrdApKR2X36iLhABrFmlMCbisV6oatKjboruNaQqk6ohiktluTAD3WR7eBlSy
p9HtWY0leZdMU/hrsD6QJi7OzGgrebSJxY3XhCmacGuwCk2rq9rkxFa0r7dl2fzXpazzSxhv5xmX
CvdKmvw4mSJxS3/I5zskeAWmfIN/jcEfpXq9SlyNEiYFKL7NGwUI6+wlRFVPORys78HSc+WK8qhi
PuNvRZH08yzo2d/MzuyEgR8x74F5FeRSi8bFquOf8Pydxtf/UECEjEHg3g21OrH4UImRTunFgBD0
WiMev0NEoCLoHxMWww3QhpAJh4bOCpwdwblHosEptXOXngvNoxniZ+zOZFJQmqWFSQGcU0fc68zI
INoabY/RnCnV5uBk5BD8sHUDrv3sb1s2zsIz7m3LOKnS1dn2nTTTISE//MkdvTEJrLzVvksjPaC4
HoW1CqoalPhGSlAjccKVCINLBRUjxRS+g/mwI/BNI+JnVW5+xouA98BEghxoQeQtNpYHS+P3QOvT
d/ts1MnIfD1oP2qusrDDaiyl4i4TUXnCO6Qo9lWcTB/akk0Mevo+Rvm8AB2W7L6q0BsDVc9YGn+5
kDRC57GaAQb3rYxgI40/IYDFIYDxKhDx2rww8uMolw3SnLMMn6nJR+0aP8xVKL4qTHPc1UmKz5Co
nVP1DCEPTO1GAJWTuTUuS2LiEABrFk1FsQbBtbTBfAyHEw3mZSkwB4Nz3rb5x9TnJreWKJEALFCt
boWF+7EvvP56V9GMtT4KiEiFIhGcKS5BFHITQbk9UR7We2ngj6JvJy/Ia5t1kNQrOwOXZ6wIfQ1O
mvAR2489CwMHLcySmrzXTIroOxAOOabG2rOpbLGKnVZOXlAhTAZMRUPmR0XBgiL4k6euXKp1DmtK
gL+VBix/npgvh3hE+37tazGk82NLmFyGpe6uxLkqI6CrStp+qpHyLsBaR3W/0e5aRJYgMQuhuUBd
NEWzPWPRF9jsJ40/wbUgyPproaBm9ggWrJs9GY2rRHMPnikh4ROTBYVEHBVrbwd+W0YfYAOg87t+
r7TMwFnXHpDWXVevrxQL4yqCN5/rL9oTyslCui/VHOrliZ1ii/3CnUPqyRy/lHzNhcmRhQB/Hp5A
fEa6tuDbopVfh6DwXbV8iMgIc/VvPuv69+2SbSqS9Tqd44OW7SCgdAEbJotEvsvJUBkWWNjp4WWw
VNBM0bc3QxzXn4ObLtQPMoTZYrY2bDRqA4damY5EjP4Hf2hj1xu8aFhIe7+D13QIxPooDgn3AiAe
IuKIyhzoJcREb5P8sUPzPy773D8taCwxD4gSJ+pK1CjLY9vJYSB+9aUSJ3V9Sww9rjnCZYu+1dTo
AlmKnt3aTFxtp5a7sj72fAqoZvaNv2mdTnEzRWGCLRsbWAsJq3UZwB2RW+q7LGWOf9or6OAAGWzF
zST7ggI7nsgU7bvwN3c61RVbK3WGAWImZGBNJreYSFT6MrgysCTdPrZhbqQ+gvL5LJh0RGYdrWsd
zuGPynw0VE1nDGdg4nTzCJht2svths+vwjhTUXdLiWtdbSwlYXYd9nUdmqspmZG9aSIQlzoqmxU+
h9wnoZNJtYFUjy3ZYHsUesn6C9X5Yhlc/ygZmgJ40qc9/mtwtftdOlESkHvph7VwhDO/cJuMWY9l
Wnj2GqcAmaNi5H62NJcZj4P71w6Gzczd6t9PVBE1UO0fs/ZQmUd4+41gQDZjFbJr1gs+OHCbtB6H
7asYsRXraz/Fxxi1nz+tz4/zb+p6XMLAQfHItjpL3xvuOqM1R34SxBQGVgGif03e3KQB8hFBJHrU
1a7wd/F0kIPOstuQdqeMpey7wVCNYG8UX1cGaL/G94CIWnTmo73wDqvjMiJUQx2W/MshdsykUAtB
24mUGMvM2mrZyGaY9WiTEXhWkjxaJaQTTLygvWMTTYSv7dMN0jNEFnsksIy8oeoufl2APy533Kg8
JN9F6z6UfVOAfp5yY4tx0Qanoebv6h4mD9siqI9oNeQiugWcyzV5OAbo0bRKuXO2HO4Ai+eQDG4H
i8L2UD4iaV2T3j7l4IzGN+YFjLxzI6sYjATtZxE4oUUufLFTsk7AccmyPWvS9UbX6sSkZIsJNCmL
hoUUs+PVcvzMJRbr+rccHnPgjA2S4l0Zu74vsGGOLDt0QQrydHfw97mFEGtL1Y3YBUxLL4SZ+fZW
mIRodrzlrTjbU7TR4inW7bsNI4dx2DXnTE0Bq535KPCuqBTU0A962BbD/r/mSgBySjqCeOh0iDWe
DgBJKEA28cePa6MFDDdLUW+rZZvZq69jP7UUOWsD4+ctfm/S7o23W9N+nZE7Uar2vodlJ+ITWhZ9
hfHwN1Oo9qKn0jexvZnakNPQLLco2srlXBkEvvbbUqbdJYw3qF6USH5ACB1jrVNC+KsgzHPfXHyE
VJjDaN/45OyG/WFg0tURU/XETj4zZNSpZXEsvrfgc8IfmH4oGSSmzXLXA9BZF17LhmDLqGSYy/lG
HpD2tDIwFS5fKtcc2rA4pyfZKylH7nymp69Vlg7fus4r/o/pi8tzE81v7gtnfxwhPw/rCoura1IM
CZ3JSGVz5aRsJDWi+bXYummLGhAxsakYHX70OA+hv0XwA7nu1JkKouRJOgrm0HQ2OKrTHM3+peaq
0yhfXOma4g9K30Jvzvr2YliFxlcxTJQV9UBp8QIsupZ0cc1LX4AWNxCJntt13RThsG2z2UkxcmNo
8gqjqOIN8CYAuFISL19b3id9/SFfG+SeDP6NVYn9XxAdztl/Hzf8yc+cgKLWjyk0rh7D1sR73bXu
sdvJdjvvb4nXcG/4wfILDgM7jgGdAl0opmi8I28t9D4mFOIJALHBRblqLjazPuL6gBcMELFPdM8x
7rSTp+hjxg4V1rA6pgHUVSS6Nv8qDZ3Zz+RLZjETzpMuw9+RX8pmwV5tfWqhBtrdkoLI2jqzdad7
4hMLnnfPxPbuqU/IZBg0xVtdVKxgk8XtGSux7OXfEvCF5u7bT1VndL02xzP9qvqlW6/CkOOrrutd
p69fhGAeH0Vjwtskae0DOFFKDiCjub+y7XXi0FhA/H+5An1W7zJlrZfZNuOaNh6DpNGWBoz6nLPK
Epv86nuQsfoFC3A0pxJcFZo2iQRYhtEoyvkmtWz3AOXW2mkrwwjHeYVbHc2TRBHEtqNb8fzTDeH/
Wbmu5b1YgOGztYN8TQczFCSxPUT+c1xSvKjxoleiSLkC7TTGHj/Mi93yMOuvDpe+VbotBf1rjhlk
cE+aaR5Gs7dA4WLYwgHxfV6gsBM7cTnX84LkxKrVa3vUY6aodPmh8xD2/SFJwO8/393KgZB919Aw
QSmhHdZAGF83J4nnSwUjqx/l2P/3yIKSrKVFg261TI/finC6zlfgnKNiFd1scjNflCTRjJr0dgMR
4uQMCpluUdomR2jwR9T30jy1AWmK2PCjEsRZx7fL5L+f485TZRdIiB/arlK2vmgV7VkkXyHnOlFq
dSvOfyjwku2lwns5Q/bacDWUEmIxRC1x8EI0+MwsjVbNKY89OjuqI2wHUDLO8DStNJUcTOW7ocCT
NU22roWG/va+RwcQqRgn6QsHKr5YNkula3KnG4Lb6Nihq9bq1864qRKifx12BFBLL5gi7br8yV+u
M6adD1Q8Zq+1b2omRqoLhgJDEOJ55NWvoLHJTOz6WkuqR4VLCYxGkoLdvwJx8TiiRDq2CAc++Tol
83a8BAPaXxgTa8WiH4d1C2NXboKMCAO99Wh8MiTrJnh/DrryN9k17Ha3lm7+8pXpG2RC2AJsmuaJ
f8E0FSupFz+FbEiKNEM8T9QnAHLjZkz03uliOPbqM/OInrJOWKk1kSPwbQrR06rNdHWOga7FiT9M
AA4hH6NxJ6JdHR1RqWInhJ2TIYVc9dD9/57VNWytZCHKCBSupCaG0LTS1sWqO/S1Abbec3L8JQ7+
nLMGh9gKhb5Pi6ptyz2H/Sd69vOP5hkGhrHhQS9kxLzPKyRdXpQ+8oGtukC8NU7J6cnsRvxZAy6s
pnYlUeLJdpC6Y9WsZgBaxdyotx8XUSouhlik3zj1h23QX7V/QKQFAzxIt4y3tgy7RsxjGV2KHKVJ
TzeZE7oeuz4D7mB1nljhJ+beWiyQi53LtE4mS9t9P9Uy7yZan496YMYpjNdgeVu353TzdGP7oroM
g/b11GPngVa06lvEZjyFvX7wlSY21hTsKJqNLtPYiT4hCLDjl61RdXGnRZApfpFAXe7dXtfaeBpM
ch7VexUO1u05PlFRUX/RThXLQCi0UAnv8mZFxjPrO8BFtUa0djp3aArV9wY+tm1O3aCfQhknnDpx
F9FYHSDYLBCbdJ6vA2Q3FnMPgOQJ7kWOuJfpjbxpxDPBe4YaKT/oDMMAhbQXISTmpy2VZwNw5HvI
zU04EshPyysHJTORHl1OJfsTmeiUhH3OISeV6fML2u5NX1aBUkuOrg8zJ9tmtGAfbs9Px8KFYBWT
B/m69IYWden3mgNiUuDrVRcb/+4y7iP81sKtt9uS1t4rbzs/XK8cQLME9aqT4u1oaaLK7Z33wZmp
Y2pdZiqct2Qq1slcEbMmlo2UxafDnmi96yV2R5Y9iPZqBT4S0EDDzUGDNMG+0/tvSKOV/iS45g9E
Z6UjZJQUa7DggS6h5sZE1TKr0cnsKSNVxwp2Qt4scFI3wSNxzA0g+FCqvpPO26DcBMQ7QkucYF22
FqAhjsL2WQXSHsmMQ2/OHd5d32M2IEa62LZBpdNayVkoCEiDWtYcCBufdfCElcp0hR50iKA1mp58
/wrbF046GNn2iLzYGmZ6/Tqd4Ziv3wPukRq0+IlQA81c4i0AQk5DwV6Z8gIrKBlLifzC+iz26lMv
TCLUI3nmM+mNtSW+hgGPxH83eAw2P89uFHcwXQnkmsqxIWF/YjFrGjUETnhZhbqMrmo+/DSq6f28
67K3M9s7pdD2g7kuf8DpUMo7R+RaEK9uV35i/kt5o6cKdKhpUd6LVIa3S86EhoVlJyVJalrc+bKd
z5uFd7I3fLc57fZ1gpxPUz1zZjGDlnEmEVZFqJ951hLwYYK22fo6NIakA9NDirHOI1rIOwnjTQhg
ogeqE94hh7oWewik1fxH3wGd8eBYXNE/i2OunWkg30CSqmvxn0TrrWYV4JfcpCj8OKP12VAfCX9n
EBt8LR3ihhLLKj0rr/EMYGMk1vdBjHwBDIYuT3o+fBPJIIwF8RPHlj0z32acoLZfkNWH0Qsv1QTC
Tfioohmf4DiEb4GiYlenArhIZ8Pw+wbXLL3Ozk8eiKMPBfKRkL8DgA+GJlnTJBa8lI25pk+uSFNe
q1Ehl87EWGDn8k8EdDpwH5SsnLGOpp/lBA1UmdGOnNVmTyUChtojZzdG/DzbPSuIYKAs/YUheGOg
gRAzKTBJmAGnqn4OwSMWKx2irMoC5xGlkGWacmWastNdbGbzOMTdbiPFxN97+VOZ7tQdbv0hOZ5y
Re0i/X/RB/28MjPPFEqe45wpqDNL9hgrXO+MdsILQqYCnBMWZiOqaPn0rsal/FJ0GLthCL2qGftF
6rmcU9gh6VQbRSI+rLWEDtr6Be+UD1ZUgsPB/n8HxrkOnUw+USBVPyT+wagQlrJHZBVmCIfV5WTb
bddJo5eaunw0x0q2seRFnFQkuQ2Un+5yIc/vBkeJ1SB0TQ3QvDUTLe66ZnRpjaVWPsqXHy1URRSH
/L5vwDQTl2i2w6cPNmw4sSSVuT437mn1OvSWijZq3MF0e4uwV3YtOy3mgtFoOCotRWuB9T76Cqy9
VvMdpv9XRtf64qdAYW+r8rrwJu18Gzc0K9JM3so0dJSXURv5VJP5fJapDkD77zVQaj76bKgHqRZO
gO596EIN8dKPqcQreuw22qU7/CCPnECgwj196fTu3LWIRhUUUpZ4QjN8Z+v7RRfejPP4F8eorf84
jbFuF1L28NjvFnXHmNSjQ8fLCvbRjQNkeXy29devMSoxARpLXrG5YqjFVYavwy4AtXz586izxkEs
JR1UuRmWOQnX/14KKwv0Qt//SGk2PJ6Z2a1JzC4WJPfHu3deJQDPYB09XUbjfJs2aJ0GJ6D4p2GR
cv3A/Cdm5vQD4SDoQzKsygTfgsSbcWAXlwg3m1XIp+Bq46GjxkTzmrKq6vjgEYK2sNONZpXPaqmS
1zaapxoceytvNm4/CKoGX45oh952flbsGpr0SP87H6NAofEzJHdkdlmom7q5Pkp1zAKg8MRzACmt
v9pZa8hObHUItuLqwYfowve9Lx+e+Df5g1LAGeRLju9hnT0A2uXyYBKyH7hKGck/1sYRdd9Gg3aP
+xHLxCscsvd3BJGyW6Tm4eAIVSn2hdbJSprLfulTwqzbsZvIr8QMzbvVTKHZ1SWOS2DdN8hHwFNe
JZovlSIRNRMRWoJrE3BF3tUBUzf7+NXWFAqAdAr3SjwIZiNRdWlUsSGswWfV2sNayqo0E+U1/wJP
tOQBlucUJan7w0FUHQuWi6MWT1eWtriqDoD1Xh12FPrSaygAG1r38UDmqnT3YSY0VGg9YlIe/F4k
x5YNZesY8jJnZr7YdXBXfo/EbvBA5J+f34T6JEJAosFOBNDlEjHXSlwt1sQ7KJ/ftyx7nZrd44Xh
3K3G8jzuxqwzkkc9kcE+2rQyTFTjsYzYr/KVGfjbXT05F22dy+S44zlTQEXuxnlvE9wq7KUHNLHs
alkB1LG+wX9eJJ+ypUGVmyeiK771G9SE+DMteD8nBQmNBaVbn9HLdwE2ZPrmJ/1KPhZauOniqsZZ
DVzNOziBonxHko1sEquQ30DNftF+CM7TfYAAObRA8l7MYoRo+KohTASPHllGJ24OpSBpVKun8iWh
HQ+3Eik4kIgoP9154WcxSK1tgnQE7aqaVAgo50TtR581pGZLLKi7oTYXxje2Gl9O2xgUGuhJWRZS
MlCw7vzBPy96nvgqVaH99xMw0bj+GLHFUnUKJg/GwHWwkIzyMnH3BVSrc7VoZ8OQQNkEXXzT5zx4
UQqGJRYaCwhv5ZEdcdzIvrGMQ0uHk8zyz3QRPzWE8sRuQZiyDVlFlgpawNbn0r1rQ62B0wArAN5o
x41W3iA/KuUnJMI0u/9n6LFz6qsxLV7MCRjKfmr/qVU75ssWFKmxK9hWAVZlUmF91X44oKk0AtgQ
0p1z/XGxuUWfr2CLQeZNwX03pFT4I3bwlbzY1yp5xrgYcZ3Q5IDR4S+ggGZi84VKjbTE3JVRkONc
jbF8db2rE/FFlFl3Prfq/uxfuOS2BwpuVehnzyQ91UzoSJynMfWNG7o8VRL3D7BNAsfMCjJgxX4p
Upz/GRxLgJUkhN7X/9LoazHz9DnRXpc4pWjUvX0aENtPOyeN/YmhfXcKfRsMcev+lKva/KtrH9wR
Ka8SaHAIxPXN/Cok6IA2miTXu5RKDwUuq1su7dHtK6mIvs2vNxIQl2H7UhXKNujoscGvdx//Ml7x
iegt8o+QQQKb+DWBezZZI3g/4Sqxiv7H9cMXo2rropT2tRpzBA3g4tGsn7wDuxZHD5ZmIXH8f3b8
MexyjafBmVOdaLLkM8tETf/xWCD02GHk5YuwT273ZOmTIEOaAQJJySEiBTF3mtH3DMWWWV5qcJCb
8l97J5pN2GXE58dIvEZKskpTTsfOsWFlolmBriqsEHBOM3fHlk0xysoTy6QQxT3ZckSbBXpVdggf
C2gk+tmpT/xzCak9jdxMWQtrf3hVDtGglqdgP9r68vG5hEgxU+9V09WhC3LT6nI0PU57u7OWXKKc
GZFZzdmB7Hd3aLtEKe4P/4F5Tz/DRipcHRdLEqO0EiyHystkE4qhSk4dDLQUC2trP2cDL+Sp1aS8
LT52ntCZk7qml/NUNU59xw860lK3i/H1eXo+sOb/fzmRaKMZ/H8nzhhKU4Bs28nr3pi2nLaF5uY7
AM9ibPolMRQ4Wc6n9ItNtPGW2NUVa5s9KLoZhHNOS30NWZo8A21H61UOsZSmEYgFd4BzTh/IB29X
ou3NjrvbSVQMGpVOYZy18zxXqlKfORZTcEejAQzgcY9pH5Mih1sLu9ydXVMHaEs7rqX37d4cxzLf
23iOX1UG1JTLJTWrtL/LX8katBmoCl9OjaUChzmztl8innIcW4hdS5hKmDWY4og+PRnEbpLSAUtv
Z/3t0XuMAUMqun5xiKs05lLogPjDzCPHYCH5OeCybz8jblUE/0ji58QdpScVmZWAnri1c4cxga9U
Q32TiquE2q6Mxon1VIBaldAwDdClN+PS2QkfdYMMfOZJavcCCnmQB+jJijimc6Q3YchEd1lRFZcE
rHXNqgI7JneXyCD3tTA30i9pF/VBUrlUCeocZ276kxPt/XiN+GJK0Bv3oTg14StxL15lxwLMMSc7
TerbtHvI7wxtOa287aip80TZNcgEVFPk2n/fbT5BQCQ84CeVsKD2vMvOTSqd/BTSDW0fc+5R5JUa
Tgqs4bTKe/gQ7p4QWrX1j1ouGDFiYk2Tzd4LZBAI3ZR1VDD93Ti1+hmQPaeEVVk+ITdM5v84SqsF
Ff2EW/hc/feEedQn5xsuVPV5gopQYpxZP4vgNTCdgBOUTeT0t/TnQ9uv9ZWqdY2bwbHgwFQnAayx
Fb6Whd8AvDd0XHflvFSb1lHyOsc5BWZheGDaJ4WtzinPXy6hryc0zp3XtO2oQfIGOrwFaJ+tlLE9
gitjEf817WzC5e5Swt57FnLz2OaUWmpL/qvhmIb1UhqEGGOQEX0cEHhnMEu8k/7SERm6bQpuWGAC
jHXmSkg5jtkGxgG1P13vzxmcEA6uevOpaGmfTo5xAwe3o0qAePhPS1EM/iX9VNH5QgVTRaEop0QE
7oLrw/IvX63w6sgBaRa9fx5aqtTp6e3Mkwqo6fs7RvO4X3mnYmtrDQev/W5V3TA7AYkbdI9LERwT
PfwKYXjGxxwSZU+WUI4OFeqEITQn6aZbob4bD4R4DAUfs876tkWpnftMoSUyClKtYhrAaQQQiq18
4QLWlyyqA1o5dFOQC1izBesKySPBI8+pWszrBVRJsC9EZI7NaHc9HP5f0wTs0xRgJhXIsbRVhgdo
m8Z3wYMjuBN+xz4uOWf8VKP9HXi9nSPCjfZyEVoE5vdPsyrlGMjzerNBP5RcsDgZx6+EUmczggAt
NuszO28TkgJCdMU3BmhilB+1saFuxb7BwV2ZJVTJCbWWMl5B4IQGBl6GwWkh4EQAK8P6vKY15LGn
ap5GcXe7c4fVPIFySSxMgc7KFybYgGqBv1PNXLJPAGfGXCSBuudU/N+YvwnPZRfHvyleBwXzmryL
3ebiwPcR0bRwRlbYWYpDgO3YLIByuSW1vHeiU+YhkaDV/7XNHhN2PqQNWyzKM0m2mkhoGHNWEXZA
pfwFyfJ+SCgSVZ4it0QWJrcHkvd87lSrnNmULn0U1TTgBu1+QnqjTUinWnJfCPNHl5z1ucwCwTye
qP93Ik4KZj/2FvRzWy6H1zRUnEZ0B/qrQ7SvThnyV0m+fm/9/PkQlVMagXxuTCUdWeYdSnDnR0H8
E2sLL6u0inVXpKJlswnwTDZGGlFKkh+tMhwkDqKhej6tfxkk3m/eE1B5SRABSZWQvXq5jgI1bkJ9
n1cTMF98k0LUaAC5i53Ad/1LZN7pQMuYrWO5Zj4h813wi/wesxgut3gYkgrF0JZPYTNPoX0HN7Y/
Mo2EQjlAoS+TEug53ZwxmqlVDgooBnYg4O2jBTa80oYu8utGiY3U7LnYXwfB5aJqTpqB3qv27w49
oc/LQoNNffrvC2t6jLkJoHnKimQTVGqMnQFg98ghBJf52PMS5mUY9ScpOeKIuCinrWuyexWRPytI
LbVYDpcMhRuoTsHcu2MCNcYNFvP7thweJJXhmtikydEw+HTREfjTwz58WfN93pov3gBELPFY/gE+
VZ9OG0S6HCZnHC+4VIx3zacknLyj4NWzkMM08p31pxhSyjUlMSVWPLVYS9RmZBv6nxmoUttioC7z
XksUjkJ3V3IJ0yH/lIRowgaFfKlhBUYau4EgT8nwA+VU0Ph6Otn7bR0xW5Stjx92pKrFNsxAZSdS
EzeOAMuSyC/8AH1o5B+mV1/PNTeROCyBQn7PIhT/BioeWkkyZQvsnM44k78cw2zbUJ+AW0jCkVrb
I/qoA8rhjuvSzwVaaLLe8jhjNbECKXBKyh1z/mZ83bSEs2m3hq/r73YWMPfv0DYxvfc57YsqLPVi
sybZp/eyU++Apiil1gTTpeE6G9JGMeowkXcHWMUw7EtehkogNADL6aN9Vtbcxbi1sMFBhmxz1d6/
A6dgQ63MtNpOmIufjQj8oIrxEwGzpyf4KjJf0wW9DoKrV9UzR8Ref/xHdLagpQPGOQqdfi1B5w8k
BKxuqSr1LEC/9aLLmyjRTYFhgX/7EjEyNpc6G3uP7+sNK2DkCMfYJiOl0nz03iLDoURcDdBg7fYV
HqF5yDveNXnz2Ae2MpPZGOLcw/i78MJHjsT0KGiRyRFdE3Tn1mZ54F4GdXTqvWJgOUDeshuNvRIE
cYvIZ9M9hfN/EgET5d/QQ05g8MXK7LxcED2K219ZTW0WZzyVxyxHHNTRYIzaOgbubEbbbFfwKCOM
9+2e5gg/9vNiObEwW+4cPIyxUvh0dnDYryt09D8xdmU08YC2cZka9iaBwcT2BO9FhwYxalXwr1v2
HFW661B784jKz20OOvRURitCu57tMU8QqKdDFA5FMTwzLvRM6GEGIBpAstZ0uriVv2zsh+u+5JrX
jsl6GwYWm2Yr4evB2cEpOXNQe4WNiZGztwFVRxY+NAKZ2p3cKDjwBJHEYgtPKImEnnSZQ+ggp+4j
3qQxF+8e+E+mKEvPuMXTZ/H6s+/nqHjTV7j9m8ilv1q1dELy88DOmEdJ/oKXF6x7sC2RuKVdUbdw
qHY768rwY4PT7ycntqrDIuZ1zOjReDgsHvmKSnqSAFgih1FU+R9jKcisjBj5Zx3N8VQ9ujfp4Snw
gIxSHnBZ5hy+AvS6qP3bQqYBRn+g43iXkhHjddtT1gMVd01QVA3u1BnYi0KsztP9e6vs9Ho4rJPl
4XlqqnUsBPS0EO/SSvGxU6IMXaYELCbjZlivdFteBnrWz7QWhp1SONYt73hzIeZYRjesowv6N+C8
16DcG5h0FO5kF2iVbJkNu/GkCb0MQoEkpcVZtr9x4Vd/2MLFIzY/yAOS/s5QLNft/aMvkFVLYQhW
/hw6g3dLwSgHpf3v0viEi4JEMjxDxARjp399RvvTfljbMYrL9+P1TZgPMBhiWDZyiwg3UC1niEbl
VoLnwLsACX9HGFqRujYgP0qDa+SeRU5Rymxmi5E12KskwykQfVFzK7rOTTK8YpxrhPuJLf0F43M3
n/oYLt+R8eIfcT23hLnwnAf86Vbx2/gwZifgQBsmBQBt4v81E/bYB/RYgy0iVRbw8CPvTw7rjeu8
hLPPDOPfCpC2CWhCVnAVMJgG4IU14zMC43VjbGowmG3jgM7fFXAf1i38xIyoq8OXT+nJD7bF6lRm
gcg+bSXCmlkNZWWWVh5lcWJf21bUvr+ELYBS72qSfI75FtPVa7ppwLfTz1qszA8M0YuGEziblXAa
mHtIGI0JSwfmpZPzilXeNjNL1bUNTU/Y7+2hjajv25JsjkXbiToGOWH6kadK0TI+UDLAazFHmVhv
Kv5T1JwnPUTOK2oOrbDAoT9O6AYt30WXtUuPDnqAlc517s3UiYcDwFpp5z2VXbSRbFbYBXEbVrs+
akwCGTGuTohS2YNIRIB2n+TpC2on11ZrbuFnidXvWbAdVYGn6kuFFGEr1ANy+gi3ATmT685GbuJO
JUOID60Z5GhbyDwxjLCsUs0oTlzorI0NAR6dbkBgJZJBuHuD67bd30Y3WgCQgDjLRJdXtp+jPMN6
TqLAM+bl2ktgSbMCn86JdZKv/aCTOYiFyliuUjaS8+lDZu4uDueaV/awYRKAW4TAnvMXt4GIjtIT
+MBRYsXcG3/Sdb4s6rtJ5ffwuXGKymfTINSXrJ8amc1P0QgrtN6BxkSOmk/33f5jgCEAoJWEYCOE
EUWrLwsJdfeDqnYBZMXWChpIyNmDDOVeY3bWhPIiTAi/KrkTLDme+9xvTtacuhriYNCWreNlVm45
usdNpVIFggMiiPuuco8PUFokYJruoXV06Dhg9MIC7dkcLujTOo+l9hzYTjzwooC3byzodtmcZ3Pg
TYgLsoFNiQNWDp4EoEBOb+sfddbaFle7ejCUQWTitazkJk64ptM6SDKxsws9bGS+XyYcES+7pTYV
Sf1vGi3zfHpIoq1PSxK0H/Gpx5yJBJiM/t7gf5odFxdivQxhiCy2JQOdfkvDUM6TnneuvKm706TF
W/sQtmN9g2ETUV2wkr46gbu0glTyyob0P4teGfgVo4tN5x7Yb0cqFD2AoXPnKPmuzlfdkaIjKGLB
ObMVm2+XLDYKeKHNlYt85Z0Vs/fpaYrcRrsC53Kt60mfhlwjdlA7ImCzeADa0ev8ZqKVwRmVv/0+
q1KzszbJf5CswD6eIzFh8E6AeiFyXRnFN62778HRmnF/to3ytgnFIDNSAMfvsePAmAK+xg8T9tLj
PvSMjIO6ZMNYR/Mts1DjNTilT91P56bImXavYwU0FS5W5IGYiyabeDEBxSN01yv9BaBpqSKbsWoU
Nr3ihzTsQPI7T95n25rWxu+ucXYk5hZ2YEncGED2t6hruA1JnPf8UIvypg0nsKD0LCanBAiWTwO9
w0rp4UkasyZvFNvjLw3+dPRUvL763y5M5+Cu2ut4RH47OpaMm9Lt8cLi85uzv0irCGp8WSCk5Cb4
6ddV8z+q8BLjypvIJRmIuTy3NNpf9sIt2HJ6iBeEJ+djmbTJY/LcuLc5pQxcdimjsuQNlbWtlu/A
m32Qse1HAAnbbzNJFdyJdwCs0Tg4cRfhWnhFPqYHR5bLLCqrqTzt6qEd29acFoBLTWb1ItmYv6Jy
mX1sXzxGZpU4UPhBES25oQBh/6jzm2BaEYR/TwPgZRyeQZZ5FUiaZrrguf/KefmTFPenzOy/njXE
91QKzawF78oVyAJJxQKQ9bWG2E8hkU66CnzM2nTiXWABpXCt13x7ehTFK2jIgXfzZL2uEON9Wuyh
Nva5Um8Xic5j7p4myG7HvjtlHIMYLZJnRo46oIrkBmRSRy7KzOc1EsTvlQlFvZ9KU14QnzE9U29d
9DWh17p8gaYUD7AQPrqFAN8sL+uucEZHU9b5eNAVJjIZ5OAbwz+JeRNdH9VI2aXVDqE+FH0DfJ/v
5aiXKTBGzSJaNjmNCtkLYbNV1wsgdAkWgrZdtTkt4hSjxKzImI4yIjQyOTZk9EkxrYKhzGfwmMRn
+IdWS8sdRT2MAhEHAb+saAYEQnpxmLceIExG1XI93W0eQ3Fl7W2BOBcM/yG3RBUEa9DORGTDUgxK
JyA2Fbz18HZ2gCv4Hhn9IMn3ZW2fzACUC3ARuihWFGEAkLkQq8PSczGJgkdWYB4+mKgiENtC3x63
E7SaHqU0HOg5KAONq6uhH2QLmwjJKTlTr+hU83fM73M9tHGipAFipeVdlOc4zSD9KmOTaz4oqzV9
pZ/vyJVX2c3ewe/fEHIMQkwzAN5zbL9DXz4glLmqO4XwVaEfZGo2OK14MCF+y3vzXE4NPYRyeJbV
h/LDXEsa2qB85indAgHBJTWkDL/hMq21+pBNbdNmUS0QyWRNP4//jFPM+t+jcDfBguqms4MGsZZ+
p11mEVRF9mkAv2LCK8P3wQQAI3zbNHCsJ8t8GlxLpWyPhf+V5QUX5U8fYSDPlgzCi9MQcDMt4nQs
zCiUQWIVszFIleckgk3uSoXubOMprceoQ5ETU+1KdeJNi//SoPcwlQF5GC2qyfxTCgr4XjGwxyxc
STXZG9Z+R/iu9rmVRh8TzDQHZzwYGV+MbHpphUn8ZlBs53rQvgohucc611IP4fHWwSM0nUOEaFpW
GGUT0qkd5MiEljaKNtcOT8ReG6pvJVoSNPypCnRvY59B18dUibo/itL9/FJCgQB7OuUz4maT/uG9
l+KIpkZysymFQv6X7clnjyVGMjJbG263h4IOvvjiEXAiGty0p4pl8Y9T7KdCnOTsITlqImdBYiOk
SNQNjgYt6ZLDttZVxRnPzTNe/jnLwVekFZExF6mXuI0l27OCaLEdLOY1FnYPsA1crECjbxu2VNuV
KU7KU9az8ETtcaXUaPKy9ZuFGHx+WB12/Pgrr8ALUXrELoJu1tIwAMoZ1j47yRcKoyKrbLHODK3t
3eW+mv50PoDH9JLc629Axwaz0G8vllKAwIMk6NtNbWJf8DrtAKNlO3lmv4HtZiZ9z3YJ7mXpcF34
iLAi7pmVEQT049tTnreoEKOvIueDsN39MQRtdc6tV9q/Hpv6r8ggVuJWW60ffQlpG0bHorNEU4Bg
CHzzWamifhLBJg8IpXU6wm0CkQj1ueLDA+g4HxX5XQwupAna4CowMrNH4CdAQCayDjEeDYrJu+Qn
3/7m/XlmGeIOp+oomohdnEOiJUaF3aXMFIE7e6Ex6+MagW6+QUbrqT1hgC6OLDrTiGhQHhemWDGK
Z/Ayg95iApTGT3KmDTtVlR/BdpV7SfCEpcpvy9KtniXTlV0Ih4N+pL5H5EEFoPbHp3H6CbPRegB6
QvA0tQ3OKnBkBYHBVpNg0R+8id+67e19q4H7JZ2oYO71f4D1WWMRfjBS2rsL8uk6FHyE8UyhX4jS
8C44sZNHesJQUbtZB409VQ/PXrFqs6uhMSqjl5DW8dYZVjgoNtjsZoRXratML5KB8l2VmUh+Z3TD
nd4INJx7/kjyCphtQhxuBvJkpakR0+y4Xx5Li71Afmx4DflQIua6PO+GvOg0utPiBpONm1gTc9XP
HN2xkQlOgaKmcYxbXDRzIp22pjmCiJ1q5zMasjBNRjGa5sPFRyyrU+tv8xnkHkJ6QSgNI5AdSm/i
PwxGn0CKLwKX+jMgXIbujFGlCaIp9hqxhAD96iY/QbR4K8X2k9AUjCBD1GC1PKlfR8zf7/T6lnDc
/vzOm8Qx4plXBA/fEjds1WTZdCdJx2Xq96uKZo3m+3yuJFrl5QZqQOSClVqNp8Th0uWYO+WCkk6i
Tbny/UQl4MoT9KHknvz6e3vc8YxsGLGZe6ucTfgXO+lU28iRqxLKltUWvtyN1p21atoidYlmdG2Z
QG1uAeCcDalGSbWObIZ1C/OC9SD1RHhPV172gFKm0mmIkfQl3ttgZUJTGiRC4uop76RXydBeYHOX
QsvIh0jsQCDrc1PFO2QsaEJGDs4cfYDWvjlML1R1r9pSXqPG8u+PsGXgS1Lrl9N2TkJ1kYo7WgAQ
l0jve58hmZiGATRjZdaTgU/iadf+nKZNw3ADQd6CSzNjJqw0pfXhc1RlnynLYTp0V5cg8DYgevmA
aksY/6sVoSTZn/IOuVGlFVENVTg0CDn1RdwrXczSsH6OzGlirQAUj+SYqW4Ln/ZmoFiS78yfEw1f
2erkqYinXuYBTg1qu4JdXjrToED7dVhg03nCVli5bGmzkpoKuu55zvs1anpg81uZPeMrmRzZXWqv
itbJVjeWnX++gcTE0E8LQNykMgSxyK52A2HuFhoImEtwL+Hm7jDvpvgoKxs2fobts50xcmcga9D3
z5v8QwMYmKAiG4dGz3bj6V1hNEwiNX/9e8vjyR5MLZgDXyo2eU85m0kC5D1WDzLu3ckxF5d6XUX5
VFpRgRB7lMzslC345YCRbZahDI4LiPf3eQeYxdY+mxM46xtvS0BtrGj8cJT1eBSVE0zaalzW7cd3
J3ctxgNx8yUAK5FQdmGIZv/PIkxvPBgN6v10YsdqXkuq34iS09kRpYkgd78h9w/EGs6qwl7+Ewbl
SoAVBLdE2mcP13mUEyYuyiuxbgfLB9jSBLYD+ys6S865ynVwTyw2MCsd0vRBGz7znuPG3PbAyHRr
0RsxEjj+LklmipAHqtR0cd0xKlImzvhHdPtWQsu22bEH3gt1ISOBZkP3tO/xgNbfsGQzon3cu1cO
EDgUVHe5VtCuCc1FBlzDhs41d07bYrq3VoProHFJLjgw0WYCQBYGAGcp3G7fN00TrL6u+6n20LxX
nvsmxJp2HnmXxD45iT4ZprD9IEIEXjlNi9I2heoDYJe7hMMyM/AB/yqmZJ38jcyz8P6QxiEzauF3
zGYbLNwtV0KECGb7r+sa9uPWp627TGkyAjgMYRkTjJBZph9AZjyQQ+HQ/zqeZZNZV9QSvY7j9FZ+
Q1+1YTjLrUVXX/Ii4O1X7hLqRTxy1mEFvA40eS7k5Gyuz1zd6YTUbxlvmLLaz+EZ4rgVJ4C15BIU
+tRucUWHkmDBRJu0m3MczSPEoj8i8+LvTZtBIbIAnXHs6O/nJK6v2F1pChNG387cneqF52eBPrOl
JKzfly2Hqy0tgc3wji72dxCiFWnuRkGWOrpswVP2BtBWu22DSbIwPnXX2DKBdoF09XbCBl18S2yE
YfAyFibNh1BSnW+ga8xHKVSkx5u2r3HetmW+yCt5afIaCVpUGIvtEEjFBD8D+T57mfhZWAMJLCDT
t+4aPDQEyvje+Fk2NSt1aM1OW3MYy34XQyafsE3HLHAjamPtChPtTpZwke9UzvFHLp4SejghOLY1
Q9PHyiqZiQ8uyoOd75AX3VUKbfqXOmTainWo+LsaohQaYt2HJQjgOwTARGCYM+K6Dz+iyEEQIeYI
4n1PAmoByyi3pSXP8+1Je8xpnub9McYt0bCoIdokwSusFksoTvH0rYdM5TUSo0p8pPlmtkDIYAGa
M2H62WOyQTkWBSAf3suw+WrLhl+QDCKX9deLetZVXUimVZX2buvrh6P+oKcpCB/2tXOZPhRJEKFz
+qDkHd49KF2YE6PzMQ72zXDCewtnDWetQqMOXm58A8fk6/nR888lelPY4bYyaoL6Byd8Hh5Cltvr
loTi9kS+yHm+j3DS4NrYLRoSNKHNonO22J9oUBEH6U5SXnDlMeCJsza6hKsmKVVu6zYlKBMO/+7w
1SkmnXrTXCQG+EuKGL4F3sXe6ftQu6IDA1N8ZLTbJ7yTRFpqdc9R63tfGUQd8FBmpg58hxKNkq4X
KUcxtgdKp1lRc2ClufKWymjL0t1iT5+lD/5g6S3DlvmKAgiuVgNifxNYPyAKJz4MMp/0AUTI/nNB
0bLYHIRP/4MCTtM6FMK5M0kvzC1T8xGQOsCibvoU1lQ3hcPWjOZmiKvmNK++O01nESb7nkfwpkOB
2Em/GuSa4E/rMG2MX+6oRxNrpatpOcGwVc1KGwUsCkC4Ekjj0WCRpTJ/jWH6ssTcTY1T6hkZFUKt
V+amOyKLtTEhBwij92HvMLv1hoGs0EzLx9ferWxYjx/3NjeD4HkChu2DGguKyFywIOEtNBZz52TE
H09YwkmHX6T15Vzy3jBorOhcEc74SNwkLyGdLN8zRlXc/5l1V6qBDWmprubsEC3oIhtCyIaL7Iw6
MNGYsySCn4wvyjcZP26x0kVLjnywFRPy4QKsNW2jbXATJ2TMJxE933iCYUm0aUh6DYF/aK4eB9XL
Q9ZBqRLmEW2zXdAuA3pfIGISoNTU28NGZ8gFy0XmkIlLZxLBVmtPVRmtzG3UovoS2/qXjZ+2fWva
Y4/AdlP3o4D2gwH0847heC5dGLJWra7al6sbvj7sVegcqI49cPOIMvMpUgda96pBPiJN4wLwzw4R
e8c0vVxPMho2XF3J2+7sxOmkCT3hyQ818P1KCx6P8fD+offWOyapP0Q78llZ3NnsseDDR1MPnJxm
HHMcM+CeKNlZmqJM3BS9H1Gg6ByTj1W1fno7ceog2DtEF1eZAvTFBVJQWE8a5ZTHiwfFyy89Se1w
dFVRoDcBg2xNE/+tVpHjxcJRCqA1YVwaZu0Aa8Gdyp3mXivCmhsJc2jWfIaGw8/GXScYSVIyhMgM
VWLSCC5Qvwi/sBDes2RdHmpwGtxe3gy8e2rCDMSF7tCj4L9PPjcznEwYYH1fnz8it+Wu7EBfowK3
Sp9T/DZwjeCJcBLP83ugsBn9LIs9frR79exlNOAcOoWCV0uYLbVGv9/r7GaH3uifcJqLdNLYFezW
+spfAZKwV99N6ppfNBu4kSEMd/OKW4X/ZGjQPfu9MIP3kNXahUiE4etMqQjuB1fCFHmFzT4Jmt2t
8Ep7o80mCd7MAqQ1DRwLNDo99tWtZuDta+DqQUGAyxzw7TrQYZXjo/CjCIWjqfj2v7u95yYto8D+
BLGkX4oWP/hDGtvqJ0WxsEjpwACQ5ayIhbzon33WdhkuB0ViCOG1ibSRsKemPCjABB6BxspJ4YfE
Kiyw+av+HPH2Ssr1r9uniCYbYjXIyDLdq6XOTFMhgkNoVXtqtUtvXtxSWxGKlj48Pan/+wyDfpZ6
kYL0GI7D2BzVJ6n0rK/EeaBL5gm4A564LzlBMHBTiq2Pn1C0dKknSxpA1bxdluaQzzag5CC5YNBu
kbuOnNiJTAb8PkzLk748z11Bya2TRKgZXMmBuFehcUiPsui1GVLw94bohkaUZZej+z94LYYh6Wpb
6bsXLagFhVBkDprl0Yks5oGAQUwyLCVCBMQ7qflOVFeVsqdpMMqYx+tL/DCSOpZOJsgQm2mp1EJt
BzhJZRauywq4WziblxQYolYFSBJXqo8hyblUz3TS8O5qvzvjA++1yIjmDceUDfDWEb6BjAZMezsh
ah8R0gDCrtKxCBTgaPZzugHHz/6yzZgqGt76d3E97yA/jcf8tOAYuTvCjESYOHbK/PHqQRpeyc6C
2f6u+F/VM7LGsw+wW1Ko7Ku1QJ10az8Xr91QjyNVeOC5RnVQbO9wbYp43LA3TE00r3xkFCOIz31d
Zvc6ofXkGaMmdpmq3FMRNHVFlUzTSgoFYCz0FHXdLJXcjVySuPrp9wkxA0emJRsaUCED9tise0J0
NmGsGwRjStfCqkj3q1okLzxNZHWJbfsVGeY4PqVHHWYJl5xf4j3n/LNMY8a0b1NRnW0aVBWByUvx
cJKyO60iwY8abr4zmkXX+Jnd+BDv2Wcgqwk1xPMqrZZuvNkEwP8Uv+6nPNZhyci7l40phrouaraO
xFPQ3XbrRQxOTHa9WgxUc31sdvWGnT0pgA+RL0dLghowrutA4/0188TAog4lX0+AlXbxKvZayzHq
mx5GjK5JqMlR5vSwV89ATtJ3dHmYqNNRY14UptwiLur/PWNhr6DMSk1BDwfIbeM7e3Uki6xJnYut
bJk5DwoRv85M1HrFt/d3aVcxL4p9HiMwe09J26R4OHRheyoVtETI5RYSrxh9DwLlZWdsL+xhwdbs
PzyYjOCvjgcuFnoMyqg/MEsJ4cton6z9EH4WLGxdgAJq2k+5PIkwHEMVNj+nzDW73VQ3bhE1VSLZ
8vUsPuhnd1c/vKiXcGWCQ7SMr38ldJQCdvoPwvQQntKVKm7T7yK9OSqxty4UWO0XHz/OBoj+lweC
eDKUiIECx/4dFBL6+AccZJM2eJ3JqoZUAXz7EuhOd61o+qGirvu+dr+XRbSRNInJ1OSNzcODmgqV
FAF3f7HlCfE7xQHzzPrjSfYK61wzN+gqUfVWzmVCCoFFn2TGodJzG3iaKvFPB+DWlCUhSidfDiH/
YCzYmrBfh7W8xI2g9RaPvEFfuAEsGUQ3WTZ605J8aNYkifkMamID1EuBqgqCeZL+4Yy3Heroi9F7
ZEjmYZE0liJHVvQCzElNLduR6ygtNz3iodLP724WK1aCYmAXCWegq9YmHU6pWEo8cBcYJx/M3M1/
Yupa6opVgZ6ZwKb8pQYYM64kKUvEmEl5TnYo0nusRf/vML0gtTAlR+GOgoaCThm2Aj6vEMhevGso
0UybfM9QVRpK5nk0BklSneFCWG7YWyoNP+lXqjZfPjKVSycdbwau/MDNMQrvyoTIbzi1k2O3xEfq
2nz4SP1dNZyQiM8pMm9804LF8vsfzH4MMZRgnuASp5Zm1yY114BMgD3yZlNYKV/1r0Z3Ez13btaJ
bnQfpzKRje3o8SCNnM9aSf87ZOdwC0PkBDvNKcBMWc7MOZ1FtymwMRFrKecOyW3rcWV0/Ih7zk8u
6J+GMHNFdlt5exC0fb2qtD4NSrTwcbCcW8gg8t5txKmnwGZ0Pkz12ihE2+fKu3tjR99g408ZjM3q
K4J9NrTz0+Zne4LRgLtUPHq+2/YWZmlPwhv7ZNjdpv8lcK9SKn2SEevEr8G4b/59xy6J9BzP8b2s
zg1pQrxxPqnVRPleHVVfTV/5ScyKRRGE7sl66Q6C/cHJ5JQC+pZuOkmlICOo2pE3N3nhbYb82lqE
Jf+vBvESEy7AVu6S92HkO/ETmuxAVrkwl8r9SOmZ3a+/+8urvt1m1DCEOzZBZwyKoOvGGTJtLKh2
A/aDERxvoFbBZDHwJKI6QA/KLpyzhEwTyyt0RmsRna6tx+eW0QGW3mmnbWi6r8awQff9zPD1Fe5k
3s8EfhdIq2IiO9Y/dIKoTVwfytuMGr2CD8T5FfETL6MuU8q9xoXS1XcwgzLsozDNlvgjq2MtVezl
SQ/QjDT2pLy3fCbBol+629xZKbJ5zyPQY22EU1q9oJQCX6R3AJ/0g5EUTPI7c44GLc2w1FKTWqt9
uDdG5O1P8hYh3KPVX//BxZq4Wmfui8tcjQuQlftuAHpigcMToQcUpm5iVzmDW2FF+/H1X/DHmKAL
6FxXwcYI3skkz/BLdTK1sptLm0H+2NZIh6gifEJulhnQvQrr6jixEzBJEuMsK9LkWA7S3plez1Xc
GlozfRyfKXxguY/9cFWnRjYE1dMlQs8SQa5YZ9yw/QpLeZgHd9AsQYlyBijmoMG1c7W9ccdxkJ80
81gHlmMqZKQMq0qrciV8zTCKzuGt7XnkjJToHalzXiCEy8VaW6lacPOpAFk/FQCzNB3PE4Ungqz4
65g5rrse2hK2js618wHlI11FpXD4IzJhyay1Y8p81r1fzBCnGlrdR2fmsZFrXOaj7YGXEQK0hj74
FjqgNQekLooCDykEf4X5WPRCxKWf2SdINokGl9bjMII7jRY5KScxo89UqluqeE8UUHsktq0KovVd
cnszSRCT5H3VNlTcTCZxyvpt4RF6Le/6sSTDvFc/zXxSWU3jeRGvtvorytSGK9KmWXSccpgXEbkb
8Q3qTmlUDhZLMBhf7bR/MNzOUOVUEBT51WKfGkg4IkFSelKsOh2AODPPG6kvqK3WjthbUd4vV307
nfXxpCVDFsOpQ/QHOqMcDfnfHr//uA+v5Tp1IgtJP/Cz9bYzykRp5YGJJ3ksFECgZtIDqhVrENxC
1Cz7ZFY8kGJ+Mh+rRv6mt01BUrxW9pQ6xD1KDs/UYEDKfV0JzLt9PWlU2gE4LA5F71acUC0DbcKE
72bgmtkgUvJ+v5pawSXxD48zGFUplMElpctYVOyKWgwbN0HaTTb0aPfA2am6sYd5OAkdqDX1wrih
RxITv6moBmyFuBqKcaHykGyaY4cLKV8PlZ1G044TkOQJloo5M3pksG/jeaLKUWI/w0cpDSyKc7Fa
DkW7qO+FgfWdCXXyImfC9OLjWCqNTRqoh+LO9nwvu7B+dOym6HKOcjENadYfUILxPVjlOmmFCi2A
hLrSOFQErXpdkyNULJCwruoeesmn9SKhbPRYysUBn1oYlNaz66fP0GpXKc+4FLXsFJ13IE7z6tkE
8kyl3dTFm6AJaZv9fe+1JjOIYOR1Q22vHheYmIMjqkZ4Rf2MF86+I7aCzcBZbMQH49R1uW8746eQ
EIybf5s1nQg+b0QH+3XuUwIbCO9uXgCyKn/gO/Pz16EHgLxzTr9BpYemH8ASMx2xrki8AWlz89kh
mtYMvaO4X0zaDMjHzXqsrrr/FitJIdR1keeHkdZ11lSWbQpV79I8gB6aol8GyzXEgVuIGnrQRo5e
GBRIsDBuUcSyeP77ddqq1jE2YW8NFUdOSGCRIfaZ07DL0ElS00lnpkAR/FeU+4yaPhWPsPaq5Gkd
xpS59tzsMLAEr2YFvBfe02l/QKK6AmYK2uOm3C6ryP9b0prge8QLpL2mJxb1espn+r73GtnsKqDv
zHEf0CzTcVZDfS9DrfCP2kCeOBpzRqRywQBulD81ZLoXZ2nH5i/kJNfrXcoq0OWm0U3FaIPALCKE
67crx3jBLNwt0gaasaIl7EhWrR3W3XlKqpjZNoMsegtTflBldN5/myVQ+WNjUU4rJHcw5EGhFoP3
g4Efg9wUA8QyaLCLDeyvuqBbUS8mSUhcCvLV4vXRvvD9pxfbmCAoYEahf7e5hDA2nzb6U+Yqh8O6
hIFLLrXuF4SDnP/7kmIAbYUyJejvVDdqnRtRVDZsh6CGs/lL4/xTKFO5UF30a/TjV2rmJWYO0En1
GaIBJC2tS2UcgbwV17rCp2EUkMd7eVnto36oToHaB2+QVd3fVsD0XXBicVy1yKifkmKPvEKG2NYa
7B8XFm7RfVxIrNmw5gPHd7mxoa9YHzUwbX7792L6yKAb+6DSAle5+9OllEruqh+PedizYd0BLHgc
+8mmInANvMi9CaQ9cslWv8ZzOWIC+4ZV8Ref3Qf95qMQCnifOVAR9QKGju++3yvo+XsYW2Edpbad
dWUaWhrxqjT7BQQJOUY92mxxlN6ftllXGq3SuLYVb/yCwWyd9rAOry0ZFCkNV1zN99IWbKxoxuJR
ak43boYvNDvVkGqRCRc2RsyxQ4G1IBKua/X5N4bvYqpoB7dpnbRi55vw7CvPIwE9slFuy87Az3Oy
n1e1ynL5utHHS9h8rzcecGxs/g3rtC4y9CSmeLQmKdty+d1EiPRd5gdFEDIZCOHkXttzH7DYKUSQ
UUcOVJReqZUW0qJySGdE4xQit4gjBg9z8gqYX4M2PxhmlWsAoxBzWJnQYICykUwIkqYhz43hDfRJ
ymNYqagt8ULC/VZ5tHVwEqSc99F6VewaHLnsMqxAOIczCllGDvkRBXHykjzCZDiLDIPUewmMBSYP
dkoxMourXGgB3DeCe48nHQAlof5XNZtrR6U194PXMxQCIFCYeFCECIzbXoa0dFUJ/7xRtbNTTPN6
kfMru6HheepbVhjEFeHTGxFxZLo8YcxDtGOfAV7hFMfMvYuXRcyrWbsQOwhPphpSWSMA1YA/yP3k
4/UWGhbVpi59KgtpdP3BAAE2FMD8KlYFdS0iPhaMPm6Psr0aAoyag/sy+6gno+ShGQ+NLCnwwSjz
WANx/wiGlrkOZpNjrj7Qbi0EogMmQAhhclTjSQOylyuVNjbGhDIowmp5veFwSYLdVZZm2G/ytXkM
+b2yvcPO+9vz2HRa6/UrjvnYFFOm6vgzkU8+QKwp/EwSpJ7qD82KWpevaIC0uBspbYK0guzw+5Gm
rODidEFOP3N+vHQglYjAH2zMmeqc6ffd4WipZObEXNP7xxjfTZayJLKaIOHOhVmASruMAOXPYoqV
/ZqQHWLlu9lx7Xh49yAL+lQi5gYXzxsHm81SrjXLmy3JPYUBz6s3+ASjOhyP9aLtHJ1qXwmvhDXQ
wChn2m9JrfEVeJcENuku8aZrX4pu04Pye9zX1UVvWI5bkPVn96Nu6GrKjAHydsfXAbIFaC1Ignjn
wCFuKbFT5JPxQWDdpbxcpsweemAwOSFUCXk3ZqGom5DCzEvUYnUk2XssH8QHw+oV5ovL69t/aQBI
SYGYwstr6oTSNBYCrU3F04iE09AguaZ3IIZnanmzqWbvQ55GsGjrm5lpVjFDvv1XoXbsbW9MtsJ2
Y++DFGgsPd3YuGD5NhoobtJdfzjTw2ms+SW4pcTJ4X0OyLm+revLiM6fTLdZAJiSyOrux+ErrhFd
AgakB/34vj8DOs6aRJX0/JprYtJ+eM3zhLxWg5BKBs0L5h0FoNKmJKASDjJTUZ7x0m/9hTeMdM4U
9CARJ04Kla+T9zpaHE5g/cIZlCWWCs9KMT/c4G01SadwDduA0uPbF8JDm/XS+yQTrpbdzdX8lziB
3Xa9o9Xe0vC2qfTZgWI+YuCFxsoP1s4j7BOMdvVBaxa8ZBaEan6jBqPg/9AQivbasn3ItX/fs8mn
ZhNghBAT6FBGRLe/NE/xf9KG67Ecy3x19gML8FKH+pQEagwlXPKjFEe39rdv2ZD9nEKyFkRyRz3r
l85tRWHt2SwWi3KSiJgPrTu4q9dFQN1fKZgFW7yg3A2bB5yE1ej4gAdgFeuf5LlO0KSeDH70P70L
2SsvdWag93GpW7q6OE2tMPgSJsDsNZToGnDMkME7llyDujLF4GijDwkgDMlOzkjgelaCtSNcVmN4
jQW6Q7vvU0p7VeTWmDE/Rs+V1ot+oDvq0VVq47pSvtVRUioTaddTg3WEc35eKmLG8lwISMMQSNla
mTJB9Tp2u/tvQGRIDkuhpChFiJrOgBeklaHVSH6eQZmyxH+r2We4GI0tVW6YCSH0x7MfSRNxPu0a
HxgIKUqr38yy/S3+ETXudJ3fDAWjmscI/XCs+/WONnDX7ImqPOdxtr3DXwE4y9ITFs9OlrLu6Z5l
7ln1rdhHk56GPaZkRKj2TPQM22ue7vFiihKn2tqRRs59NkCXXjwG5KFzi7gMLoaap5D9AOZlPxXE
hQAJJhK7udSD0NcylOkW+KRoP9Owe8H82153L+/Ud6mo4DRxqRh4WmoRzE6rA1ENlgYgLSvUBLP5
+7IThKzo1bi84SzQ4AGveJDILRwb3eEdTmntpl2jthxKl7NOORmK7+TJwbU9+ZasN30jj2VqfWAk
Q/WCd4TEX2zYkPkTF1Wsng3LEBUsLrP95CqRUtJ8E0ZPYOCKBLTA7Zglr2xhhQpBDFAwgYyA/kAo
zvZcnXqPVhHmn803avgFT16VD+5faOw7MyHSglkFvMKLZE5yue2AYIhCozRT3htHul+6K2Btjx/7
iIFPA0rQrzdul2V6oeZIm2muU9dnf63Cs+S1T59zRIzbefQnJVuLruInKesaEWfe6KVl34L70G3g
nfXF157l9+K1foNKP5EnovEGrRYGgcZp6Ga1TvsqivZ+Z9lMaF+LeHNUAiSw6dWyb/Mi1Ybwo1GN
MfoMpNdMpUHw1IdnS2Ksyxe0DEXZdhIb8Mcx0DboiB4+rXsBhr4y9NPL4dDBqJeY9OdBU8W6SZUK
rvuD0E+PPHdprCvrO1OuSLagCiSsZCG5QwmUHd4EfhXQpsmq643do/c7Z+R1PCy5fX2IsW+0ju+7
PPe7Gn5RekjcJcLr+B4hhFN2C4HBw2CjOm1CqWPHUSdcYxQAeUI8/Xx3+hTrG54QNK1c2cJMbFDc
UxuUpWsUz6EGpdxzpg9p+jYU5w2xte0IrOtqinpUEobEuIC5RIcLLX7zhI6lduzZzWSjTR0n6/1L
kELUhwrEe6Qv85ijg9tsqxX904+8GSOOw5wMn2nAMQP0vPSkau48zePJIVQ77jYk40JjOMPoAE/Z
LVXvuMRmo6Cub50Lgred6ZShOwHxD0h+nKpLdEzXCEqi6nUkFFjcM0FGrPiCX8nxe4zlhnRZQsJN
6NLCiHIGMThiNRlFvXXYc7evUbHNsf/U8gt04UlCuzw+zKbqGl7UXcAj67uNgxzXwKNMSHZNTwfl
YP4nqpOt4h6NUk23JfshgbcHXXK7rydzZ8DpgmmAJ4sizDTVTqmvA3+gHIGHU7wOZma0xmOamMM1
P773yh2JULdfKpnB/uOsh0T5PKELqIgJGIqMJ/2FeNBWDrDmVd7MLG89OLB9umIJRaPhVTQSv6s7
IzW/S3sBT3l5S90zGb0gVTU5MeoQYKQaYAyXn09w7jMV+Il26V0xszGhuSGcBD/qNfNrH4lq1BXE
O9eVTKoKTay2KzkrZd/lclU1a3L1tMdmtiY4mggo/eMKhI+IFFGiRQ9ahUa1O7OzLZ0/GUadsPqq
DChcEu6V4ve35q+fWgnaAVOVj00v8CYJgoAIJS/3fsAZHChwi+U7bmnxnBxZr9IisZT7nNo6gS+/
tpzFgxUr3FchxyFhvqHyAQPh63hJoYYfiMYsvdu414tJBvtx0GZMhL77JNRie6LZ+pKO0gyYYgei
ifWIMBZwV1EgsiXf/1oXdKtV1PezLZ0SzXDFPwNcYyhZB738geSDYYNTZFb9e5xXGWvHdirvj6Cr
DLLbF+zMAhFNJ262fFMUzS0G1DDqxc/aDaitk1wGPBqjHfcrpmDKO3p7AkYolIHd3cQaCdNgtjZ0
pD6IrR0l5rMFGqE3LaL1LMGil//p3f99ZRBtdt3egxs9QvpZxDCBNEOlF1b7jaien9c1G26zH8Yd
vurmPSMwyLunc+WAOS8gLGyep1xst718gp6kqE+k5agTQaoeQPK6cb3POKdYiQtds/Zild41B1go
PPqK/QlyO3LwMuaLAxznnL5TrnR9+Zw67WivOmrliD5+tLasU6VnyyqfPnPeLSnhxUGzl4Ch2N2p
qLUWdxXrCIfdCks9mGIUQQH2dbMwIF278RPAicgR2XKDPAE7houXGXJFJBtOxY0DkZZJu/Y9SpI/
DVnxFN460xVYoTJgwdxpcKa9Ktl/q9RN0nMu6E31zoL3nZm72nbulPg8t7oAiGwOky7Odjc6MYeL
s1z9qBJVEV5wmIdW/mD1keosG2a5t6dYIRp+XexOyhaw79B/Jv3p7aXbLvM4gXzVMFNEsc3o7CEG
QtZaGesgglqhU8wZ8GCTe6ZXN4b983INB29LoApmlsfGTbnfgLBHNjMFgcmHTDHOD4huUWSURpiw
fcaxQrjXh+zLfIXP10v021ll1nis+NxmN0wN5FQuC5DQC7BSa5v5EYZQlPaOIBnJSmERt+s9RYYN
fSgwKRem5Z7L58s2kGDC/p89RGNbxhWLQ6/Gj/UBPMCJDkAD/RXF6ASCzKi0vOb+aTygnpLiu5ff
I0/3IpnxMpRVHrwcC+1F5SMaUVroQl3ajqBF65vFn1JPH6QvbZcg08sW3c/QrFl2FrVjf1C/94pf
ljDLOKVdyiAVcoOb08koQGJ3tCuYKelf1WKl2tHbdhzG+CT98p7H+0mTbcW1IGcjaEcWGiRhrapZ
T+xKMdqTitWssXh/ke8sLgMgh9D9UUBwWoJEpypWy71jLmde1vd/Bw8xLINqPMJSXXNHukz4dCzd
pAdBuynQXoRTigI175iZsfkPcXsoJOMBAae17BpVg1lNqMbzVDMC8KSNBvzVn65kLemksLDcUHQ/
0ZQLS2shmTUshLQoV5mHz/LKFdUWjL0PGSKo9mAAR67n0ESl9KzbqemSbEA3AXb0TcQ/KoYjqXWn
/4CBIqDGeEtnt03sRUOq74T2WCN6JMZn8jg6wEkyS4A4zX7zwKcH/9KjJxL7xybIUWXe3XFXajoF
Wcm3rLk9zTuS9WUHe2AwAoAafROLvUpVB4mo0AnOnBDFujYrcZvCEhIhLN21MX4LQiF9bt9yJfV4
cPL9oz8g728lm0n/NMV55yIVaaXgaiLEJEm2RKRK+qPGBO4YA53hd0XEYaW5broEocxjdwTBR04Y
dEPOX7/qZStuJA4nETJvncSLIieMnhEKsBqwfLJwSLgSbtEwSMdBC6ibL3f24q7gVu/8m6/SLIm5
1uhs02WBp0O8LzMk/3mbKl9qiOMQsFKG3mUfVd1g6YrAt5Ft89faoCyqz1bxflmfdxo2eekUdj4Y
zgvsBtkUBxbze8lRpejyDNsHipWVVLlIQxk2OeIfwrqIpkm8Ka2G3ryH/1mJoN3PYT61ZuUni9hK
wYbF4qiT6+Q8guSZxq5QFkU7gcyUeVmMpBCc+CiHo+SYN4938BYoLFqGOfqhDXE8u/MZVeb1E7Ur
7b6hytX72cZrRX3SYu66tVt0Tu6nLHW/e9zquPryV4eVQDLjTyrKfXGwheF4tDMS53Vxci9zRvE+
entQ9FcaxEZZnL8cB+Q4xjmBYDYOZQMH5pbw6m5AJi//RwWfpIIUw8qXYQ/tlCHxystZGWEv0Z9y
DbgB8qwGfKlr/mCAr5/Xt/sMH640fgWKi2NVrjCJms//1ssK8IqftJJEW28GrMoNSoBxec6Q3yuT
Jues5SBie3mOueSoF3vELazY+jNgpoCGNpY4YBQpNxC7Dz3ae63T4faKPEoP0wGhzatNpDvyShnQ
t2jHC40eb7UiJ3WjfbE3u1leX58LFJcnl+0olsiR6J8i3KsNn5lTbibvKFjMKGK/zBMCCZYrnkam
C7RyhVGMJgd08xiKLP9ar71fiZzHhRWxX3ZgIZOPz10pnCxETNUeDmBOdHt8Vb+Eo07KrKAz2Zsu
8uOg56nsLeaaFBXiZPRwvNrhgPMt9i6N1yMQNSiB1mqldaxJs82MYu/ZjRyMI+VPTIQrS2CVPzpz
5FZiDG0aha39lkfM33k8/KMHuGfNXy3J36g9iAWVrAb7X+3UggRxuEQb+tgKf9l31Hf/SLcl2q4a
aXK8++j9pAFnrPMuM/4rTi2WfD29wYyN59jN5HOqM6HOovaYHV7Zi0oIjlw3/ZW0SfQUMeljNfZf
Rd/6mnX7Tq+2ZexMVbU9U/3ph/OciYGEjXx+uIAZy05LpEKZX67mdS9wrHivJBZTSu2jDlwWJxlv
ujkQyj86GTSFX/l9Z4Fn50DdbCcowMaDDHmV8SGvYX/cmz9obsPEJM4DaJvL655glfL3LGypiNMt
r+44QOwP39Im3AimDqrfyzwKuBj9H1qGUBh9rJ+TcpKxA6KORuxI4gh09Wn1gZnCTJ1ChKQ81MM0
NVk1sTjFVu5Z2G0lTw3u9/Dx6XHZc7QnFoXEvQJHdetFNJFlaR8D3xQ69SDOcGX6QFAjpdkxvb/v
rH803kW/P7Mx7L65vqZo5OcU1yKjlesBe2XwSMQS8Vfgaixxhjs0mSxiRRJGJYrdu+ZCEPE0buOl
D7RG2cF6sgj6k8n/J0V86t8zP1mEOUPyQ8X1OTcubetEJc3Sh8PB05iGLVbaL53dZlc653UeWF66
FAH/cePSBBZsPkZi71JxyZmnOp41HC5Xi3w141S3yAIjkcd8nR16FZNGMbem4UrAzStYB/jA4YaD
taKRCDA3qdim87zHeAZ6zTew0UHZNAZ5M5KXQeXHYjHhBaE7STpahlS+zfTdTyRumIEgGY0TLXRw
3TzMalYO/YvfZ0hgbRtYiAhBUiloXxhtVZdpzpV/0yyXpKFgN2jyRTImk77a21gy9+TfeCBMserl
1UvTla0JnlQNbLYZep7YPCnjudXvXRz3hRezXPZktWnEfShU4vaC/YClKtgiIcqDuozO3gOnBOEe
RiZw8b6d0RAvt8lHdWT1idxZrF4LBXTPyydhAqm9lT1pZcNSkyLoCNC/ofogedGz75IEYF2bUK3o
Ad6hdnH0VV7dLNxiJ29y/S3cqUbG9dmpKwefPyc0FnNmj7tBMwfz53EqOwkr65WGhsxg/TOOYDHC
lUzGoZf4ihvy9U4FhxCLBDmmib7y/tn4wwo7Xs6pyXP4J4sotV0NdGbLjbMCVGseIIJV1VOhDeXN
gi1tEEvST5by09YdW3MjJ8nfUmjfiwfq+8VwtogqV7lqWDO84a5dKF8bpvNbppjaLI7ZjPitk8+2
dklzazZvLkw4yfcZshD+f1vjNHy6ztpSimGPZPKqxeJZ+i/62un/5YF5mRcR3I+LrxGW90iqR6mU
kwIdsEAQmgA5i+1gXzac3MAnpZ+t4rtMZRn6K3+HEX9QDkN/LUMBh3dzaQuNaevspjkIVEm6408m
G4SfGoBbd5lqzEfeJb5AhJ25K0uLT75foyOp4YNtnmqf5iZv4fWExq9NnObGwkb6tHOE/Jqv3ji5
R0YxidSWcixKZfkhp84+ewHy2QYvn3A5NQIBd10HxlBh91gqk63rS+VrsGGD7EmTpzKwIfPj3Z0j
3viJVhsyMeZj1RndGyNTgnrI4kuEjQTwddq6s/6kmKmWNbWPriN4DfKxtcWjkpX+aQ0aWvH+liS3
7WsQzt+wCFI0SZVcSapBtH9YeInWaR2+gO5+a26zE2x7fxEyNC/tbgyE3AMk76cuvc1BXYMcToqs
YTbP0P/LI52j4iz85SZsEK4XtO9YmXH4iex6sxwnIuHznh5alZD3V7sWChh5VOdN8dzfN0j3uxF4
QgO2gq/ydQ/kfVGnDf4smsGW24yjNtV2ImBJ2KaoEeS4HbZ7oUu5pOGafPqe8tcnLFNQQGxJfJN+
HrWdrpRwYl71WLDnBg61pd3YkXoB0rcpAJ6wGzLP5aHJ8qeshcuQxLgRFZ2Mgs9EfI+BlqsfkUXo
REhXOJeM3bbgatXZeQ+shZQvBkVbupy/4egooUpVQcqbuNE6KhqqXhEaBvsjAsoZBHSJ5JWFrbvk
XFn3ppvHhWMAGQOwlEcEfKyYtEpWGnXUBXjj8epfR6SZQxhbxX/zflNujpcfnBZgwMo1A9Kfbi54
hQS4ADNGHp881IpgYc6TuZVdrB+hx17s1GJ4dAt4/R3atAx3TBYzKd4hYZW3qbg9Gwp5v56QAfYE
PlDOlSeNPDjDXUTWk/FvMYqSQvdtn3tatCbDiSHTh8H94xr6jUp0qQq6To3vGC2LMFhIqamsCAcs
1YR+TdcatHRrgNCTrN7voq0a54gtya67uXGKIg5uxWrKUntwKgUBBAxW7e6iCVOmuPUr7wxZpk/F
VWQiBjnmB2z182Kr7fZd1RWJDLmelNlFKKP8xJbakUqmir43xrxh9xFGXWXXqu273DX1xYl3uu0W
Eu4oedUiGun+bskUgWnRVpoZUD0VhWsEmDg/460201lUCOfHzNDf65D6B0Y9q/R046ILrg/4dIjo
D3Y4vdsDdRkGoLOh1Udw7Z6fYi6x8aOzCPuSC4GamMuQqoB0giMDvMyCIDSVOgpM4yqiaHyQ9zZ7
z62OPdhQdGcA+Mwjyyeq/4i5pgo1i50I8+Qio5MOh7FsKshkePxbO/iUc8kDoK9ZlXLKt1Eq7SUZ
3drm16Y25eZSaezoGFqBiwa0lDyqyjqebzoKfM7yyYrftx+uMCiWJh9WeDg4EUD733wJtY1ZSJ/s
IwAFV51x+EmOVF2r8di4H5DN99rQiNMSb/u5Yy6yIizbDyhAOQFr7NNEWUuDaV2Vb9nIueSZTv4c
2CcM6MnJWuWoO9mNx6lDOtcgQMYOZK7834XSnFEzVJMGADr7OETEk2awNHJdS9P/R+i9aivuzwEZ
KaATd5AnQ33fHMxijGvWjvz3JS3d79EpHWKGmAP/fry+fwK4C8DJsh8LMi8GR6M4m9pyT2cm310q
D1FfA2ubdzBEtKJaFfKzZca5CvPJaIbOa1Dc2ddPMSLX8I6lU2TwiNV3lIIblzCyplS4pLz5aPWR
5TRKauzRFh/7Fvf8WuVlAT8+4M190ne0R80l8dL4t0fauzEcW9LdiQL1LmhLyjK8ZNTvYjzDQ+/w
WPBD07DjLVZAk1qzXkphjBo8pPtzUdD7M34gCARKlRq2jmKvqBHuU9CfWKdyMi+LrlUgM7nGu4yC
HcqpMj4kgUrrpZVQgtH/E64bW7um9m3W0NHBDhIqhyOFeQktG9jdUC7ZpCe7O/0UVFibMQpnT57N
V1hMTlVIA8xTiRXPZ658oqfinPO4tgYhk6UIEH51L2U7FAx5W3BhOrtQ6++mIrbayQhILacW5Yf0
VcKnm0ENArl0USXuKOwenoeN9Nnu//muILoXeBgbgvUWEmoq/Rpa5zwwirgbIZo5fo/6RFXePwZf
jcikkWiVJeHxuyDXpUix13xKfkY/h7GGy0DVFeObxfpdS6iQcD/miy3A8/Nc+cDU+OWIKvwxBEq2
vjEDODVC4t//f9mF3g6UH8hx385iDy4/rpvnZvaRk/y43lrrELOAQakuoqd7MohjR5obFM7etznr
/ztpIeFKnTHEJtIWwqKoOCLC5uIce/G93chdETDmivv7eBwNotCrc/ltPqSTZqbfLbBAf/iKHgaN
T/i/wWsBkSctaBDv5PHK6tmMSQJg1adOkHjcQbZsl+CDkO+vmW1iNMYElwUapbyTo+7PvL/4t1Cn
urhi+zp0uvgHlPQcEp/DaeFtwtHH4JO1B2BVTt5eBteRBtiizDmeNCgMy9lsmw6jg1kJsIHbN3Xy
V1FXeuOxbjsri0Rm7ShJUp2XkaMl7Vvh5guwcNr7VX8EXdCI3JZZSu6wQP/UFhy74pGDO5gym4Vm
Xf20WOZo8tLRVjkSNETsvwlDpL3G4MLqzbHtFdz8GPMVKD/MycEZkor3d0UVW4MoK+rw2x3J0nv6
2ELDqAUzHfs8735Rm1XBJHzk1Z61hLAfzhEI7Ep3EIDx/Q1rPJY+4ayUfdLdBAktr4MTvETGvIst
4M3jv8eoxsQrTTRiG70j2nTaVEFQ+IqfeUV7EkaU/YORcoY8Y59FOW+Aet5SaBI440obwXu5D+Yp
z9iIn3Bl2FAz1w4XqJlZQaMPZ8BtWMt9fyrV6nAz/wM707L0uGUrofrWqn+VHYpc1cndBGAuEHm3
7N/+r0uDN0Wl/cuEQEpGK8qAXRRFMd0pHLCsO+IPbN5AaULjDRB/qn8YEry98Ol6A7TuuULrU7ps
mfloAxC8WoxUfCv+q4pu4c9EX+BQYlAx89OZ1B8GcixnAma322gRlKZetfSs9l+HdJHXMics0R2F
MHyLkQRd3pBJk5SOaCixOns8qIqyfeOeatoeCsxJkK7zmf7nmZWa/yhB+QmzoL5u5YU+78bFFDGL
vtS4fQKBQSnXeUhixbxTEJy9eAaWAZ0QGGhdMqsoW9FSTv1WY8jj+W9AjmOpFecqz8JBjiupWHU9
7CP2b0lIzVpVh0a1qOBmgQc5IUPDuCuxsCWE89TKfD0AcbODQY+hAfFE0jqiRMjXe9TzQh9F1n/F
gvsCUYFZHbIiw44j/1y2KBI5g6Ok/kQvYyECrqEZ6LeOY+qgU9nCE2uruQTd4G63RWU+Yb4Fed/Z
nX9qzvVU2zXYNAPgcUeCfmHBQUFPItn/Es4GTCEKZQaMrl30krMFdWJMKNf54rMQaqHqJ5uTJgyZ
+i+GByB9RSuv7wa28GMX6SRKXMfvdz+Gk5vL2Sf7vYQA6dgoNWSIflxXvmpu+j3SznGXmENVAemF
ex3jLj1pVoIpH3LvGBeSZlEDV5r/XwCwnVBH57fvQpCMKZcWsY12wrm3Fp/VC2noJllFbewMNVvA
/q9wLmSH2QoX1InpZ1rl3v6et1eoLT1pBZ/rzXnOMrnk+Bz4zY7z9zwgvXEfbCc70pX+YW+vJNjs
KmzdBJFjAEi3A8JpuD97R3nmR7UMgSCVv7quUADmipdjnNnw2K0AhW/nNdEslsKZLid28QsllUiC
OIOVqcSxckFLf8Oa5y0l/y6s6jSMR3u7tHuMJjn8Mfbf+CyEZVjDx/nwfxMTPbWrbgI67kEXZHRy
4T2ULwSaW73GcKn195UOS6HuYnsY/idh83tdsdzlS6nHZIExvnn8g+V999K2SMI1I0zP/Hwfagl0
FMVbrKsYyGswPwNVtjGpI7N0nHuENfJR1ufq/8mesnBdGifv9zWiuNm232jCbRsdmHXRQo8C7ULQ
i+RqRvUY8CCQ6J5GHgkW0B+4wr52BvAo5PxJsP4qoedWsklJCxxmuuHE6TJrgQ55aZVby+rvoEiW
60f64zAz2UFQgjf0Ed65KcfVjMLIcA6B3pA46gV9YmjgcJPQxz6K+8/h5DI2WUq4Y6IBiX8ntlTo
nP7wlANkHHXZvZZo4xZ8IolzJeTwXtqicMRMn8xybZt8LpMMBakKVWZ+7HrZ4Ikq1M5dI4tdCNvX
xW3Sf/vxrAwfotX0RoX13pdN60SNedaOuBpCxwWzQ0ijX0tORq/r0QSs8+7eh5ff2xOjnokuBifj
oUiWW5n3NXjxjNYbvVZwjNpMzpi1Guo0l2u0tjHhMuYPDMP1IUrf3dAPEGe5xgI8DZfP3fII0Eax
F/YjbM3MnZMF//fFp6Us5LRtqO8FOUNezj1nq5F1VX9rwgCkWUZpnsKphtrzyVBZ3a4BAw4lw4Si
iYLIe33xQm8Ww4SYPhnqlkUujhhtZgpHAuppRxmKfjVTYwHY8O3xQaUboviwkL6QPHR2QYqdU6IJ
DpEhlF/b4ivqenuIIScOvyfbGhJ/W49b/ALIThijEklqWckhaVzYfOuY/nNMGGJoK7pKWbakd4VD
O2UE28Z7dghM4RfiM2F//Bdqy6Swxskp3XmX8swF3sZxzCHxew1y7IiuYCHYZH4lHrjoGIBXT5O8
y1W0k89xuzIW6+xCNiZt0aGjZFhPt9vCXUedGk2inAN3HgEVYy7J8wAfM3l0jODCZ6mPdOeVcMxR
Edmd5j3CcQIEr7bNZTQgopFu2AuM8qQzuSoWFaf4wI6Q1uuatXfrnaroySkhOli9mLGZ284vLg9C
m88FNVuqZKjNSsCqZrNVvcJ12u1CcZ25f5ic3d+FhxVxrQdpCLZSS3OoMmQ96zMgWtQGjb2HyURQ
INIgFtghEuJpLPAdykpg6B/rwmAZqCSla7qxrcM21VML4G5KH3Qlp7azaeL2wFDmzwH+H4FotKLw
ch3rPziqWvbCvWcwI+oEKuYmvImDpK+yR3cf7yRQ3mEyCdZ0PMLPSOtCfH1lCakaqLRdrcwcMwuN
GLGyzsNHXnG6AfKvGThAeKqqNpTQmf97HVicq+msbC+NTsBDF3jkU8WZWRNCqd4fuCyYi/w99xE8
AWOvzTL+TR3qMTwruf6qKEBAhgXZ0OOHRJlKDhAJupkHZFVMtepGzY+uPr4KLOu2uKPUF9qWbM0c
iOsg8v0dr3Q7Z3Bc7IxyX+eDwETLud9DvmqCPkz3L7ssRT4EJWM0bzb4ljDaVV6mlaE8QW8tv1hs
zNPH/aj8dR0dow7fhBChuV3Uoxu0T5FTGAu0KEiCdWK5SRyKAPAsc3Pv5MlkCisvTi5be2u+EZXm
YqNMEjiEU4nhy85A1ZhEj8+PEyvd0X34vn5avGmOSXfpdWMAirui6/Y9BHzPxKzFCesOFWRV1gAJ
zNH341uoCLOTZNpvftKXEWqFjGQeBz97rs3e/nDVWhUycvB5Ks5MXvOb2vLoxS+X/EADqxeKTwZl
xWbI0Jsz3k03FBrs2sj3K4KI6MlQ88RhR4TcXVzNHUDvkBHZLaY2zL7WoPGS87Jzv0me5wgAX3gY
jL8IaY4Tu0X+UWaKd8V9+9TtaB1UCPN8MtWWaPTD0VN4uv+xTHyxcBViE+LheitEvX+MX+C7ub0o
gluFmg3AxurYl+rgliPMRtKHShg5yiSnRDea69kWNNzZemT+Td8yl5kZ1ewQPl3mJx+KioHgnipD
HIwdxaGO7IBSft6AbChhWk7QdS4U5GP5O2gLjBKWb8pj77kM+qKIwx18xnz4zJ0o3bIu1nhiZH2/
x1ZW29LQdL/Twyzw9eX/6zt78n4/AseBqhXsTeROkxTPgF8GKhqv7hhn6+LlMTdDqykbJfyoHP9K
i4/Ao252dPScFzgJoZF6blnH1r77okvCZ/tyo9/uNzbQAvP7wAUX2bbYCmiO8/Hd2Kwu4G15RUTx
dbL3yszg3u8ZmhAztzVHUcuHd4wU5v0o/MgWLTL+elvF6i5gREvvzV47opiP/3Zrs4D7MWKmr3U0
vTOSADCwTXcx/ZCJ8U/OdUtxIBHLtXIy4Os/QI6q4RmLWkkW5DgHfSFZIFjCLfr4BniJxWy9BlES
aTd7s91I1OPaLaAM8bJ/QxMjjhJUYKHvJDyBAq/6RKkvgHtXt5jdpbmYpLWtfyI83ZYw5A4LI5CD
sDDWxzduY2YJ0gk3FuoGz/IMffNWza0OFGEYPM4dk6IN8bfxcgOiboZ9XgYl8axse7VgpJ59J8wh
9BCvVpef2axE5hzj5WmL5RxrElAcX4RpPq1uG6dXV8IcQjZ+0Dg4R7j+xRjuIDKEE7vG5xpOZzNW
mRDPV2IwC5F46A3AsDdytNDdyFwTW6qSdie9Ykhf3a5/VuDZB3uMtrC/q5R4ckBhWQzKKzaphbDK
n22RqXJwvj5zinyGnmks5pJedKuPdNkBnYX55/SNBY/Zpn4xTfWEEQ1rtrofU+sM1lkbYixIGXZL
NWoHZSwNxfaRSs1XUltyoz/4ASvQxRNGDhvKBUqIZUswG6JQ5fZoVDy7ESW7xJ5yBdJkrqYDP5RO
0klkfnahq0uCaRlvlAB3Mwd9LwmAe4PmHyFK2N6ubtsKmmfYDTtGJkCV28hqRKapykdffLJkav2O
p/Fn2GMEAI/iIPY9568dqTKDJiPLMD+L7mOi34yOKWeCcvZ0Rz5yG9ZmW4JlMab+mvYK0asVstVH
B9mFAJ8oSFVSads8wxfzrkMCG/f9EpWTqb5cRxXaXoXjei31c6c7P2mxD5RvI/qjNSMhxUF6lXQ0
y7Q/PdVRnLSN1zUQSnt3pX+9B4hgXxlzSurZSvGvwl2B10NbPEw92BfG4VoivSL/5WeWX8dWo2bI
gv542DtR0W7/UAbiW7X07/XycvX6g4PrRusYBJNZ6haIrZ9fdMy+Os1rlSBkFPRfri29sf4d8ogy
NDyWwOWiFYlSJx+3xNGQQfbotR2wTl4jsRWXslrglY77YMXKJb4CJ8Dna+mJBvPLlPgqiKqge94O
pAdvlPNv5Ds0EEzCCOflPDevkq8g4syWFfk66QnqQvO0zzIZl++Cb/xFMe7lcNJcJEIelgWxaQCF
ZzUYnk3+7gDbZ4xBkSTV+mdpQGZ9kldM0itiSSg5lY62sKKPdvVVPGBsMBFjFEDljirfp5+EpaUY
nMZNVAEPEOnO68QLItNALdzYubYZV6SmsgX1YOiz17SVwobp7WzDxM9CNOlFhEHP/otdQbcP+Qtg
4EHnFU4sel60WWEhnP6xnszdTCwgbnjv/Ys/ZYc9J0ysCgXymmtkqFWjP8Xsr0obIQDRF6gu5RO/
NhSi6SsBnNSnJsWoFzDMqHLfjmDAJ1eH0Ef+caCBt8nP8S5z6Dgi/fkY05VE/Dm30xHdFKLspXIz
CxfZjgrmu3TNj5rUSD88hqlL1JLIR5CdQCeKQVcGCWB5ZrOGGwJtUrh8e+RmAMqLBUJkSD/mozI2
Q4Rxk3kKYlSOpkXo+Sv85sHegpUzpJ8+8QK3kDW/TofvXyncnjHVj84YldS5tJE197J+vEzFD1C/
vNByDRgraNsosojbkqEROmrCFTPWsaQIV9FZB4xlUTcVsAVGF8oGJKi5XSUgBp3il98yNdw1Kdgf
SBKG+VfLvOkPbQiQIkz9YJtIIvJoFhTeSUFpYHVreSpAjvVQVCmMuCweIVHwNYFDwWY5dGX3WJjp
kImD1FGt6obzo2c/4bPbKoL1qKFKNycwRjOpWgv1tHhBZgNh+mw/WWRK+l1QeC/pqkwyCkTfAxXQ
0ztaO9Lif9Ybxn+2HlPMBezDOpUDBIbemrxWSb/Z7xpq9OB78sU+K2VVIhRLZT8GpyOF+QrlHr4M
+zRIkgJUDKkAC3LZ58ncj4acYGwUn3JvUsgTzUyvVZBFwOPbesL+BzgMnFUrbNtX4fUUgZ+Wh7Ft
Ktzo/mNqCR5/dwJOLvtMhX+w7rDAT6wL6xFxehoRaoFYHIOnW2PjKv43HKtgmiNimccsocND81BT
au1OS4KHYoxdA7Ou1kXoi6dfke7Gv26v1O98Dq3KRHmwuz0BJRgX+ED12KL2CmihUFjVdRGCZ0Z8
vyAt3tKuKZ6iBRi7AEJ3/hCmbaKuybwtRX2Ng0YeD2/fc+zqkYjfzcZ5eh7KoxIcd9FcwbB0870n
z8m2CqKiE8FwusaQVfIHjvTHVq79PdlfiLTrJX8+umiQKVXPGP3o/RryZH2N/fXdDTm3IX+wT7ji
1nqOopBucuw3vns0Xwhz5roeVITWU3B54nzonThq52J1W2pxlF1f+gm9NcqCrBc3U57oJf7UNJ1g
7tsb4rex/tAINngWVNHvn6UADrxUyae7G9JIxZ3iTxHs+zUMCxdoWXPVR5jR4cO3MxGwAcfZK21Z
8IljjgfFUY1Z56FTPVQcj+BJ5YrkPXn2go5wmyev4BztrV2MVWFw8lsrdHYEWgn/eo+plI/AOeqG
DSxoWHa17XdAgFRllkEelHsM6PsYimaGFIcEimdPNI2WwWfKi216nTWbYnNu/VBgMKRMRhrgtvn1
piqThu5j5zjga8+OhSu8ZTeh5G3kSJ1LWVlb4aZZjg7n/K2y9B8bA93s5ldAfrIJeusOXun/mKPr
ADLuvchINj4UkL7+8lxymKDTG8KRPLdp+S0XMdNwxkmgWmM89JXxxTmDZpGGO228CAl/8QEScVUN
bpIzgtMCiN4TdnPvuoI5ccBYW5O22lcazF4Fdu7SqKYTsZi0+Kd+IqKUQp4gyBf+2DEB1w2uwMfD
grSrSj/bMnPYpoj4+dvR9+zV26IMxqHwrhsPk/5WS6nQbPDBo6anfxFcnRANjj8nOjGPmEA55gPm
8HTO6Hl47LjWWQDYV30xIIbRaW5mntZiX1kw90Rc/LQDTXrlBLw2GM90OjVt0aEojbzA9AAdXx9+
wHL8pSf3NnD/OsDdfRmBAQS9ow0feDoFxvkcZrgyZdSjqCoKJnOLLSUwBeEqZvMLJd+JnpWculZy
uXmMS8wEjscxmWHGGdTDZZd6GRRCG8i/nr8QMWesbPZEDRqUopsuEE0cuMaWNnHTRSS6Dcys5eSD
rTfTkKEUI5rt6nHsAQJN30D/nldwsRaa2pI+MaIBSQcPElX479P6u7QlyVkmNDQNw9QyqMR8FFd1
C1ba2ojMg0EQh2Ted6f+08u1rpQluHZ6GA1n7lIe3+4ftl3oHkIS+t99fFojP9BOWcMyF5qH/vv4
WA0QSIVH5OOor1XUVn15nEgmKLS+m1S/NuZcYTa05z+L271J843Qbq540tYbjs7cXCnoKogdLAtQ
wJ6Dc5msvvm1b8tbDn5+9QpEstDScbyCQTiR6PdmJ7d9e3qL6Fvh2C/nddPs/0kbLoCm7BHANCjt
P7s5CRtgIE/rcAblmrDZCRVziCEOiMdrbOQtj/SmaFekgao+jkW5jluwGfDmpqgKleBm+g83rmQR
Chs84iUq+J4hpVG3v0NIvwp4O7hb1n5cYHkhy1FrMHTDI62Dvwwz6wNdanJ6fLyvxLaILSSZm9Zt
DBZzv63OieZHhYVRtL9L5a7VQ2JAfQkEqPO0tvA2ovSbih4lk6lLwc951OuFOU6zqSB94hZ78ytG
M9zI6n/D9WjDBgwbAhJSb49RTCXc8LazbjipF+xgQttfZrjL6SsuEQiF7W6LJaYXBTBdZCLSTOj6
F4uL5rUDoX9dpS3PP0jTPGHeCJCAZuxFA2cAvJaNKayDHGOQxa/r6qIPc5OCyf7wE6qrDq8g+8ux
8KwJ8O/wkktWGMuah/RPdd5YWq2N0/wHu6Lqrg9u08FSvCifgXuXqw/RHRkl/jIpNxrR5y6cTnbJ
kFs3y8zPmM/Uu6m2XJMZEn1aqVLS/kukCIFLHv7GK+SXeg2Kjsdz271iL4g4H8bcYnZS1Ym1hL2y
pFUnHz9HaQ6FiLmoKTulbSjBJ4neb9cJt7h90PobO0RKyCmmNxCSTBcdZCVrh0Scrx5aRxvg87vI
kcMQ1OIKKm6Ztc9YvA5LBDQ+Ug1a+OR1uyE9RWwySSOkS8X8HELLUEe0bDG1uB9NpNK45sUw3W0n
5q9QXTHuhMmNOp1U5Y3lTHD5rDiho60epVCelNa/uWkVHUSgY619eIlPN8ddJ05zlUjQpdxSJqoS
+Oo4MiiKAM1zIc2Ia3b7F0BB8s6wVfeyCz1cXPuCacz+RKGh8AHmPxipfLqXyA6i+rUSjJKn63jH
BKhMwscLFuBwXD8sgBh1fBaNWTc8/XgEiCbVU5YpuNkn6dfGqDcn2hP/DynaedpqVAmlnIHHDpdH
HYoyi69T7F5BedPP1RIUZG/1e7PHjBLyKdgi8G3fXkexjkL8RE+dDC5x+akd9ym0LzbOdIqi4BhD
U68UUpLfXOkATLt8wwU//Th87NL6HdJLsReeIhv7ylKO57CHbX7ygfJyN74Ej3eBn9hxOe0/yLKo
Utxjjcnu0ER8JfZ/nTtWJEoSU+vGrnvBnSeSyaq+qwtAaqxbR8XTgbRm+fKKmsn1hZTHryQaMxnR
AQpfgZ8VzIYh942XLqxn8pWtat7NRf9LxGNr0aKFg2ZNMqDDoQLv0dzBrz+ROPBF67+7WdEjfi8t
DriKwQQDfiUqbu7N8YpduF6/BZQ/IQqsGu3vSBDMj77RMCTh+hMh3a2GOKCLDuTAOj/VVgDLLUpT
fHGbCM+Ubuq0a7IiXmRaN+MJO6quVOMNoeIIyYx7VvSS5CUUgNfHQKnRQ49odpe6tZlmpIvkn8pi
uLHIq+nrY6O2hEUywE2utePewIk8QJAer5X00CLQ8f+qLpsiknUTlUGEX+D9DtpFgrXw8O8nKpbV
SqqTRTAPgbRMl2cTJsBcYag3USXCqodU/iIiYrFclyDCjOFYx879C5V8PoyRYPpXiVLi07Hwusbh
qAxGHMx3W+iXjeW7C/oBe4meJ/qPdBgrE5uND/y2vJroh4Q2R/RHvqgvQ+7xX+MNjsyz4YEIB+la
HEaRKMy7GSNmcmsHVEsBNN7hF+uW9ubZZdrdtTKHeIwr7qOQ7AvpjDcOMDX5xvLotP0NgKMCEPdO
EscefjSFABwwF64IXWdBd4J7JVtosjnewPzd4kkkU1LiNqMWZ1j65P9yKB/8AGTvvVEaZTHZLnlX
tqRbROAZ3oJaAU+FyAh1TmCTDVPf7At3DMYTmNnrmsiv+2zB8954Wx2jGsKuF3Aj48SQ46nMjj/2
6DjfYwEFa1s03G1ZXoZrl3KgxGQWVvtD1ulHr4kPdMxNJDfWdkQnK1c1E0k7Qokbi9gzk0BgECyN
r7loq7swdfCkfwDpFnUHsSeNusNBYxn+SpCGiz/4tvK9BVXT/TatudbAgq/nIqWS0oroVTlOkXJr
CVlw8ikslUu3llokcO5ZjzwinF+XxaeMH2g16FlDxIgFm7X02FHBT6fkNincfcqC+Mr7zbb+llrO
zdrF0P7sc0zGkGXIqtQNgxw6vzO+BcwIjoDfe7wQT0UIvMOLBSChVxUGqzlK1EjgwFlPwRyyJFmz
AcMlWUoFTgxdmwmLBcbCcU+y1SihJwZ38nocGq7j8UaRDqcxZ4/1GPXGZc1Z11rPdFEkbp6DqcOj
iTV7LHug5EcRFZPK3WDZ17dOCgHAYWpHIYc5haer8NISxCx47Aa5Jq4Qg4TdVU5fKW/YDO2B2Zbx
miT3ZF+0qZIMrZdRBBU5kPdMd7Nkr3EG7sXlWwIK66X6oKO031VDt9Wl8rGyZlihd6EtM1WNxs3A
ocyj05x+oYkXwkyiWJw+E4XbJOtx8DNonqqro5BplnvwZF5yX1LjF/gAmgKT+bNadYuVWqSrSbJL
c0mEQGd9x0Xau8udEuIPOu9DOw7J1X2JU8PkyGYQPorNgGzKD74bQxpUhMHtHS93Ya228e1gWsxV
zA/GQGB8FuPEhEqDPRHBiVW9lhUmrd+5JJ80b2OlfTlnjEJwBaTgYNtPIGZrU6u7AQtNxeLaEsf1
kpSGZfg7WakagCzUL3LlwpSgO97DMTGmdcH5bVeossm8q/EVSwHHWC38mHbbeH/XQBmdpm/eNrte
IL77s1i6II1o7eLCVgo2msTK+UluRf+ly/OA5zFmAE+1ygqPwFqd1+IvunGZ9NCc5tzyzc+P4lJl
iRtFjqebZ3igxGaLNPfIFhspoLHtiGAONDaC+xvJl0jCO/ZKd5/UtUdTALFsIiS0SG0puvDHZMZg
YU0ugMV4Ve7YAxY5z35TGNMWLLS+u03gsowhXJ6xinXeN4S70pnwo0wOzUxsomR2eB+nqEEmx1hX
vyasmkACuHUvZNNQlvHzkaqUs586SN2Z1iNn+4AMmpbveJgSIDP+/ElfHwzKYFwg9plwWyANiT0k
WuOyifmyJMVkrGpjOyY/oNN3/7Jhc9RPvvzSLRLgL4LUaMSc5AR2LoH5fHr5WNSiZGitnXW7da3h
+iPP+l8V6A+iAOVpOdwZDAiPId0eNWJepnHaOrZBkOJx7zO546LpAHGb6O2Ib0PY4UYhssrsiSZb
cA6/tiv6nLfLJQbfavt8eot1EDeYv1/JfRtNXrF/C7z4X8yAf/euycDcHbCOBZv62R910lRzg/ls
0/ldaE4ICeXPdxYmgl4WXuVvVYJ+5aKQF3qFcdk6HszPT8gJL8Ne49Q1wFo2+7QfAr9HL7jLkDPh
zeQ9F9zPB7ySamqWqGXsbPVFHnvwna/fAm7dOGAqgUhuZR9agxc58jl9glNWI7IdzyU5JSVpJr++
ny9CtDCbu/G8PUnYdiYvr0dc/yDceBpIE3xfevWcuN458h9oAxQ+EaRyaY2R3KRZ9sMduL9mYN5c
gxcnjtRfbc+Jg5trMonJ7h7FE714hov2hCyrCIeC/XGkJK3OizV+9QhaZicqV/245ylYaoJv9S+/
HG6NPfPIJRHyZ8Ep5C7pXA5r71DsP/fov+gvWUVwR5WfdM1UaZgbsOZ4RKJvNKpbhrHgChJ+XShG
HZy4/A/0HXwKy7l7Ye7FsFY6tOjU3ObZTfmNRSXGDk2wjZ05Mv5cMZl+O3bnhwMgLuER3c4e58vH
u4YmwQPHZrBlHMjZkmaugapA530cpF8HnKhU1CIIw9KkwnNQe1VrhwC8INmaEnHjG3M08FYP8Gaa
d+O6GVEgMQUu8PfcuhqOQuFQ8+V5W7c5XC0mqlDCOMXLWdYEqHbUdal6saYrrtiXESocxOZJqt1l
RfUzCnrlomZCTAia7y94VumxYc3veUc5Gi2eR9OUexSQ0vthi+pNBbZG9ZOBHDhUA16LZnBDq9Aw
xdTWLMjXpjlmT1QhH1s8EAJFPyKA5XTC1q5HTMGaoz7VMnKz8SLqiUVNi1y+MGY7K1a3R5a5fuHW
HsNEwuGnAILWyk6GNzc5xsVl3vgucjkh12QmpVS90Q8X6l+ldAfBA1p2qk0fgKAoY4eGAt1eITfj
KZYChv4WnPjmeO0HozGtAxQ5wdjncZcxu5kFC8SgFc+iClMK5yrr52mIG6SQz/VxLAuk1RsbzO03
XGANJWeLnIkTOMXT9lnYOwH3/c4ZOtXPuH7nT+7Kbk3EvniowIAnmERKlqOXcyxV6EkE7gYE8P6/
YmQ/XhusmBSg7YDXYLnJgb7bLQ0aoviW7q4XeMKJW3H9hLSzDvWp2yB/oht4+MYAXIKSEeABEk/o
hHQ5k8O06a5p++6YOP5vazh6V+2uBbf+8cjOfx0pHGrERYgrXyWsRcL0s5f6VvlxBGvFl+cCmYD9
qtBN76iD2LpS2EW2/i5Wiupbg1OUbkGcq1sYBku02vH0ErAOj9Em95Et3JLrQAUqxxN31YVJ30EF
rO+1QQbUw2/FjvkfHWkIhEISHFUGFaIr+ouA+wEtBsNB4Adx/PSHoaf3gxP7umrvCYx1D6TfAOHm
pcgzq/AQILy3zd2rL0Mq/8Ntcc9jlvG8HfFUucCj/o7g5a9YQJDIsh/ZNty3WapaUFDw+TSa+DO0
RmuyBBquwXDeSfRx375DXYH7sbX0fzMhMZNUpqA3T1XwCGg/7zle/sGh9xF/udkTJ3wShT5tAJqT
vwv4JYS0ICTPAFbb2lVr4sJlvC++r+bETrw3a8CGz+WcNLEpP1i4moQOye7YF6NC38wVd5DhwvNP
e8kB52DxowFnG1zr+LMJq+7fKaATo21C6v3oRSjU+AEqDgMnvZ3iYo4jDRz3leGzvAQT/tZ30APJ
MxYd1iT6qkuhdycF08xy7BCvPtwCSU1qgg41fn9xc1YfUK7HTxeEpfJSruSqGk2lMQFPmvC8CJhX
m6dYz4CW5REccL7u2ULnaKYwl5YsxLzmaLNCleIV0brDaxSxHK25qNFg9pIvAGO8ZzENCRLJd0DL
S2xxitKDIWtG68/AtM6RrKvsFKtVxRFp9btOpWEUN8Xz0eKY64K+S0vlyceAaZ4nmZIXGPR353Tr
oWqo6FuXZhSpfA9pnCzKpCnksqnYOeOmIZB9GoVQ1k9hvpsu/jS5QL1Swni4sky9xOZQCP8d1CD5
DTcCe4NoJSd0CYw7iQilsbTk2ZXe+0Lw88j2Fgr8ALHHIAhjtV1PDVcbRMeApjGa79xiMdaI/z74
+GSSQkJlZiTmTehd5rrD6s8kI52/ST0NMLwmJV1jwq9Fw3V0Pyt6zkHkDRrmFF5c3YITfojPUDTy
c3guATRjT5LghBvNsGcn2FtYwPNtpMKUDtc755KgAla2YOeHO60ojHXEXMMaLyMLi7GmzfBy82CV
5/3T0uP0qz95Nj7VWCOgJo7tDmfhKf6OHG9PV2iRA2WTkOggWwpF/o3iwYFZ1EKyEKGKkBKYyq+Y
5ZZYvou6gD+zoMpELkADn0WEB6hKuv8d+J7jKGygFeFRh2m5UkpbMBCEFmUe0b35newJJ/5y3izm
09xXzhGEOaKYAtAvOKCgSjQUiMTPT+kqqOox2wFmrt8YCFHalyxKXgfXarFqyG9WcUBvsZBhYizc
3hqkTiQARN6qS8wqSMmeWNWYm05WYerWqrlzpF5JvGXx/mjc0/ALhoXxZGxu27md9PhrPgFysxRN
PVN1rpc4ahkPEcvqv6ZzD7Yc7JFPCh8P305KEL07FtiDH2zqOp3ATlTpUYiy3km74dGgNAF1ujcg
mU5CvtZ627Z7qWAOHv2SIcoJ3OUhjj65VDFe3R5x3mLpbxBeXgffzeM0z/9+Tip1zFoYjqK0IbwT
+bqVMOOEroHro/wjWbKuol4pFx7+eEBIXp0p7yEfUdNlR5/TwnzThVQ8PfbOqHd3GBFvBjwvDjS4
fGvmF+CU4QjcJD0O1+ybINtdSXnSaFgkOx90tnvg9DaNAeDO0sKbD0I3v7ImbV7UPDC9By5MiFJJ
OBaxvfuexzKpK4Xs/CaqPuWv8IhztC8CZbReXIqkYdd1DYa+/UjX7GoR/wLnaoYkLWNEIDMjqin3
XFESoiGi32N+P88rj2oXGZvEvFjxue9KrhLLMv+h1lYeNQzfZzBUbUX3TZi7QSgNevHc02M7duHf
tgpYUYFqQwjWdinNimSckZJ0uKzclIIb7xoKO1xzv0XhUnidcFiD5twCOW0HoBs/en8JpA9jybBO
MHjT3C8NtxhACLRrjCpQMQnGXXAlozbo2Pmwk1/l7Fcgs2XPlCm/Ktxdt36YeDjsW1mJADbj0lWr
j91TchIY4pjkum/j/lpkNEgSXsIdpLz8rfPRc0OdPaErbinDbCbYXoykcrfTiJzm5xM/emGBbP/U
9+FlP3+wXs9DiqT76gxwm65KsLoo0HXYdgZIkFjcu/8ISg/5BU9pDlTV996Lg+HG5U56aALV1cfe
aMMa/2tAkFOdq2nGk7wj1VipT75L7DnTlrCQNc7p4HP1xdGYnv+1h6FyPARb20K2hU+qtQ21JHRs
rPuyU3jmw5sX3O1V7HUxi3ObVqNI8vhboVdwHdwyY7VT4GT4b8uX742qXXlgj1MCeX0tl5qZtYn/
yh0w2mKx0T+RxE6a+cAQM0sxmhw34Wwk9MS3IpeRcubBnsuh0KuxCsxURRu2qfd4dST6AJ8wJe+q
XI4lOZkSdWxMq3TUvXe5Unk0Bi5RAf5VZ/jnAO19rB86cQTvp2+YoulJPUXkXR/T3t7acK73R/yc
JZ+PxTebVZbg6oZ2gGyX8gHeyfyk/A80bgHiOQyhQE8mmf2UZB2h3jtY8iAuGILi0lhuDQPhJJjR
aAkEHst1hyzaA2dTHqs91Zg6e064ktytEVm2z4d5wBONNH52Uss5rY2MH3AMMIcVrNJCf/yVta+P
KzBCGDFm3c0IjPWpSXTMdkvTUmjWwBco9DYFUOYmQWbDePtNP0+OhEihRP49DZC4aw9Z1NlmzLmz
2x7FnhZibzbIaWcmvAHUHwEjqCeqnpNJD8Hsh14zPHuuZZn2nrPsI/gTV/kWF+cj5K6pCspyCS4v
NeYPDryuvfxlgon6Aby/DLy93xHkflkrbjOpf+SAjs7sZLDU0P1ASqvdfwLv7Zx9dvLIj3oRiCqf
9pBqRm/xqHJfqKCeYgoMq4G9qPEAhU4sYl6S6CDKub2WyKP+fR6ElR6O6Ysc11S+MmUXUFTG/6Jv
qXFEU2N6iE8p5McDixku9BfZBT+GcNG9RDx1Eh4TuzzwQcGwDINJ+qC8mq0hYL1TmSgLj8x47QTu
tYa0kUNZErnwMU14BeGfMkJ+w6FbeumnO7G6S+S1OABSnPEFrrlnNpdskcNC3MaDWpKzLGl3CwaF
/xtRTn3JSTD7j4PbWnGh88kUqUF52YVRqvLwnHdDwZvUD5S51e5XVdrcJnZVMBXB6VsVWQEwJLZ+
fgP9LqBQkfF3XWO5sIw5hLUO+Cio2Z8lV2+HuXlPUkrROSh3o1KJ1F6grCaN5QiM3T70JVb/nUgO
t3LsrkCTy3RiNauV645UoSSpYrN+3FIaFcwMyLgQirUzfgj18p9hxYCaFAJmYsufemaSRR7TbaDG
e9PqzlLhf6kDIZSn011cTecOC4XQh2QmBMSx5Nv9DzO4v/3vSzaiht8knhcg0XSdVVRM7mPCdsJA
ggtKY8fvRpP9j9epBvMwR03XJ2PeAj5e7QbiN5/nIQDWxHMbZIboz6giAhH0xD53IRIEEkvVEp+P
J94NAISCsG2psJ8btxguZkikVR+7pdh52DCBcbyTH7tfnjElUGgu7bvxFxXni5kouJaMW+OM5fNJ
QczlsbZ5vGtbqYKj9lFsXJkDcWWmMNO+0aJ02YouimU6yfBdHeK43E+ZCetSHAQLJoeJtp6lGycC
Cpswu9aqVw3iOxLFLi8fmmNUUFa8BhuFyRGNM1zcROGGH7QCkZ3YhXbojPwpG2cKpAr8Oc7swrCF
DJ55o91xajGz770ZZUE3TP2mobS7qYPb/0e0KVAiqhsljS7zfGNdk4YRax/ofcXa0yCE0pC3wEAc
Yf0DSfiXhOCAu1HRayJxAlxRn689DlPwkEgMHpZukdr3vqqSmGCV58cHTUBnRPBXSjD17xxtVtoC
BeTQwKHXCgUprWPxtk8rFhUz1muo7CGYwLfmmLfqgg1hNHjJk2yU8noHSPeujCgd98ItKYwD1y4X
bG8Mk3o26+8T0/tSvcfyD7czyKPdak7gJtUE+yNnJ9A10103C5UDhZijY6ZZKIWOoMYRDVnl/G0I
Lz36xHJ5gymo6VdUPZp11coz6ZIxCuyJff+swjqvJ6FLi5noUAAZ+i5d0JM0AX6Ty0Amq82sxevZ
tWQpihVJiVZVH6P1O9jbNB82jifd0V6nSk7fxQj5BaajlY3USxWi00EolzcAZuAwIm2/tGMP4/31
h2UM3HXjEJj9Mb4JsTsO2CAmu2P78kacuSK5gOEg+5tZttaEqgIIWPKdASmyUtN3XIObuke2Faw9
ZEa1RleDesfF7b87XSDz1MfexUE4M3Z2OqxKlO83O9fxLbNk1FsjcKEeNio7i+W2pVigDPwk0gSF
0ZU+i7LjWM8DG20jHg1MNxs6N3COdCNqp/8fe4Nd9NO88/L6G9Y07+/b//dOZpJGmsviDQEf2RQu
Gre9nSt+IDV2duKM3IzyTiuZsYgZvDwciZhi8Z+WrKxVpZ0m2iRPk5HeB6LZDHvpOiW8ZSdD3yfE
kNQQZEvxeeHGK+cYd/DI+ozo/f27PADzxpct2FeTBgZ0Yom2cDimwGQewMex5LuVSVHI1WZOB9vB
NEng3FG/wDYw7LMKQ9tT6Y7Z7AF/jAGlhKiqyPZdJVi7RZqCqn3LgrejZ8Heh/FVKY40jrPt5RMg
7zm4KhJMzmkLhY/NM8oePnM80bvHVtuQdtBV5+8qXKIV5KtomsNEsGL/Y710QCPFWZXb7kG8HFDa
1MDZ3KC/LqWDIsklVmQnoJNZQJNYpBL0FJbXwTAEATJhbgoItf9XXet7UKRMsmQOppXnIMCeKWiy
s24Ud50Rdg1rDIetLhG4/hfB290L5ci0YApy9xsU3slOq1yVT2VZ67vneTJFrm8yRcf4mzW0+/ot
JnVp1lywR3JM6vlqJLJwz+U5xhzbCJ4y3B20qfj7YGjxrwuPF695qSWGrtcYzHJjJWYwNlxa1cfl
XXk0kf2TKEFJkK8wAqo7RJMzTcHoY7vxrg3sgkAfI5ywkK8fkVNKQ4lacPCifZn1yNukA701t+cW
d/pPBP4/MQ335klinzuZEl1VbnaoaIVC9gDzLBKK1CaptXCkKqFyctiPjwGiKCIvsmGilPQPnZ30
C6BAuJJybGSXEBjx275y+iwZKbto+nbiPRJXgy5p0DT+2CZIWYe2yD29nB1O3Um08oFvHQqrsbCg
EH65bhEo09Y/NTJhHF9mFzK1Gqqfe8ExxYptAps6kKppl2g4I/T0mLKDBLsONdTZVfEOeuO3UpM9
UY7F1JZ9FUHdgvYHILnp5fqj+tTIus182fbIzH4XAP9BTqh4l7Gv1+1/XKgIMj8QM0ChlJV29fio
lILyVfprS3hC0Yrn8rUj9+I+O7KbWl3+m39EGD+jI+QMJVop0Do9JTXMKViIJ5LX70cIX94yeFOb
Sd6qLu+2BH3u5E2COD2grqPvNaB2Jgn7KfZAbsDaCwmn0GUMeWp+ZqXMIDBTXmoboW5MwFS1y1o0
Rq6CgcPhFsZHeLnbzLgVj7SZndYjTs0Nru2ntV55YjTDSaM6mU3fmK9dwxXsnxfzQdqZekMe0zJQ
jAnqlm4/fH9OmMHIr4Xc7pyn9EAmGD+W+EBxteh/BhHq1MNaLpqmF5N81OgShM4dV19OYWtz1Yh8
uQtbixyL9kTJPb2Z++k7T1TFpPfJRMOCvWDXrtzogLnbyL0kdwb81z5ITMO2XNUZLUmKXYwDrFj0
fBbqM+Z3gEBkG/ftlCyZvN+kiMlIt89ufbtqHHwZUVH0WDa/ow0rM4ipMJ+kgePO+9n5HIfWO1iF
QqEWFEdhGf3wRD4Eq14VLAcefoKUfzGz+Vbl6cF1H5hNiv6WNe/2TTOwBdcmaMECLQPDbq2bXZWR
0uNluwvz2oksS5CkuK3RyL3HX8P6Uhw6YjCU06OGR61QziBapNTDQOo9U58MxFnDGCi0mkwiKiYS
oqi8amVjY2XDj2O9/hFYf5VVj/P4vFzsCN2bwZWU53Tc3qF5a10kKn2tGFMxEnTUjn3c/ABjeSGq
mEhoh7u3j5PdhgSYl3ossa+s/r9ahVGEHpgD3c06vU6xUqbdwlc5WLVgyo4qhWWAPK9QBp2FuBea
xl4HBdx5pnKEwdf+hrYqQHLGiJz2MhtAuiQUsgFuKLaQfSrRGxAnQPkfYqterUPZGrujbqCxuJ5i
g+dB9Wx7kpv5B8UDGWuOvbPg1XTSMkLXLJF5ZvwebE0tifZYQlJ0DXStl3I0pffCJiZ7pbWRnWkS
3NvpG9uHoWIDEIhWlz3uJ89RkfFK7nr+8l6SVT68WNA74h4VDlHj6opES3LslGkPsu5wCl1kw2rM
PS3qXzqHlIpqRPhU6hiQ/wp25kciuzrNDikwXHgi9AllrLZCgT+UofdJxJl9cKLdOuxR/3scLfOu
puNJXE58FhJOeOLb+Pfa7OIienkYXft3wb0yakCKly/A5y/ONlirgXX35s83kvD99T3N8y+JkJvI
j86glBv/MuJYpB0nT3aNMdKy3LY8zsyO7jX8bb7eTcCpmaJQ8vfqBLdyETLM6rz9nMvDU5zhk/fb
RneulCjuISJcwvbTO0KGIgyiE/QYqXCU6fia2EIyPu9fZ2gSCeW8B/q+gqcNFLX58pLS9HNu3wF3
cIsNiUaoQ/fNNcPvjviK58VXFVy4RcbsHwVeH8PaIW5xbE0GnkBq6mvr2iNuhw3OQlPH6Ii26UCA
l5zykiW34kvToBBwXbp52mYUCV3HTsPlU6v9Hu/kD8pKxWFpQ6tBRsm5dC8lxs1Ytci1sQDGz9Ie
Yd5S6tSKidzWdVRXJ+N7jZbt14mN0TdHmpUXUiwquL+eL5Brf70NnVJosWgVFvAWl8BnNR0Sdh7G
MTDDKiJA3TA/v47SjLH7/29y2NGrwdnqKC/eIoHqh/ja2lmrIBcVPC+3eMVcpsKFDJs7QDxoKIwF
G6pMeabIlfUkDrk6h7vDx5fhwJZJ+PQFz8vq3WL8BW8vftI1Vf9QpPPPA2WzgVhKX4+K9bTaJPf7
vp0qStbrHTf7Th32AG+BSEqFPIh4BR5l3keVBGKQ05BXJaBlBKBojzaJD+B3EocA35/IJ/PhOYmY
PGqs5BSPCr7rHdILgF9aCEmgS9F/CQcvjVUEsDCUaKZlID2rs2906sOZPW4zN/n4w14KgwxvhNGX
mCflHhHIZS6+xH9W/z9W3Sqq2BC4U01SF8i2oD7yyehtsFweSG7Ws9A9XHBnjPIqD+0Z8zs+An1h
eMLjHhhXg38Ft3+rY1oA17yXWXUHLd5XBKmD4cUu/4ZWWAg/z5kqZKgWa1iM3GypZPefv22qSiD8
MYF9Cc3aQxMRbqj4T9EawEBLntpTBdN3zTRQuKOVAAkosXrPTvZFOiSPVgJ6tbkygJQ+oNj+ROnL
PaCnodZQgcURmRBfLRjyftWG3AWqBD4Y0JtIvrKfCQBUZIYjuJkEpdl2wq2fT4MhyGBw3pSgSHje
QS05Y38G6AxHLVsoOXQ8wed41V6Eju9R2w5D0Vj2mk5z1UXddhNmSLD3WsV6bTWU/+9XdH60G6lo
Yw8FVdymQZi0e4LfV2TbS+/4+WUWmEzhtX/csgb13lJgNMkm+rxCoxMnxprLfYlMs5KlGQqCMVjO
vkUVXr+uGL1mxyjhOxPTlanv9LIoN+6nx7uIQGH4b+MZ1K5lxfFgoImzH8jsbLLYviJLTuYdIcLE
6BUcIpQw8mM4x47AWv9oG4x7I3oEVCfTwYhIRSOb6Zd03j2GxgyQiuoB8FR/UQBxCHlqy2Ln18ES
PazoE62norOpS3GR3zCGrTvPTm/dUvr4lm5OnfKMwfzAmGc9U0sEQ8zC6R0tj3CdVVwjuOUbGU6z
iD2J54D7j6bJUqBTzEUdZ/8Th+aeXY8hIBkKt3OiQw7Pcuk2k4chGjARVaGvpcXvDpL/HMny/OqR
avuj8RgddKD8rb3kPexE6VILKlle4Cwcwhp48U4VEtE2HcWKY4d7n8yS6zjmZdMbyg/TfmdPH2/4
h9hXMm8YA62ma6gXgTROJ8d4LfUMVFm/cviNj54luDLfzosdeiZtUtjq5jWinTVK1xs5fSHcW4TM
DhPtUtSFAIhNymFMdJPnBk6O5z/1Q48cZCM0jUfUabICV3lwknhnxGRe99iRTknPxaczFhiTdA5a
y5yocc9P0gRumT2JfXsWZObVxwCNYmhe9o+00iV9LYU48LkARZXXS0wlSP67A2fGcBsuy2lIOWYQ
jxwhoxca1u4mWl4CWkWuqqRQbC7rsbX9j3XFj3NPo/lwVDkStxDMbdmDfXeI4neBMNhDx2CxIv/f
QDLjcZNWb58cyWwC6Oj71IlaDMyFP1saJ7fjam4vbp103wHhhRx9+xDS3J/iHhpQSGedTSRHC0Qj
2BUAABuPzgBVIBb+tzCaBKrhxEg7to3NJJ3pjZ7uVWt4BgauVnuQyEfQmxYT8BhBIMTSg1bDBt6P
7QvxouHTicmiD4tENITmqB+Wx5mEzJziZOzWi2h5mghKGwNcP3aWz7+L91AT0wxpH/wyuvFMM1A+
4Fy+rJZLHUN/PF6d9QV9sFrk/t2u6ZCFgsKXSFT/AWjmsrtn0g0JBoBbgodBfcnxcwbft9SKKSB2
wJgnMLDNE65yB5u78PgovGplEmSNoyNPCz3IzupikyBuCHfdhkLprOgqB2NQlzjhm7o9Onh3K4qR
PUTHdFgvu7Z63QvU1DN8P/LrmINtSg3h/bzbZTB49Wz70CMYS3AkhrqgGB2/rccubQLinPz7+53d
wd71x3b3x6OXAu0uErNn/GAB5AiH7nBCcW9wj3uj4vntBS3pVY+6tVsI9n+gZllRpShWykKklzZZ
uoU1w42NXFwpr55NkvQ2bINQNJZcwNvlw9I+crfpjv9w2EYpW1mZ+na6oKzj9Op13P75iKrAolQQ
+u23biVhkQfFUM6V5nO2YkRCsfUuyO1NqJYTD4Yp4IajAqzrsBnArut7KRgmYNm18Z559x2qVqGE
JN8t9VcXFxrewDBFg80tYgL4GMZJLSW7gX0ZeIkknwLg0XmZ8JmtLln2drWbCPC9uDerJy1Tq2Vy
Qua2nxXnysLZ41yZv2LYQqN7VMsJ17AgNCdbIEaCQ7UZRFYCqu6JMjAKMWbVwWb0HSDV5qp7rXpt
4JUrNi7yGQ0XQ2XrVeccs8r/8CHthIwbU9NFN8HioXT6ykFVU4342ZJY/g4lYevJrEjN7TaeGkm6
Ilg/Qlyetl2ocYWTTQ25HI1r1lDfu6kbcfSvORdPDVv/yVVn0H0GnKArP1wc2WGwCWzRYYu2Js/m
VolRm2sUsRY8/siC9veOxGHdqVJ1m3EtsNRmzVhGsxLS5GThnuqSImRP5zUvnqBcgUXwgQ07q+b9
ZwFko4skyfaPX9eNJQhmbWcWhaqzmUxttvpIsdEfi0c/SWze04avLca8A/3H3ym9sQptNsKJS4pc
BNwvu5AQS1fGqx3R3vmrxs6Mkg0Oi3695uHZWtOWpxpPSP3jerBpzi5cTY+6VUS5EXgK9OOHWCek
ZjaOJ4Xg/Htb5pGTPOzvjS6PAx6p5OQY+FQuejd/CAqFT9X0oRsKIVVy6VfQP+X31LOeH9l9dDYD
89OA72Ny6/8zyYXCgw29md0ItBmyF1xPF6lXsqwqb5WVFt8zugDB4JNGaHUeDYqg1oDfb40W5UkK
z4qQ0f6kQvrFMEDf5+6EX3LvE97vFw3KrrjUaas8kVUNHSWB9ovZSoycB/eAWHGAxgTtNUWE7Oz8
EQ3Oi3gMMZp5TdPw0a5bpdskE8nRIdh4tLeCt4P3tXDxMFo0bM03UfxPlouBTFqdjch8bF3y5Na7
rq0+DYV/BouHTJHGy5e87SLcgBkIYiTX6z/vSJFE4awS7o9oXOcs3M+wSMMXHWenw/SbQkObOF6H
7zZNL2uM2/hkcUPRuTZFob3l5Np9YOgz3vHLZs9FMKQFac396LeskpUulTBZ6MIfPo/3k97YqwX3
3vahn32KrljBeHm9d6BbfYPeuAsOPzvJ+vLODietxXgtIhKFUaA2bMZ8+7FioK0FwBGkzX30Swsr
rinM0cbZh6QOiKxK66Wvk8Me1Kiy5+Nde7HhzwLc5OdQVdGTtp/tC7YG52SBSKByEksMdPeomaPZ
VmJ/Nk2y7r6ZVJwGBC7FjntgaLr1JECrn0iP0xq+GJpWfwMdCHxskTOE0le6Z/lEzJlIThE8CK41
tb9LgHzmJdOlECeP2o7OXodZELw5d3VDEWK2FNbRHPKCepOW4GtbbzXfmU40bTHuXPa0LSiWJEpL
bV3YAv3latyYnfbtwb7fBK3rZrCYQEn9fc3GrlWvTWi/n/zryn8hzbfNLrydZ5jdHvb+80qWXzbn
uBsLGmSBFjhlVUk/N6lWBh4UdexLFoGnjS7agEY7ArqMAiXaghymU628P4iubqsZqv0X8NSxiDjk
v1bYp6k7qy5RloIpt+VpBdWpCy2zj7c0c+l0i+cQUZlSQq7hK+QDsjXwO/PVz/EKzemuEF+eytJF
+cFCQomieodSps5bg16uMlo3653oZGWFdZOO70lXXetFSTQbzOg9NxEFktrB8YHVIN8fgGBXrhnx
iAvVRQ66N7BTfiRSmeQqUpUTEQaQoJ8SAkD0BuSJxSKbvdO6Mp8U6xShrYMxRxjpBkoMGK7afQ6r
NMuY+Qoyn+vok4eqkrY70FHMrqX1nYRTzf+9z83y2u0tsxfnydssgyDpb2NZdPlLBwaFXhHchsHg
IlsSp+9lIfk87kf9n5OSte8gtjmrSEktdiS95mc+U6QxUxnoMNaT+FcPE6iAJsDZxGBqh1oVVq/9
VlxqHV5ELhkvNW281o1HeC7vwS+SZCubKrL4nNU8rNZ8RR3bIPTZyJZpYACZLxHDWF++kG9w56y3
u+sWqPs9537Pv1C7YAy9m+CjDE8OdKXOBPgwjKTN03HBao/Y90HBp0H2EPqAF60bfmKOVEY35e7n
hKtfn5m13DstVmU8Py5x+RrgSp6bSiajrJrSA24rw/TqwtY1RuCOhUROJbZuwLmwMs4dpho7yD+q
zlAT+/PXI2ulBhrk2Wu9rqvWKo2H2WIUZRHZjLu7lVyaOGDE7RIFLFqhuzVNDvOpVprVPIiUnx3Y
qNL8EG78DlPQ6t43qHSJ3R0leaizQ9QMCWZey74N0ElPmAjbxQkF6oDR3fLoeGLwzKVVgCDztElv
e/20VTRc/90tdURrYWWIwI1xsdULWPlaG0k2/L/ZxYJeKqy5/Pheqk4sLBJhCOr0K0pm7KMnl8nT
r+MMmI1Ui7jyhEYe6rTSwzXizt36sibSi5qOVmcXcSzTCbZWlv/YNyYH6cvQcMbeRKqCCdRiOKbN
MnKFLmFEjqPIzMnKm1W0rMAQCm5JVOTzQXXnIoBA5HtD9izI3Q+VpN9Xf04C2Y1GVtw3IWnwblj+
XqLm7mBSlYayIO4JlRd1xI+EvMOxvgdxCfpkvJXTDBbhaTq5XjIHU3dgCsFwGTKtSFdjVNz/12Pc
rtke/6l7HxrNq6UA5MIhNDtIRHMvazl6HOqm9yR74eQGXZli1X7BY1G85OL24yqSvPK1hsnVNg6y
DqmuMO29WjSesGWW3uo4sXjaLQFb7L2E9GsUJCPyHphc7EKXaXWGueTNVDQddHnoXqSenupSXGtl
2pvS9oQH4gNzwsb+uhSKNl9wByvDurWRuXfxY15MVwE5E4/TdBk33cPQc9mKoZec1jHREb1QtUEO
PRwKMUIv/uXIZ3djvLgBAsQNgv2QB6C29kbdgjcudAAA/O3jvHgdBGcpiwo23eSHdYz7ec1dLSMM
All+/vozgxpafSIz+C1rVLW0F/R58CzxCna7FaazdA00R50O4UWIDw9cd6dvvrgASpG3mDA9p03y
219kiJolUHG9FYbUlArL+c6oZY5PQnB6QXsDmAJlbGgAwnLaqrSyjjEQAqqsYUfVTpSB+VtuzOwU
IrlFykHjwI7CJeopzzslXCXvJDkLdLEIXeDxoMJ1dRWdGlQ96WRzgDDAJ2gQEnLLpuqHwz2jWKHX
Uw9/tAsrNpTIvIQERuv1qNnEXCwlheZgiu+j41xiuWy0eDjwCU+BNrSsJKEJFGogfCG9PkyYKql/
T4rE1uVhh3kKekhaeld29ykaKN7rmPwW5vFOpaWBTzLeVdARACRjXYrh47a2R5zckJ65LrArUoJV
43L9LMtcBOluSEQJts7nvpKvQvYumH2KjJKxoJuNe/qDJlSEEzXZROgGhSbkC8Y9tm5EOen5jdkl
IJhw17klHAkhG2r3jYiee9/yUtGLu+IrY41CKMtoRddswicQO+mNWd4y0Do1u6yGzSScrhbjQ1rb
U3Lekvtel4Gs2IqodzNTj6DmFScTLG9pqdb90yBaz9QqjCG5h6fCIzVnRRu4UceSK5yJSxrGX7MR
ZrO8qpzwKOYVMq8aRNXVZmBWLD6/bK5GgqN0kXsZyZ9FASMRwqReuPHaSJVVsuXZAyRyyzQwgNFn
BW/5WvnnEs6NmCVOrLAUCFMyh4zJgcm9w7FKN7c3suwnZoZQjdpeVYj0dF/FMuyONfMKImcQwZTk
6qBPIjYr4ykO+Hr/YlPeJIN7YnbCbslAfm02e8LVpRiotYOClOC+i9xejcWXLa8SUiiUbW8Sv1H4
GSlug/0N76A3kYiy+kx3HMrVSL2TnvWSOhIFHVYPO1ee+lbrj9Tfk9yfh4kIb5L2ND/+sJi0oj+6
MYtj8bTK9SPJ9cAtPpve5lyWcspP5gviakBobjMcoqa6hcpO90V8e0v7lBRS0xr3E6+I3kxgGPIb
lAQKT9O4ntGNV2iFNsF2IVpGBbaL4wS/lf00KFYo7BBqEqkKQIdd9HYX02dA1cMQ8WBHfHeyQgUA
quWKMSB/U7CmqzihyxliFDRy9kCm+mpdp2XsYTwr35t/jUMO8Lj6gHczuKyBA0SvEXtPvVhOY5BO
ZCob3jnZwdCOAZbJCMQePClDqYjkJcJREQR7FTs+fbQWelvOYXZn3IZZDJ2qbHyTCQd92X/WBrNk
mZHwaRkwWGdONQQxyChSp/bqwfoT0xr/fL+7qHX5vxFSm9cjK7Bd6AzLZ6j4jihaw7GG524fW6aN
GkpX59xH1JNKujpzyYLgJvVhEuF8JvyKQyhYnSoD8BSmcptqr/r20kcHK/et5DL9oqfXz4xvif52
V/W+qU6OB2+sjtlJNdb8NivtB6tSDMiPbSff66c4+qgwMWbkEvrDIBkL5dRkqMpmtdw1Rgd0R+H0
j8Ef/9j28KKZXrQ0QFmFmHb960pGu+erIMVRMpMu0BYmy5qImKSm22DdOx4NpnDQgDLaiNx0G/D3
AT2pdSYYamm37pWRJJCX719MuHX1SJx+hKDlCouI0NrmutbIkfP6mijn1b0GrXcTd8gboXmoGRiC
Ue9YJ77ZIQUv9xg/O1VWXn6J9MTu4OiERILX7T38uDB44+gjABQmuu7LWot3yylz9i6RRlNJnNr2
VhMnHOTXiflVAy5KytXtn0m3h87rxZnDcinkxR213WYdyyS9Low3o8cxl7fzDd/umw3wop9jM53i
ui1Bkh5puF4dYxZLh/7Ygyjc3gXD0Zvll8HJl2zDvPrIU1OHaT2eoA055WqxvmQL4Hcu0+4AQKEW
qqL6c2IBin6/Ws6KO1MkSms5MRlO7B2QOi5SvH59gSTW67dyCzAQc3tyDoR/Gy9nNVNNEP51S+mL
yhe8Vw2wWTuFMPrwTEwoqRbyJRe4vqQ1AfzGIIOEEC1zXgopusuUqbiBEullTcDvnH3EfB1KMpzm
Kb4d/VjYrmO9gvyFNFxlWr0UhxXIYcnye4dAUaLGOeF2Jyu0pNHKRjDUTrLKrzRM7BFXJpD40oN1
ISCOSH3ygSvOu1qVQKSkfHq34CaEEUCntOImeEAuP3Jhbex2dSNvaS8Syxob76ILqfrayHHGJbaT
0oP41Wah8Lm0S/K0TzU8XS79erwhmXxKViGi3xJl4lDmc2n54pq4XuGpKe6RCGV4wzIqr09GFm1I
8/DGALHHURF5yLarBPV5rzrvjYzIsiM/siG7rISJHvU9UGWlfpVUH8uuzdFIuXL3wXxNpYej2AeN
QCRkAhQlJ/8jhmtnOyTZq/gKoRNnlWjV9TgyDMjj7jR6alni5Q3i4I3FJbdNhuoHgzOEuqTknyIw
KE0vDXhjwAHvZBDLk/jgZ+uTXv6rgM+tO0tKTrBEu15TyIJor35aCs6GTC++Zugydlq3UO4mK8/G
C5J/ZHNPp0+J3GVJv2N1eIU2Mz7LSo7KsjuJxTDav5ehkkfyBj16E6PCLlQ69+KQBCnXOH2EvI26
bNyBDb3iMTvJ29wCm27UVrQ7vEdfpvmnpb8w4LggXXjDL3YhbIot4X6QW1/H19BzDs2G4ax/R4HO
KdwHxTFULEFxd2ncRex8xdTxUxGWRU9k9U/k5Z+xAE1N6l7LKOfmjhtAhqllVXQeT8rVjTPfcOgR
AwdIfSgyEYnZXbsfA6TUbcmpDfrYWlPxmIa4KX0LDhWNv5HCR2WA8QajplRlCtOUFPhfKFny5GmE
kPkwwdQmGJnyIlC11spP11ob038aUgJAPmDqHikc0lMoUoB4oy26JYiaH5Xr412qhxgF3tU7A+kQ
W5fxXjoT2g4DxXE408tYQ7gAY3g6Xry0IgWJ62hC/SRx1cfvAznefJWKd/Uu0nZOGNbpa+5aSDci
tIoxu2t57cLMJJa9LavSTlHqiVCSmssNMsMhGl5b5u4Fyqm9azCt3+h/oqF9NftL10VbrDGGtCfP
deReH2hgNZbOf5a3cyln2nYNYFeRxsUGftI0wwVrVFqVWYgwAOaiCXdw5YUwymmKK/EsFapMw+6U
ZsRoiZDo8ftBNXwiam30vCKZaRcTwwoqjkhwE99A4AwvlddwPYUe0Ese7owVp7VJ/BjXmi/LWXIf
EafYoDkkzSZxUNqo4LSoZya+VT/XtMHtdHJArMWzt9u8fZ/ATDJ/Ap0FJpsgzjuZbHXsuhNhaGWS
5Yfah4gxPKuJrJcpFMBlaOSutZdVqorAfLOiMIKILitvm3uSv1NNFN6M9wyZmR2s4ejuuPawTjqm
LIRTvBNwAj+s7BYiOViHH24aXKToMmv97eRJ5W2M/K/irxhMyy3WhIjQS2NHTVpwDMTOLj5W21Gl
5vvDZEHCO+sekBeVXgovIllnUQk+saIrxUnNEJ69H3F/Qp5i+WsWngyTl9py1mGub4IJyNTf80vE
OeiEZ6pfukQNItPbIknpzaLACf3eq7HxWJAc5xuvuhjnA3iycWtM8qa759JS1al9l0yXb1FgV7Bp
OS2XoJjrP6a6pyc4jTu55RDdbi9Iq2gtL5h3rpaOunqepQooTuGh9e+N6Ak8US3aJoPdrzESBpLl
SuvrabdIqt0Sa1kYJj9cvNva3B/CYwqPF2YthgoNGGHCzyj2kUyDc6fIDBifM+Vp2P2jl7PwxtH+
aGq89KUzQSpakAMVYF4mNzpiAp1ZAvYVN1t/TRqmYKDNRFMXMumytXyU01MI5kgSG3vKYfQkdmwY
YvSPcWlh+3YCDOuNWvX4/IqTQrDrS7cP4e66WG0z2L1bxPgdZln5Xkgozfdn8ewHI9mWtjntyC05
yhHBf6Llpp5kmRey+wQXjm7QL41ITrzIrF45lhLYNyKmvJmukR7lc+lPKruuPGVJGNEK6Bk6x+rh
864vQZgACXXDxY6bwZCO+TJL4Z+9CbSO6I/RP+80jv0rhVArkk26ChPFGB7oBz2erwHLo3+4ifhY
vH0oymAEE7UfzK/Nf9owtSAwpxZHxUwdNf3ld2i1YNuE8MKIqq56ADvnuwL3eY5LAsZx0cgbsN+E
vBXARybgv2J399CNtQjHfDpRYEZv+sLjJVvG33IVk/vZW9V5cOJujp62Drysae/lXikStiEZLAMe
lKqgzQng9+ihhPwEQqnB1MC43RvAfW6n8fDDeKVTYvUg7PJxzQ1MegkatXvoA8qkEUqUzECIYpzl
wgsknnBYLChOAhoQeYGXnQVbrgWwVz2iODyMe2dmr7+hthtz6Upq5m8ucTtFNmDTmeHLjO34JdAk
zXdlJ0ZI5PwFZx/dG7zjynYe87C89beFJAGohD4egEWOI+mRufBA7TA00hwe7y23/nb7DES2Qwgt
c2Spbq7JdeGX/iQuxSBsiVD1hEM3zuWSGCVeqPqycFUIxgvoCGTFYfODhu+SRP/FbkszzVpdMG9b
H5UE1BjcfH8GuL6b+w8CPc/uzXaPWUgK3pCKzI67fn5mYmhwfcgEYc872Bfjurfl9vo5rpIja7/1
dJFBwn9c0KDJ19Wk+YsI6jaLhk3f2Vn6G2r7ku8CTKDUHTIp7sjpgZl66+05vZH7jwfrmU13P/jq
jpgN2/cBYtqi4XbK52Cl+9xN7F7W+iAUQ9QVd3Bi9l+kqucVpOlDwLWHY+UDLJnXh3/9GWXCjwFD
oRPNDjQRqJXIOC0natdc/awIw+CVfmk3cpTPZNXmgf3AhAOzDC0Scpb50RqlDyC7Ni4MSlO9dw1v
yt5AI5wuUMbVtcSNVfp5xkiLiW1UdvfBqRfEEafA+Yc7CnH3pZwrGLIeJ0/Q1il0538p1ojlWODu
azVHw2SxOT/Uctw2oAkjx5+URfxKsVP7uhh+wzwsCgGNBBb9IMWA9s+l1fxwUh0rq39SolASs5SN
rjtHkRhxdTn5YqrsvLQNGQ51dyzzLBPav/1+ovwTIil0cwZDP8nhmc6GN+M4gAw4kYhnZJyp3ohn
SV9M/ilontVa8kthorNQiuSUySZD9GCqZCvuHpfeOWCI7yzYjCsr+hLX9H600SadSN9QQhx0JdIZ
xW2c+fDNGV0NsbpxDe5xcpOZf1+5siVIGqKSp90QWTAN7jVWwqD9pTPWSthQqQ8NF4Mcyl9VE/wM
6fekRkGvJX4Kr2IKuj0nvRJ4wCGVTedshgiPAqBHIsP3bJIIe+z3gNZTdAfrt4h84t+sPxNLrw05
fC8dNUsJdid0y7qbcO2OIUDlL72BzV7JU13fTCowBYkfpU6YCbd4LjSnDjZetqUBQfiCnf/WbuYM
yrBvWJCJ16MivhUVBPCY97DPkb3RnYdAVVPkX2RYX/hD9IwC81u5Ho/zGc+TeKTCU6vQ5T3wNPsm
+9eM3sQK+tCWWExxZo/pY+PNIrKyC7VMex/vcjElP/qv3oFvc7xcC5RnzgUsvItQBTz1muJJ2J3M
x2v+6OxhH1pA8IwmSuzpdQ6+NzUYOgCtjlcH4a7vMmY5Z9JrbuTDcLqNjAtqX8dFKX2yJZ4cfJgv
WVuVADFV9oI2N5651pdayDqMx5mHOxYig4fZxMwsIIaQEiYSHuF5ZSRFQ337nPwmtJoHlJIS0b3R
sQU9iGypJJYng7J5rHLfItNMwl9OZCQza3jPDyFy6gvPwxomBEBJJmTrXYoEk4yo8AKq18CO32Ia
EQIjhsT0BREsl0ZQ0Fv7qMo611nJ1FQ+3zfI080wOl/y5RWc/HzBuebnHQprjUiZWrdZJSDV4alc
XGalE920mDGMzVSInqFJPpKQaLG2sTc18Gl9SO78//fiaUzr1WZRNCJ5aC5jnB6R3p3od8nt0c71
xcfpKwowbNmCg7Rn8eGr7nhDKh/X2AwaR9bX33dhkiy1aaUxh2H+R9/CVWNapuuLxRYAJRdacj/7
ZdXSdhk8Snq1bRsGNvm2+y3j+abphyjmLteWlNmPgwGK3QGULCqtV7SPE5ZFS6yTZFzdPlkiY9LW
vIuLuftV28wh/FlEwh4VLfps4s1RstZLK1SdRM/uA8xIQf8uC3RxitWNuXsAfVvSvz/NCY5mYQMg
4IQVZ1YRE9JD9brH5u1itFb6R8x93/T4w5bbmp/udUiqSnvGf2oA/jzm1pCC5QjbEkO7nYADTEJo
NpgSUg/eNkPnZO3912oYmpkd0cYQ4RLeWAVtgkpYvSnTEKt1a65SopijVoLVRLztpp3UZg1wjscM
dib6glkxi6otuTdmWURiiiXh/fODX0nV/4qb3qRw/MFz8gPIxdeoP5QCMpH25JJWxt2+1Fej4Cvp
5lUpobaxCafSWss60wPNgIIL7xLew+glwyLleIqWzZ0b1frj9jMJFxOEB3CTMTjkAaMpjhcMGrJC
R6fBAyEUx00Dlcngsj+nq+hvfwkwmktjpSm1Fy7fUGkIl99zrNpEG3QUIL0WP7Wgs8eU4ICxtKr3
3Ji5Aba7JKYAlzCAoCGnX2ednVunXvBDy5FpovrvNBdCbU1VPPRXqmecsE023JnNiw7tNMFCg9o0
0BvxbrpKbp8G6G8r4jT4s1N5DE/AWElQ3gGTg7b95ZFYz9BzbdSQGIQZALy+MGJSDE8sGFcuzuoe
zdpx6Y8UiPCcMe4dO3NXJ4pJt3h5HVYsl5PHbiNPJufGRHKe62yysoHzSxo27uTbm3pqCGgbcNs2
DEWz8tSN9h3D5KvaO2Dj7UD62J+HtecRfravWS16BvL3BEUKWvWk+FAcsznaT2imTi7UzyV2dPm+
7wYY8PVJTuK+JGOLIOjXUIjiCzhuAidZDVM198curBOuaEBS9UyaCDn2BZjnRptBM3MJKXsdRqBm
O/Q7sk5Cniuj9sF8lmE/qJrnLYc1io9vecbKaoOVkk5Olt6EzvKt4hbmqeeOQjGRtHb0n9KbHlNM
IDHw08RxDEFwTG9aXJbhIwLyROt90ZSL67TCx45lTVUogdzWicWxhU5a8eak68gyhR8eIZHECgVd
V75k96J4giNtE5RpXuulC3EZQSEKd/KFxsmxoqXVRtqh5zGbpTaVwFSS7QgDhnMitmBK3iixc5kL
71hJ+j4Q5rSCwT2PM0vLl4iADiN8XVPkA9R/yEemdBMg4rzTdg8V92rzGwzVYSbHJBENKxY003Ur
JE1nkoPRs+WrwQAwfSBeEXF7pSzCmznH+qkIXkYbAkdsa+K6CIJHIgFDIgADDkLJCaiZm6TZNV0Z
UkHYWOqUme127+SoY8yPPN1MegUiv3peuYhgtyE7CnT/XRI2GLs+y1LaOGIP64XE+XtIvBUGrknQ
35lNrdmKhXvSmrMtHRocvMpLvSeAaZYptqCYEXUyMzvK+ipa765RwVaZOlU37gO45tgsgFmxPMzn
5HSasrEgNC/3mXM6E23nppAu3jVKLS9uZqTC6uON5g4aeNgM6/+nKFig+Jr37L/8bofeST6bjvkq
J6hxee3j1kGZ1RGnI4wRtuUvEdhwm2x5o/1BM3uA79PEPGgwelxWqOcoD7t5ZTO5Tw4ZW5VSr4fw
aqmnaRl1WWuNEKkkgBNSXsY40o3viQgu4DlN9C8KrHcx7V5gUvgOb1qztMRvDevcwlDTpKsrUn2N
1jw+Bn6F3PF/bmgHTLYr+RbUxvk824wSkFg2/nY6SteU9pQwvGqSXi7i5TRDWL0Z0zH3JUCoaxHT
Hw2pc+vwpg1Rdwx1aI5UnAlpXAnyjIngTuWLokCUr3JgU7Fq/OZWCLkuc1B9mQ645Ks3kj8CSNFQ
svwdGJ0rCo+DIGXiZ1siWBSpCHnqNbF+Xj4UUp6tceKCGipf6fBCBd/tegZoqJ5mC1g0zQrR3aKk
jOo9LHWcyBIWxUMVJ9MPD5NyP5a4LFWAQnu/YfCoPeUBCPigj3Nw8VdGq4mOccrSyVL9soEv8bWZ
xM5yF4udyUUkGU/7lkXj9W5mP7kt/+YPUyyLTP17FtPMLJmdfiQg7eecZ9Gsq/Mb3h+vqBufpho9
wGtNkkyDTVwU3OEeG9bKiqAe5nTd2ia1M7CPo487Wl8u9riIN8gai2MD/vNuqEbhlNl7cJeuK07p
rk0nBPsIbeV+a1CM0U9WR7765nXEbH9kf8OiMmJpefQ7Z1IxgSE39xOtIFmKP4nVySTgNiIe/tqK
T/IZjpinG90zzNvp1zmKlJB3gMaHCTHBRLntnlSeiwPDlrJxKnNyUxFau9UV72XrGgRwVL40PxEz
hkaoJtUVO7E1GT+t4s4YE0iU0PuykXYf7PdBZQMEYAL3v9Jnd0LnoGecS/KRGIwo1LLmgOTR36TD
8b25VMDsfoAGZws/QnwDCrWechLtOVaV6HVt5QhW/fW03y9CJc6pLRpZM7TBOPkYXif1aJ8L8P8W
b/DTF9UH3xx4+XKt4RoSP7m1JVBC2fgbBP8TVSW4m0KUujwImh8HO+fi9fy5YtdZWTn8tVtsuMKT
mY4gi8Jc20VopJXmj+zNM2BExVbMf1MhpeB0/4Ba0zkdzl5qS9B9solEeOEGL/1DLyL46W8TI+vo
E0KZYDj5UVyklRRxk6S3jaQPMulgANqjucN7ImouUi639w6DaXkqd/qMuvoJdel0YXSUWoSjujse
zonSOtK2+Ui7sQjgYsNhftF3uxaZT4WpT6nUoepR3TinupshrGKhYOr63SmfEfX7omjMpEA034L5
dPNTceEKOlBOzQnqhOBrabJJ4ZtvzT1qV2rgQiWkNnnBjXwpOG6rjZzuzUHtUebvvDhpfop3SHT4
fhj6QoP/TisgXz5d0N0evkFJgS5xef/UHwxjcv7RXhjcQEaXnsKL+O3Lq+8/kArdoRiA8OqcDksd
8HpN3ELmwbI8AVvg+XAdlPfNEgMVW1ieB7K1uU+tXcwlz1NL6RPf8kFH+DA5YfN8lgHGVfoA/LCn
+7lY5fFpn0P1T4ikh6ZFoc2tqakNLDzWtS8H1zkz6Zrrx9q0CFUxXZHP7hHFPd5UK+vlsOAURc8W
HK42c7syj+HztC0Skp9CYuBzpmUf0KUAdVU2Nooj493WEZQghS7o/9IN+/1fIZuOp+2QSgyoWhTs
W2EZNjfNGrrYN7VuwCxNr1IeBE13hjm+aIgGYQpmWwd/1yEhKyJl3ANA4QHW4ggyy02ptV1IzJhJ
wremr1Vy6IyTGYeYeraHLX5+pAFntMCloSVBNNSEX0lSfFNkGnndiOa2PZC8a3Y1i+WnvW3BzMKj
YroFsH25LhMesFpp71hlSx6nEZAJsi6zn1UGH01+lqb3yuTPYc1qNMssybWFHTIrzk54AUKThE1o
0aTNO5sHUu+Zn6m2C7LWoxMC3Ehs2miIfuydZFOcEKOo0DTTBb+WGxd+chUuXa+BbEKzdbyKE3RD
fVGruiGTqm9c+VkkrrZqySA4dIjCc4+pGTKPecBK2j/5fG7hAYytNnKlLr6j+ZGwhpUO2rHkLov2
+b3yZ3rHRzdfSIfMezPIFPMOL2u8BUyKtXftZKWPunDeWe5zw9cegrotazs/jOufKS3GOo4QbPQh
0eIp7Uq178gGTw1z6BSMKsmwdPw7C04r6Njzc+zhuvnHtS3YUR6mWZYwUlN/FRtE97hoNt0FV+0X
dRCuHVsaXtJglAcohspEIWd6ZF+4RZcXXe6tTuWiWi4KJ91GXZU0D5bCZlKiXXgdslw+DGwNNq/G
GvC+XNgFI2nBSXI8gZbMEf/K+3GiK0hvIca/AxlsU/xDr59jEF8rh87ZXd6dJ+KWhb8+pDc9ZZpK
kOmX4Dvg9+gXPzl88yxtyezBru+0OxeIyvpxwvCWM/oBj++QYMhIQVBWHj1H/SgW7sm6lxMxDzTZ
w1yUO2bjM0qs+uwkK07oyXHV1lLiKH/aarTYGa6mohFEuKnYfY5fKBN4j2pzfDhBVl5SuJvH7FLM
2kjAicnEMa+x559jZuEwF25wdkI6kjhPPqKy6I6lCwcCXUS6e0k14r32MDaWCzRnURy9KnHviQqk
KZhA/aDGq+ejWvvL9J6SkL8ox5WFtH7u3HaNC87fg8kqBIryLl9IeouF5WX+jDjYUZoTINg8Gslp
v2IXZFfH2PCIyhsnqechkVS66IQrFHYvy+zcRWnVqooQSnnKNzr7WiVafQRj8XTeS9Ae0do2ZyW8
San3YNXuyoMMRDP940luY4hH4IID6tF3LV0ubaSsLuwJgPafTuMikCwOA6Mx4V+L1Wd9CIKtiTt5
Etx/HakXg2Aqtw2uEf8yCBwXl3s9nGyQemdNx3fLvif1eJ7L/nXRiSlzuJ+Jj9LrQEbQ+2EIQP9Z
PXo9oh2xRldxv0hLzDjcIh3lNWCNSsHczGlR1Hfa3Fr0a0GARTbdi3lIH4XLWff+9JDXwYvV04lm
mJswb3d/uRl8kyVTN+iO/Q/fw8Zd7OEozDXlsfjoVAvXNF9hOI0pc7kJmEWyaE+CthwP9REJ0ZIv
Ak6/y0eStFbLtCzTHAR/sRv26BC9ZA07u44tzQ0QrDDu+nHKVuItqX2UVA3NvPf2J9Al1YJ6LpEa
PLqTO/9+BsmeLAJ5dE+v82ef7S2NkKeOFP4dFFsR3wLiSTKbMGegfvCNgucPt+OPgGhHz2Yeq25e
Qrq93DWxovU+wo1hr2IJI3VcXVYUHnsfs+LNSrIR+7geW+TvH2zXZREwIsFVs3lxjw+Vg2l/u6Ti
R0TD40qBNoxOi2NmAGVNzRpcR57CLwqkifno4hnjrYlJraVRcZNBRXIOkI9dHr/E2WBI4kqxiWVN
fbLR94VjlVbBAIVriOPQiYTOCgDH92edty4E5K74Ueuc3C5M0w1cD+A+9+b6Ok9RgSipyZ9AyV1s
0zVmOSaotxDNO9Mcsirrr09H208zUP3PlFrhDTlZQnVt66Vh5/vvsKBDN3ZRrWwu0V4x2bhwl097
dzMSHSAep4Xf3aYJRGGRihAg0wSKRzjNG24kvydk7eMP0GWUxPjPoDcANOQM2bEdY0PHiXXfmpYv
CrJ/nuKTmI7xcmXjJyQlimx3t2urE6rwwHuw14CQ37nJuGxupV9EuLkFDsDNZgjDLXcyGTu7EI1l
QxpZ88iFlA6yj7YM5DIlSEFplx4k0GQAIaY5UAHtlW8giVJjlGIYEdMVkVJoONGuSAXRRhojrxx0
qOWnjErPYWyiGsG78mbodMuMw4SfvQCrT1QW4vM7/IzPMzx2a/F65ItITNMFJ/8un9MF+3knMtN8
6lRLsKjlv8NDzK4PzCdOsMrVUjpxO4TkdSdwGQqz/FmTyee8EgXanhqLcVDmNxQANn4lJsdv2BW0
JuUu6soU7tvHaHcL3IdE2qvwOegJTjx+WmxpgTXpelOEGqPwcPOWE8mzz6hUHfr64e9MPcLjWAH4
vwzr5HHMLxnxBbQJAc4aWSnFVWJiLojVLHI4xOZn4FET/OL+AAcgxwjUFJEqe2WzZIKDjBxfdZQa
fiVYIsWh/pmxIFZLu3IL/um+2z/pdxAJnTk/sixczu7RBMPjzWn2TEpi7cC4zT2aC9muFZ7PZH2S
qp9gk+HLHuql0JPn2LFo0WkizTlLsjSIWlLFHM06eTtnN9AYsnM+rwwrRC7coprFcYQvJAk4IC+f
NweyH7lfxzo1w4s5i4mRY/peMEL03J9kgpcq6l/WzGcSqFDGsm6dr/eKU2GDGPoNgAEWv/TQg8lD
JzkmVBB3BT6gCfYqyJP4cg6rs0zQQ5dPm2D03Apf0FYFA5Pjn6ZKdCED9IzgmIrzM17JZDUoTZ3g
gZcCEp7HOlrzMlb0x2/eqrxzDR2dKd48jXl7O+3vGn/gz54TP5lie9X59MINPYDKUW3zP6c/tlPQ
wcct6bCoAdB6oNLUCQhBJyNRCqRbGeKLWKUc71bESKHaaZcYCb+at1vvcSvhnLm87BEDPTUQW3t0
FNZlItJYQpGQlJbta8YyIUlQebZUQrZuizklVMH6jN9SEiEnDh6BIi1yhiXQO7vnxSCWH53BTlIC
5Onf+I6Tdx0rJzitCAFt2oCcsaj5XVYLUZjSWLEl930aKjgvj8m+JL5440CfgZZv3CHB4KaggTCs
z6MIYi3/N/6rETraQBJT4U2HEtJeEgMoLwh7VckYscZx9BNd93PVQ4v4+i36lRFjbDN7952fEamU
1iqosJPCQCNkBzAqcH2aQkOAJT1fdI83F8yMczYxOXGmKfDcF5cJWrgzce6wboalHDifZMS/Upen
X48P81ShIp7OlibaSm6OnFpAbzwB8ILkDL/AviPZvmcQQ5zXeOeQWLy4wrkFTgmQrs3kglfnqozD
zQc5cHjvvEPYaUirR4o9QaoM//Fhx/ZGPEf/jwSl8OYu/cArWgRwRIHudS6JeVNcod/aE1KIxiEh
BneY5hAjyeRpqLpsZvQngQZ592YOvPOnafLawVNj8Jnv+80ddi9jZwIKqx4z/0eXFtspve/6oHQ+
gHUwW1qiw7a8bso8Z46otrjGDdAsjuPJnIfnioXTQYQAFPIfER/I59M/XQ7z46MAsSqMK3PT/eB4
0L8oZQY/hrHp3pxUImYuP6zwJn6nkHWk+ZXk8vsSNlrLL77qv65jaVeie/KGkUSCTe8x9nR1jynR
PDPPKMWYzLkmGsHCngUbelKpCz4o+ruqfC2oMPFhIgo01HeVk3e84bOYBpMUwN43l0AdIqUUljUP
0YGvCNgz9zSPn2f1VN82QPXbgGM2m1ZKDI7Sq2aHvNxtn59n0e8p9UC8dS/5+mj9PrkHqGqFk4no
a3E3LqOpzAX5EqRPj66yGg51BpQwas3GH45ew4BKr4Sd4URT7YURKzihva/w9jYA8bT5ihom3lYb
9XdbPJPQ3IXWOYUGugy6R6JGCDmr1eadiOB6TYKHxGHDxEd8Xz0GBsKxhMN0fpa49OmqESZuQJmX
VgvA7Mt0vmbdWq5C1C9/avp8/NocPgdAlaZPNExtmH1JSeQkNvC1J/w/Y19EWq8EJKrONb0HmWc6
zWkSHqKKRhb97/jQqp4jGDXJ7Y2Y+VgIYbHB5dmeJhIHz38lxNxulfw82IiFWXwG5vfFx10nk8Qu
DAsj4e1FUGf28fKMOoODYo0+LnwdAsTJJqlotfY7amLoKO8WcG4OvhKPTxngqEj26iP9UXF8+fyH
hTHiNvTex4sSQ4jgEWi6LeEnr8ZpXwyJFaMZbe7L7q0B212w1TbiTGgzzdly5pCxzGKogiIp8X8Z
R1mlc6X9pNMsQX5jbp5aq8enrkN89icKDbdPGSJoo7i7M2BfarKr8Fs/gMO/zuRQivj/W6lcHh+M
zVznEwqPm3xz1qQWZnMWEtKBa8gK4hJscNt3jcs7f6YAPkoivX17zmmkoFkFCP/i8wV8Vofs5GXt
h4oMv0Tyyfci5ZVKlx4nJkJM1snwwAXWXwK5qtuAOmqQBqVDIOHX9NEretZpVtMKQy5WKyRR/WpC
gKpyhbOmRRiV92vO5jljjvJsAjIGj29jOHN38BEQKkR3HRBxBzQp7zRCWOREjAYFHCYN7mM+EO7j
/f09rymhA/azIlswRCxtFSxtn5zBYzQEukRl3sxQiwGzCZN/kQFaDzrfPKEdYOlvoYElrtNgRj5T
oRCTCO3upAX6zAPVuETVX7bKgiLCwJfD2CNeRozaahWBx61uACvBjwNWgsyRoaZFBhGXxM3MYb38
HQqUrK876QgjAAJP5lbEOU92Q8cNXFKV78UNo82Nrqm8bpdFg/qILauX5oUwacds3osoQ7bpRyOu
f1XdHMRFXkXYhftGfyO1LNClxLDCQn7GmZNB8trDm8dr7llNhwGn5dBtGMRePfXvjtKxXsYH3uJN
LYEue0tdRod9OyLRG1W/M11Kk5Ii60nXXFyS1YLjab6qXzDeycCOTJd5ewFzEbCJgmUe/mpClIel
YnCcR8cSKXPbAU2HSzS9nT2yhv6huZ9c8BTcD/xT4T/UjYhknIEL94Dwe+uLrWhHgyyzADbJ5DjP
OaN6c/tWdR8j+PITMGFFdwDSDgTmPuo1uw3M1gPg43rWq7jgM03IWcKyXHvuAou96R3o0FbL0Ag6
HJgQ9VYZO7V7pu5Cpv/gHNIvLAlYNYdEqYkvSGv4p54maPfOZk6lNFx1fjYJ5X1/OYTxkeTjR2fg
vqMmUUYjTySPboAZR2J8NYj+9BhpCqZNHeNb0mK6VDsnJMJ8gNSxmEBf2cPEhcdPh5BlCQlh7DkE
qqVV2CEIBHbVJ8ncQfMzqtn3iUYIonE2rIgeTFtvMh54xGW7zRN/X6BqKMZ9/dSh80WLz4YFfatY
cqau7N6IaepS8itvXkRx+qoZNd76cLNyqcxmeK+s991VWCXhVqzUEgq29FfozCLjVgWrjgywYsFc
Jvf6L8sozMlgXV1BelnKTsVSRixkXXQwSXPyfQvHRmf3hLoCG+ue9PRIN0kKevY9zFF2XglJW95s
TaNWrKvMyESA5TyaWEs8dZS1ImTb+fb5AstND9EpNCpWRrGySvVVvegqKiDeS+z7L8U1jOcZvmYG
txpzPqBzIn9G8zki4f5+nZqOpkn5cDttpnk1Mm9N9W3ksUc+fV542zSAd1cAwsANTezi4m0LSGRL
tpAKUp1lzFzjagee5udNpvkuuCNdNfwzrpxo1sENxOFxmYdUVkceJ1S1Edb/Pwfa0QYjg7YZA1SP
L6jvqm8qLUq9lh9oAbJGkk25bqzid2oiiufEaDJQ5b47dIL7D2IkdWIyBfYHtPCofRpJ82C20bON
mEaqU2tF3P+oswfsTi5DAo9VKNd9VSMh9YlOhBNubbHu8P2T3doCWhjPxzMyClsEY12pwZoZL2mz
BFymSNp3GhIrDuL6RG3+ZygYDYJm0fDgHzw8s0ro5N9X/tZVsqW9gesXSUdWJGGLN6HqpvQUkYxE
no5ogubpoRCdldF2a53nuMTE3R0yQOwmlQoPiErCyleSZCgfiwFZsVmiTnHV1H+NCaEL+9Dbs/9M
oMitdqIblDNwVVoIvgsNQwi0oU5YEIbcIfRElNC1+ZOrUGJb4UHAWMB1z4E8XvLSXULkSUFsCpOr
z8gv+/rXuTB9j2eRzeeiG07Axn0MVcNqdsYE0SJJ2Gj5GNSHqPqQFUrRcLo/BvsFdcTjuCE1hUFS
axv2B12Nt16rj/mrdgWzpi96X/976cdvB53gH+UDS/BVLHmd59zSJJxE65cDnJ9qW7mV8anYU9mQ
xaOJgcD5jAVL7uVXfdrUdbeG4/Or85OyBHPOp74XakK5NSjRIeSmadrEvgC08SpiK38GqkFIEL/V
FLn5CaR1gQ49aA5mhlIg8XNDyydsErLa6AmN+5Iu9N7OEepSNelMXW9sSZDGWUsdGVmVkUnIwNrr
GeWyZ+Gz9yDzw/kMzckBpr75O8kdoXjT8e66cJyesYMa5fzJ6zp4Y0Mnwiqc/crEPU0XTY/5LxJn
Iv6QmZMKZQHtyEuYUwLI2EkKyqag0fOGaO0gD3oYG9mLfyY2npvW+F4B0AQ9J2IH2/Z8Tj4loHFw
QaeUNbMISGS0FZbu2Z8xBNBiCVyoqRUK3DmiVX6JJv3zk2q8lt1+nSoz7X5D7FKElLpaNNO4hXD3
r65RgBcVVYcAKBNbtBh8I+0qzDGHGjMACKTQaPuia/WrjKY25NELa91XalRgkOuKOYMvaVVohfqX
lDtx5/N3JsZLTPwZu7rMXOf/iUQ8hjzAfJ64cA6A2+IBfvp0HQoYtfomsmeGh3rzCaQS9xJHZfya
fbv1EJZdT7anD8lqEvDJSgy3FHXw3JtD8FztuGThLKTOFptGIN0P3c0JkMkInYtBG2KVWLy96MUa
ve17Q6lbmKh0JNUzlANT6uO0fIR2NUIYNGUd1MKg+VmytUhMPshOWDvAdTSuPmAckokhZwiAYZwR
Ae6JxFwtN8sce2vJ2RREoXE3z3gCwNN3WL3OzV2AAPm3cZLTb8/pOxyZqfEQ8b3ZbQyuz2ikWutf
AT9GrXC4iyszAe4Y450suOOHt+gT3/huSpqBuXtAq/bqTlSQu/x5gZGu4bo+zxgkX89byIKu3aqu
bBI2uhICu3mpvbD5BZFUr2QFUF8LK6wTErgV7eEWni69xe5ed+CqMEJx1MUWIhAjDUoRADeUmJRD
CfgLYDV+dzUhmB8GWJon3YFSCNY6BhrRN7MgWlutIETShxc2Oi2ukz3JPn3jxhFLJDio8kMPcXmm
Ep0K+PGLEsCFC7KDmDBHuCcOdCMBVZJkhybRsP5qCRZxRRPTIc3yIUAl2lAuVkFmqlLKTDaqeQaJ
xetiSLzoTxOr77ZpIBMRLbih0mBhZ8ILC+QEMaDMakQ5W46y3BZULSpU+7uk9z49+6j6KV/Fo4xk
iV6CBQh59T/RiL7aJzrraU4M9zlC7k8zWjlFcCyLxuWkHcYytjsbtwMdCsYpqEN8251GzATq1Adp
z9zylE2cFj5MwJFjmlAxcEoymEAVoUf7eXP1rAkim1hP5FBE2QjmHIa7Z8Frz17Flg7pQ3Kel9H0
K7iIo5Cmj/0xAOueVnzENuEjMNL/62PuthYTh+QKz2mGDFb4VuVqjzWmr/4z1zBrQErqbva36//W
2VAmGkIh3TeGRTvqCFXZSAynEEagRP3/ZVbqCQ1V1ZLb6n+eirK/YUwgteyi3jgbeShFVq2WwUfk
9V+IBZ2WF1MkAw1+ROiEpbNIWeaKeYhrrO5csEAU6pm653knLE58sBvwWOyfq9CY18d3Q3zrE8Du
749E/YoLBIWnzK3r4YPH08JqDa7Y7QtMZyOaD2t3JSD/3olUj9r9GorIyfgiCeqxdEFaalNpjdkN
5py6GXIJpvR9I/ORucWSppnWwwrpyHOKc+6DCjsIAi9x5uQs5zG0Naz0M0JWxx6HpHupwzb/P30n
Uj8p0ER6KK2QGCqAGbjyKEqK/wjB6Ot8rvAKa9iO2oaGzsdrMZHJJwIDqR/YHtuf2D2E2LctEHkq
+P2YOtw6QqFvjZVXHw3C9tSb3Yrxyw0Da5EVHzQYnGGXU/thEQtmZ0Ak0uF1h1/tZF/r5bltxHFD
CzD5lnTWwDr0KAFPt/YdT+VmoqJro7G843Ymy8+dWotDL/jN+o5M84dNng7tGlMxPaPez0smmp7G
md5rYrNYtpk2rLj3HldrJq2+5B+AkVLi9j1g0+9beRdAxCG8prBcjvyYmi+6qsjSEZ1rIkqHKJlI
CFI4lAwmC8P3VXj08pEjruDnAQUqCxkwooqbOL9M58SQ9xdSOMOsZUMVUxUP8aGH2fFoNSW7lP3d
g4+rHauQje/luWVrxCtAzdyiSfdnqir4wHJsDvIVCHX5RVLjAgidJQa8r+1C6N7qU9c/jhTs6jfc
oyJz06VhuX7/2L8YRWedGbcrXEVgHDITfe+G8hCDe/h/xss+kP5Ak9XkOfKrU0iVXaUvdQj8bVbJ
J9JmF9KEu97oFFFGOeU7mU4vZGyTAg0nxw/v0jow2FfgrRNuZRIQTvwJZzN0IPLsCa42RN4H36vb
tISsu/dfBk9fy4iAn/EmSplV0Gn554LuMEttvFNkCzz+d5PjouVbx6DwUfCU6InZkhBisIf2sZ/j
ZlWPrCaEkRrPZODzFrzGp0PhPhwMDkECbm+/7D1ZtAIz3VQw44QJxx9tHQCPgnaax6Lb7PeogZ45
2HijdFscsjCdLcAjFcyW0I7b6/gkvU4I38MY5K+m59regr7ltxQCK1nsm8EZuCE2J/itzqz3hpQx
KnnvbW5I4OAYzZ8biafPXavSQpbR7kV71XVhvTpjMh62t4HehUXYQTH42dg37Z5ymiVDuh+lDamF
2VkbfXnXLLu9iueMkVQYzwnS9pFMUvAST8b932IwK3qmxfvOz7uUPxgUyvOAKURN3wdg7neYRZ8z
6qOUqt7MtCAo+GmB2cbsYuuyw0LprOPLUduNKgpJa8eJUXxFd/E5K0VMWzpyc1B7lWlCw5vbNij1
iQ2cRktmHTquJGPAjUAAA8ElDRTIlh93RZCzvjAnBNy+EKOdiZXy1DcgdDRImC4AUFVWQ4zmaMih
H9zlg9iZF+j07ZSg4T2+PkWTgU22dgxa8OKSjeMiZg9mkyAKneIQ8RVHTEeZZZTjdUpt/meuk0wH
f7rG/VutaFq6Li4hjDBtLKBeHT0cP0vhnfUxyv5nqDhadXcZa8+lZk3wItblX+CIjY6UqOhbcZAP
79gJUdk9hZ/Jnl+OR+sgY9c3eYS9D2ml2BgonI12h+cHM3SgyfW0UApJIPERMa43s0IiTzfgqckR
6gAJUfxC3qLpr4xgErXntHeha88B1Uq6YncRh2EAdlTT8k4MU2TOR10FsVIcMnxs0cHVtETbFGtO
mYOuCNBPYcEFTXWm4zsSi33LT/r1JFhYmN5n8llOL1uAs7TzG90swEmcy8KAekias/gloZw2ZuWB
bdk+62OO0IdZX+uattyK5stb9GOm3Qbsrm6l187g3osrTU5gIh2mKoIglwXJfhmo3OVr3XsXdHc4
Uol41OrJr0lOQscjsm6tbxaYEt0Z2WQc1zXVdyy2cONjrH9krANspiShTrO676gQrkCMDTqcP1o+
EUKeT/gzUgFfu8Sh0FWkJDpmuoPVZDYbh+lSEUqOErXbIJzv5U7nPmrEh9sFLm4re0NPYCBZqsAc
7g6IJ1M8t2kUDydKMR/IlGOxCB+CzF67ZInEj+9W3oZUKteNVLOZczkqy6DommSH1xerPuLlmTSf
3hXgOitju/+0nUshfsJVDOHbhWKe28kXkuvKYrtRu0M5kzYgxxStct3+EWchOWtOUjBSDOGdqrIK
PbCBYorkXYbqS2e7QSO1Si2AKBpEj8n7Vhl1KkqrzDTV2mIIQ5DRjwy/1JEEYsbI0Oe4tQe60sZi
RpLrzvA1OxOmXWEolyLXRtu8SZTqiKHvC9qUKV/8PP8o3yTebCXqNsHmatyS7ICgOcvJJhsFggoQ
DErIOM2hzs8ZVB49lBzdQK3O9cY9x5DUOT1nNZflaELpwCSkr7r5y3Us77r9I1Lm63yJI8HCVk/L
U2v2HtxY8ntFoF9E8AeNH1hySPfLDyiKY5RoaerBcu/3fjKdiTJP+UTGdDCbGdYdElON+k8nCiP2
mU3sd70h8tEyYd88Yw92t1ohm3Ge3yBrXY4Cin5vjBPt02Su2lsQx8YpgGxRD9ry/OzH/gvtbPO5
Ls10WIId8LCbV0fJj0xIRgZJIkWhpITRr2XUjmoiL/QLhN4zfOWmS1oGZu3skaimk6RTuNMKoi7Q
bKIj310PPJyYjsXrkIpwSuOKrFBhe7am3naECxg6QpR35UcEfMUk6ZcCZ0x4PNIp2C4MLHY9GOpv
mO1BU0AtuBRIkeDtvmcFm1D2zMfPhtwl+qLT/2sKFHfMiBXECKEm9FkPFW3Nw8jhXR0YTjZu8xuY
XMyyl8+/eIkVe4g53VFuaJRUq55/YrRmrdO8L5rx5jwtQPTBuyUIM1VUIDV2CRAoT3uhbiLwbY5d
+EMLZgmNnAXbup3Bfzt1RV5IJqaaVn1iTG217GTQ88feSOzEaE9nYaarmrkfyHLjbpQcmSDLGzvk
YF0TGNk6d4Ab5hj31EgjkNw9+bVHdt2fBr21rWJuaF1FCj0qL0mNBATUcolKzJ4cEf3fNmqYUHMg
47vHpb/D4Ji/l0RxqHQ1zHSYzGIXDISHZ6lfazArU+qkA7R+tXZgDeKd2tZ5nZNFxbbWiR9uwO03
MljKq6dtUivDOoKmSr3RA8pKYKJsXeBVDlW1h0zi6fd+v1+YHMD2QFBHlNEUOQIc+9ol41mJQJB8
FSp21YmRApdHYRYAwvOkjNAZnnaz21gmX6gwL8Orzd3GImI5vMgtwN9XoALPmtPIq1p7UQWL0ML0
vxN4Oaa25cLXOPSHufIfWdByd459x4r54cJgzieD8T2G90FzKLjiPeuO74pBSwMOuv9UovAh9ra7
YtrNdOReXEms7SWnkswHYVx/GJc3+MRJW8aZpxitaE9gSNdT1r88uJjOoGYrN1MN56LGkmL4mDzM
F4ad1Yg7p6rDYpb0+E7WnRUCldir/Wr5OHqrGFkU+ZwokIQum5l0R7KIy0M+XBHujlhk1o8bKmDk
dJrl0R8zWRSPnlMR9nuhlgYoD2xF0RmU4kYl78AzzLaN+M9uM2phcwetbTDMI4j5ToZa5n2FkY4n
tUlSEpc8A5rMyURNahsRfXqDdsi2suOJ70AyaS6OknqosA34ZMZyiKDT6pccQCHQ4tQWLDMSBUwr
Uxggm+hZC7xYRNBwjR7mL6eFLCfHlXI2w1K5pZZrVONyhxu+nM5TjXGGDX+eKP+UanxwBbNTCS8C
JwHanlHcfJxeFPH8dqArwTl6nkrxLDuPE0eSg+ESo4I+i4u3vhMfqJ66leee3B1+WNBJSI6Xi9Vw
B+CimcXPWPBgvYse7Rk7MFxb8PFjWkWBpwsZ4idAmZchiJWhNOcrPSwtBqAIQyjnlRyJ0NlMLViV
Zv02UNJTBoOGrpvmaD95BjEs6f1nU0NDlwfY96+NkQ5RwnmfhiO06OgnkTw1jTjQwoim59Vz9tVK
FjPm4+BRwO+J/3J9nmPEI9/kclonA3tp+KhPH7ujQytLznTiWRjIdspv2hue+rrxfMzWYEK/Xvzp
Mkks7sFijJkH6S/e0dntb5HPVfbDRaBnM1vEcVO5nPkqiNjtX8yIcDLloz8VL/meT0YloKognTIy
XvMGPK6ZX+FxFqogMBsCAV0H7uNP97ee7h2o9l2IcjQXchb/uODmk4+5mgpbbO6uPvjANbjNKjEV
mTZeajiHaJhhEmONaRt50kQ6X1Fu3l0c19LrsnciVhfJLY6+IhqSeqFdpoRmpKPkjQdk1lQ2Itwr
6Y6XL85NGqCBa5/E00WE8N+FH2GH6wxoweV42Newx/vxH1Cv7VHab7xaEJQ7Ttr73GbuFmo/sJzo
LqT+uNDYmLLP5AZ+J8+At78Dy1DuhgcxOWVdoADhTRQHjrbiRy9sW/e0yuLk9IKK6fZJzWuU4zw1
ErCD1DOkjKksLW56AMruvFQc4me3XwfAVTprNr6TdkL90s7vvmhcGcfslOnzp39d1WyENQNzxmmU
VCgZsdfZeFStHFilaIrJIrnqGRZ4HeU3XGurY+jLUzH9BuGwOpfShXdWwXUascnRLPF95v0nw2w8
wyiowjKCciQ/lFD+2isjFkrjJXYw89ai7rG/K3/AH9cjvITx87pfcU/MXs3hJCwVgrkrG44UlLY9
qaaxkwaN6RTB94hoUhbXpWjAwll1BW1Wa4E0TItxpmGj73U8kPUsmDGzjgaszCOYdqY2ODZ9U0wi
1zH8y6NPKKaM5WxN9rplpffOOkm4fpbdrl0TIGwE6QDAOaYSCEY/4QYeBPEDY38m5k4+OaQPA0WH
IyuIdV/p3lcjyDdbSDIWA5fd6FANMh5GODstlAXfM8ESzU8+PmxIEB/UPgPkqV5rJmNrWbQerhyS
3xYYEQDjpgpQYKMoXvUcirBA0fymOWdPR3CyAw5XSsQuJU5OoZmBskjXWTUcib+cx6v8aYRGMJjD
DLNqhjJtJz3rNUonSJlh/qnpDJud7LKHvqNz8MPykjnZR6j/ip5LTuixZbCZK5DUJB7KyH5C1pso
CYakGo9570d/cg3HEZdDD3l8+xmGsBYTI7wvxNID1OQ95u6SIUcVTQDrOWxc7vFHkT7s9ImFXsVf
sE+z4ftrt8SUzysTnIlZ5C5h1QnSDaMA6/ykod9F7wk3yjLBSjvkU8riCh88qivWAbR0cQ/ukGz9
+L/P3KSNdNDRb96qlotRGfCGzqnzCFk4qd8cIu7Oa965IO1O/sAZoBuuySnxUGzLNa07YktqP02P
UQmU9BSBuplwgHkTBk9m6cimszvJiC2o50NWu7kCRtAFxYpkj+t3iPtqavql7P8NlyCQhGkuSy8s
aD4VRkhys4B015Me2pMonghxYgyZh3P1aeykHHkVisez00Uosz4fV68ucG4ytEK9I9cPpHYph8Hw
NHDjdUduRL9LGSzHtUCZKSZg2rwAZ+tI1hB8gvFEkmK8uNQEAqFeUBfDwpR0M6OCLWa+MMtzAc9M
mpn91svloO2ufg8/KqOeTw2pqdRc9ISczoR1QvsuRIuiVNGpSIKneLCCDjKwOoQdzcSM8/lCGko7
Hr8Ol2srBR3Bk1j4X/+e7orkwHgGHPbeRSmumA0Fh/K6fukKBPlX43g+EIk8vclp8J2af3ZAeo7G
jo4x4WP1FyljU4LLGXI3LhJ9VBUxfZceGFk0YP9Wfe7KJgW6oz1BytwQabxwLtxa2V4wk64aQla1
eChmti1MADuZIB2LTxapvVetsrYJLnWWxsJGdhYSYTcDEPxCQscbvPOSbtkErUgbwb4BgzeSmc21
EB+/7+Xuy8Pju99+1XBFt97PHPHZM8Py/pAOuAmdiq2TnNffHzOtSLEHdX1RT1xWykqYEJH8B2Nf
sRCa2WWbYuqzS2EyaYY7hza7suC8Brph1fG7bnbG7NfY8M/3oS116VR7x0WApk1w1Pcrx2UL6+TX
jIKVfzTXVI4M8wTdW+lqFABOGLCFE5MKpOiTu8M0w4+2JrY67Pir0Ofhaqk4TqVCBHRge5aD/FTp
CH+H1XN8Zgb6VYLzn2yN8Zg7BI06YZQL5bd5dxyiHNSTtH4DW4FXGSmryvSxSX/u/OihMdjnISMz
z1RUTDOtqcrvTZm83foK+MSzFEPyWfSP20MhYVpB04wMmjRqOclQv/iN59lEtqFgmFAMF3mM6qsp
kR2uMTpHGC3Npqn9ojIf9yMNkHhk/0UcZcDMCsKMi56bt65pSpClFfuDDPcSe+uijJYLibG7jX13
uraw3O3BOf1QxFxEUAUDh+XfOs4G/9o3HK+yzTRarpOp35JFm/LknuH4cRZkV1ifr+0iOEIGJHPE
59w1aEVj7l3eN5eMQy+1FimDAfVDUZfypBXKmOP1O6PC/CXaFTVY4JbpdBVgcbK4Ikn6fhGv0eN1
/KMvmOe2k6CkPbw7ZAOZyp1akFVswGm7/27YMncoP2IRgHzF6lBxTubm2B0jyz6Ik4vDvfPu52lV
5GjQsKw77gUzL+ydOi9T5bXxUx4RT6IxlCnuOehwjWWqX7qYMXwewHa7zjJMZClZt6D7f19QB5pJ
k8kdUGzMz05jGkSChbUnP5olHoxqawPEpDUniXiYAup8jL8UNFqZAG4CrVwKiuQeXpjcWNso3xQS
PMuU5o9DwHWQl76iqTq576X2IEBsrotilYWl+3Q4pPyLUkZnRskYVdI4YwtPgCmja6uJsnTPcaxF
oDn4ycPVg1GLYDDeZLn+H6frPq9zQkzwBaiNkvCK/pj9FpVYVb30IxP2DT9qi2LhjSSquzVsEYdc
8GFQByiSf0VnNmSG0GAUCMQPqpaw7+1zZGm78Jpp8O2HRpT7P4NN3muO2eD7csjTC0O5yb9Y2lzQ
DfOCu8gBJmTYvIq5ITZejxpqxmi5RlyoipALUCU94ZrU4A/hSMKacXrGVpTb5bQjyrtAqXeo4QRV
lBBQUoTLrCelayOrGC0u7JsEfsi5gTazhjowuv8fiDV1pnvkXevqQWzIOgub9YsMo7BAumQQeHRI
61MxkSptahbjcqwZWfX9sjMsuiMwzs9SAzgNf3pcxCQQUotcSJKkjqecZ7gbrXYFH4/3O/+SI8qG
BgnlgE5Lh9FM64PBbsBM/pd8D8ibaGuED6u6o5gwtFNrGkxxihW+6zq8p0rxmaWNcMP14b9YAq1I
redWu8Adr+XAJgWSqs96Ge9y+2dH1wCeKWCoPM/pu+FoDEow0NiFISih+w/DrIM269HWJ0q8HSQj
tkIChY7sqvfFX4Qib8UAa/V9UDpEZFqvOktDBo1R6tWPUYZBx0BiBD9KCBIPMLoHhiGbXF+WgZ2R
YSnnx2hzAyV5bSjh5G4qF8yeegdtKrHEhj5SFXTfCrEzy3WetHpdfTMfWANYJ/63t95B0VvgInPA
taS08ERdYK9uygJpGZ4MlA88OXgp7Dt4IKaTZwsgLJA5Fn4R0QAJ+wVQktQ2jhkbCOEXg/6Sx3ST
4Hxp8ocBhiXrD4c4Mza7CaT4UCkZdWxX91tG5d6H3HOGSsu8/c4Z8jBncH3YjaLlCGTTmiF0dYlr
JF/WiEjoW/lMHJHr5xx5qPsrwD/oU9r38oDAxMupVWlcbznKddOfQk5VKrK6hVAIQlcdMf/53an7
hHvpKguqHOKH65R9ZXXhrOJ7RxLTdvyi6qLJcr/0HccMSS73eylLeZj/zIg32Dd36ZZLMPE8Cbkw
bK9M38ISionVPZPy8hjmESmW7z1VlD5j7WMpPQ5bkjHR2VtCQrN+dxy3fHIhherRdFUS+TGC+oDw
kpwf1FLacqlTRpB4lLE0TciEovT04w06SVOJDkiE9HVhPjOAHKwZhUeRG3XlSMzqVQg8GEN3BZ5p
cGZgz0uNYuKlu8DXyjdZBXeJJr5Lmuv9caBwP3DtYxouwOcqbs7rqMdXWthXE2169qfNgu0kKp3D
/ROipsnB2H/mKzVYseWxouWu4Np072pmsA+kdK1lARegeRJsg+ZByIBJruEJ5qnqCidVzuV8F6A1
IZmX17hXSeKUig4H8Qayx5WuzpjwYWKFMZ7GKl7jCjA+YKLhmjlvpC2255rOR5Nx7qeV5ezgm9sB
dl8ziTaKUluc1F8Rv+87Jdm+dqu+czzDX7hvEQUmLPNOO6hS4ek2cN9daYexw724Cp47vI64EKuC
XkRQFL9myE+2reXbBaheX/uUlBK0ArzXnd/iMM32wgoY/6H7nEe7qY9Z5iIvKDxzPDXtFFV5on3E
9oLzyeangFS/B5DPpy4F3CmCt4xDFRoFthWwEIWLbjThsx6I3Yu7KDJpD+eUEbAb5a49MP4Bir29
0yd2oyahPXVbC1AhMPx0TzeYOZJpo8VWJsHuMjYBE5LEsuGFSe4KGabIXNxdfcm66yBX8p76JZSU
9StACwYz5n3xAxtzLdjaH3DerIpX9JLlsAFP00qZeX2rmGgfO/da523pjcodgEJW+49uh/1+/J+T
KWWFafkuSY9e90TAKskao59At31Km1zZ+M2Yp+0o+vS/5OUeK3Ysc/Pf9wzpqiH6bCbpDn5xgPrS
ZWpJPO/xX/mAk5NfPekKHTd1NpB43bZ3RqQyoekVlqlBDgZNTEBBtrVs7iJgKnTLNCgSs9D4Wwbv
S/NyiYQykT9ZX0lC+DomuOdwTxtEAdBe5n7KND8+03yF8vze4qOZE//3s3gTFal1x/DFQPpK2s7j
W+1SCvBO2nvZljuLHzwhTqM7EJrmp5mPZFx7Ey5vj3z2BBU7tnG+qedM1jDTQ9aXxaTvijnA8vU5
s8/CnFDkiVbfUN4uEIm92K8c4u6sEe5hJsuCDB2Gv2errgfRMABv23BamwITeCctyTLLx3zf8T5d
U9DKBQgAFWsmoHGwY+kPf9OVkURqMp38TAB0v9QpYxjpjzbGlSqfJFImqcGv7VOHyMYibr79mIQv
HS3IcxprNJ3SLPGQ4X4J+nAxvormOkLJR43JzDVvY028WI0gLywd7K/rkp1He7AXyn6oBHGonZdS
H8IjU4keLtfgofhZS+4Y7GgH89rNNswrwK9s11um7uWP+5VVpo0dpNrZjBZlSOxhkMCP1hkjNIkk
6w5DStWnxzRYUrBvx4V/t6Oxr4TdhRcP1RazeYk0k7C4fs+Q8Qfa3EFjNVbHqojXtG2SXW5wbnui
qKm4lb8D9dDvW9creT+jcWNpRG79PYtAIwQDEH6h7cJQoVkMbbY12f3kRZjj7DEp3WtyaIfh1o1D
ZhR8Z4vz0/vKck5KuHzQu0nsng2BPGvdNyqzS+Hvkuufl2z56SYPxDbXZoN6yu0oqPciQeZRnrRY
gto8cqTgNVhLV1vIO2eVOs1aBfaccxgun+s/7yabzhru7z3RxZ686f57RQs2Aea0oiJUsXZBoWj7
kVdoZvwXK/Jve9QiBDT2/fNBtTqGPF+uqPx1oNGxia8iKczA0GvlF9OA6dBYes/GIMeqSNJ6oPoS
t3B1lMhQY/uAMP1mmSmn6oEHJ1c7IALncmlIpRMn114Jzfi5o3LW3NH0d9MZazfjChOaWyDpoqDb
O7/iWLxE9UNFBcOTuuI0Yt48AIPm+S3PqeO2eqmo02BTr0CX9nztU4m2OhTvYy2FcqaMfZG7yjfe
7yDNmhflaG2ZxYRFvgB/+ADASBFSUMHAYv8r7EUPj18/52GyT7hZK+bg41bjLRvWT4FywM6E7kUe
05euqw5e1ru+EG5SeO8RIO0wOi9DpFSM6rmVrgEN6ze40y28N1NjMa1AlErVh6gIjpGjtSGHEYq0
ORsQYb6no8vl0yuLM7hqkfyM7HvvqW5zuJBPqqB6CuT+Snb/zqR6r8CY80PV6RHe4j5FnWcBLmSL
MrAgsI5JOCBwlnXv4cRJgPuaGdo1ImLZynsgD860iPJsck5H7F9j2v10AunBJxb8MSEIqiMsOLL6
OJay2k3UTaKAnfDD+5lRnUyby6dIRlFDfZIVzlto00+/vwXfJHh/ZBpxW3iKID27AdSOAZKVoQHD
NMPVD5iOhWHvjW7MKFElXRiYcr67tp9HHdFm0BrCac22aKPBLeerNJvb+ejFzIETobO05DKYTjrv
oqZmtkAWbuEYSrxgi9kWIjdkA0WsiqYSrc1llHvkD9V5FbauhVeLQ7bsXz0XFnEQmCUXrehaQQ8o
FrVGGvw3xUqXZELAZbabj4LSYIaSbfd4XbRnGqE07/9SkhMFnyRmbDR+ytQS0OIPKm04HCsWq1VS
08zddzXZgDKpsXc5xMBEew+hFS9CzYufZo/IrZkUzgyaAINATXa9FCGoRTVYmBKy56WeeHy4ketg
o1IQ++KopRWRTli3sMa6mZ3R/2fBGqkolnMc+HlXuIOINfnXov/sh03iVhPl6Qv6n27TiGEMymNY
KnS+oc8L93cy1Me/y0di6eCPMZ37HxbZYmVZw2bRrtVG7kXh1Xf+0c8pyzG3ciZBA/sFmEes8aSm
AH9s7WwwUIaDuCE3c/xzyQDTifT0f8Un7e9+DQqludx0ZZMag1+uaX8YtMcwn3ohlt6E7MMDb52k
m7PgVKx3xlPxTscycCvXNWaQ/hmvefFGwRp1XuqSZYknIIt0hpS5s7+Bbp0Jhme4eiCYgjOq3Ylz
eW0WrZr8Wq/JDAQCCgf1WvgmOwnIn1qkHkFr2Y8MgxrWEeetgmo8hjgmqsL7Slf3+4AUkQd3GVTs
JkiCqoCnZfGgN50lza0UEBpcYfKpjR2SQO/KEZQWCByQwUM0RppJCVybeE5ciypox6F0qlIIZh0A
SH+7THJ7xAHAsLjk+5wZK6JzpB+cRPsihhmsOxvUjT+VHPKo4mX58EwdDYNYKqW4OWwg69s40tIv
T/kyfMksvEam7Nzyu+o/LJlqo++J9yHULBAUUPyZI9M8mgMEwAW4+LdGWsM1bFD2trIh8I1CVy83
X2Ghp0izMMyCiRFuAgidb+EhoxWonsU9O7ZHJeSdezoH+Z1q8eADdpdTx8K2WGvcDeGnR+ocZYb/
yaxmvvEAYoUnLrBFjEyrpYs4jd051eT/tz2a5536eNHKh+fCPZlvtKJbfK0ffo8L+46cen6E9eC8
WEKSy5CXNsRziDqDwp72TKS87lLTyEgV0XxdXkP4jG9ngUF+SCUnFyaenkvo7VU75v83opo/vQ50
luSCX8K3bbP65GW4pDKgU7iXqKnIaIwq2nDoBYMAQPXLJDTPSwiPIPRN5fhJ4emTBNIItUn950nY
ibaWewvzJwCQXIkDoJwiXt7m9IqYSakG0yEarVppAViBSVICoY0txX3FVNAZAGDlkICF6Q547Ixn
UILmjJnlQvNiH7DgHiK7emN2wlS3ariDay4CgfK7KZMsjz3VPytcr08gcCBfCnCJG9IDVWIgYkgO
wokHLHxIs1p/FhK+15v932KGNY1fV1Ky+tKVEgZHbGhiMHSqrS95NIPEfQXJgVf72r98HrF7oUO2
NYDm9+/iWoWxDdBcQPG2pI+93jSRwDL8Sve8ZfylvzYFdcLjes8QmugCfG5KrJdLjJLRfYLwW00W
MRGq/tZdU1loLKXF7JgOE9HM1o0TnvET/HX1ahs488FG0YP3VXC3ax3fGR7YgRBp5KTewQajcTz4
BDW/dMuTL5Sl8rkVJxviucUnWXKwyi8lMy8/eHbe2E7lPH+QKS3DPGhW38TKZHOYQO1RnPD1G0PX
V7B7aflvBeApo8vmdyaIHRBLdsYzKLxVOM7S0vKL3cctOb+01b4nH4323SaYhZtcI9YpgBc+sEor
zQZcVhBAZfpRcOzNHtlxeHauFrxYQpVR7J/KkT8i9YxRf9FqiXrqcGXfDqlxcFMQdvRDw2e39623
TUTE4iTFNu2UetdJlgjWmbI76xU/fGPAifgNyWYYJiLwJ0gYtq1uzr2aSrPbYkNF7Gz+aZL18oTM
HgR4qmSdfkIlJIFa1A2EbvCFzFI0wujcFB2U1ZoLDfzMe8GGwiIE3S3GmEyy3lIj/j8WqXYSBi5c
s6laF3dS4BcqRHmpKobtS77/asl0fa1vr7bCBjTSWJnu5IXXVB4gz5KDy7ZNCmv2npngX/09JoKW
QxYa9GGVcx3QgG1xT9O8iZh1vDsQz/FV9HdMudW5yN+y6Pc8/MV0nvHI5Vrcb1+2tDRFfuY1hy3r
UzmFacIt8nw35ysWwryw+SMapWnrqY9RrvY72iD8PuKfZaeXs1SoOH0nCyKdEUQfZfWeDP/Bbtma
AmGSe8HGvX2lbkD54DHOEnFrYNApms4T7U+jr6VMpea54KFtfP2bNbLD5PcLNdFiXHBL7tskAvzn
C/Gzi5whzgvqHbdz+3Fm24KLTp7ZoUvUV1a6B1LfKBCxqtuqY/CKp6rRIekfAzHw829KHDz43mqA
pr65VBK/advTIgL/tiufxEc5wnvzkUjhTwCrGPf8Tca5YnSw1j6A8ThVI/g1JHDgGzn8Z+vssKQ0
Od2NgHKFcORgktokRHheNI3Kq7OMzhTZTEiwh+o5pd6xnBor8Ewgxisv91xJDyB8466Z8tqj623g
W/IDnYnJWzAWsMY1Cvdfv55qwMT6plEuXYwLO+Bj0S1b1LCTqoHgGimecKfAFQj0GD0NGqH5F/Vi
ioiEF6rO1FlFgCq/iTn1nBaHB9hLBFWufnkQg+H4vhh0455UYI2drNEiuyPMzNtyfcxORdB6LTW2
M/8kmDfbPgTdTRqPCdDCjp1ARdl4w4guahkk60rgnY+Ileyf1Whx2B3kQ66a28YFKFpUQp/9ktzn
IiepZfm2N5pSf6HRgGEAHSZzdYq9edicaxAcTixiBt8UCZTfmGuhWLJ7qbe4k/sXDC1VT1aXhg4N
1Iveg2Hqb+JEWSsFDvnmwgmXnkEfhQ+YqwkK/NLnD85hQziQkUMlrQp1ppzP1sF0CVLj+ZyWXroq
Rgju3PG5iWoz917rZU+rR6h/RfosuMmSnPl1GdWn1hNWP4OhJeiLJPUim+JR1CVO4jw4u6r80jx4
2APPyS/rgHZ+HeuC1sAspI4ymB79XQrLJUHDaWbFYHIuVJQ3nrOqVTlSbeyniPd6rwqctfrNmxpe
V448Ba1gNsxD72THBLUgq28tnwCgCpEiP3S4gQiRD+5F0tn3iyHzJNmXI7IDkCzOEzMUfkLYFZF/
a4MJrv8GwukMbZNPNbcbq+qXlNcFefZ5kIZ1z6px0jffDi6pbwWeTest0K96lvMIuZHFiT/FHhWx
kdn4asVkDWplY6WSMRbM+bwnjJjv2J/5sQPk463tjC4C72a+UjJ/vQPlAy6yjde2jQX18W71CUhQ
fhWR4CjAH8+cwaZnIxG0mtHwxd1zGS0jJ1J/ttgnyX/7qGPwJaZyVELyzHZ1yAQUoiWkuoVH13Re
ltCNDT1xgtko5LbjZtY28hGu5Gc0dCKgX72O3GnXkwVPzLPZcHN1s21Mm/03E0RDbrijqooUURrp
0nSVCqr84nnjdaWZzRcixBfW3SrpdVC8WiaS5onoD1DXCEKzopbc6509Pqaol5OTq36eKs7jIRsk
P/h1jMi2m/nTJebtfgxDWvUpxVvWbngTfuTmDXWHoDyoRSABbnOhcVC/unsBdnpD7CR0GcV0Gjje
M+/BAMkCy+mxJakZ7CbdLa9qI3XlIjuiaUOKivHhnc2wNPZrdKatz8klp+x5UdiD1uxBTkRz+5PF
Yvco9/wY8QhTkc034chHXI2Z/cjwAIrIMJ2wXYQXE5AI/9e9r60sI7BCWyNVO0CKw6Ol/xrOGhaL
7biLHEx8nPmpzoHKDMigCwyXiO9I4KWq4XL5LaAHo341rrtBbTOZCFewAKvd4BnWGm3jqtthTzn0
kAdPa/4ZqmN4g5UmKpou3ugwp1Ixxukf8QALe9n5UX9MUAZfz7PqQZZZjuooHLzzEPfcrxUnoqfp
ktzX/8C9HqOXUCzsaUiMSp+MTvtIRwiHYeRL24laRMYvv13RfbJs646F4swe1q0GvECs5yYQ2Xz9
9VtNWmE/Cb4AIubS/kfEzYBrMcuuaHEMU4fmtb8wo9KkX1TqPGg1qo5SpdKnTElBxNYwp6vDp2iq
5VqJ0WDIfLiLLW0cpHu4N5Qe0Dgah+stsjlBcCmnfGS1OW7+9PCcx9OEj46PZdzznojY6jaSHYPe
vAwiK40dhR3y1dpUoWH9XFk0i+1vpAlQFJaWbEa7gdIK7GJeD5bZWlsVVvhl9/xNfpV7n3wq5e1V
z+p0R1y2d/Ji1RAADv+inmrR1j4BbnseFNGvpcrHmB/4FWa2QBWRCiL2X3d+6Dz7dqgukZEChO7u
bfri/KeeTKHXjYTt35xLsOJuJlq2qOY/7bbp39t8Ntlj3waBhvizxCuqhoqBfdxSLE+wctZj2EGh
Lt3jwP6fj83rKobaM/FELcF6MzV8fY+Px6h4dxhQIElIyAZXFGT8O2VEHZGALNE32S4li8FVSR/t
nxA7Nmptf3ROAkxBVrr+oiO3eYWELzJxZtzMs5s6/vfJXIx6pUBcl71/+a3AUo7w+OLyBCsBBPUG
dXWvNc+nwMpTD31vBG01pFbJjX3C249kZjrxeO9wgdEowk+p4j09108e9TgaDhezFNvv4xQAHI8H
Zjp7ED6B0E+dHYgG5XIazqbZ0HCqQHiG9qsXFWlgEc1ALHF8XtsUqG4sBWMqhMagozY86eXwzjnt
tDJDsCATDiE5y3t4Ywk3HTYNLpV9wTn+Ir4JpmCd5ib0ASuXP3cf/hiEo1BQjOSgE8ZSzR6wk+Ld
GTNSogXwlAuBQsAiIJP8W6Z488SYxsWfqgZEAAs9+Wqv5Lidllq6F+mre1s/whdKnPMqupq15DbN
r+TKr778QFwEZhzSGZDheNm7nFt10dxalH3P8UYbb2g8oZcuVHoTBsqDxNyjnPrQLOmPTYddplgV
jcLQYFeYsTckQXmmW91atf6TibtAVVGk928qM3VfoPe0ijmmuTZUp+LHvaAv8qSQOLw4XS9pHJ1D
9a9JH1jsfIDQNkBTNLvfczpb4smvNMVXgZHuSu7JyPUuy4Xs9n3aq0OLWCmNLFlh7E9DP2Wz9BQ3
N9nnQByPAkqShfQp7J/X5BZNucZplfaZU2+rz2c88LmDKs7wX49G4jkR+c6jYSCoLEqc9z73DMyf
JgfoHKHlpSlRggzqWTRJQQ8e/lf3J90D6rUrdRMYAtY6tA5etvtSafcyZvNm6NyQsWULLJstd9RK
0QpooQv8s4gKFJVIAxz7hsfuQNSNWtD3KtBSnI4rJ62OZmdQ4SCoB+/2mbPgqBsmAG1oHFUoWczR
LrsysonfjCDMUwFidUs3MM2F+rtpV8r8NmfWeJJ09N3HuM93nnqqRA4Ifx09h1kLLMK9/amih0iC
ItJjQ79/J76MHNZYirPi6kvv1rlUjbT+3SrA5ukWdeNiF6r6MNOM/IqAwm0jxamiXNq5OFIk+/3O
ZSFtrkzxXALH2c+2o1G7fULyRV7jC/WrAiqofqZ9CtlNjFhBM3QDzgJ75h2MvpCac+KQR/aV73YJ
jiNc0e9mleXHPI/5S19/E8Biv2A8YYHi0anUE2Iru6jv1vX/1sxXZPVIWt++RTv1Pk9IbY0m+d59
6/alfb33Ys2pKUnhHc/yD6APjPhTL6QesCNOrUFLrjJVpSG30pKjq7NCHxmHSNPpg3bS4fd/7FG8
vYvmHSbeizjPKPODqamSaQq7Z9+R6XuJ4s8AfJx49KnChWZCradDvPU0+gaO6nLIg3wQED3Kcpxv
gN+w38bvk5u/U8lu50r8At0v5bGGhaGKvl5YbOwCcnyYHkOiiRKni+7fcSX9ofqWvHUNE8UNka2f
ZAidOGxEYn50YhTc+qKcbY6W4+zerQ6tS3y0womwSrl5WZcmx2CzRwcW5UUSRKRSQeqdXqfoK+SA
F4em/O+7fhRtsCyx0x1wud2jHWjqllzOizgn2l0wurMMo9FmChcdMkw075lyc+olWCoznkzG9BGx
MXacunE4IQRzuJOPFs9P7w2brWJ9hKprxxrs5jgAgJRfFsn8nLjBXW9f+m03zmfjiAWlZb7tyeIs
BFt8OQy5HoMpytKJwPva6FVDZ+6hG48f4bJPQ513qNl6NLN/82QY37kMPmcPJcA4zf7wSEBDA9P/
cUWPTteTwEit6A+OFN073QuQR2Dh9u2BNQI+pRl4Lhw1r49b6Y2NI0SS6hNbwLT9TSLHCT7ngNDT
yLP8/0SBb/gokzmb/0jNI1Ghp0YW++DJQyc3xZH2YR2OAAC6tBAsvNXl2uiBJ5A/vtdQNl63v5V2
M5avehusr6zqfJHb+5grxJ24pfPxdkHL/KuiW35uzkYSW60TUG9IgHjEMipo7GdO3ctAOh4cCRFN
tzRDgA3/q7TazldW/SH5G2t4RwGkGKCtT5xtdykINSyef01TSrOodxKhl1YnMMyW2aB0MsTN5q2Q
A/163neGKhriicqCw0ZNtPS2NfLB25sXD2rSXIvy2oyDsLUSbu9xx2xyg6hnxfoorMq0eYmDArYJ
SLdjpLcfHvikVdt1Sgt6ci0GCTPQr6OfR6mbfai7k7y1Wkosb/c1JI/CAGkWLRGMMdpGd0ysShGB
8TOsg969Uwf5L03jNhAzDr0m+QmEW1K8/OL5+kLZWCMpKFu52SCqjvwIBKQXDwLonVgJF9oyQ+gm
6xKUFklCygbILZ5sMzXSo2ZFjWpMUCP5732ZjVU6mak0rlu9qCGND7coRI5YlRDgI0CgVgtrlKwC
Vr8L56ysXQ9Epx0S3BLJP9iFGdlHqQg/ByxJ/DfgiGYxz8mFJrALlKiDxK6CJZOAv2NHye9mNA8f
3dcONbJ8ACgLTGYSF/p3w5rtGW5RvPZqtf6XyAOhF6q3okphsELvSxHWg72vNld/rsr/BzrYKRJs
tph3p73Q8ja+qtL/SPTzo7ShkjGmDwVS0ynmj1o9Z5UQnb2fPiveo+Pga5tjQry7cSjlcNCwbO+P
z9zppX2Lu+x3sdP6o3Hy6zFN1aumCQlCAB1cG4QePdlZlAifDRsZGjrZMYlIazMip1slgkJ8ZB9u
c+CN19gPhDat9FjzGR7v3nx4n9XXOG3XMLWRRQUelJ2Yvr5WXWRvg5HHVM+NjGH/ZDDnCv8Sjj5g
7tCAunhvwG3WrPX4i/0lNKj6vEiH0FhlI/JulV2vzGIkvLBOT4BDjy6OzI5BlLeFOgLPGFQcnnvY
KwQWY+TRmlpAPTbZFvoh+bf75MrWwWdCIj6eRud1FlP8gOwATXIZpbru6sBJ36KdPFPmSVNSIpCB
eJAdxsVclxQKM6K13XrJ4l9WQbLPhwiocX5V/MS4swrtze1998wWfkLyHeVoqj6mvwAb6vz50Ig0
wxJ+vGYQ/578FcnTnnCgkFOfWeCPdk7/KKMO3A9g0BJIJjsUnLpfuPF/5Zy4W3QX1/ivYY57LtLv
1q6t1lWOoFh9xS2/hIxHR60epgpssPC3DBb5JH+kRpmCvc4BKh7pswSIXk2ST6fUdvPdno3Sh5/i
xw2rcQ1w529lXeqGcfZHevC+kjkFbwt7QgLEhM0gWhvu17iNcvX8h0rNTuoBLYkxZU7QG/W4U0e/
xYhPUvbxfNdSMr+ZPPe2kh20WAy5LvyDCCNAo0JmEUU3fh/dMdvIJwghilCDu/kql/bYB+uRWBZS
3NJcFyeKECI98JIcW2IaHJZlWeAa/Ih4MFCyYE0s8iIsYrxXsr8ZVmXVeFIlany94CltQN3X2Nhe
0QuAz5/IrOdjpp/7ObXNRx+TQLobiLr80krXxDgTPEyu86ItWSr8G4n+mjvcJAvrzdgoWL94WdEg
8Q42NB4a68jQendIGynGliE+rvsPo4RYuzSyANm4ArOK16PLfZAZrDyeV8QmyO9OO8fQKGrSvfZH
ZW3fLH32zQvMEZB9MoPoqPBliW+BxeMWW2gWUoi2slKuMBZnRM5Zs0njVOfoq8qQ5uKVqc+AOXAV
9EN6SszlFqIfict1FUtHtWFjcpI71lHflinA4lGver1okYrfsNe+SKeu+mBcbDrvRNLaX4W9dyjp
LlYQ+KIgGHusdVb9J2lnH24S/ejKZEqkvbzgciCHVf1+jvk52HEbtho4Yd2DJDlIYv/U2sSq9pz/
PuGjlQmNzDD/lPAnOCzNSdqPAHxX1Uq5cPn+UpXr3dJmJLJfpThgQzchsSNxkxhouVnG4ERoz464
I6I+zqSg3vknuXW4OXleFn37ZaCtm4FDXJafSiRp+LwpX7BImv6umy4zT88oMYTQ6yJa3EPh7w54
REc49wSvj1wTC6XwDk/K31SIUIGpTq+Uu4Wt8Ade5s1RYU0Jws6CzP+NgRJAJAN5dgMB7J6NmLNs
5ou7IzrtDhF3a86f6oPFSXu9CVs7DfPYrCgQjg78REKYCWrLWW4KApvEGXy7BLPM40zf2rIHHStG
FeusvszL+vKNf57S6RlQw+iefiIDCv6dUX0rXqe9sMLZ8+CgsJ1R55Z5gAObpusZ6lTGpeai/YB/
JkGYeMWYaQuNJpTp9DzclN3PKbXylTG2u/tibqAQVVigOhl2SEfo7j2q/sekja2EQCa4Lxrcx/1j
puP8+DVGGNWOuJZr0FFv6MxBeyFdvJruvMiuCpcENiUw46yZ/D9SQazz7NFWNHn9W2yzQXaCCRA+
yvWH7clmYiq4Wx051py3STm5NYyjWSSxxlJDEjJspY4qb4JlK/govc+4Ry9Q9HhrBaWYftKPe3aF
YrJ0RDyLvhlMSMWNqxH4vpQ5Z6LeOE2cdgOrpDK+H+Pk5OSup11xW1Xeu6wLkUbAQsuBfTtwI9tB
49YJzmPyqhZ9EWKDeqaWRY4SzNgVBGpEY1zFHAC49rVHuHlXRN5fDELhG9VoV4Ppqi7y1DlwMk59
NpHhoDM3kRK9AqHeYbhJQFnXvLPgRVhyg7kx7cAhoh9gqNi2ehcXd6JDZfQwlDkj/b2QHoDR6eR/
/K1DziX6FjharB/ZMJ5+SlD3BUUqPHf4HG0TWPPAMpjqD4pJL30WrmkmRVy9otu0qy7vyX0s0xDW
mxUKgsRUDbxtG+9nL7+qVdGHKlDDpfkppS5Bt9+1pZYQ7p5/GJCAWDqWSpKjyhf6DneB+x1PCtmF
R8Ra/pkEzqDa6LHpRFkb6u2Bvz/XuG56OnfzO11KXMltmtOUDOHY5FnJRXFGXQ51tq9yuE/tN+UL
ic3Za6iNpAafcoszDznQCy1NSrYJ700Iw3NnYMD9i9hw2XhNxXeqfSn4Jb3V4FVjFvML1lSZZmWU
0XhtmRCMCeH+QkCovXmdNbk9FpEbb/qKddTS+017gUIpCd1irxu+556GDik4R/LDCiprVA9e9sOL
fjGbEIvUobYRpUmofy05C7GMsPtiKbotdLlK6jar+TKriCyh1mYmzWKpAvQ11BG/VpUs5DL55Dit
VMdrPOQDBAcjLER/+iMKiSnZyi7aNJGdXr5K3BhKTi+ONBmDseWmz8w/YECG2Y7sDPV72wBX6KQG
6PaWjSMA7naT7D/voeB6QWuRJG5KNMjigx7Ys1ut0v+63SHHWSSQk9IWb0Rjyf/R4Xw1VnzpDkQm
mw1j7YBFHybY1VG7itjd/jef33a//k4deyijvygH9DWOqeQK2ctPPKnf+RE1sve28DXY1E+asv4A
Gl+fZnw6bp1lznN+TZdq2uusSTd+Pesu6HiLVssKg1I4U4bUO9MM5j7w5x6TSHfKOeUiM4T1R58u
lqV7y0ohPgyA2urkWDKFXabGfTjQLMtbsZlLb87XG/khEacxzgFIKssRwRp39GjDNb0WsMg05L6e
BvLJ/CjqpFLZa/+lyD1MH10QkGPYtoMyilYo5td9nFvYqaE2H0vikLMd3QqxSvY6N2ivHRUx9bFZ
edT3ORq4YxBOAYPXfbGipyMS41KTTAMAWgGrbAwDV3/eAuPt484olMp9jd0CE/okMdagkyVF4Ix4
0erC2itIJcsotn7kLkZJMl6Un8VRhrfYhbSrd3S/MMtFX5sHfxx+lfVSUMkXhsz6QGR1oZdmtn9w
MjvrQD/nhlzorRdCJsaDqkkayeRQVpRgb0+ObTnKdOlb0oulTYLFqFODPdSAkO8S/CYPXC1z6/6g
R7LlFyYniQRIUj96vaIjuwFSTKokJFe3PHJFdNjbdS+n6yeMWCLtx1p05AaT/ifONNVIDMXhGTiY
TdYZ91ZLxT5quyCY8GoDv5JN+N/UR/2hy9Cj6oWVCcW2Am56WjyVugvwNxBwuee7TC3ozDfODRHF
6TPgu3FGhgmkS+Qhvyq7KTbqv0NxKYPTcqfmUXtMhrQUnlaEavbfzloZin3iKrDMtU4bNmi1O2Hy
bKYwjK/UzZ45Bz+M9JrGn+hiOToI3nDtPly0YCktT2m4NuPjOqz9bzu7V+B2tGBE04smy2VVRMaC
ClZmPic2rEylZ/okIgXp1XOej6u37gtHCN2kDijisD7LFsVZvzMVla5t9R2jRXilne2KQH1wzhVp
7foGGRegYvmNjtuymPmeWxNNINkH27m2H1gCLESlS7xPJuSo5g+nOzSAl1mRXLGANc4JSP9/UBVK
vEodcAxrDTWqHgL193jMAlNtwsEi65rv2VuvBoS3bu49efGM9/H+TekQHuKylt4c710lFRv11dIz
8Bw98QhGNGoCnQemgUyHDh4oxlefAkX4pQZTVZTz2W48XmgGyeP3xJE6pNAGDJK+wXB8nG4d9w3I
ab6yao6s2zQAy8wthRnOAelqzxT5ZSVcnOLyLUzJpfnT4k5jsTNAvbHxuZqbUfTJKZsHGfyWV9qy
BqVQ/WfmZR6Gid3BM9CYEL+dYjJJrDid3psIlBA1xXPXbzNtrZfnraziQPqmGV90isavzXhWkxS2
KeIu2LQ4OCdQJ3v6DeoYDUka26NcBRBppDiIR6Pz69LAAQPO0FWLYLsYaPkRz4CwNDCI5eO1nDEP
JPOyZemorRD544WVf2wVj5q4LCTFhX0MXAtcfK16JQ8IsTOFWn0iihCNIH3emWOiApS2e+wyFTL2
0wJoxHIoP5XtMq2rM9fazgre26GXImkJkDmJW1WOyxLmpzjNF0IZaeGfjoUM12emsbPO+XYQurer
nTUYCW7h5PloMc7Av0EL5QTIJvLTHm4IAlR1gqM/HmfiYjUki+oikCOlHPXkhKzZZMP+XRx65kfW
+lFQn3zfr/VRLj+WK0XB1xHPrhR1IZpN/A6iqNZv4Nq+L2oIMHRpTKOUccc6KAy0EnpK6qLJBqgY
zTqVb+iWVlGOKCly/624B9dT1Xo2GmyCvtgsO2r3nIuDCoclFJ9A9FsvPL4o63RuC8dMDUc3wxk/
GR3zZ0XKxp4lmsOFh4FaZ/vSt2w2OtBDfHvg/jOePoC3h6np81g9ju4W3uI+DzyHTz/ywi3RdHsZ
hnGQJvv4xdoO9f7OfjSQDc5M5JcO3sllLtIOPn8YgpRZ3qt4vy/u3kErmhl4mIKDlLS4nvjYGjV6
KuG5FhHsEG+lOrujvISlFJT9f1mBpvG6noQhKm7xN7uaMotFYk60oGuEKtuo4Nv5L//1WwmvJcgB
YwKE7/Fia/wSBAvcflY4tHc9IoQTO4k960915wSbSgiot1OpB4GYGPUePpV8F4Ho4BttiyScJ9oU
8FspxIMzS8z66hcLKOEJhBudcJhh1QoMt1WRVmUgbKmdDAfusvocUnirZmBVprgsKHa1b29qbiFP
w3u9khrRaT3fDXsOWGP3cq9W8yF65ggRUQYxRZKCx6j/UAyCOAwXRFVZrgJueM58PY2DRZdKNvBS
j9m0VqJD8k6203tAv5pbq7zaA1HIA17C10pq+js2/G9or3heiPAJLbw4fLLgItxSu0MCuF3FU4l2
+mHQk+aEzzgab8vCLuWY8P8AxDZnPjaLjVU9/8KTUq3KKQ55g5Z0sAsH+MLcrpTXSOFqwC9Z0qrv
PsSdASBQZe3Hf0+GC7ezY84XxLT50k8+obOdhc1l1D5S08hfk0dcPNjpxx8TWzB9z83oxxNdCtZj
G5nPAylZMpruZr+4LP6LXuG669rs1wqHovbOXW2/FRHWQYxJqFlQxtM9LXwemqDnbpJIct6kqObc
YtdQjJUF87kAUfrwvrgz7tI8afrJoYHcbLHhPEG+qvnPVz37lHXV6ZVtvLUgLghaaoXvbm6XMAk3
6Nh4ek3Np2/eRVpcALdbORmWUzymIe3VRjZ9vx7vNpvD7AzaDLfWTvsL4q0Y0he6i8aClk+8HALg
a5XX86/+G6i4WighWfrZVkA6tJbAyk7saEwVlgVKRx6lLUqNcPE/fRl3ayAidfiToTtWNy1hNjjt
wxyZinj30iJBkZWO3kMM6x28CCg6UNutzbVz8hibNTPBRhMybI+5JghmKYL0pDMBEvEKu2HXXcmu
ph21pTUaegXW4Sr2kdn/pl+j90pqdj89MAMFm6tuMx3r3GMCfrCgAFJZgN6BKgbkHJKMLQ5g50cf
Wex0zvyovYeu6g4bAU4aCCw+sM5aHRKCTIPFhtbKh3by6EdYy16UBj38Jt7OOgQv6zwOEVcIpaP+
f9FO1eDLLJfy6JdCBOMgrX5zLn9IFU4ntNASRy3DGclpYfW+CQMALwkXg6r2WvZM2vQZ8AT6ryjo
m1Zn5PTddFIF9FTx5PYdcOaa1hZi5du73hGNEQXBoOAjW9Os0gDGAhMGByDeJymqC+f8MDa26qE0
DtPkd3rvpvY89zo2K3Jo2Yn1lsjIhZ0gdA/SsYiDB1j+GTMT/D7Y6LukJV1nA0kEvMS/itNI8emM
Q3+aCV1X36S3k6ovx3NjdME2Rx16X8xYfg+zgFap+SFIS0RwBH0esKMr3eM1Rr9EKMEBxpCraHAa
ukAmpXw8usc1+sXdv+2edspGWmT1Dbwq5YqCt00E6eJYFkGTocoQ29c6hWpkhnd4vwY7BKv/4T/C
zJHrr62aP+bGZL6VOYZqv0TVOgJR6AN1X6LlY1fmhwbj7d4ON8Viq1i6COw+GkGu3eqScN4KkCCD
WRkHfprs3NWEyj5hL422sTfPlBpdlcKk4zyREmIszdHH7yMRKAz5EvdMIiwWTOn7JhX66jAOi8xr
9XnHJ0JnRx0tCJLOzN/JMGOb1MfEphf+DuLDWSF9+2FlK6cpDAPd4mNZppxxluDf5ixYdFb1po/n
DdvKG2l0h3ZsEWYGf9zDUqXujeyhK2IRKGjGtWRVbeb1WtwzF3rT08C3Mo4bYmQrmZ0CvhopStH8
cPKBowLMAnqeFe31ZcejzhiX/CQKyhUzif1wh7MSaCpvpGCCynRu4WDQdS6kN/r38TPWvPntjjbZ
tFv2tM2txTmoS//09iDW5SznV4dgDEP5ADugXkLp4vtXTY1AiFBuDJ/IYfunc13uggybwhS+yK8h
P2DipdFNNFHAw0uUNJZg7nPE7ig+I448cjgFnBiLgPwp3oB6oLtr+/yLpbI+pJ7CJsGxESEVKS01
6xuvJDBqvDsjTXk+cLtDLdU460R5gusowpauQLpinBQ++sUQ6oGcOTIdPmyB7p5p0XDIi5DfBsiC
nFaG1M38juPXuYye4CWpcTfFF6cPQ6zIT6GeIlzvCeEqCyT7zNgSfHfNgo7Nnl//nrgaQ0V+4cl7
1/9FCKHL8aQnw47Zm2uBmLsQVTYIZhWaPF5ZvV7H0VpMlktUcffSpKa4PMgNy49Sdr9ADK0xI0IV
32pth/hOxzJttwBMSaX2pk+AM6fZt4dHn4goxUXoYm5y6RXnc0LCwc1Df0fm4RoGI9RLwnvip19K
d/MnXwUy+0apLjMgodjdv3+l6CQ0oAHynQut1o/ZhpJS+pb4zLkhzPyt+f0N6aUYEjzGNV44w+A/
CUgyvCFOcKjdrD5mM/CcQsAyBrvVoUpnxSjGXXRI/t1MG67kB7Lw3zdsw6ezj+MPAB3WLcc0gX2S
PS2yHejG/LFSmiX247pldx79hiFlZv4GObAM/zM/KoA10L9tomcpvoXxkxY+5EE4o2aA9WriDV9x
iYPjKzsR6mTy3/4Cc1DrAPH61HrWdAzR/5lhtlH6Z574razM0jXpXpd5pzpfaml6TNXs6xg/X0Kb
rwbbWDR2l6PtQ4W6Y6Ai6ZMwpQ/blGf2z9C/qyxU2WhKAy2PG+bCWVJzqUfsUA52H0NJbzHSPc2l
gkL2RdoyfvuNErnQZ0A9yxesV2pnjMSf0AWbB2o+HiFI+OI0NVSFiy3G2+uE/MO9DtQcP9v8TGpe
9zjPfYr2uy7IrFTb5Ow7XXcMmPwT1ZF9PPmaJzQN2bxit2uNMR041pca7N5xb2e8Hp0iDan+4pBz
azhZOXZ8MU3TGdp79qVv8ofxnuKOIZ+FdUeqLEHlGUgZm6BxD1RuOl/P1iIqeF7uiNx2jeKFXfN3
SJKj6G9cJ5zOEYO+rxSsT9XguhK5QGb5ObKQ1A5JGKvmIvhsAS8nLX0EMWp2/uAvIi5nExKNuBB/
dZSJMB5EIbE6+r/MNQri4JcLstQ5vop0SyITiH0k59TISfw6iw+TbtpEJLiBthOjfrWaYpt880rA
V5ZW31ERII4g38lDol+1Y0Wb/RjOGztDuVmkPhhxICPzP0V0iD+5FwwAU7qphakLuHCAZCLWVl5+
suRfcUbeAzIM8kzkg0YWOAFdoMeTjgxhg6Z1JnrvIECgTbXKDURZ6iNmy7qvXo1nzu6iBvLD1zu+
Ap0PSUwgN94F4RfYvUsZ8eV69eI5Gl8XnoPLZk6432BccLJZOxx/h5N2SipBv8SopolU8HltLMeL
aaWTd64op05gA4P1tOeqSnqJQBZqVknix4ufr+2knWgjNJ0Misvfb7oIPabzdRFNC+uDpouUcOQI
x9RiZix8p5VWLyEYuVDzyDTGLGIvHFhzDc3HI6WtoDgBBpAkWgsXSw/567QTq4flDVHB+ntPOGIx
9qSMsyK9Ly39TVzAdsIWBKQ8bnetX3HaROjJkmHOcr+Qtpg/vaPWkzYRp+QJKwzVcljCXtNFrCsg
h2Zb/2ltoFCz/A80uENluKKZiK+7wnbROgNPhvsu7VlNuqobZUsWa49c497zBJ9zwwYxYK7gezU1
WA7BpMEAd5fCBaJb90MgNlLvmUu5y6aWN/lsG1+HRYdVZhpgreWm/r9eiVU1y9buQSULhwumShAy
aDo/OqE9l15usDMxPVGsF1yIXhBRBQQ/UfP3btnUta1HQP9umsflSkWAAIdT/Ayq3WwTnVrVKHPj
24RF7BzWYyPxAsttTYjXGEPgvJ4zC5WhlVRiHCyN/mqusHm2aL4L7HB9ELgF+fvKyZ8d9+GjMJRa
CWMQf6OdW3PGkNtmec7El5N7rryju5fvg/NphLyiJsvFbV2tzAIUnkDQ6pJHEgSUVwBV/Nh4sXsT
7w1rE3lrDR+8gfV8LOiAdmtQjuqwl/2nj3rmvrTIv099ohgu/2zPTHkl1qT627BJCQhCCzXepoxA
IMwZKV5u6m52wbeF8AONAIz9i8YKWgHVU4XJ1pjDmi/bFP6LyXDd9N2O8wlW8c9f1fY17Ypj8HUl
cqIXEDM+ieseEaNREIstQQGYBb7kNoFcEkCt9Oa9PeckF9HBt/ZEOavz1KLtxMmPp7JTs4IpQD3F
DZg9iNq0/PDgdbovSpzoKXk26d7MvsqSCb7gxA7/Uzh5Gem0oghge3bm9M07Tdy5I5bjZuTKA++L
nskZcjxo9vHe4HleiNVo5HALr4Ws4E6m4vC4gETA2rXwgErJQ7ttTsNXxNvda9ZFZSdhQ4zasO4U
0d911N67++YE5kBA27cB23AP6U0F/8ul1dfOZyPRCdfmpvI5vxE5PPnrcDtqrjpGuahyG5O6GqBe
lRaiDH7qDhxrbqdmzOMWzQ+5Am/9fixHUg7cinNebyVOM+TnYHd8U0+DOHLOz0z/OOHhbKmQ2gGk
6TQ5gorApRCZZIP8e7G2zgm5Gw+VuMQk85czgGw/E2WTXQGYp6AlxRuFyRbXTxHF7DqrftjpGN3s
1UnYBxqsCmB40Wq+U+NO3Q+c+rQUBr+70S7YqgqPs5/tbARm5YP8wNzm4Oez83IGunWsw22WUNEW
TzOgzybe0J4Czl6lKsaeIolkd/JM2keaYRUDm81Fxiy89DdLR3F4eCssRdLyLfSltAoTFwZlc4LR
sld7Do1XVAcxzGztdvo4zrevwYquyhx9+WKjzhSY9tcJTL7DnwBawrRJIrMe6/qGpQqidBTd8KJo
edhpn0aTtmlsBl07N0d782MGlf2glV7M8pVM4t6i/aZrRH5OqjGDtCSN4/ZStOCUM27i1L61X7vs
W3/4TGspvDV1T7arLu46zlW7tjwp5kJSBVLzPKhKk7rNp+dQ9IuZ4e0fos87+0utqfPUHECHi+/V
5lsVESBZeylxFEkYk1bJRRYQu52TqS7D+zDn1HZWOAS/sdFDQIwKH4aAJXDw2S/RxhJbnRFY9TeQ
zjrwiRGPqGZ8NkEhI1mZPTSK0C6HJj26/oFsZen8mglWbXMjYH/xOSwbQpQ8HK8xuMyHadEK6Oz2
ZNCdndTl0sQMCxKlApps6KZcygwRQ7C+3oZPLpjB6CEMGQkjFcfdVUqx+ATrM2/XHrwiyWnPlMv7
+3EETWQG0ZfD1o5N1z1n6Ao/BDRB7Fili3+q6sNkuvZSPlH+jwNDAZT1L/qe6vzKTcRdLQbZ7uHb
Glf3AVJwcLsBnmZiaVmjvCIMCR7XnIssxD6DPu3yDJMg7u9WiFJL0wL5r51Et3tZm4CKSmnKh4fL
H5YfRZeZcXwBRg1e08DeNcRCnQP7dYAP5g5aoipsrAvNqE+V+Npfdv0zALefmmtUJie3neYFUKiz
wy33zPnTmMNpBAWSRG3oEOALF2RzQ3ANkSqWILTc8yk5WacWIv5Qt01cTSZG5V1WWKH2rKG9/6Ma
UzAMqVU1nJdNhXPkkF3HU7uS3llCB8Iu5i/nBuMv2hWxx+AF8fxEFPbBYYg1vm87vW5g501NJAb/
LElQsG64uuudIbqe7E3AH03YC6kguazGcGgjyrFrb+RkDBHO6GwymCiUrTX7ieMFoZXRwCC6mVKF
FzKc4Jng5wIOernBG4RyWwQi2NHWrIIUk4IMpqX/vtsW7EWxYO+fWoigysp1xfG5nPywyjPDXNlO
6QJrm8WB8kuwRjCJqOq68uBL9xdvqbJWHRz/DlmKOBYDKZGWMybheR8jx1VCxz8pF3g00sG7j+dw
F9jYJOI6Nn8dqJVji84sTPLa4X2qjKKoRFuZB3zkf75mxD9o6MrXXPzkQMcWZKJAKf4vkwpDpnjT
1RKEwgSYbPCgU5sQO5o8wymI0DkksKoND8sSmrfTx//9EXhGd3VYFPX7U/rso3sLM6rmaKlXftda
ym1NvFKaWvf1iryViuKMg344SMgZWAmFzJcqszs5IVXHJ0qhCTnDMt992QFolzAXnMh1ABxDHSWG
LmTViQrgn2ACXJhVGXpz2sGlKVC8egwKTkDcDicuRGKVHA9D2KpdjPCrHK/UH+/DpXOUT78Vr8x7
452H2dmTtuo4TL4WUsoqlRyPtYb3HMMzTzwDz6M1CkRF92WVVrk2K+5OSsgsvCV9Zvo1rgrF1IMA
EDjYcYZmOqg9QOjqpPosk4yYqvhH+QToUw0Q5JshD9Lb/Z1nsTmELNxYqlsF5fEwE/AqqQ3EPYI7
PZNaK/kvcXu3oFoJboiKf0BBQai7Z+kZRpqtNR8YIw8dAD+aXXbxWNCizrj/CMEAUa9MWkkGPlkQ
EkbpMK1C0KSN/Zz+v2ypJEhmxb1tk68ZoW6FcFV2BAJznPr30Es4oOm2Ub2XLv4p2N42LNcNvdsp
CPcQm5MZJT3swjbv+tERKcfyyjTgHinp2TkAmGM5KVV+aTY6qGdcpRLxgsGi4HkwtWGUIm8rzZm6
GAYi6M7nH94Z7o060PryJlzVBSHSBwDQvdXURUw+VWdvw47t70m2NDWBbGYNHlIKaDbA+KB+SsCC
xEbqGuXYQgx28HW4F1+l20cPOHUjruCuXFo/p5XRqYO/QWtc6CcPAHYL3wdxFuxKVpdKUL0jXfxg
MTaJ7AfT3nM2IqdP1HRxh+1OqU/VEoUm3QA1k/WYYd//oPbsMqbHhVHNJAsYKKCVWFeiMssYwUBn
cdrzEdR4jjC1HoMwAYz5vSbbrdbJ0RQhdxnJ72bnze2Hj6HxiLQXmkx11b/1/9M+qITYCH2CroWv
JLqRxgntAfNo3eC80UXLqsQEw5rJwUAvWfTPe8h2eGA+mNS2D+h5w4G47Z9pqHR1Bcx2B3/v3lmk
WNfmTR1NTsdkZDDUW/tbX1aHB08n/UWS2Z8tiCQq9gD0/3A0sQvZTunxlVLjtzfXMlIHYVLCyowc
/JL7jzcrS8pVzOvrRZfgeq/1NN0MfUSMhjU+psk8YjV2Uk3D0KbHVDVghzXUJtNnm8ARzw9z0n2m
VGD2VRxaDv1KU41jXDG/6yGGt+MlIKvTpPvVvSiJTxtIQLKoB27ay+EDHkqDL4mnqKSQcAMfZyb1
2pJcSLBIOslNz4de0P5S3RFi1F2Co8ZsIRPrPTeAn76Zl+NJAfWV2400olkbt9/GoHNYiOTWSyPR
EWK5YXX7u3UfkAF+w/r/zwh2f2URWPHUYGpWi+f1T20VT3Fe1wR36VdUC9S11f/Dglvli2EX0MDg
KrJLP3TiTx6VnKmIOV/jgFFQny6yK5PKkDG39azup+MShL9q7baBPBul/7ovlhkvjgU1WgYi+Rws
QcrOnV01SO26MlTK66L5UY+Q0GpqeBY8SUYJI9ljSt4yEg0vcldHfj13LIhSuEI2BgPecAYlLVvb
3qVAqvPWgA29fbQn1No+VpHG3mu5IjxQyBf9s5L+pqdZWBT45gOFrrAj9gNNOY7n0xyfn6ZIG3uP
rvEF73PxckFSTgddQ4asNXSDJMaew67AI0iVn+scLD0xe72gT9eCs7EzkAgvwn3LldG5TDfGunJk
5GStT2SxZtykL11823uc3PtFAdkM/k/jHogNqLJS3ISiSeNk9s4Vq3bblBD3fMcVWDpPo2MaYrEs
cdKGZiAPxjJWWgUh+2YfkR8BAeZqVetnaxV6t3Jq2hc/jGWlDbTnJEvHiAsRsKXby7iQSYwjr4dU
0bHvxkR4uoNAvAH2q4oSPvpuI+P3LAfO9HE6OmsvxJorTauwOKzrT1DYbQ+8w6btcGcSUYkbj52S
EcOYHqFnA9CIhE3hj2FJG954fYUzFihkRUNb8ixD/pPXRTXD+S2h/crtOjk7AyX3AyuBr5UortF6
hOVNHMNPEe4+806Mzf/suYMlhJpAT8HEx8c+cDScq6mpHcYqS0vC4EY1wphRV3icQLWiBnP0WOuN
IGmMf5HyJ4NmIedkynoglTEuhKCdHT/ISj0ezaAvB/UqiujELtnxjtoXucIlb+SOH12WJd4ATfKl
d5YtsEeSMJyOnRro0X/eUepObr5kp8u/JcXO8FN0EQ2SKDw0kwJUaHViDmOwtKtAfMEnXEHCq53f
j9keY2NFaKF6N5+esunkK22ifyDaR7W+wh3ErDpSzFP/WgXPcfDDMj46O9K09QgvnUaAE0xs3AyR
lR4wfDMnA58dWTZr0IbiuWmsiA3X8gvmmxYMGUUN8X3Pcg+gpuBkbmIZBH1KlUCqnUJVEo5JjhhN
LtmZCrbmbhgF7bDxD6otC40bJdxbjZiOUbxJUtC9v+I4Nbv7kQMqcC1yGci2OHndDpGEmepmEqVj
cqLRXaDwdqYnVo9H9evMhEuGeJSN7QE/tahcuiZt6Bya4ZS7+gw3CR6Re5nx/XqPybaA2/1P+KyR
GKvdN1fLzR92i9ib9r1TAgWfLXWV46ZRtvG/6OcWwpiPPliM3CdYy1IN2ES/zfrxJAoIRVGoHRwE
PTHivju9tFnN9tqUYD6b6EgzZGLzTtZoiMyzW9cTlGYOYYh0T6Z7+WksiSeqgvR6xOaxZUsR1bvD
WxzeKdnhgh8Zxs1ULzsb9XdVkhAvr1sQ249D8p2gyGDtoklQe3fQYSHSJ52b+I5HYIkPqg96SNGe
79Qrbdq4eIfVBJ9bn4dIlclBJgQmyHGwBtVSIbnRksPUJoSgpA/7R3/9pvf1pIp30RhXUzrnzRY1
7gr+UhS7ZDsM/688V3DI3is5gGekUolTGKl3aGpnwb9lxlg2KCvyyjjPofQeMPte3dAAdFt5S1Qr
2lpDFJWgFJ+zzLWpv+gvGA3yyecV8ebmAOqGM6Uc3O7ZXFgyJkOQp2vJqGErMcloZyr/JbeW2nBJ
1lRbryTCgAJehfmoGhMXTw5LFYxNkhfC5mOqC5DnT2/3LSJr2s8Eg5yanl/WIgBdXmx1waF0ufEq
u4aKpG/a7CFwn6/XvSXwGuhHbL8wE6J8/tfseGz7jyoV9bL+v+GzU2FlUdi+dBV5i/tQKKa2hcxg
0eyPC7TjzvVJ/Zpf7tVWYcKbr1GRBcKpM2WjkLYp6T2tb7AXFuwwsBQK1e9VdC03G+GwtSvLmix+
tAwCbcBgTbvqZ34G3HOqelxe2ROsu7w9TTe6k5rQPxU8qm0B6cX21mawECdnqx8k5uq5Ngce7hbg
Y+bjWu0OUSjdslIzftpAHs+Fcm3gm6IbEGTcI6nHeYXDU3s+crp+NqMj1Aggfvtw5LnEUePkDyP4
X9nThzdmNq1xXqOafkMTNsVprcUzWTDxKBKMyUUR0Ws5HZwFIA5LZlER61zCQhCTbHCQu4l7UV4Q
HIM7THDME9H9vNYFfsLomC6pUOu7dctAwLhFwHuXgGS8yTZ/ehE1KLbp21qBq9g3IXOApVtbmqIm
vnRi2QNZsIAEKVpOOWWdUKyIkhqrrXUQi+W59BwY3AmjeKPRn86nwlAbyR0ju+Jc/QtSOKuTI94W
MQ86romasvzHW1DMfFtxAbxxiAc/sJylYd3sDgb1+csFQ61s2DGE9OxDUIKS9Rg3l3t7aXoJ1l4N
xCWWhdjT/FuiQvpPVWlUaprILadZsstYdnXj0bmuYSffAmoR1JZ2PEK4y6XrPcCs44zlgthQgLpt
LJS2Ur//aHbos1Zzvcs5ce+SUx0N7RJmQUfsqhaPhWTr6HvcYkGuWP2o7Gk4Z7ZHzTi39K5Xmd8p
nab544SKsbo2LJe3Circ7XbenP/6ouWpXMah2xoXmK0dW0Qwoewklt4uX4+1rTlhT28wm5heUYXx
P2p0uUZmlwDl/TBb1Uh26J2YZkY37ir6WVxSuULaMNDbCDOAjKtz+hQab7UsrvybWC0zwo4w5JjQ
JHSWM75OwKnyw1osxTRQCEcM/SLCNtma5vVXQcWTtcqXn/MAeM7gLDtDKRutJQxmeYXrBYJ3be+d
QKQ6hfglFT2gOdmPJx7Iau1lgd/xYH2uGfj8ESjmrtG12PGcU+vW7vTvocfJaTnlhVG/UDI6gx2Z
hxJzubhP8LpYlIw2J+RkyCaf1PWA46dzvf/0pIfRHxqTSG80llSOXaAJHfMMgEnpWxptbxPvALfJ
jopO3Wb/7qWhJTSdJhh7CtaGx5j88dGFTH8+gSa1DsKlHJpTDEZRHZPs3jsH/J9GymIVFq8Ylj6L
LZMS7Dx8FNT7eeh/nHfOfj53f+avvTOQ9wqPRJYT/bHXhJJben6d4iCLIOQlVLS4Opzjip653JK7
WQt3H5ILLqXr//XRQXFnSuxH+znTEmHnw9PwgRU6yR13U8w8846PGliMRW9F9ePR9jumR66hdb+V
m6O3uJOhZ1qp8x5MmO+KyS1MhrUoAZoPOC1NgksGCUAN9u2dfjqHyjuAwxLgz29adyx84oyQUmD+
WdJRlCVOKh1ngA3d899fd3BiTfmFpMPozPHxrSSzI3pCeFopBHnp0KMNQjgr8+JOH8E9tIh15jc4
f82HRoGt9+TgMJOJ1TGdQfLPLitf3cJ2K3RN3LqJvdS5Vg6Q9fGooGcJ1i1Xhybox7SCjU3sF6O3
Twboc1gdQskftpbRqs3ph8843gbTsiFy5bDQv2SY7tgAhSiY9/qfrtufxtR+jJnsUhNSLclKikji
71yXgMP/Opk3uUi+x2HPnIm09WgALpAOBqoVTsZNuuAfCqvn+KrpwK5xJKpHgpl3z75J8lKrXyLK
z5bwOHlzGg7wR2F7p8vK9ClqH9UMlVnrgQSSb91VsZjmS+dDCDw2Y+wvLzfIiP5nEoLbSSi7Ch3d
l7ArfLEKdQLp+KSGdBLd8At3/wh20B2ixs3xZ6VJ/0gKk7c27tkzK1NykjaOA736n3Un+TXWQim8
wOudQnWQv/8SNGjEUBLzBry09g45bOhqScIizEQdhGhFB172HhQZ9yd8cuylF5mDUTs7nw91OebA
XCGYYtnvKdPz/6ytFYvxZaJUmdxSpU8JWVoMNzAH3XGswzHVA1moF7C7Em7BzfdpvlaEJmVe1CX3
PC2wqNzvA2+a/HaWZxSGwTH4H1D4wEWEjhRfxmk0xA3Fy7eoglVgnQaTvqRShk4CbuUWUAXFfAGA
4jk0K6g+MGmocR98nsEu+77ip1xj6uJBQ/Ay8jzijMjY5IEcluP+2IsnjYxonKURMCNIEtV1pwKy
Z+5hOaKrb+I0B7Y6pDCRtGKP9PV5w9TOeBsOzSPjS77UC00/GKn/l2TVyNWcWKNl/gb8VFz1ieFM
IbnT3UkN8bIlRpzcwyoPlDI+cOpA9xMiuKFIddO9PMMnKbe1y0p6Ll+oUzdpIcd3z8rP6x7RNXpC
G38Lc0TlaGFlemGMVMlSyvo+A4Wy9dmIebI6du96yekvgUOWlsfvsOddc4+rO7YYQrXBmKF0GAUS
tWp3wq77wNg2ZPN6bxh4Mkk6NPOCoApFUJvYT8LyfmxrysdyzcVG5osaA6J4JLBr3lXR/XQLWF9b
CfVAp1lgjrQwikGa2R53kEfZ++tkCjT9iS87Wk0dd5KXqWJPDukKregnPqLiKgorrDiDTrPZYL9c
SVpCd4Jcmf7SsyvTRsfJB4CD2VZZAufj8xMYTrlOr2xFExQmKZqo4OTA5AGE/7ZtBWG+wjXo8Tpb
q95OeSxFJR7TcXkn/GBTf4/wJfxl/4IHkvBFUNbSD4dMweycAiWKTRmQfE1ec4KvRupn4vYtjHFb
Ix6IvEZ4gVhUfmTcfwKO9YbYPo+eeZDedopY7p3dDDkchtYpWyCyFDTQ4HbmgqiKXnjJRGidVmjC
qIL5wmRn6wsXFKFVax8MFdVM1UPcA2StuneB6sbGeyHAs3QjugaSJWeI41w8u90BNG0MjTxY+fm5
rKqszo7OYS5lP2n8MwWkElHRUzv9dY/GUTP7VE5LFojVaVfoSbHachR5GuhP1CsNgKvIzdoJKV9m
lJ0J9cmhuE283SjR2TKVLt8Q8sQeBdE4e+lAflv9Y4xTyGZ9+RXG7avyKKiPmwtqh2Mjs5Avo1o8
HECUoTDO98twOjrsEpAkp/D4/M6VafeOB6ioQaehMJJrFHlnXws5puIWI9h2lQYgq5BP/Ok7wcG5
lLvrrhT7/afruSZKSe7YPazE1vlP5OUb+Qh+3yXiZxFMBsgz4KTF8NltoAp5xAQio1Lfoed8r+xt
aXczVWcT8mlrr1BxfxlrzUNEKNhfT1TLSCfeO11/KHaLBvu3YBBF1vY6lgTbyyzdiPxpUbeGnmnZ
0/tYDEdlquPMHG7KHY2ZtfUY7wK3vLgwbE94SBNT6552TOfTiy5NZPT24+LBaNsDrzJhRGNTP+ES
Cae9zjP2/sTWVbpSIaqxDA3YeFCWMtY/s0i0ElqivYu6zJY91TzDDWFKXIrfaAjBmGGor63EFVZU
BOX9OXSjy2OZ7npdlkPBiBOFdLeJ6XGeUgexxTnjuzP6OAlDf3Ov/nzq3zvY1Z/Oq8YtDU63lOwb
Hox581TbX2sYZQSPduZ5afGELYgQVPwJny2kBqg1AnVRHzdgmbw0bDuo2SWei05D67wQaeTeKM5N
/vKpA8EX7kJYTDZ4vAoHsWoO76dNwDGfeKg8buS70DEIcYHz4cGGFx082KSvfuxUm4C/EWrYmE4b
3bv0BoYMa3RJWiU8YBPOKfzlJnzQ67JVOo8INtMomXzktXLVgbuwaN7a97MvyTxQrCPB7UzPAzYP
KCpCRjsyxNR90yFwvD9MGGsEWNsOaLx3nfxLkUxxTMHg7QLiRxwTmEJCuerEpBOtYvXNH0X2NUrQ
EVdqHV2FThCMVRhNBUv6VEXNI+HkW5lqsWma4LiVkGZ9bIyHAMd4JmoxCB4Pldzf8Vzpq7T8HLd7
/Az1OGDwG7X6VI60DudT4Obch7nMJlKhXgrZm2woeDWlaCT/9DGuYIWNoNir5+PqafhlfhFB9+Pk
iGSOhqW7uP3fjZNcfGvTTPVwbBTTXQ7T1XlYQXC0pWJZZveTJTtkGEdexfbILn2plEQHc3FTTWv8
i81gicA9E3aKWtTkCgBwctgFcIqnc+oFVFR2JZCGf2Vyxeg5+3z1/D+U3L5jFE+UhO8vU631AaNS
M3ksVYLCz/S/dHW5jk72JWUGFPqOv426Kvjsx8oltuCb9pgPHSu/kfd1hjHGeaeGvA13YrBIQ3Ma
yA61420sOtS43S4I+r9Dg2jUZMMepCEenAdk/0TtRj0AhuvXQ5nTtZEGCo0Y1anze7g1yMo/WVrQ
8C1VwXS8dKmEjxaEzKRGgsqH0arfjA5N67QZQTk48dGpMKkRaqNzoOnWQ82fgz0o5OzCEjVr6MiB
YsZANF+pt0rJOx7PsTOBjExYUNDaPGHv12ZkgqVZCSNQeW5OKlF6Mu48MwCM9LgTIuN447dtD02o
+OoiDCKfcZA5r3o08RN4m3VDb9yRnilCxEXFJsfgxRxg2NzIGyUJnyh2tFnmTdBymMeeueKZVkqb
CPFlDGaobtqXWHOHlKrmdl5JNmI1M24QJ7kUzDmzO4NqM3cJMkBrERNH5CLlXkTfa1FBjXCItyl4
JOf+SjOJDRhXzA6R/EAu/trBfCGPfybxtUdGoFCtaBHkEzqc8RE3ael1Jc6waINm3wdhBCLw4wSN
tZq+9kz4M1WGbSWH3At3A+1gg6fyjrxiThm1tNU2/RzVv+9RvKaFyfZ/LN6uPXxjLwuHR5JxdpPx
bfoeCeW8mUEvjtjNI5rltJD0ZGbCo4X01dZyYOYR5JNpBdKdE+dfVV8rRK8Fsbjj+eGUK2skxdi9
a1jgEN2B2kpnSwo6Rdoiq91i4zjMtsE+vbXMRl8vIo74qG8EOK1XKk0ai7GO9b42szuVzUYFQxgY
9lB8KT3ccY+Db/CI7A2VdAN6ui522/u9fzPTg/mpIuj5xoqEjZwwuYvu4CZmCbpfI3ijbYiBiocH
nNXhQiMfkz9uPwK2eRKwt4NrjasMXWcswFcrzbVPdWY6UsImuEZiHXT0UreUsFI7Vqxoutqe7xFT
jZ47VStI+hU/RTx1e5vilyQQQvKrCeP+/EGlp6FLVOadJ0V45JgMlnrV+tRo+nS0O5APc48dntBS
9j0grKhh7COp975xH3Yp4ReMkcjedDp2FrtIzHbclB5NlZDryw+NU3+cRQCJOEK1RVsLY7OrRuGP
AEF+nhxo1KoCy3gGpJd2YtAx6jsgyuD6Plj88dRunk97GWIQaFqC5H/hV36ryN4f4NpKrVnss/CR
jOPFPhIOF+SXjwsXHAZy956Hjok5He5nLVsGhq8pqHj5BrB6v2pzqrQP0gJ8iLxs8tCXeMH/M5e0
E5ycW54+Zbl2ucnYptCYXv6nhzOUVMHz2oakDlrl8CjnuBedFxcAsohD374LR49A6p1xWa0NMfkz
LdJHElSusrKHZlkqLFoJM65qc/LZ37lvsKRr5Lcj9Yf0RF4lWZzPTcnfcg1RERwXhNAqC32NkRwz
zfbEEu4sJOJ7GP27EMlLuCLMecQYpKzkVp3DIIhUYr+jMhjFn0BzGttwmrEwrDRxWoivQ3Ftyjib
clSaXXl+5rGXlrJHQ2bi/tCjph4AJJdw7P+OokOyyDxxBCTCGBczP30fi1K9EGhcN2N0kiyZkLtj
M3vZLRTgbxXUGlHZ7F0x+7RNjO7UZRQZbiW5MFF7GEGUeTejqKq5nHe/8Plh3+HRxq5Ok8ygNrg2
M45Dyi8yRJyRMOLGvC9Sd26mbn2Dct3V119vA0N60lzPBtcJ9bJzTH4Yo2/qk/SOuuzRMbuoMrFQ
wRV76TR4VwZlXZbZMN4VE2P/nyIxUVxNY5IASgkNSly7oC36asrsPdC4Vaaw0IQQ1MA1PCtvhzhR
eGjWv7++DdcfgK8AozD87hsPMmKsJoEHDlMAPPUYGU/HESQF2VgiWBjAHPNAymrSk5nEta7rmIex
iex47bMpCYIlEvdU4est77E1bA7dWI77xLo34xfOUbIjuSZa5sYec6YC74dWUsmuYa03P/leAXIT
CqSTtzaFP9p41uc8OiF4NL+ysc8Xrk6u+sziutc9GTvc1TnhWce3YoSHT2KxoSDtvKxxTcELe4Tp
zVF2p6OhUrSIFz8Yqrjj/uKDSTQBF8byn21NUPfDMZjPqfnZHKbe4ByLi4ShSdGRtYRHYUCrGcUT
HnORxQEP7ZuQO+kCja+k4s7beU608KuuAln1X5QoVTpx3QdsLj9GKmsbm4hpAnPuBjFAZeERGaS0
H3fkJNb1XeYuw9IIv3Nwya1jOpVoWp0KrfmMFa3b3wXlqjBxceDQReeqsT9dXBMfx6W6OBRpmdj9
UvckoB4I3/n6WdxGlxLuH4kmkALqfKKe+2vDyy4N9n/3YnQI80x+ZBr1B7gGUol147JIScwFbhIA
83PPqC/fkdDyxQU+rbllbFkw0LqpK2QJJksduIbup4SwVEqK5n6u5pABv7gLR+aLB7CcSjWsINng
amUs8W4KEFSv39WijqZkenQvebKrOx7NnVyEQEf+a1hySnpUiHJeVfsn91yx+gVhNpP5MZyNlL0i
a/wIdJ3KmnXYhNPmPaQgRfeVA1887oS6wLPHiULHJOx23eZ0jjJZ9MBDXqKhZYZZ0jDlxvdc2JkB
7HAKIh0IAVg7LOm+EoRTl7tQxcYherRBkBwh5uOdL7z5AAFjFTRr03WP1Jfv2GlxSqNMYU//A47N
akhmy73KcU1vPiFe3pBBOVUHjwVxZzgR8WMjoR0wwmFF0zQ1MPdckHuupMtyYpsTiVB934yhw5pe
5HwRLrOC9cWWDGyF9GIZrLQGAyP6S4h9orUprkXYiEqbCB+WxlFXfrVd++OpxBxwqNyccvGzmoNF
EXaY4G1A06YiQ+M7Di3h9SwNJaMZii73nn/QGUKkQBYdmYXqnSUI7mEvKdjk09KaU1Dn16mn9Jpn
dsnrMPL15sJwt33CAVv9dexFYeyDsTb4pD4lZ3XqgE7VzoXeSXE5ydQiy0AQSVKq8IP9jGW80a9J
TZeCMFM7dWKE7IVN0N3Ofp2iu8l5d4dF6AVdhWOtYpWb0LUdxUbeNZZQ24x+9VdbGiOa3bHEGhiG
7s6tiBliz2Aqmr8ns71aujox9FXljOouPWXvLV32xH3XccmjYDVWm+hvQpJNb2jcO+owUosmaUI2
nQhkHtC9WyOgePN+ziRWdmWjuIDyZa4uVfQauGpsSq9thI8rQynghSVvN1B58qLfL67d8KhDAlUb
HTT7Np5UVIRYG568VLl4uZhMNA09nQzaDCW1IfeXv+JHpqJUC+jD1h4Ds5pl2AsjAS9kpMt9FXHM
x8jWplAnBN6r0wPFlYjQa87WZkUds7Hkxb36Gd1OFbpMi9znx/XrM8acV656ZCoftVZkeG9vYFeR
LIQT0ylhkjbd+HGErdFrV2odZRvAHj+FEKT2bJnttnWNkWHZ10FsfkdJvVg64bLn2TXwpvu81gni
Jz92wuAn34bqW9ZKkeg52BsyexNH0LZp5tXUvOfZAoPemXWdx+ciqoMY7/1NvFOgJFRWhPA/R6Y9
mYsVx+YG6izQGgof6mKI9OKUavkXcIR7j0GHXh5aiSzEQUzeyDnioaA67WwewIwk+5bEW8UNJ37Z
0zk+wD0mCc8kUCijvi9iOwR/QUULcpHXLp0IQXJNjAHlpPYTYv/5o1EESBTPn3vVely9vR5+lQSh
IfIVpd7FFkQXeno9VD+BOwKZNBR2aQKdteOpVfCqIUauN+/a/ihlVtYKn2dXg3AqB/OFldqbplxu
xbmH8G2n1TQHqAlmWkKj8v6jeLw4NuWhDoURg0V6w1zguII0je1feLJSKT0yiNaifrZjCpfUmaFK
e3xHhUNIc19gTvUfliFfFpQl7b5fdbM5hEfAEJnN1xzI9j5m1dt0LxSDgUDkuVeuaSZhyNML2+K/
XelVZgSimzwDHvLowNoc81N+xRudgLZmiTGhYbd4t96Orc/bNEypX9LK8ezDn9IPkuccetzQI3/v
AO33c7EoOmNxfiYPL1TMGr1rn1B5SzMt+ukDhF2L9t6KjpXG3Jxi8qE/eTijXGiXMwsOpSYCDwsi
CS4iHGal0tac8aqAlpPMM4et6+Bu7mY/T+JkHlPa3wF4kcYwm2iDr2gqSftyu+TouFKQn0MzuaA7
AhtU63LYI2886CsNPtWk+IHSEg15eGZ4hXbfiEcdSozai34ADYIqY8t3dR6RdvYbXPOIwgT4udpL
jhDRvzezfytB1NkmtjjsTDysVM6GSlylulOygPZfiA0b60seow+vFuXaAVoErGzfTVCFvv5jPgyi
mn641vyTWs5MUG3tQ33jDTtFIwi5OVPMH/C4OtF5isY2Fhcg4RWz770FXh9PzC90Py7PfNOWjDXJ
TbH9cGJ7frqdfyDQKTdmIDVCR94Y9R//1RyN/0P/JEi1AZ6xQ3fxbPa67QN2l93XKpkTCdb7qps7
80bGt2IRGvwpoiZvMH0IeUaAR9JEBwnmnguUA53ckN29aLPE/uR5cwcUeNhUo2V3nlv/WENq0hVo
qrCpqby+DCv/MIFwfWSHjdUKAbmSrjPIdNZoGHLljxBJeXSayiT8RBTKLOvCFiAKL1m5Xsm410gy
P6BGUwALDqB7TPnN4QF+eN7mLIPJyVvobO5zi93iXf1875FTEcEGPpSuswVKgjQgjmvFMDeURerd
x6FKM1WSNfzrPsPtTA6l5k7RKUPOgI6AiLGOs0tZwKO1LQx984MrV8eriktleXcdftM1t+mXgm2g
DRRKmZZgUjaH8pV+qD+dviAUlBYUGJBqKXPEY3P7Myj5sAP/oHDgKsdKnL3vWMhfI+DKgq/yN6TA
fM2w7IrX9h1l/CgYRKl3iogS41MkKYtrGMkWatT/xI+00CEH+6JQXpDJx2cCLIW8abwoL21fgXFH
dYHcvmIzx+gCqdbdwjOSRRw6t7dft7Cp7yVAbI5LcHDgEcwaYOVdMrJg55Q/NmgjLszs8v2gOjnH
6CyLJNEgKtzYT6ptGluByQvJlS364SC6XSUy2iX9G1fCUk6FLK2J+LlE/pRXpyc7JPtL3H+KC/9q
Axjv95TRyQE2BxjBDQpsjZBRw4Cfn/B5TcIdZyCkFcLxqhCVOAMPSq/h3M1zD2yewUEvjc0FqGrr
VIzIbSq0EfUeqScvRdPoEmeuIjJMUYZEMIqwWTP29CSnKWYyJDyTD3W4qn0dWNEVrYLw33NxlecF
FCDxuFM7kH6qyF384qQ+IOFzwsImiBFTMH2CzJhJF9muzoqm3dXYDwMdYCg0lSfrojMbfHr6Q6N/
lSFDG1nYzHgkVPrmeS914UM4sEVFuuhStBYS9a5GASfHIY8fdWFaDK5D/rv+VlEGVo0deBuX02ql
GesQMmJoTPdeVIy4lajkFbPicNcb9I+prHQZ1cgxeGt+KQvvPK+jiu/ZVht74BCTeqrK872L8BdX
5K3SbQ+LzSJzVtuqcGGvOM6gbddeKRNhw413/y2GKGStZmhWBgImJ+2Rv32M2uGOymsqRavd67Gg
VYinhs3oi9JdBRbtbXmI6OkcSbvpdSAqJiDklG2H9ZgV1XEcIm0YfVYnwnSG1df6K1oRmFejZcQl
QN0LMmBs/iYgRGSPPThUNxVysGAIpH7EZRbV8k0CwO/iUB+EH71m4UcLBELgOEKgRF70RdeDkmB6
fOIcIuxco7KIMWJgx20mvUHYQ2oDw7RWCIIANVdskp7rTPh220EatnsjbRKKR8Gw6dj6SYKVVQ14
GC4zd9BRv1ZQBrGSSf4FudLFV0GsxRB9kswFPWIaTo2TaoBxsCYzO4/ERNCTr9oMa6LUutoLgnVo
g6POh4W0m3UIk6+Jlgjh/47DjgvmlXFSsGiyc363ZRHlfaIjxEGjCwLxKulHT9N1rYjaPvfS+WhF
eeBEXaGsxdsByUX/ZgnPdyb6g4MZDKvjZ+Wsh2eBHuW+dImvIFjcXfTFiyYJLg4n07k4g5Uteqtw
W/byPpSPEZJjJY+X1bBOrI/IX4ci+IXFwVGHkHNZx22HyFZVSp2+rBLA2lloq0xeC/wqqgGyz4Aw
fHj7MCPc6TvLMCvA5aKVaraQxW6wpqydIe8Q+fo4uF1cYKHgN8AjWoxmbflbBwInt4QCMuQFdz4f
rKeu72/rgD/+SEVKQymIkaCvwX/8nZ0U1o2oGt5V/v+FdjsPSlDGU4QMoDTNvnPV/FNjOrDP54ZS
hFUI/CjaN/MynwgdSeuIMfE6LOGeW7pCVaGWl0Q2o5s/Jawygtdzk1JDMSmJr3iuNSRRH7HDDAHt
Mf38QqPCqF+oO/Y9WZsvdxy+QdpGZnuITIddVtl+9nig15Vtk06PriqgXvdH9O7WYWeZIm4Fekne
+pYzFbQDMbDIop/ArwNYbn1906x9knM4o6r4hEFu8m3cnp4m8ZiYe7XYS1/xvVg9/vVggRrzrX2I
tNMoK8ymXtrnA6OaKziR99gFCYQbYGrcKpsuAlHZadOfXWAK9Zf8cpbRf6z4BVU6VQmnesVRGR3n
U+tj0K9gLVXiisI3gF5e6bF9tuvsy5/8LaUWf1uBdQsjekbJNGhL34H0tEQE8vDngXiOWXW9xb2I
OScE0n1BcyE4kHkeheC1boqfhyNJ/MR94Zd9FoYYFOJSlBXPhHhuUuxsZNIhPCXyzXV6VNqwcOQO
d6fNx6W3rAIZ6EKHw99ebwcW5/OLtncwY9zdGCqD4dI2oSQWXxrzZx829LxuToonKuAE3sz+BER4
9dBcpJ9koKbwIvHEigvxW3sRTWq3C33oQrqtPls9aYigNM9AMQbmB2xb/ZoekXKyS5pSJzSX8eX0
jMJmyj6gVMtMSHoGbCi/KWLJFjaQyZjwG+PVLjL9lhkVsISJ5QBEI3TmOQqscF/kdfz9tLp42ya3
L1AcK9XMkr0/WexaU70Zk/M6nG9fhhj3HzEmSoZVrE5yQgyIQROdsMuJJwJDU60syUOVripuI8l/
ohePIxwmADRSvCpULDCH0tkoO2Md7FK+mFoBFHnodH19vdshFlm3xVqPVyRAvZgSCIBIQ1Yoipnv
Iehb35VQJq+8sqepxHGUqxdBPN6Xqw2HIiQiXEPjYznVLTvP2tlomhYFKYEkxyenXZE8OruSUTiw
qAQpwmncHfqBfBy/Fa3i4eAfKtgOzqAl6eJaRPxb3clcADakRwCgZQxlgW3YFYwzrEqq13Ki79pm
tf1lKXBVHpkiptQ4XbAYU64CzhNF/aPTLy+99ila5JKSAwm/HjAKTZIR4d/ySkMX8wij5XKQ8yeP
g3wr8WVQRQXkOKMcpLqhFV6R5aDIu47qZ/W+TCp0669+R56xEbU0leKBiGO0WpJEmaq5IMeaF2BW
/ReLEp9kt+w78dPp4kV+YzdeU8YQsAP6SvWTNPcQ+WQBv0XCZmz9QSHh1x0E+fOsXMvy1tzYuxjb
Jwcnm19b3uJHKTO5bsU/7cEYfZzG5ryBfPowEkJ+PXwDcQxrrMXPfH6ydoD2LZnzEtNItrUdreYQ
yMMXsPoE5EPzdXWBq+hasXm58jGwNcYT7+nSmUrV5kWXB8T1l0np7OvO05eiEoOfoL66+/knK/cz
/1hkO4M4p/Z0EBUeDJppbaKZReWsSvrI1GAYCD/le80eBEj0L87WRFXp0CHkOGfonS0YBf5v/3P6
2UvvuCj3aFqFFiN3g8AJel0+GUKa6Mq+9cmf3Z0PawrHp5FVuCD8CRAAsm0oRlmkLVrND81IeXYj
WH1XFZ0h/wVdDJ+TqzwTgmMzSNII9zdmqd+WsR4rgLS7hEMD7UfEG0ia8DfL/s5if7L2xq5DyQ6h
rBi+VQiKNQJj9sLepH8v9s4e7ngZ/yzZZNkUIecAHN/J2bq65kLeEpDfB398iJzkdFihqV/7P9Hs
kKGtyYEKX8cLKfbifF7IMIiVnwRkhzMQzayarN2vAlA/mKq3JySFGYveSWu3VAleFyYc3yUUaDBq
EJ4Hoh+R7ZDDrKcGKtVjnJKYDdE3/zRAtvw/r2tqjyZUXqjuS3oYj96E6Hgr9SUnQAcgl9S5DX2o
GgOcXx+diz0bEkDSXeplSoqBYQgnJYiEmq+EKZYjOYKOc/zUz+ukDuxWjxK2gm4EYi7RIYUDxVeq
3JjvNmwArTxR6MEHEZZ9gbbK0JFCLC9cFq+6qKNawEjSxI8TVQv6VBNIT6TEkBjISIg0EsRT216O
tp2BGcvC+DxD0HUyQ4GaSc39Z7m8/nTaK0kBEW0u8o/ReflQHicF7J9DzisKBBw5Pm4JIyXpRfHB
HUA3ICJsz/DmXO9aupdOZxOeP08ETR0XxmEEqlxRoAy4johTF1Rn6dAWMTtkZy1i6k/P+q8mkjzK
xk0eBXRtP1pwPI+sXN7Cukw6w96veLeyBI/4FDDEvCZvRK9PFCUcrKZhg0GFVyO00YHHfFeWY8d/
g5c5ie1DWUqKrstR12U3V1wIsbWLuavsAsOZ3DTvxDUvQqqIdYYQXVzUYJb1vM9nYS2aNzNlArrd
3COLSWQqTcHATGHYk1IoIrnOY2191X6XEMfeaYA2b+z27wne0FO4V7ELTuZqpKF+AGz9vE38CKIh
tQg4YAIRTuHWZQpjandptO4eVPLA+2NPxhe24gdqHag/mu/4EcOkSvPYxBVVFmuE84sYBnLzHC02
temHgaHisoo6uhi9gDanFiahyAFA2grqy1F88tz9SAvFw41sIWB/WznmYQpRStXh+V4ETFEiLkuz
bEGxQVa8Iv23uhsuzb2HCZHLSKOJ4JiR176j+PgVzchuS/IdaBuAf8eAL4ChRB6WouVN6EaJRybd
HTB8cMtAWmQvNzAMRnP23xi+CHHIln61caSrWWDMJi1zwRGjp0IOM/7qPhfCir6n2riYsIzbCdOs
A311CUebHwVCwslLQzi9W6+aqlm+b0qI3vjmm98CTZKDP4MvzZjycdtdaFz/tMORJJ5l0zBuT9gY
2UTxILi/MigQPqUE18rLz8AZBtqaWh+V4A5iPzB5TGzqgZpxFyBojfw6HnanuJViPSbCLoE299ZN
6EQLhM7JEW52xU6qsAH/T0+0JNTcwTTTWqa3HCtmLoo0VNhAXCeFSnVxnvIPrEdbGLXYw4zOo/GF
qif6HUTkfwuCFsDpqSUaXWSuHUeB5hfoW1Ttr3v4g5g3ocqV800e+KAk9aACeGC0HfY9NcaGv+23
YgDr5C5+OUt5KAULBLJ95aVoM+DJhOo4Ot7Kw0twZV+biQDdEIJSaOM8nR6tAm+r3hpZVqnZ+88X
k9xLybY9nmbQytgj2e8wMEb3NMLz8hgV/bVGpgFsO2XJrzQP8M24f2R2GDolHdExj0Vt1cfM4ayn
dXE5ZsRKe+MnhAeCf7hWLhR98D1cy1FTiC1UaoIMc4YBvIv9fLuK7M4hlBWGVMEMhQUkCOexKXMx
dwbQ4tugI227xw8LzorS/EHXI9/AgD9bPdfko+dph02wlwlkjRAMC7HdhDmmGWv7arIEi9QMJZDI
fom0LAr0xCt3S6gtz1PB2QmJDUJpyqqvHkrzOaZu0J/lGozNH5j1QaXObpfY/3D2Eo2URdMm0G+C
mU/cEqYjkuGq5XiRN6hqDSu4vWoYjjR8bnheS7fbUJzhz4unuGT8K+dS02uurLJBXAGnOhzMK+Th
82YG2g0xl4zLZ65zZX5TNqbMIjELBshq0KTdmpN37GQbt3JHqBxhcC3wNphu2iBB85j0c7l5CAWq
ADQWLEkbx85veYBW/YVsplVyhBOKgrzt9XTkk4qGCH6tMZXWjfDha1PKpgULE58T9ZT4HU8xxLI4
Uc+iZc4er2RX5nzjbijyIlqGqjKwxYvMMYxgZ4vUvRUuLZBrhfIwS16ZFFWzz8jptX4TwG6sDbFi
pQvIM0ztPdn1ohu8wHOQfi6Lo5TLaqKYckq8RDnXTejmtzk7cZgvr+H6XB/2LmSeFpkE/LUjQLZ2
n9d2XiGd2KQmA1vHbFMONa5HMyt87PyCAYx5aLxS3G5w32XK0iXKcdVYZ1/CHnYCZYRftkuUuH7e
B1378l1h+/yc0qbUTjV1kYdGWa6dt+6hSOj2bNxmVylWZKfasMqjI2wJoToQC1/kFJA3krbXmPna
9kk1q4mP/bk/I4t+3uPZDFFktppfnyCXyTuk7j3m2u0n8CogHcOLuwEHidq3aor7SmCfJywzeJLc
Qwg22U/ph0gxzuSwCv3e8MTSbAGkqoK4v7hWDlUcr+uFbFx4dUgVECT8IoVLoumaxm7dW9jrPrMJ
2I19Lf9AMRp6IAIErBwZykZxOjK8aU18N/D2xTHtIfYHkOLtNk3ZNeOzaY3FzCewQYiMAuyguEIk
ojNvn25SbiBL9xaCxIvLcdfs4Jej9JxzeAv/WgelvokRIkDjRBgG4A+AFdNT8HjoQH4VSNH2EuLy
AsmcBLJ2QqkUfxXWts/GgdcI8/JOdU0nk38lnKReMUDl0WUZdX1YN3nUUVP186zxXJMw2NKO7xPq
71a4kgWmG0mxMedvcPP9viGaPhVKpmNMSTwuViIjoGzqET/TamW2y73FxEgrmXy0dm7pk6/QQ4eJ
ZbFI1hKhsetokk8N0lrsjvRZWxSpAOlpQjJh/T4NZaw8eqRScLKpQ3Ul0kMIUUmdgiSsreHoVeou
FrEnI27htMPjPmq6BNoIBFMh+10s75PiD6dlQBXfr5wSOYlxtSkA8lu1fk8KFBCeU7t47YMhtL/l
RxhO9b52nVda2XzEoB14pOXF8ygb9/m3kqwUJspqLjlr05Rfcl7QnN+n+lFqK6IIywTXix3aYiv7
8bvL/jx9//iJ2NRpco2f7dOGi/z3Ty8IO8CjyGT3WyybtyMuIqUjxsxbPZXX5NWDG9Rykkai/W9O
QEkZhRGtfUyGbKFwNMgRB8/XeDEkCVqe7CwR0CGGRq/gZqXP65uzQ01MgO8+XK81P/EfpwH76EDp
FMqjGx2vNVGuZiI7OTUaavlDsw37O3cDfkiH3cL4CHZPYSLCpgY8TnLDVTqlXjA2q1mgiiJ34gxW
KtyXXw1IRkLJJh1avC46Nh4dDH7k6q/U0Gir3+s2CBapxwTvZi5TvRx+Tf7bBBudVhURUsRlXvRQ
1oyg7O9MTF2M90V1Qw+XeC+8KgAGbOY6O8qFwlig8cj4bfuLX56wKVLz4CPQPNChw5x66dHrIHrJ
N33dVc+5DWVezqhILbEs9+S9jvNl/txzUbhlNpn+FVx/zaqHSYvSZRudka+/Yf14+COh2roehCEk
VXHwZ2DEVbKvYI/Q1CTSkizZ3lF7v6WSklnF7Ax72j4JnXrmiyIP7pLGX9obaeIXtXrNd7cRrDm1
o7/2LSXPRBmOZqtXPqWdfwScEhJYjyyAIvrSm+Dksaxwd8wq9zm20Vul68Gxsiet5dmOUvbFoztp
LDh/kvd/3gC/7GLEnR/K+BEytvNX8jy8/vqv0nKMIi9oRIx7oLsXR0l0kRl1ohuo75su70rdbOOy
Bv6aUPPShnozILOSBX3hOBIBgnv1UK6UYFJtomYE8OfQNOSRYKLJGhA7oqqBHCaflofPA6Rsnz/M
yhZ5xjY9qZXiQqXPqgdy4rt1v8VvbCzrtxCNoQl+MxlvvDbKYVv8spCQ9p4aJlZ4rQEmdLefBCJm
FEqgjQppFmeih5G0mRbXnPDlONySq5K5suVBV70XWYIGd+rFQytSLYSW11OGzN87uQLPK62JfdO/
j4r0lzOR8VoNrtabMsir7Rv6Yd43AAwLbkPqLyOEAQyC5ZwhZRHLSXs8ASCrKTduSvYAtncDaQUR
B/ZXHBKyf1n3xPolOmEo/tj4x/TFqFRV/XLQYoXpU0sBR+ai62IUiBORF2HNaW/QCPlet5cuVdhI
BBGiiTzYOD7w5jTWfBjMnvbqbiL/hnYBV5M4WXiBdV82r5UCGJUGvOEsQ1hOZ6PTmcR4nNHtezEv
l5Z9yngQZFjSSkYF6EzQJNz3qzYUJhVX9v0iOeZ2ntudd9yBDIC2Jav+XdodxDAAeQNfWKx1nq6t
V6H+R792d/JQtr09kep2OAxvcqFf6RKpBGSlpT2N1J6R3ohgHULQa8hfhNlKs9YvclP3ybzSPMZm
8kBrFgwhGym8525iymIYTat2ldEd/LhSa8GOvVAafMvcyL6yXSYu8rye8bhD86rboIAbiibdoZd7
9xj1kLkl/fb2qXzn0cmTguMxBk2oud6Z/tqAiE5efyk+CNJFkl4EwaFLApRQBnEODJmMSAzc0i9M
0TiNkmbb53W5qHEsTsgzTGMBeE45+N6nnVuduLcv01vtS30PjuXXw9Rv6SM03l6M1lGTwOY8mdwV
s/xdQi2xNdhHqmA0KQT0uy/XWuTv3vQmtA4rsCK3AQIs7MDTsoSKpT3t4cSDuj11ph5xxnRqGjsV
F2+2iGYXUtiP7ltmpxOzGo0+dtgOQx5ufxG5AgmjCx3Q16TBznhstpFRUKihc0s7QiyGMOxsfwt5
2P+EH4RmSQUHvda4FBfkKYfymGGuFXq6wSah+mbOlmUK+KIk5+YG+SN7e5UO/w0RvwDhReI/tgfz
1pOXO14ReYGYpAJqgokgOg9Ow5lMzrDbS9awaQ8uNcE1kYIZxBN0D//sZmf7RisvhS3Z+j73cPlU
C2SbFM6chMLtUu3MC92BBOigmhJiyu07nSrEQ0qnsQwlN4NgB8blPXIms+Zn8l6tlKaSjOwNqzRO
qxpXnMqw+P1ywLSQWH134jeC3IGbjAnnko4JiEukOxR3Z5O3B1EfFJpfg/b08T9OXSSn7M55k2lK
bym/tmU5JqmadJEmKBbZVf39JiCjgtO8N23h+kX5+8x1+PIG49avgIGM+8JOECjfDxXdGcliL9FM
EahbB+H2ukBfWKaRFcvRCRX59BFWq83va8R8Ak7JXQUl8tCOoapPdi2CVYRHySpZoYoLK5H7V22r
zYnj9Nsqdd2Io8n18PTcuA2baCxa9lE5FdrEru/dIfsKS3eljYuhidHXoNDLaTSId6JaecTqDal0
A+ubaA+vTTlbfvCG8Kv2ryM8raSyTqpvThkFJp6j0+7TpSeHOeex0RtqI7wAyvTxL2QwIgY0SyMl
vqnR/ep+X16tHFLB2rzW9OPC0UyRdMt//rBvTHjx3TZLhUDH2jDXoorKdEYqRkLKAML+UoIwUIKk
dE0xLDNtXEpDTgIKbRM9R+vWtEZ6bkpTdwMacd1KJPupEAMnFniGVSHrZrq2o+xvLAOSnfi2RIJE
ZKvAiD4jA2dadOQLPQfaAbD6+ncR8KtGI2i16mjXa6gUrqyR0xlPQhErjwzlIKFj3AOxAFcQTBVK
oYzldHEdo+WnLomBq7AgyB90AqKuFHjaY+5yC6svn24+El5RAROscoyumqxqkKG7knifPEfCrF+1
C4mXzN6Mb3dUxs4atJhuZ+n6vz1t+Nph4UqPBliwGqTRwaqbPv8SoBPWNZkVYLIi6WmVxIpjwBQ+
sWowc9ah1kybQABVdiwd+ORsBy7VIb8l3RPVR9E8YdLIZMWc6HkEPxsptLzfWIPJ4I84TACAUSzl
QIbXlQL66TgYU3kgXgC1MGYsLabxq9a69o/oaAySPB3l85iLrM4FEOqw2yB9qKuEgbB133+i7SH+
U30Bkb0+A3QfgwQL3yBIBsDvDG4wGfln7WnwacYQalhgr1921FQBBCen+DicOmxtDfprqcmRhWmc
Xw+fbvJzqNhjtspQD1XrpcY/fAzO1xB3HYfpUYLOhPZhSlfiZma8dnQoe6lqmLEvLeRAZcY+VBeF
a5syuLN3foDLmXwVKH7p0ruFBVEwecFV2/RVVJQdrf55DwevUpCfcqz5K2HJ+znjgQ6yPCXYqxhy
mK/BuES4bO13qDpHtrhNFcpfN/I6tO4bkqivIbKuvcobftMijL+/298ZlEAw5MhzpHsHjsvTu5VM
RssGyziUIqWmit3SVHpGT8eLLlC1eEkqQUjJV+65ghyiqd7CPqQbn1JdouqiAVfLH+lXs4Dletpi
U9YhCZUmGgs9BOxrxRITpFMzkQdarCBLqWUUB5hkU1J2Va9sbkwfdXs3ZiQGzx8B/eLIN5YGsMD3
XYGZHzw004Ckzm7ZWZs3IJiRy0ESQCRTsRaRzAT73BKUQo0Uqm7yi9244qyPhE4wp+0paDdgNDcA
yzuAMLceZeB73vLdcV/eZ+MjZWt0TKYnx+RE1DPJsj+LF2L0Xwi9SALJIWzAQ1B/ZDz2J6FdtyaD
YdLtyChNLUFialQgJJKfQIagOHrh4NqleBXCBkwq23o54zR5S8J6RxO3KL04tzj2pPjFIAe90cu/
1HOSP/yzPSdyhuXwzMnDf7zntapl+DBk3lb0AaKDet2GLq16K7RnE10o5RxfpunXdQZOZmyO3uNQ
nCV9C1tWpQeM3hlqG9Ec66TGvwPuBvkztOS0a4SPemaL5si9YdeGPv5y5AFWxLjwWkOIWR07qujf
o7WcW99Jg2VLLLuorHIx7+1fHPe5G89swniN/vr/JCnZs7dgW/Q6eU5XIydz+yDf5ahKC3MVv/Lb
b7gpQA888WrAZGo/guAkeTQOHNrBFiTMrpfYj0zl885TREwzoK1nkcVy2hbhj3/K2r/HTRiyMqXx
/gPT3nGbZyQ1Wzue/fw6WJRwmn/V1lKzwWNsfypZTaGInlYpHC+Cr9LwNd8GJUdLX8b4kP0liR55
ewTxjtl6rIdxLtYIVzXzc9gobBhMgDnDamM8hUx7weV9zQrvklFVnTdh2UjLSKTOOmGo5tH1+XYb
CbkgYVrFErneiChnmtGAhRBVO1ZGrMTTauOFIrbOVTTWG5Vn8m7HFpG+gzEvAqEI4G1uqolgc30D
BhJcMZ6IRTCx/UjbfnZOGHbTqhe5FTsoRUzDO9P7pzx3A+pJ3A7+nYbv3E4OLafJX0OWxxuVjnuf
OMlmfeLd7gdE3AnBM5x7cEfEuT/3nHIhdpA5AXvjYxbF6fJcDb4rbhgj41YmV4IbhGo749o3ot8b
aWetdnLv6DiP06mMfbAfXmqA8sD/o5DHYj9clSNRpqVvuruyqiwoNrcRPf5rPvEUk6clW06Rpuns
gUqU0T6MmILaNw1gRIWWEfAHdnsYxxXFzoppRXKaIYy/AsWiX0wvFEQpTwC60/YCWrm1wkrG8mtg
XC4sLl8nIhD2sst0iqu+3xB2tkohMDyq2q8kFv1DFLtsMg+zeLZq1SZs/dJ62zFODgo84hSpBxsK
Ih3JpeTXkXOZSLlNz/Wupv0xSPvaI6pzbHntFXmxH8kGnCZtR/iev9fDFrvGy8ggSIEn54xiLk3z
xB2spuHnFw3SPZQ/KRmtCMNwI56WTQ+9OVoVxETNlID8jVBjDmtvkpS9kVg/LP8mZtmYmWhFM+QE
d/5u22U1xvNJtI95IuQIeIY3NiXM1IG5C/yQ0GEHacTrohE52Kn8THstegMTIg7zWIqxTSfXFsVC
bB8kOuI7iIYv9R8eSkuT3etfOs8byYxkfSUwRZDKie4TCUCyiIYa/Anx7RpH3M6IeakXtBu8KRBa
lECu4kBsPRJ2TaG4/EO0pob0JbXSUXyZh91rjgy6gREOUs00RuMKlpgQtSmNdzYamuszeKjQIwvz
WL7LsB+S+IydUSpL71gvcNiwdKKeoBLds+E0RytsGTmqpe9aKkUWM0BZczo5DuAKnrjLoteXWx+I
y4PUpVpXe7C5Dvt1NNm8JTmqJcvd7QoJN5iyitav6Vuh16Mu2wVnTARGbV542dszXtd5SkQV413U
3Z5oaI/8fBIu7Rg8AYoIYjUtq8qBksAAe0zBoUBGUldfZbBBDNcBYAjbHvEa+1Zz8riQBq0qqvkv
rk8O5xhl0a2N1YHiUPDCvbpyugoo7HAFBk5zM8OM/NZRH9ClB8gfDjddJDL8KJHrfzA3BHW2vozV
dQm7wF6qQnXfc3ILpF3TT5aM/n/T7UyntbOg/iYgug3Ra7JfhRVXc02jMQz8Pi1DBkLttAsbqoEn
mvTWHT7THymbYKtK3L8HAnpjHvaTk8/Nu6TJl7Bk05MYaE/b3NqF4bnFEVu+IVWCd6eVQuIDm+fp
SIWkYBjhK+ka9LkzaMnXw2QkD6j4qNDxV8WF24HlTc/Sd3+PQQItaGSEeB/fzBqQ20fLUL7+pEW6
Qx9YBHWORGqJWKRQxBCtu6tW0KFlamdnyei7zVVvrVrFBLu0OMc2OWsp115Sia+Y8pNJsgbBjB6B
WL+LfQQufcIJJnd1qDQhiuJn3ahwU96+5PXwjkNz1o5jIkYfU6I3+jSzY930dpizuW8eWQRyCKxJ
0rTw6brCF9g7+JjQ32M0Mbg7gEDszRoqHFQe7oI7DLoYFbYdydD3w7jxsiX1QOzk5Hs5+mvcjcTq
taB/p07PEbTqgltMMXZFj9CBcw12emd+P81l1n8PKPM4+YrbAhsqy7+rpje6GY5sXcc3/aK2lAfe
25ftOx5MwUg1EKLYkxI7sjUF4dkIOarjfgNJ7cikGVO5nE2OIe47sLglrFPHPKzO2RszYH2e+vLL
zhvLkVYLlKq4jCYBNXGTDXch1nb4nbMmql3R8lwXPcca+0/leconQ2D/jSkeS+34uPo4jExfyO5U
i8FyYDfnSsf90NhhqEmMvcwqa0F/JxgNQNxzU6rDoA86N/+N85QO3QepVqGZrtSqcLAYMaFnesqh
ZqlBekQEOsiFQV3mS5tZmlkacsdzmHivdLuHpZLdDN3WHzsC9A6Cbn8HEsvhQlYIUOZp6dIG8WYZ
eC+s1iGiJVO4mvAr2YNxSrmwts28JdqKbbCjf0t5GCzFkdtLNbn+ephh1k4jWaWuA6zGhIGBPaPk
KwKwR5n00Nc1xDaeyKUEToUz2V8IcWZg+PIZv4yeWzXlMpJ6X92031beCOP8KPKFdRtO/JmGjAS0
R1U6XsLzioOdmQZ8B5pW6B9YBeytzhZ5W5QdqcMKKaeYdIBjXvZgWpRffHwQ+JIIalgvzt7VB0Do
NpWsv2s+rN0k1+BhamAoZTGGmN0jaSF0SR1SES0BFDKs++6/q7RuKigYobYVzXaegs9JU6eR25VT
DMzGv1v1eKANl4L5oXluC4Xi3BPxddoEMlZKWOnpI6OLG765kxlyFytZ/McYEa86+yHxRPF8Fcec
d1cPjEcVncEllvll4kzSopoCImbQrTH8/IFYNWR5I67Z7XP4acP4e+0qL+oV5HqjaiODbZt4zMtE
NGPkYNe/bTC2Ogqp1cBFdz3pLRLmo3rg19lIDylbwyAR3BrRYkTV+8icRR/9cYzImeIg04XChPdm
s3fkrU85YGyYAyHkdwzCL/0PRA1t8Od4BMakmHXhZJ15e1x1j2ABiBIjLXT91+53cspreSceF0Dm
WNOl/kWdOyVp6uNZsoQMUqw9Iz5+XoBuKKUNarJeX2qM0tLEnuMdxg7NG6xDu+Vs+wiXQDaQrFCo
FjZ/LLc9Pb4G7iWmrovIXRJ1ro41Cy1O6c0spEHQb2Z2SE3GdEU7a5aGJP9jaPqUZpnFPuygSY17
qn3HCAZW/CX5gxvAneNb8HN5bu8p7WKbgNJBuGqWCJ2gUVnv9teVRtOgGKdQ2zVHh2TwFxueWH00
2aCbonpuRtixlcC//qybUH10gsVb8ofmcp7A3SMHws7F84h1IX9nrFiLhawLFNl/C6q4vSFrV4i8
ezxYmL04qRZdyvU6O8/50p39CvPf6ZXfn4cuJ/XE2L9sztcrzYsck0rZ8xIHW3ChWzfnnV8ftx2t
uCt5K56/WQMRlmtvpM1/2zGkGO99Ne2AZPAw2NBDNXdPxjg7mUq8q6ydZs+a6p36JtqnQrE5pk/j
JJbs6MP4a2zNBi4SDyQ+GxcaC3nPl/I9S7v/kIS/1xscYMncbilRiC56pvn9KeYRF14xdmjmig3e
q+SrY64ZwUHk24jfs3RHauXFGR/wtuoPoBcgUgNdzC615TQJZz5QpOFv7vamwbKr2cDMi1VygTtI
d/YJnb3GGcND7CnYVz0UH3X2V5UvFZ6wuHUQ8Vfe/804Y06FG1G1dJ27JqOoFr7Oz2mKj5Ugy0RM
Cgq8IkuiKHqvcL1lWV5A0yT0wFgDASp3Z7HSOrc8qJecFEnyvC+U2B+2JGhDle1jyDlLIbQxy2jp
3t7PMei4D3Na39F9pSxo4AvU37Rq1jcBHJ+R5ICuPTW2Ycfz8xlWezozNMPbWB2LXI8s/WS3wRQ0
y/DXbK9DPXSsZ5u22DOhlHA+viwq4bfxdz37vAMuuFcP8U4Sz9bQh5HYKdTNSYwQ4fQ3kLga9ueQ
FoXS19eoudodqIwt8HWr1KCGeayl8gYPqpeLIvG32VxPAi7V3sWB3vBZ7YG5KIensDBmg6Zyx83G
tbKbzmu9UQN8ICG9OE9UZ7eJhpUdTg7r9d96APoXmLOWaH8XDMCumiRHy1Zj1enVcdVWzz2fUFwM
PqBDU+xIUcp2p6j8RQ7FPFAVuQLc9RS/Te7aKcguvGnT4VAbODWX7vPUMQngAZcZHSysWI6mPjWF
SPpg7sCwMOAJPv4p9xma4Hxw1CBFgu+5gPlWN7aSNx89OChTy7Mtf/q4WDnZXP+E33QOk8aPvPJG
6xr1XvBnCRzvan6JuOPC6tTBlnO1wq0N4O4uP9YZ1dAF4BSc/0u5cu+Zm8WbVTo3qBaldUz11aYS
yAzz+nSt/8bsNaXCnGG4XlxewtXgt0LQpEhD8E/7gJqhoAAtYU/H9YsbywNum9siL+6/Z5zs200w
5kYBP+prp0KNsMIJkX5gn7W0DI1g999glbZ/4HSj/WWYI63+hIxBoHrIVIh6e1OY5xsKBI7FSCLv
hPJZ+qykUB0RmCEYrpCQry9os+EgTlq7Eg+I9sAqpGzn5gtVhbN8m2vhi/z57B/N9mcHQH9Nk3ui
nwSZ7vLXvfxU0GLfZZSe067cofbWE9sf7S4GiJ3s91eG0xGF8ju5Vguw1N3OfrHjU5PF0GK1uGTv
Xy/9LBxaxb4tgqylF5JDPG2L2nqa2UWS02vganZHoUFQof24jL/szIy7ge8LIux7kXhupwFl/q13
URXaaVAVvvwxpfk6zF2AuIZPlyf3fh4Q74EcCfCWZqiZvX4zdX5Pfxb5tQccg9rqBG7Bnv0UGDsC
b6d9uSAP2IMwhFoxiGbEU5EIt4FL6gl0mVAJEL7Db74WzsW72D2SUUReTXmqlIkGQddUEezR7TDv
XYsJpFhERfxmpxSWLK7IsoMu3yKfLr132XqtO9uzo94AvL0zxaJ5XEhkkjGr2izhOYPM3fSpJu3F
v1xEFIbLWrkBqC/Kn3SW3i8XqPU9SCxPfvqpOfQ2U1gSxVbbXi8mBAtkM2ySnAYcP9JId1qxdDbN
G99qnoG5yas2K2k5NgdQbyFw3f0E82mVPEVzkWp5ExCEpf/4B5JwqG6PrdBsPisTnfRQtYpZifpW
CMeDgCIQ7d7eLP85h1NWeo/S9T7dt3mbe3yN46im1IRySb3Koo/MlVOYIyr9KAG7IcAWlPcSsxmp
iKCnc3cntHaQzeSBrit9zkfjv/L6y3OJy6z1/BbeaCYTSVVxItj4QZT48gMTtF4lF2+9BTQrC0qD
g8D5YOxjqymH58XKWuNaQZNyUzW6Dmr9MigxZeK1RD2LMwOwu28xTByfiaF4nPYLesuQvLulp4Rn
vZkQBCycvGKAdo6zQSC9Sr78T2z5myaRBtuOFvDOzTSOP4K2v5EIOgHRqipF8snM3fYG8qtfpAli
kK8uKX6V2nQyfGaDvIhLE07g+4p0beqqvn2ErwiFZnN9Zn6Q44n5iDtHgXlLlnbQaJp/ILkqqLCQ
FBjjrz758vMQaYhvaMZUFJV+CLAuJ0xkkhrcF7JxrcA+aBSZ4DvicttjuK30doS3FoQQiBoXW6Bo
i+jHhKsHwnBUSkJg/i825deH5RxS41NV+t4NGYDfxtRLciFbf2gbFHkJbBrraLHjWVc90YU2W9kW
cSheSgtGK03uzu9qhQWJnCmDZDNE884me7ia8HPU/qnAgQ/8zzHQvma+q0URrxEH6ANFwxnJji7t
mYNokzSMCWYI7cCRdhH/sfMnoZOQMihpoPUWvKqw0r8sJXOQhUdumlHqfWzKUCj4dcJXVi9zZTn/
q60wS6MdieGTEQ1MddiDyNGKTsSN1gBycGAfjgL3WUunYdutDHvy6j0T08lsFpbftaHJcxbuXt34
JKmgU+XoeI514/a9NgU3JUtzK5owV2J6ek1QwcDszBIKXOMY+gJoKu57w/MNCdsiPxVN+pJhX+wa
w/igoX1cvz1xZst2+enPAwh9za+1jmjTLHkMnwF4ZC3XjtEwX0hlmgZUtTcR84d2t5ZnMLIyNCZe
9jI2LeAqsN9B8Jvf9s+lmCpbhlAw4R24Vpg1GGC+gg4nVlx7u8s2jcV2gFyw0erfkiBEfnXbezDK
+oYPFA7C3kvZm9ooo+dkr/ECNv+w9WA5364N2w1zghiKczhTj5j6VVb2rejcx7hGMWiA2ukWnDhq
v3r5u4UdCAP/s04NWY9gbHN7j7ibFnkSMwyLFFenUQ8ucUY+LEIkHRwHT8oTZGGWj9glM8K1xHKb
9VEr8Puf/n/eLVEpYlzRe2kmiQ5K8M2ZI1GQG/6Rd1hvW/oqFowwlLyUZSNyT0aRkCE21OcUKcm5
u4czR6rN/ew9J7i9qb4lG8JgCcoQ+3C/nqoKlbPgC+wZkQ/h3EXoV+8SEuRghfuqgzAAKfS0MOzB
+xJIoeAzEHh1YsPCGJIYQBGtgLHPNfHJ0NnO7HVdMYPAj0QlUH22Jf4IqsB0772Z6gkM1v7UvW9H
5C3KkyoV4gt8s0lHi8wHuEqlpvcJrxPU3cVIRlPpszcLR3X3LjsY96Ij/CaXXpFqTMDugDJSfz2l
2mCP/8pDlbT5PWRve6dh6d1GEQwT8JL9YXiIQSa8sLfakRsVDXSP8D0wWNQIDdrlhq+RB8B63sM4
+gd/r8kLdARMHmNx5RiPr3CVXme2iNep1UmrQz+GRenXtC+Tu5UPcycke39WXCIaWjC1u4zj2hYF
xCA1vyVX1bqYPCA9wro8M4SLxu9JhTd1Hcbh0Rj9yRKZzC44aCcdaqp35BmpmBNlYOhgq2jAsC0M
pdeFUaBNq6R9CcQ59gGNNgqWM4vXIpkBvRFvhdf9D1KjWgIFfog4b2J1vDbXZ0kMC5WEEs7ENBgd
qwsmNiQNcCvRfJUQx6jZKCwkPysuq041hcPvK2jumTIeCzxlPat8bJtRBMtEj5XmTCdxdWYzfpjJ
GVwKyIbJv8U2EGxNQxh6MKdjeJe6SVxx7KUXTfGeIZ7Zm4FbqpUcIrpEKnlsWk9iDgn1Ke2I/kcD
j/+pSaIsQaE4hOFhrLy1vEHRL54ruvMVOXstOa8ptSRUc/4JSJ/4zqGPKIVH0Gw34K/w1n6MuCSw
YqAJDLzMRB+HNcZENuKAN22LjmbPa3+eobeFG1ZT2mWytKt2VeMUtuqzu/xLVab3x+5crai4xFOa
TNqfjB0VpeliyWEryzANGbc9s/tqCAlVCMFqEt01XMonGwdlUbo9glozmh6pOovkShyX7IGox6OM
6aAhiEqmGHmybjTO3dGScD29OkynXWzrbfA5GC8FKIyzZgNoi48eMFOYfga+vFn67KiOPGgGjvcE
QIou1EkFsfP/BagwBbCbU+t/cAn2ah2nobjvMizq62yyPRefDu1xKiFQ8uQaC3c4k0ACJqG8rJxl
RWNojj0sV9x4ROKSGjKqOdzYZhBdz3h+MwpNLxB2/O+PWIqufwlrNK7okdOt3m/s6zs7piwbytPC
4PB891GtgGDP+5X11dbsvT41qvXgSKbq7hyXdXpRiUgG5gmQGy8LzXWDtSjqhc6Lf6sndWwgtDut
eBSDF9FJgrUikcAVexz0ODPO7lYPajmjOb9IN/kAmY1wHmZ/bisOaNDQ4rlkLUsJL1ikeooJvQNw
xLGS+yRIgPUFrpvK4E97mvj4E69PnE/vNIzHKSQBTptr9FR5GU2Gg2Z0QZeF8Nmwo0T91WBXnOCl
ztr5ZkrpnRSCBUteqC1Z6gPfosFYRZjbISOS8YwuLMNH0+9bPqM4XT41eyy7eHgW3Jd/KspeQavV
aNzzwL7VPw7yQ2R9SspVM9DHw0HtuYO30lhi5Z6Vn4KVFBVXlsSij2TDCCs1EcGajb52fZWasr9+
jDZECUeyUN7w7r605e/zKTaA/IcUA0qxw+n/HvXITKrbqExY1XEeayAnx+MNqbzi1m+F1/HMgJ7T
0KH+kqZDlvUJcXh6FXk3RviEaN9K11s9pbgrpiKyBvEOqB5oLlGTwjq0h08tI3rAEMVhELF5VgGC
ui9Ojkzkpkk7mMoR2qGOcgJ4Ag4mNccsV6kT8yU53OrUVjke6ssfBKjcvLL+K+J9kz+8xv38VbNN
fn1MvXkcXFIYDX/yEAioSOwAQPjuEe3Zocu0HhgSyXs1cWazVOD+1O4vg++Ii0lKGL8caSHilovz
4aD2tgnFJSbGIfdvwpRE1vldgZhRgJEOxwBrZLzd5JwXwvpvifz6WY0teosppiDlL2qO//MeRKfP
9NX+FK+9V/FWApw8GlLcVnynNG/KTIC0NOxYc2in2Cl7oQ8wGmQHSYc6hAs1G+wm20r4wey608kl
8rlqsWGtEyJjamLuUFdSlhxsWhufqIvrCVKrGO46aioq50KM7IJHmzJKFln8GMxQ2YaNnrgFHf9m
HG2n9eeRIi7nwPO1j7tky59OnOAMfDvNUVDqCPKLpqr+0Fk5hq3BKTO6IzMEVd4Foi83Tjo5rpWX
Zs/sv/0z4Sz1vZgkP9Lp3lZBwHh2z240N7KMtWIsKNS79X1bUeJT5sD5TDA5srQbhppA72eJaVuO
rW3Fm6xtIuBdeGoEIzW5BSTknz4cdAVk+EmmIdosHto39GEFpPCG8nPtH/ZQSFuxIIj/SgE9tmX2
N73wjGEMfWNI7trOH6I8u7EAkJS076D8G7YiR4ISZfHBsa/VfxAUoW9r21gBn4EYsI+ICHkkWBA5
x4wbIc3C0c7j+ZXA9c58x5JvMPvZbhLjFNl2JtOZxFTRcaiIvIFG4ttZ1yGNRx9M4/1/K2jm7g3e
2HjkXJdZ669nLc6hAe+bLH0mav49YOt5Y68y20PCLevZpLZnwrYEpnviO7/1Em+d8gU4EtP32Dg7
jGQ8T6KMt2zI47fvqMkV2Q1tHe48y//6cGVDzWDGMLSHFVMDkhj0sZ8IKFrmqRa4p5YCvRJOXJxG
yLdH/R9xdqHHtb4wYcrYDuKHPFB0kjaU2Z/ylumAGdq+ihRiL2QU0rVE7mqa19381gw1RAJXS/+9
CkGVl+t9YFfbl8ISbW9bR9vLbSX/ob3UUIoZ1Vt2wniOTakQpA5pI6DnvP8Lj5YBLsxuC3Xv5QTw
hyct/9mKw29Vc8ZVtapg0SZHmt0uG+WHmZSWs45AwPpTSK2zJCaDzrCp72dXj7BLkw4BAw/ysGKj
xegW7YGfgG00Q71gC00js4Z/s/BsbR7d48qqaQgNHCYP2CUUGhClgFegBsrYICWr04QoaVKrAox4
om2g2PgtIe0tX6zilYVGHKeuAp/2QMyw5bh5KQ3NXmGQBkiaPKrwMaio8QQOfPixaqkGjbY9gjb0
psFp/dtkdfSAWTKqYlI7/y/jLn8fqTNfXPg39ycOncupwz/vN7xd2hPpoIpOEdvafkPkLB4XiXo+
NYnFpPUPeTV1gscQenI8Q+SeszFtSjkwPvEMwcyq6iDfkGE+H9n3gaYCS+lLpEh/lovl4NUU8PUS
2NJiixur8RR0mV6K7tJzkVQuVtXDLPNlFLNS5DO47n9YiR08VUZaJL8+9D7ItMVrOWaNF4Pmw2/7
/k3wPw3cBfooSktTxqdOKpIogB+pFCCbPRZOquUXliDvQ/6SRXe0JhwNa5srOtYRRJrqYTY3mmWy
LTnqcj2IThW+5Vl6f0/f9hp0qLHNCRc0CsieSCEYyngAMBh+YCytuukhrap22EVFFcRzcuz+oj7A
LbImrLl8GHQ7oZDPtYTRAG/eMkfcMl6wf+I1E8guLbFoLetCNAkB8N6Qr+lEeQcWXDujZnONU2/O
JJyclLqbrz9OhlgU3UVsfbHQU9VJHCLJ6N/RJRW+JIsjIzkkVMcsPVIwNOHWx7i6cmgt9uU7LIFd
tsOepkP8Kpe2lH2TpsVE0etr1DuwdtuA745So5vTUAycRxIaJSKk8JFEvdPZfHBIA6HjRQArq9Lq
S95szKp4Sr2Z5/oJ7GAJksvI0zWbWwDRSuW3r+eEFNsDOad1NWkQY60yuj1/DkjJ0CFHYJAoqxXA
ZnZSKDLX43GvlqeA05mBsX+AKq7Etq5CO/smZc5L3wngEbq78+dziQ97Ve3xClzRfwHMJq1U37B/
ReJhA6bFkyplSmW0MHj389muctOP3gEdXlq6VzavGfhZ/PBATYLCx/kiduWvx15fOhCVbRCp5MUh
77oMgGx5yeTgX6DJXnpSnaMa15H9620ACbgfFOTLBQ1i01TcmApKRwdmcm5z5HceKjkPvmHCPCmI
aJtLdJ1ljXLXQ+ImSYTh/5qBQMj/4ZAPJPlS0QlpBcjbxwCsQD4SKarsxcarJacbU70p+IaoM2ZH
HdHFr3e5/O7JFACtRzi8iDTt5POKYLW8jG20ze+Vg5Sq4zpj7TOicdJlVU95TZpMRDBbXTfZQRjY
NLTYdoY+lPNVsK4nKBZBTt79Cv40NIpsxeI+0lU2QoKdSOMIjajAGBjSKLFUgHguskYW+UmDPVQo
vDbPZoivtK3tW6OAHG0SvDQu+hWNpABDhDvK0z2WXcTCNYHOb9s7cL9fzzQ72hgaMs7iuA3nt8cV
SHPb8xaFE7PggU/GqD2mqX+50z72V6N8CkTMeEnkc0eGqDlmjqEZSbs7SqDTPAXCw/1CGhcTCKLR
cwFioiTEold/Ii1BTJqe/FP1FrUCbd01cdt8P58cC0XZgU1RQUC5r84EQruaqVhCC4aeZ1Ae7wES
zZ3a/9G2h+eBpTQTnRRwYBVZduPtYl8sVWA9VpzjaBtcQfUHYwbTKrGSyDcmaZ7SAZfO6sa7KIus
cF1n9aoSiL9knD1i4DNWxqo2+HoUEgF554nlH0ch7EQ4UFhOkErOytxFZsZmwBiOdKzjyzDzx4b1
gB9ZxSaVAjxbgzioFdVjRkuAmG8DczTD3nfQpr18MiKgRUFUwf+BA9+n8yWz5ZnFaGHMlaIR7gCZ
MnTh1KWuKzXi0WA4h+6bBAc68UWxnZpHaKfMP123HE+fkQD9uq6vai0Ji06uGiFOPvXJeQqAK3jK
gMqmPw+uF2iCO/rlbS7/K3HX+0jp1hgi9oHmDAgXeNuRlhRq9HPLQWMaOybSY/JuFG2MHDd241zB
R7lM79lazi0p59/VjuyF5oSNz4lEaw8p5/tml+mB+vpHwCh88wZdNWdaSxRQ+OJx29G/JWaR7fGI
NqaGc4lt5+7oE48is7lhWSMHsqUYSBcx575OydR7ngN/T0LUrUKotbhZwIRhU9hCi7Wjii272bjM
/vqQXI/ZUXUZSAj3LgxMi1A4UX4HEX0qn1uAA61X5LN7xb8ceTPN2Wv+uKi6O043ZxxQ1k/4ZhIL
bGb277h5mPUoVX2ldG2NOTBRdwV8MSN2nlReSoWtb7SaKFZlmScIor7nvCIfmH79lLL7dBIf/UUb
wpTQemuBBQrg4QlUQe8WUoWtPoy9VnXuVPJv1RtLYueN7AIgc2GRrbd4NIsUGFP+Yb1ShV5bBKFf
vZYpJkD5j+6I9bKnrtSLmSMRaRE/H0RwJNiW9140TvIjExItw7hgbIyKu+Mm1ZARmMWjjpr8CGfB
/vypxzA/D3MdnQkMg2soljh2ZxF9rWxf3/jbONrMwVgpk5BZoenXCOyYckw6uiJtAiyXmVQD9mGm
35JsgtNQ9UjzVck0XgTxfWW+Os9LsoNXVrDa6lwRNpBKTYoC0/AmblrCEQHdb2lWOgbvFzfaCGrL
OCUVPwJC+ENsNe5zyyFwhQTv5OaXENgNmHNOySHrXCW4RQSU5uMUbrkAQL+yOBNaCRuYT3cy8jMc
iypTlzEDSwKqzGS0lLL9U3WOP8XtS3MIheFQ2efCyhKs7i72uR+SE78i/UjplpnJ6yRxT0rPjZqk
mk08xNl9dCBOrkmVP0mgMbAyhrUslb6tngDcHaoDJ+EcKvnPdDTcPlAn8pq0TZXuBgfNvCxfeAF9
JsCWuHyFJ6LayjsgAYFkZU+AUzH8Hy3VR9ekCLujBzeTavcEA5C1gw0HJicn7zaoD2xvjBZgcCqD
CeEKFSPQ2K+hlMnBxV4RyWnbGWYd0FW2Uh1VRim54d7bMsKHx0c38AlylUUep+XGKcRd0fgzKM0Q
exaHmVLJxfBIuts/wBuXGzt65n3fEo3yu/x5HNHo72pZu1k+1A6R7UVHwxVDSG2iQvscwI0fYStC
ig0tSnvKXpWLSPjiRmAwM+lNjjj0bMPufoYacHzc874QJVo73N20bp7PBR+vcYmwlgnj6GjYHbo5
O0kylQWRfya/2hP1BVpvlvFGKgt+nT8noHb9CBhzZMPSfkcrEAoyctVGp6yxjkAlVxnJDTZt/t71
ZVNye4TC8hiWSvr09ikEMjKhllWxx1oHbeunMg7NASeUeIRLemDRYzwXqBKpq+uvHPNYCt9os/Of
CgI6T+IUYPDOZVUGkdsG4CcjQQ8xTftI2vMPuUe4GfXtordTsaE5Gh6U4JhDm8x9khBSpiI4SJjZ
A5HSV2YO+oal8XRJKfni+1T6iBUz5vTykTNyJfgtrVXoEm/znI8TRYLs/jeg6eJV+hBbH8eJh56r
pOg2PXdOIQwbH++VfxSspaaqpPOAlnisyOJeZvvpiVLz4lc/ETNfT4ZigeRTP3rz8IIE1nQ5bIww
98m1SaJXfUApTeAeVPX9F6yEqIQTtEdaSAnSQjiHoK6oicBKyzUAEEuibabHbtRsP75fi4+akju5
zw5jC74EPaT+6NMaKIZ0N+19+U6LzRqbJcZCA5zsxuFFt78fe+JRk98wD3fQwK648St2NTCf9imh
ecNPv1SDZ+uL12we6SjLzKZG/cq6rkklnnW6xyiNs/8kigeu4m47iKUk6K5N8YWWBhBbKZYI2oNl
WPGiBIqunklibazOe7Eqr1uQl9S2gp+HLV6S1eyTdxC/G1vpeXRp8tEzar8QVoFd+XqOueP1qz2g
YDnDp6/SwiWxs107dHFUyXEueAI/yFbJvh3cTlb9r41waLmoXLj7NsKgK+2EfBZ/zo0xPeR01ARn
7/D4zjoPT1nZXE1Jc9CP4g8Zabm+ji8brk1iau55hX6N0L829HfmIFi33wTkNnft7zEki98XxL5I
/tlLv1YsTIdethHQwwCBGnstdSiNTIbXA/xeli+uCriMVDpZ9BBhe26CqgzlFTT0DbMFmYW8ToCE
PMawlSXzHvNe0tzPwwcrvpL8HHul4nWiHlK/B8ln95dmLXUW7nmdCTMoi5caHrmH0UXIsgFMFBK8
FW7BbaweBWWeZySke1m4rvj4fhzptGvfpl5DRG9UmSwMQGcG8eR+ShwDZArjkk+R5Lv969Ez64Ak
bGnoN3sPOFIDgdmuJXGwdLLKR5nIAVuDUsUeC0l45G4iDku0hgSVeZg63UJHmBAMqW9FUmCU6ZCx
55up2LaNuHFRFSm4kQUvQqHAyRQcN7AScfbjKtNdTq2igkvl7alN+0EnAIjH0eg/xlpayMsNkbZD
LOpgrjsYtlr0BEYlmY6Pfved9GEoFGzYFbU0z0qOg/Xzh4Au51lI6RzBb/3JM4Lzi1jLI7OF/KL9
7UYIkBaQBPD9zja+zU0+RYDoTyLgUYd7i0QfBx3ovqGaUyg1xWJO62Emr74dmJF1fVUrrbNJ7yll
3dPUOiEzINxdHjsVsP1BgClM0OVKKMPeCXxKwPBQaGZ8BkV2UwIsMA2PI1oUszTlkr4acacZpQTw
ZJtR02N9IfKQHghmYBqEoozmuLO5U6jbh65dg2WS0AGQmyJ2WM4wT7oBdr0hsmpmPySFP5tqbXdK
shBCUaHn2sBOdm4toBWS20CN/dOmEWDuv9/wZz96A31SiWekc5PgWrtV9LBTdzoTn/mDvGABWTAH
ss29rQMAXbMtA556Ntw0aMVCiMGjtKPrKxraEaeFNyYCAYc79m3XZINg2vmOXz3sOIG710wmNw7G
eKoEemhohvR+TLHCkwiu/PoyY98YEEVy8MB7zoF9GxRMJ54TsV5/r0gZJtkAVR0M4HnW4O8ROVkJ
u3lj0kNFhVQFLTAf+KhK4W0r7LO1XoTohmdquH17a8iDzSeTAlLRJq9NRFv8cH1e9+B+U9i0ee9a
1kc447m1lkoPweSBJ3XZKvs4S6NNrrcvaABNj6pXZwQrgftEjTL6gVQzo7+Wb/XCek9rxJ6KAKw8
c7oHLt1So97lOE2qXwaRmn8jmA2jMSyy3BX5ryqjnKYYnjQtwxN00EBsmkaS1LaXGlDM5ijWKphz
Dr/AEiEvtSFR94BJSKiipP+MzW6/6/Yf5no+jrVPpSDQ6qYAF7HvPs9E7s9+aZCqiw+50k+XO5B5
kc2WZPNgOxKAmWS5Lq1XZQLXTYrPYQHMfqPabUNxeHdLk46h/TAcT5kKytrJx+NRPglKVt8nvEtu
uNTtTFRRy6OyI9nSUP82AzfiRCZQR2cXYUbvu9I0sGzuCY8a1N+7+/lGIAL3qc8vg4xSval8lhPF
5rRD8W7pQT5Y+yQ3xpQMX1II5LGs6zpcD+C4xM4tjnIbPmLI64oOms0fGTSbiLljvxWeUyi84Zo1
GwLOW8Ag+WCn9KwpcJ5FS9cz+suDALxVUK9EcAyKEkraAbxRNBniw1/eNRuZUJsfrMn4g7F4oMID
5rOPDee9Wv+HV6OihTpOPUFMPxhe7HcJfvSAh0Il+ryN9hHe0Gko1+elu81ubWEg+1a89bnObQeu
d7yv1ej06jPYtL4nzcybhOfLs+vnYNxnAeD2unTpFogq4qcWzOTRONZtwt6+Dt0Vc2gBb+vjfxhe
MGfPP7GLtMaG1mYkv9A0Xm10V+svzzdAKm4RlZEf1vIWMdLHF87ic+M37F/faBpK6Uut2hlJJPKX
KDHa34K4SDzIgnXW1/bi0cnc7+3n9Dn8d4Va2l+ItGg10EXXOlqZIAzDBc2AAIErc6UIXN0eG17W
gNDBEt0cOPf3gSq8vGWyIi8PBBoMk9bKtRCnmGlwFTKj3sP+0JIxPOP58SHzYbxUL7PlBShC+ttc
0Oks6IZcgMGivPbP+Zpm0koIGg6ySO3YLNC08UGESeVo5EpJii9Vr+9bXl4HBe89b+xPC+t9gM/2
FIXCotggoVdD/WgQX9ysTEmITu2PBGjic/NoJtxPsCqx+1wg0LbwvcDUdyPrwYjCdQR7Wp/nVuiX
+ABh9qi/KWxlbLZsicSyKXykPcmoUItAIZtyIwb1IBs0FZ9Rq+kmWIfPQV4HjeCUDpplqjLUZ5dQ
SccZnwJi4Cew7SS5T27mb8ATFsXqK8DeR2DPyAEl7l7tABSrHTa54RbllYs/lhm0mlT1CK+d6eja
uBk0DUMD94A6IRwB47P+ZoPv5JfmcXT/xX2hbxsQGlKhzrNs1dW7Tquovy41tdFr4PCPwEjRr1ES
qFbUDEoM58IrEykU2VYbgf0UPsQH8RuocAs4ajLfKTIwUVZbAHPB9PDL8Kw2Tar84Bep/nXL2Ma+
YpbBATni+mdPBLUqDQMMJ+4ZaIz3TxnE1vggrlS3K/JqUDX/gJMUMU3UNIUyBOMS4ZCfS6dCpKCS
StLNME/XIm8BfynEZKCi7LB+6NvUsFEeOUcIW+MTv+55raMr2p9I5FBDXdtQP8lOBiWvMSPKehFp
fH+TvRCliBmwhalhtnK+jWLGmuiz9iV7V1FX55wgZuuZyjZD7/TM7uqM5KpavU+MMIikBifCQD5t
CRNkToEnDyKGRIrVHdReuF8j3atSdpfzHbUJAn1m1fbwWqWv3VcpQkHHaQqYNuj/g6n6b2rUFR3D
bC0lInbkaYZIJKtpY2FqC/HePGyayO4Fi4fflEhUtaex/6L5r8e0Rk//KSUi6bwIfNg9Q9PVtz0T
S48zPLlbacZKK1OKDf5xExSXnxf+vVjEJQATjln7gCy6GADB7v5hqd1GPajDLvUum3alA1peX9sI
VtwNlWEkTzMF4+QLQuF5i+T+6ZKSl51kduuo5DKa1mgNH0e6X8ACNUoUHBq/Ofbry7o1meVQilsD
nu099vD9EIb4B7qPlMfF1As8juJa+G94672ZjbewJ4XN+LqEKPsMmADdk/Wq/GiaaZMUccG8KSym
yHjIemM7lvG4g9HUE9OayYHhqek5KqVDjeh3BIRue9F22vPU8Vc/3i+2CgO4fHjb7w2wXh/qc1Qm
VjLlbmNDgWlG0z8LYH+tnu2RdT8QnaPmrElhhfWI0tW2OfQFvoUsTJxjQRcOsUrQdL+uzeTLRHLN
WDAJh/K2LwoKvwEd4l1k5IhlxaLqXP85CkFSjn1WLn+75V/4zPfmw1vN/y4s8a/P/DBWfLcyccuk
tzdZ/Q7kvZ2UD2cBE7iIVSnhUOMKG/UxmS8pSDNR2h8t5P49PW4hlh14++YA1oMwNd2OP0XSFgz7
zkCrZrgWdqIn3trYM0DIqbatFWtNYL/NLAsz2uxlBtIXQH4lJItGAczYvm9mvtjaDDhWle/PHhgb
k9khxD+uWZJpt2wTZtLAstqcapAw98Ng3hY3mmDmoZHMVsM2RzEtyOUEZMlvCmezo/stqvQx14dO
/AdRYt5B3jscgaBX88/ZItwT3BiVDbi8d4PprWruX5i/fBcWXqLergavss4bzOr+9y3v59xXcL4l
HCOjsNr5GrJIUQLnP1JDC2BFGa4YDuTaJlxkNmxLG3BCgx5AJ2z0nfkBiRaouE45OehkmFFC7rdR
XkRZjJnEOa09nMRZicptHXJCrJOkW2z05kdVzl+RmDav1KL6zRgxbpM1qVduMlGjAVpoc8jaVb6I
BBtJUjOXYMDxaCwfAkHhdVcuVhU7/T1RYp/ylYYd4cu0MDXNcIvjxt9MyRbZT2EZDpONQAaJuf2p
xDlZvLfBF8MVaMQ8tALE/Tsozi2ggDEWeOy2wRldDK0Mt2TeJq+ZENETouWy+y4r9oqil4bsApAl
HubDM3Xxj4Io3V2Xr7rRTbkQICq0Dz1P6QUI4dycY22fSy3MYQBrTGwkG2qJTraWlwejsNj/odRG
TCxAwQkWgkKy5o+HbVT4Zq0Hk1cwIVbfYvGDD6rv6zswcddwhPB3cDHhDvIkzw4L+cByY2h87vw1
Y9GD/OnRLHoE3OrGKawOxdjRiTDWJsL3ZKSCXNWaK24rC6u7D26HGhYg19AIP790+8Va/STDuHjw
WCZOOb6BJi1dZ8OvHNa4zWVNsJLUKylQ+fI08BNQPmaA5OIJjPxRGQOjRZ8r0eUlBTBSFpRO1lvD
cSJJZiMBsDQ93xo+fy4cTeGFdKEZb0goXvwIuEygtm56g/MSNkU2dCgdXBD8R2/2QLPeD/pWO1ya
+8y67FY9vV3fjyU9p5oa1tZyCcSYRbVbdBEoBqGgK/2ridFJt3G5vj7fPRGSc2uhXM/4sKs54uaU
R9kmdunydV4DTeomeV8XnhwMaEoJuODWyBtg8TCUVebKdh5tbCnTfp+xm9eCUvK39gySrrqj4i1t
usHOOh2Hr40LVKqXS1t4sKXqAokeLv/38KAXWy8Gfb1H5gNXmRq7hpUl5SnEv0Qj7IJQnZpB4Kyg
5aPef+mSInzssIUxfLK/6Y668QLCym9DWpt/fVdxilLtXGL0u9xBQuTZP5FvMrzwkw0XEJwN1EiH
AHQyB6QbJh/wlKfuxby4vhNuSfzaU0VCvyJI4ApGVruRjuuZrpETG8w/aUAx+GabJW6kzT214GKY
Me2WMK53wWczH3VOjG8PSQV0dERnVQBDQLuvMnxR8fvaWZQlAdwUCfWR6a3p3ZFPY8Y44hmAJs4l
3T2aKwJC1PPX52l/8pL8oSseIAifTLijZeD95Ga383thquSd0nZ0jRxyamb/0KyVNkWk0f1DgJ9w
qDyzJjygCYXwlWBmYVPoe2wAeWP/c5p24GpC0HSQHXzJ/HQXzJyklToy28vXWY/55t5CN14EnBhc
XT34qHJMYin9NnyK1heFfudbtBMfCNYyjbUdKFbmu7Y+K85zxR/bGEVLbptgInhPpRRr+qJtVanx
RzMc0dCCD13tMNPbKWecJ8V0t+ktHDupINd/yiGH+OGNxeP+PI7qWJNiZJYYKzYeRXb04nBUmHPx
BIS8mOn/4/w1OGRrgVmUNlFpwIa5rlwyMrXN0Xe/5F6JJCJ6AMoqxLfCGK91tTVNpixdn9hMQkKq
rOkKs5h1pRXmFveRD1jCUZ3fQuwV4ItvDyw02T2GpI61HugTb9aFxy4xjOF/RGJpoAzYck1L/AOZ
JaWKfXlAHgNiJZ/c6+O6dv90u1r5fYkC6inqJOHhw/TyJ8OU90xhxcmlj+MY//jbEPANqmqC6QHf
v2kqlKu0cJF36TiGeS7i2bi5HlNZ20Z/1wnWZgYqzwzvCip02DlAcrU0H6JyFwjS4JqXPpurcqhi
/BzQJwAMoL//kPDEcAwlZjEETbXcTWELkXSrY3MIOMcPPd6G1BCFSfGz3g7BPDtR/b02DbLAdz5q
vFU4TJj65+FqSE9kuKZW86kHioNa5axhOkYhzuBVZ1tdoCAKEg8MFKzf/FICHcSKyKptHinJ94fB
F00OPjFbJkD0fMNJBYGWJjdiPMrrBpDhT5G48C6xKecVwXOSRCpkkXhqosD8YsXqp/6cuYsh+fh7
HQ1PhsrWr0LZIENE5WuRhfYWAopA/Vmd53Hj5j9jp+9PaN9oZJ2IsF1vimeWUzFcoqKNpDO+zuY9
4FAxXIr7BB765DTe6ZJ44xYCX8qhyt6Ndmbdp01kFIUW2QYChOSqlhSNM4pe7ExnNuslYX4zbSC4
kshkVU2utGgHQ/n0jrtCt7kmDzrLhExJJHdsJnOChGNaB8JbQkaOXkvnGFjxR+J+rNaOck7JzDY8
IezwjTWW8aSDEG0c1MWGeL8T4Vcgdjd9sgrbt/GiHAADQigyKdA/l65k4lRR6w9hGnI3QqAIV9gZ
PTOhIJ+xiSJUUffylO3yTpd9+QQ9vc5qdGz+KGblbu97pQsLJh4UYrkfrJ/q5zuL4nz2q3NczQxc
bDgte0Bm/tz5QzgnN9W0hdumgP5sUWFAfCZfnDIniKWs9kBHUdkOfNgboJBk1Qi4gCcngyAinhvG
vuKLS/XuxX6zyJ8WzOWKhccGNS1WpIuiSdm4qKORNuSs34WZ136CcMCNjIBKIyqMsOsuL/rd7uS+
JMqeVzVZCuYsK6/aVGIQ26ePfwvGdLA6yrSECRAFbkeozuTNH+uA5lDF2BuQOQcVf/pxZBxVJEAJ
aPDcPU4lvvaoPMSCkp8JZGbXK+EBxPO5BisEbglPvUEvuEfjuHqoPvifTZiQav4YkLDShTa8CbAZ
j3r70dXs2agDBzuWX2mcAt10y5NbPCkiieCHn2KWNYJp6YK7EHuVV7BR/CGO+yRv6NFRtTqaKnf6
f6ekt2IQnULTxAUeRK1u1Mu2mKyTTV2rgUMiHfsvI65lXHZKb8U/ryZjH8Vo1BOmvc5ipwX3P2Fq
iHsuW6T5DeaL0UDkKBOp37GqT7aeS2DqCscj7fCv8nq0vGhB3wYsQGMttHUWbSOTNpz/3F8E5atr
trUtJIN09ZQK9ZWARjey0lpjtaW6BEcaL6YvWEmfFadFDUFMRPwjJSwWstx2O8sWzbZi2cmLNOZc
xTKrX3qNr4RLmE/IbbJGBJaSdHrtBdrSQmXzr9SjCMV7mpO+p0WOGI4hWdKMfrMBSv7NK0ZGR572
ulpP6PPrAi+4RB1RPX+5FmSjRMDcPyh27YacXD6hMjlQdXCULqClYgv0WbpsDjkri7VN2pAlugiv
wVbfTG6LWFZYjwcurIXMDzuHpSldEVBjE+C8wlUeUtJtLVTle9hqtzoPbE3mdetzbEJq061aIFf+
9dlBLUVIEc/DxGl12NZaPYXSGbXXAEOSqAKd7QlcMFLqBkrEV+91xPt0D1PxZSFqQ3JFpalrvv60
Q5PJwZFfntKiCkur5a/Qmwc/1BNtdLl230/2drDVDLmuTee0bcW77d2vYCwqoWlt8ArC1Swjpu5V
Xq9HQQyBXqT8HJTWOblf/ya27nyst9oLKxjTduw8EP4AjW6IIoxD4fJ6q06Cvs6GaoOGYeGcHCsA
kZ59H18bM8kvDlvfdemT0KzE8ATWtMWnz/EpQg6pk2IwE2Ntax8GleQzZ6PSTO0F2Ftqzupv6w/8
ZhtkDhf1uihM+8a0HgpOtyrmstHqktr5Oin+A+PAfUFtcdQn7LPKyR4VYNlSGbs6yKO0z3QrrBBJ
4Ub6f+JcLiME8uSdGKSGmEf+bT9PPIH9JaUPo/jSADtsoCjwqMBTpcsXmIkoo+iw78YtG6SgIjxp
nQPz7g8AyH+pyQqUGUIzeDlftVfTd+NZX+LJAQ+rnxGwTJ6c240cvpfmdPCOn0mJAIFGpaIYfgiU
iGdcmJmINulrJpHbL3GcnqNzJkdYLJJXlVvulk7/r8hKQ2E3/ZX5IE2k3ZS6Gep2k4dl7kXrkzXq
UkjcvMQksdHDaBVXOX4g/P2XIlv5t0CNY56J5IPkFgGV7VBzXaYpV0eI3oOO1dSkie5Lx+9zNdGj
MnPhIwpyCibGOfCitUbpQAaQghwrbwSjW+LZlIUgqzuVUXavJes0xTpgHZZkOninziDLzGHTPiLm
MArxbunKP1Jf/BXEXBdQ0koEnWyny4FXVJXH9AfBU48FKtzqeYWBKoN7aQn5qLHez590leWANjcd
lmmUlL/0ZB10Aa5zYilfyyreYj9WIa1PMbCzQ5FZ25OSPeoOQg8mBBBGCNEdzJwIXZu8GLSrYdMz
44NDpJZ3mAXaPqCKuwVD8UK6jWyRG3w1rGFzcB8oql7PYNQ3K1jz6BvAugfvdqQEyF0m+2vhNzhb
MXUvlnPmjnK1aK71bDuuz8PUW7Fbh/xIhl3nj05rfNYYDER70G3yFnlamCUm2QX3OIxVgoRwOaBK
++0ZEU4Skhqg+Yp5VXc+pH334NkhZmXdPOW6sI2kHU80TugiImJtescTZ9tTUUAnPzNlhyxLrwF3
naM93T+CCbEJLHFhUG5xKYeNUr+CIu1ybZehR4nVT76YoFqRrjbzuRdHXx5tlrPtcip1QqMmh6/Y
uQ3iAJ+hIli1mGYBX6Aocci/pL7llLpvF1cbj3Pgml3WxzvNSY/hYdJERVNrBLuP1AjpL7L5JXGC
J2zTYGMyxvLDP+zBaddcjeJ5pe6z7npDku3F3RnacmULkX6zBAbugMPnLhbFtGSR79leW/RiFXMe
LFi9UpFK8T4AFkvQr3oKRveSDhFDRwS+kjxqO94vxKSwbx/jcjAt5qgDVOR1+QptPyoxx38VqJ2r
tiMC/I9PlhUKDt23fOJTdJYfxuo02ufEb1CJ2siMhzl5sxHK0VTW2LPZN4hVTwb5I9S2N5EUh5b3
jOYiQUIqvnJ/0LZ73WwFHQGFjw86W46X2H29bTTRRnUnG2jiKxsgwfUsthNfdG6QSCwyJ02gf/4m
SvARi/gBj+Hc8yOgi3bcShdONQMkMHUW9I7NF5kuY6sQVdTMM5VwIJSAzqaQ+3LeSjdAtaLPfB8b
xQNuraRiDpP2J5XImoyygmVYeyyrxbTug3XOhGB3cUYfYdzZAgSlUiwd742+wiiS4x1p4IRe6suc
xRgdXjfKZpJBu90cnIrnAeLl/9ncvDdZxsMr1mSSLg8n2ZxaytSEh/JFT025YUjr0AbQnC8SHVEk
zg5TrAPSRB78QBjUHXRKBtKV8ptJD/hQHgc5xCYHp58y291QcDUV8InxF1rLG96UL3MzoL2CyGLw
C1iPKgJo98vpesrW0kPFowD7jDCQFhZlJfff1yCZ76Umf5YTTG443T9cHPUPkf57TwN4MZZ26Z+O
6zx0Fx0Mta7Ls/PO/BjYXmca+7UhpbbQEGeoq6J9ggg8t5zRgAgWTWxaiqh3lw8Wh1vAQuGPCJbY
l+TiGZixIynxbjKuSsMZbSCTHPqKEk266RYCzRnDExdxn9Rv3kK90aALMTQIEl+1XHq7SXJJZzBR
sh0gC6si9V9jueUBYiYYzQHutEr9TaoSVFAUZOWuhsWi854raKkpsYe42HAWU6bLoK4ib2xqnWgk
bp4ynC5wffrhw/F4koskn6Utop9KFwrMmO0cSxsEmyLm54ShHT6sF995pdm7Gziawque6XynrDR7
auQip6G15yKAwMToavh75GKX57ahbwrOiRk2IXKoq+r0VyTNDeid9lHM3atdU2Kr//vpVbKWZ91a
Ojm+sWt+1p8OHplZ4Ki2UoeWsM1NbHXB0AMGk1VtKt2/hqEFfUqOqNZWEvkwcqw91Sm+MR4buMYa
QxssYUdPeh9CRUbvIJv1V5EWgxr9L/dqKxP4iG053RJ+Lyp2u3IkAXcWlqz7M2Xmwu/R1pZcFFaU
yYzRfNNUi9B8lJ1MNPAxSZIfX7PBLSYbUIPjp9KI1FiT16ClRKfaS6JpXCROaUhAjsbLvMca1O1s
U0J6tf1KKd+4Mef64saS92wkv5LTsQ9WBFMniI0UjU3Q+odrf9YaJWxvEDH3b48XFOVj856ynJov
ymHr/6PGsUZSU2Zw+l7swiFlKKgqOU7MkE5KdVeThkt2PtvJQEqAbJojaP6JjB0g0WGgOCnT1FOp
aKzGJpvqSHAmFzqTpiDbW2HLBfPgdbwNyTqb+triT5mpQi9U6VrrxK02NkMj81ugiTn/s/AI1Xgx
Fr593Tzl+1yRvFhLnVaykJYoPjo7cm+mLaS2BXZqhor9uHii9G+qn7Oz4cWgWbch2IaadbgyRxlB
p+L2IB6BKB26LVmMjLcBlpM51FKDBp7uqukpVmTupZ+TE+hVH5k7bNhsJiK6q7GEXfNrwoy/q1k2
vnYzGvwIlnlSZCIdRFXbPBzAGsFA91n8lRfzmIyHpCjMFhtRYEpr7DAZBuu3sNWPGV9ebR1zGgPs
fY4aPpNDGLp/7NdDb2XUXHHeKe1q/Q9Oj550PmpeNVJWGK4Cc0H2FzmKpgrst8kBdu6+fxHdYpwb
VrZOY7TAVsitXTmeczmLTd0MLPgver60F2tqFZDP4zIxV2t+HYGQBlj55ARv4L+yvvM4gqPooZg9
saKxYeEvBFfnYo9L5U1CWwgkjF+yYxQWu+fF34yTYbiEyu39SUNq8z/ZqT6GauKLRMXyQXGpvtU5
Fv8Oda9wDUa0L5TG6OXe8KcVs3rdVXMKzguNb7EsoXXOjBJE3cuEhWiU5LV+uC0jB3caz3FKAuCh
UorTUNCARDXkiH5cQbRVZbGa6DBlkUhKH5vococKF/j0cFu6a8RQg7/YpKlHM37rZaJWdRo/scOf
33rMV4kyFabJG4F5ec6TpD0X7o2ftMpLdWxh8Py9McJ5rUXneCvuUVCheCneU6xG239qqVDYKPlo
JywV3QyPgz4bnAz382C/aLL+D7YU+rhM4xw8vF8VdPoVhdFqJ+ap9bHRm3mReiPR+Aq6Qu1uuVMV
AuJqeM/t7dfakasv68CsJDbkPVmdgdDNPFFPcE9ZzgCjI3OctcYtvKfduV3bKMPgVq9d8bVdahIB
swQnZZi4BtIMQ6wOPo9xhN/9CUXEtMpIdrhIHUdCqJ/jX9ZYlS05/mjKFIBzrHyNU+Gi9DJU7b3q
Zb8pPRWIX+ihcVFfeGIsWK1sPIGmGw4MVKq7I5xpd+z9FDHAreU4/fSGt4vQO2EHvcSRvrhumo1C
kly0xDstVgoMbh2kvEwID8Xwk8bGGldzeVlZsQgMrMHdD3HggDcVImqzTFPdxL7uTq/2Jquj5c6c
Uc9vJEkEFODpvpO5HdUpXtLcQwRAsgpYvT7TZ2J2msC+YOtCdF3wV6w/WNSoRMTGfyBHlW1RGsCk
36WJUtMhTaSpQkfN8dRHPD9dlmAo5wcNpYfrl4+qs1sVwfi0BqCaBiPAT0O+peL4tlYCc8rDb0jx
vGISPriV2+DrKoQV0wYg5ZUNBd+HnsrVZBSClBYEQQHCc+qbOahXYYWTNYNU6hZhmE7B3NggkWQw
IdX8BW8FMzwJ1IppaHiTtT6f1Mq6sMnwLFnc+AKvWe5Ng9W75raAf3AOcFk8AlWHHOcFTCzKfyJj
OH9PNbbrmKlzwA9zi7aPezzjIL2EWesFsyA0ry71NhnH1alvRROqeHlknpxLUnNBJvuDz9fjMVSv
ywJXaPLMxk8vEogxWy4letTcl32l20BpbU1ak3RC5nFAtn3/TwvhyHgQMGDD3zFqvcZiMWfu54ix
u184jWBVxkMkYQqRXrB+LWe7CJnUEEvHh7GFB2xQ7oZADtfbKSwH4HWzhwZLDDM4vKhv/QzQF/Lu
gvisdsIeRr0NP1U4zfI2b7W0pKKRSZklnVhitG7cFkIgfJdsRgdVmP5RxRye2mqqO/f9IVJrweRV
UI25Ks4dACBzkf5+5ovvsrm9jJ7SMFPT3UsMg+H8sKF+icTiW5wbiySf04VZrT2goUeLTn9oWwdo
4uEFg9A3R83ehkU7wzS7NLe1ttrMJWKjYXzcov3/PZB6M1YBd6yU2Pfn+pfw3fJzPDTt+NTu12Zs
fj5Zh6bLkxUIZEc1F4NAadzqTcyrPFoQbR+ytRt8RZhEcQx9ifnjH5Sv049f0w3h1GILfheapNZn
+HGSndcdFMkwqSb7X5NSo5/ILIUDNP6CdzCpF45+SnPa4dy60lczumsuCVO65YHTKbJRFiRp/sUk
zfRIqqX6/T9JCUQdXx98KLfz41r10XpMjZ9dgrcYbBcYbLIli0rOT0vtjv0zg2GpLhdQsekGpYo4
8hRy0cKMMG+zcgMr++Uu/TIucVMFC8eyzjkcOie84NBDpxCCRiMRt/Gm4mda4WVlA+RMrc85LJxp
wwREhSLDtl+rJngXd8/GID7VJ9dbW6JFimbKsncElNbgqNwUqQ8fDDtWYtBkCBX6vnVQSTZBmjwC
mNU3AXUtfU6g5KsM3oBVzwqxt/qvUcc2B2NvNgrf93cw5uGxb59R9FDXHJa/FTgdL/1Hsmmd2NtC
vMpT1/jIbDyPoYZ1bFP/wdt0UAc56Ow+dfjhQHkU2GkVuCVs9Ze4XUMM+/FsdhkB3mnSY72+hRSC
+cfIlEDq9UiscoLvKc9ju7gvXW565+eLYpB5nf9F89/4y8mMW4TKnmqvvXkTkTUl2hv+/q5TeIlb
tg1aRJV5DubrTSWBixmvWpwPmwfhZpYD9G+MyDo/nGbsH8/Ya8KCL5MqAduK5oq8NvrlSCfjnv6g
2ARmPTgwMuOZ3k3D4V2csT4P5K8vCpi7U/WvbzJmfAweF9o+E/k/5B37dFUSoQy8bve2s2zbTbeq
237OJwzfEAu/j1Ej3QJ/l9G2AE5hEe9zDr0OznAfqhi5OnQJHF58K2tRuHbI9TO05gCsBRyT7yKa
UtKHh9KtJONNtJJzxpe2HrmEWQnibWl0pOwA9Z0XoHlWxrBmjWOqNSBsbp2VLXdjYKzNJuq2xjdu
hJdekqg1F1+/4WwGDOl7CaFNz2Qkj3EpkP+KLR6PiPgOweanHLuzFPKOCzX1KqotjzOUr3Ic/yIz
DGq+R7TttSq9mrsRgjzuUj+wdDAgGq8wDUd8fUlsuA0DaQAbzMo3Y+sbR/6zuIRWlvfZ3p7JUF39
p4t/YoptZAfufy1tnKNq03C98To8cjN+5G1NTwHy4YnMvfN2KXxx5z2CmR5zC85iocJW9He8Afu6
RVBHwZinQmS6+NbT0+rKYoKlq9I+ZpJyFw15SGLkVOx3TByIUX0UZDuGF8AA1Y34V/vhvGnFPVbT
ObH/hi0lJEvvNc0PthFDbwEshYhcakIIGjr4kUTr6y5MUfF2o7T8QSxpUxXvsxyDmsBv9K04AtPH
tJcZ+Dd0sC3SZpCJ9zxPV0zb/Q5QLuZqMbfYh+f0w7MkfMC3tNZz7GQpPnKhDDrtXcHselRA85/A
jhLv1MWKPouNVA/U14qgtN7AAWgmNsEM1oFZ4h1GYJBYdOSvZ86IUkrIJ+wSe61Xja6ot6sftFbE
6bOozeBFbj43q/sX+T4N2I7NQwY+6GOHj0Y1JCdEJTw21Z/GwjwFEyg/Z4HWMRY6siIPFWSTOdWx
Z+Iz+9cNmu0MJSrb0hDjCRiiqnRDfRvmBmJzvYZUUcWKKit5ZP2iJpNf8c2MLkhoPXOI/U5tQaFm
kk6qTJENILxI5ByfrPyT5TU3/JiteTeISrQB5mhkhUPKwTJvES9iQZDKaywAWd3CUdeeBDZV9RsS
joXST8zBLPyliQD/ZtPKIneOV1rE7J5nD8t4V2Qw5zkWtaxzD8Pndsgt9X5QstH4CWY9UGXjAtzN
4/pcSSpq0O8rVWVg01kCcCb0IOsaQ2w7aEunAvZI9DjMiQcZ/qwS2isSOoAhEdBAZF44JbeJ4PIw
JW27mVFxX3dMTVpCQ6BVVHGW6wIcdoWXloj/IUN6ZcejKPBIP48rbHh4vL0HXShrKMTVNElPW6a6
lUYMcfWDl0DFuNsxDeBbhsZtDlqPeP2HRzIl0Ch0QABRo4dSXD7lQRt9gsEz3g2nAYiFBpt5Lhn7
xPRnasuRKZzKNgmgcdvq0YjJmUprt509RJMpLg1dJ83+cCCyUR1ZnZnIqz07R0pDRHyZSgacuv8g
wppS9HaSbiH7/11tZk4J9OEadcabQp68SIT+1B+qJvKr3z2xwS9YHKomerVbrFfYQw9XFb4XiWkM
+j05VYOec1Z2wpplQZ8SmZbaJ+DbBrP/Gn3vutQfvNeJcJs3mxUtMY4vYpzqMiLG7XJVyoZ6GwZl
5ITUKtj6MP57H6K+qOwlMi44ZgX9BZlGg81E7lZfUdH+BGzGUeRCVH1/qP00HtqzU/HfNrjuEgox
GrraDKQT7KdXF71lY35F8NOw2XcYfQkbu5h5Knoj47VtL2V1o73CpgnW3UyXbp2myfko5TFHF0FV
ZKmmsbt5qUIg5Kq8SGbHKEEDyep42ucVe/uZHildq/UjZwALdE9weljon9eXyeISlMGWfHm5jgWB
0tR2O7hmNXCpvuRD1r7D1i3DZyZJ+W/LiUTJbDXBAguwX3PYXFDn1QEBz6rStRAmqRj598vqNzOb
4Rg24YWm3/DNEcX6CjZ7BEgFF1sMHM1mAVXeXH0qj0hX8ht2YPVy0eN4+ZouO3YRduawaNKhli67
EcV1S13L8N//cc2U8LKpI90dn5PD/Cfygth15x6PcgC+tHZ1zpNGGBoPwJgHNPNLgTl5Lgl0TmiD
utyCtrhJ3UjMf60NLm/6dG/HO5uWOPmNdaoyHPuzNAI8hezws//bA3HUaOBwmxC5onB5E7CVI2OX
yu3j3vK4Fv7H9Y7oSRViln168xkumGFyfSgCz4PEn6ntGOS05SPBblp+Dgmuljt8jRKaFltysJUq
2cxO+qx/YqLhYNcVeKAhwR+ZcHFEXMkfpXhu9+yMlKGIr5bVTpgaKUXTQl46ravjjQDhMymAXORA
aYBnH9pSgxVpap/x3hCgYtBmhut7l1CUy44V3zyFtEmnJisK1fV+h09eGG8hRbB5oGsT8wzKqtge
NUm/xZHS5R4zCpYg9HTKRNkDXdCM0gVrYvoZ5/qEdcPoV3Nzve1kJp5m2xLulnif4/tisyB19Bzq
A1UpEImzgiUzjtvZgKbxDNjkG/kasKOw7YvP9EoC4lr6pfjsaqtNHzsjuJ14/7t3VODmvl5zoEK2
2989H7MIdzfzs8EK3TYWN4PnX8ncZi1R2FEEj9zr8BuVeqLmm0FqSTE3P//xnZp0fNzLPq6E4oyN
sPZfrVbKVvt47oKZUHha63LlehPOOfFn731UN9QTE5uXPbcpc5hAv62ParRv+apJfrIVZuzgfEiq
y86KOde3HNUQz9drdwiocSgg35r2x2xk0enPmYMpkOAqcXqSh2Kt+eQeeqQzZBnz7iym+R6gEB3a
C+vtzrgx+ez+a2Exdj9qsXK9OjsbLrJBv5rdHLASjs9vfK132ArgV/0gZCasm4A4gl7fc4lrP4Be
hzi5yqPn0Bs8dodw9ygnqyqEi/ktU7DaA5MxojYyaHx4qyCks/eIHvNjVaKjQ9biR0oyiucbvr0W
xLW4pO3JeJ9At5rW+msxoyVbEuAmRB64LAu5+BxnNtd3xtH+HvgI06DL/udZYlVxGMDSt71It0Sr
4rMRWmWAVs/UiSW5186wPLR7z9Oi4OD1sotETs8voUhI0GC69EkBZoF3R7sMLSjx3Fwdx0/1Au7g
a3eoNTcSSMz6no7s4h2HjCutACseFZWYY5NJPdxQi1IN+FCiWNcpK81XlJbSYA+qPOG3nduMLa3r
eATfOvCipzyFnLnUMTl7ADwlgnufAimk1dUd3B/uJGGiBRRtb1kn1air0g9XPXKu/6cLUXHtz9GM
WeI+CvL2WrJqlN3XfAeM/P19wlm3hxmlwXZXctyckDgzQfmCYwZeQ4l+BVOpRVsZSBFzHQixJvgU
82xZCY6VIXhvYNpwCjtHIqPns2QHo8mKBqshaqHRdK+oQOy7CoLk4WY7NJZeHwxKymbYvh4M0pZ/
yUPl8cWB+gocEU1WOur3ORXU0C8rueq21Ll8C6LQNBEJWEWiW5EHrP4MQnoVbJzHWw2PPEcaMoIw
iZcRvDBxN+TTbPGhOcJ6WILKR5HqKbOgMIadYDmDr7KyquSAP6LHThAGxwUnOFnpfRDj9mk1Q5fZ
mwSJAKdGr4VXXX1b2VROCQ3Cgbd45TLZHdcd4rckhBEt2hc8XDRjmVkOq3UXxVuWc8X3x+Ao8TqA
mDHhnOfjh8graC81Njsk2YekIytG1110sNia18HbdIOZ0uU7eFL0TXGD87AhioSiBPQwQ2ZAn3Gd
XoeEiVzbZCY/723yepjy3zw3Gmidju5Pa53TvsfE/vr5wNzqng4GFDiyybLXKOuDTUFzjlmUhXCR
NBD9CnpacnvmIk9IcvQXgYZH9n5PjN323eTiN65kBmbYJLsdxl4kur1j3AojrerpbWbqDrvWRBSL
mnvXuwaXTaNVg/bPZhE+c4+qavPMqfhgJF0NsZyBwLnH8399hjQcaAsCLlre2PXMZ5DxYLIJ/oNP
vvk91qMzr12SWTIS0Rx6AQZSmyX2SzrJYMzftQ3Q/lI67CJ/p9uEpjmjjBNBz0FpfqjMpzvmj1FB
he2rnC+HGF5HDS/KDAmg9D2gp+k0HfnBDJPGSoVaOfhuDd8LLEc2ZHUe6UEW8MhlYryXMDEN+uTV
y12fVd+n7rwxc876t62per+MkiDqIkOOOktTuo2QTkYSxqyvLlfj6LC/bkJVFrEH0dY1X3mCZBEw
ojKJCseQWW2MGYMALKPo8nMMFz1YeEmkRIoMZO/+zAiUW3mRkcyIExZOVyv3c8RIMg4eBNZ0nS7/
g2HxlsYOy3Wr79Wplp5W+0m5aOHyvDyViU15Uf8Ygw6t/qRvaJbSX2lZHhoFvskMfkiztXEwKnbR
VqWo0vuO2N9fr9GmFKI+y+VQoanc/gGP2WQMZiXGHXwqaNRSoGXyelVCQ6OeVgtAa/s+OCSA28fB
XZxIrt2zibdcz/dYu9npgYVJlhq2S/qhjhF8csrXnKr7KyExoxUjlIZXgxDS6SFx8VxqeQh2iw6G
dWZYsHf4FXB1iU4VAP4OKzyvnIt5fz1G5I7dGUVhw2cDy70dhPmrHGfa6k2Y3zAuwPIlExDDEg8r
aw3hwaM6vtZhRp74bbKLaqhHpgCy/+52ui/FX+4GTzNGrJyGtK0hVFbsUtf3J5Lfe57hLYRSvYaj
GBBRKiTYdN8z23TRNRpUL7P2cjj6LHBY2ZpcJGe/64It5h1OStfFcRDH+kF7Nn181ztCrpIO6R/B
fsWQGrdH5OGzSvZe+tQsjKIgdmu3dPz7LLDfQiyWAQJcRHbKCifeW+gIahxSOtE+DDe4HB/Ly3c6
LFu3QmyRYRUGw7+e5oRw8Jk8clqYe8XVlnJAYlxQJQMx/tLLgx5mHOA2vEKz8wQK/GmO7q4+b0Hb
rBdqjX7hksaEqQqe+gCt8WEAfx6zgliRUCCgLodnx+c2FaWmUSWE/XKfpfoqNq4w6Q/bbjdKpwOw
J6VdObJsW7Z2B4EXPPCw8SkW5mH1SxxLVs5IfGOk2ylb8cwnP7sLQvCYItG9XsW6GejXIRUvisPH
vXcHnXIsCc2gAOz0iq9IJRwlBLz8YebvhRmADnnbzf8piyvPVgj4WXNA/EArrpIvJtWcrDrglquG
M8B1gKYe1PTcReoP77jRFMgYg9q3NqIC95gD0TvN7s9pcuvlMFKLSRaBqmd1wreIJLS4oJgAaMAa
4+sari6PWRRHbVZP3F8J08+Rquu0H3tlndt2QVe1dBSBgTV3oeW8i42QMonZii+9y8QQR+gV/Qms
L3+8bMDEbvyNvHCZQUxhqsVQLu/l9Csr6pI8hO79kVGC5uTzKUAnMVcGltTKmOgqrHFc0YGtRHY4
rXTzp+kUX7EsC17Hr6k/23BHZcEMRw7h/HIssUOmqcAmUfRNbpDySo7kCvvNDnbRaxPYBRDFSSEP
Wvcb6E4Jy5dyg/h4BMfbucKYXhVDRkWETCPWdVugW4JeZcNiwdpUjeNXzv1QQAC7gOxfvRoWhS2L
rpuSu1fnTFrpl61zgrrJO/M02pmuV4+TzCagHVqz/yP7vH78Vce5viDuodSOYeLxXLFqnhooKc7L
PbOOqI4xcw5EWYini77pmvsi3eHRhm4zfzuJaboOxsLByhTVhbeWecN9IQTw5XX4EY0mK3jW7XIo
LpLHf2xspdBwCTM93CNONQ0YvPBA/8ZWBWLw4i7wccm/dF9B502ZX+8i3o/xzrTe1cNLhaYLjq2f
LhlJhxqTCKAJOI1ratQR3rTNT9HxrDp3/KSC4FSAbo6P8jmLpmgkK5bAEUVZiikPmoeAUy5qKSUi
8RKx3JPJlMq4goWKfOBOGBQ8KEtbqB6SZDLzDqWuk1lEa+ARrue2eNzg8gy2nrQqnbh+WTVECvBp
qJg3akxBZ7ooqadQwVfEu13onao7rmv5u6SjGpToP6JLkks/I7DvOnA3SkUSCZnlJwMS5xNsLdiO
+O/Sx4fUeQFCHFHNEztQIwVWZp9IL73pR7Q8kLEeqJ3Tu2hMPUkTF1UKxH81XpDRMR24fGobADFE
qTR8RGSrhUwTW4Yb//gHGPJlWJsNWXvQvPW+Hhm98nXFdcBQKkzi2xgUxgTDS77jHqk4o7bgvmJP
+1TwWDKHia+SGDo+SAW+7MKujr5rhYXxg8KebLobyYs4qDFPJetpwutn3qSuZ9VrxYlHJUky4iSu
VPVE00a/YsIlr+K2c9syKiCoRdwYGBenDQERnaOx5Fg1SMbM/LgbwvHQQbbU/DRDyZ7rwDoLLdiu
LZuWtykDf7Fuxh1LVGNtz6Qjs9HlYmuhIHT3EOXmD4PuUR2sTjwnO8+9UE4fXPsLBfp+69ayj9I/
CL0hFoQewhIkoXrB0roQjtuyxn1GZoqjJoFPtFD46cTq76PQ2h+f6DpCFbypK8Hk+xfx4UbUuUFe
nu1+B3vmvp6YWWgekWAYFyK9FseW7p/ETJD86yUlWYM0Tjbe6V7C68bnydcOtvAsfcvlMxJyRC7L
JOqUcbO/BBw+QXRLpU72NGYxpDzKeREHP7/lFWLfo61r9fw8oxCI69ZxHlHyeJ6AOqni44ZALFOn
ULSIemNS4eHSb3xUXs40FtlFGzuUgSqpWSWLrtCnhxrGnA1m5FfN5q+e45Z0HV5mylpUvUVkdCtQ
qB3K+6YogccZUC61qNtHWO5khy1JxtW1VeUwJ0XmDlwJVLrGC61KzwZKay/I0NMMoYq4rWoY4Xpd
WaGhBLQCckitmKByOmMWJIn3MQf1C6j2bxdmmmXJuWzH1JXVZ6MG7V8J0Pt4x9OJyqzDqrorD9gF
E5YBQkFcHRc3F5d3TvoTQTjHPX6i2Rz5l9R5yrmJH+vWzieeax5cTWF4iw/yoEZh85g9M8Doi/jJ
UaNsvWbWgA0N/XucYr2vUMZ+W45KrHryhAMEkjTyEUIzui1rcxvd6DQjBVm5r4qx5FlLhmvOgpTF
C1kFe56VlyU4hrJigq5Jx2X7i3FqfH/6atUBtulrJbsnSBIBwJinTTFroEfMEVm/VMHK+YZhua8u
KSHXPY1v02A8q/nbSw4g3C04CYI2AX6yjxO3HpegOOsUnacj6+jLoKuWeM7W2V54CZMI8jDN4DnA
YzmPVx5g+aHVw+ybC8Oy3tve7A0HXedHzuLVpwYWzmZYwiXChNhuMm2kgHF04g9O3EEu7iVuPYaM
Oj4JhRSAFU++pcKiRKw8wLfIb5ICpitCxHCsC+y8SqgNDRC+b8MMMMlrIqKuoHps2xHpwIQYQRn1
HRidIX+dRq0RLm7+Tvp5G9d1N57k0VTqZK/zBSrR61JNILfSG5d+MMCZytKVqXywDeJJwmte43di
kdnSwS3vodxnQUUwKp7aWDUiDR8lV0QoMN/KQh1khNE/Hff5Gt1rmq5+enPZdWIdcPd6uVW/X7x8
YB9Hx424ZV/VmiDOvkmwG9qZJIL0v6aPkE9Kx4X2qz8XQJSfxCE0MNRSNRFuarfZsFceMPJBj5ZR
2wVn5sOoBJdjz4PsNjbiH+r54qXO+WgNYiPIpjyry1sGYTIUx5yBx1AYajWjXMH+JlxZzRsUAmzD
gwfPom38Bj7CdzVahVRqdtgAqUHdc8KrnwUQ2CuOTgS9k6kgtU4f1sHdGMBxv7DUoYocvdBo7uEf
oLtKOswDd4v8HWLJS2U/3J3NGZMPyd6mY1najZ/Ipcc3GuAkGm/VD5QrB6NpPj+ea4uDzr3CmT0A
xTXTbxJ21AiXYoiKhJyNkUy6jJZ8ohBFFS8Vdgj7PtVZhaIns2m3FW3ygLRFwF7Mm0ZdNH1EK+he
ZM59gTEJ3uLWC/cHxhgltsXB+tnWU/zVwGD62UfaakXiUJZI7I57n0v3WeUwJYwgFuBXDDC9qewD
iVBAk7wUcZIZai18KTv2dz78MMKJCLIHbFrZit6Yv7uUy+i9o+ZYrt3c9qh1+PxA9Te4HW2tXEVG
Hj6BZBgwuzgRdG1B+Kn6jam7hz7SpBQ7zlj2o7HfcEjZh0/AWMlBPPB/S9yfncSa9XEnlSXpOLKP
WrIUXeJAMWxSq+u1k6sUlm2Enjr67kOejZG/ukClQqbS5RP5659eFDv8s1U+w6md6+yx6DDmNXlg
Jj+7b7jnD/7Kx62RZpfrhfp2EiqN7Ja6xaaLjLhy0xCmEDbSMUtYP4hsl34cJ9KDF6oETcCT8PCp
gFXp12XmWOOErFoZXOUjufyDxu38NUeqSJq54ik1yyYAmD7e28Wk1H+rOE6J+Iqelnsra+zrUOWF
aN2GbtSynVkbq5C5SkDOd35Clvzadi2dmCurMX2NEUe6NG8ce9IlB6sTWbSZX6Qkm+7s3YZRi1vT
DHRa5A4azwd5NCdZCgWKzXWsvAZgywPc3ODKoeO3JLBfiBLNFV3BAvM9fpNX9LC5Q4LLW1YHWJfX
Y8Onrdt051Ud2Kco+rCIoG/KO6D9jmBWeXGJDbNew8OHWxPADwtQim/nIjKhLC756iQe6ic+GU5s
2IyeQLL+O81I3rJXqRTWDLv81St01VtiO7ocFM7ptfB4u7sr+jvI8ulJvMRlHtML5OxKezJFdmhe
4v3ikYADJaqMf7a4HRDk42FdBxHw2SmOQva4wY3bSgaHXwuI2gdRzVbTIK3PMlW8ImpLUqcTQkYx
MozCnmhY1/vrgB0WAEVo8gm4vgK2AN9e3b+M0jxAqonFBAp3B517pz/39vt+PM9+VR0N4oUduJpt
2TMTCusFUv+c/FoQal974MQ88G/s+scx3zL+QBpcuMu2h07b/0mOe5/WfGgsUjimSLHKnA0AMJrO
nGjne9AfTzg7ExOWpSzxJ2AHHRqTiucxQqp9ybTUMdZDuuOVUrsN8SDaPP6ZT5qYzEd+S7RK/Ec+
8RwebvYoYHDOMafPHtQu6/Qu3qW/8lInbeyVIefZkI/atWtVJNaBIGY96WL8NUWto+nEkw6Wf014
0/ibBHsQFLzgYzq9/gBHcmjKlefK0Tu+9PbpohfvJfefwUqkHuX4gME2bl58/5A9qxNz8XMe/gL7
L/in/tnfNxHOgDxYUYlHraB53ICGTAC1JbqMErsOMOfwyH0jd+UR0IXdxdrlfMWoaVo65/kLne4l
Jt/vSdeaMJ+fm7U3lWodmRTgqEe2eV8gNz8QbhtElNJ4LJy/Xg4MUt+RINO0uewkStatLphIuqzu
spENU37M38RwxpChPecG02vry2ZJQMM8D+JqaDsaDF8XUsjxHwtiFDzuThuj4OyKY86ZjjfYoGre
wLEyVBO7Qyt3otWaBpN4y7OYfzrTiuGILIGzqd3RSM82J5LhMDBf8eHepeGqTOzdjfanekLWCLZt
ErdVmx3j08GzyVwWkY5Uc6lTD8oRuDI+ZJPSPH57bQt3HC6DE6PSINvP5hjRTXfQtYyt7RGy7zwb
zAnxrJfp4xhil3LlFiAUNRSPUMxN+CplTK3fbZFPp67aYox+3Uenx/kgheDEHTnkOCD2Q7MGc47t
WECZXS+3Oj0rKsQ/ZGMqOPeTPonNhRdOXAoi2hFCSWAD1PXB8DLBY3o66VzM1xcZda2436HkkVNK
3OtVerETWhZbqa11UoQMv4EOfHZthwdGGN1/kTnUEkvcwSgt/qttvD2ffhTAByLsBk7+susvFrLN
6Le52mg8jKEPVKX18IF2VPxwd94mKCTix6pCxVrSgw0Oae4spBGQU10c0S5l0h1/f4sHPb+Gvnmk
fegpXD2bYSJrp+QZfqvNF/r651D1gQxAlI9Sq4hpOUrVOyeH1bLn2MGiAJpy9BP8JFzRab3gk3SP
RmQLKHwzXdJRR6lJVPgUWBwvQjTH14IJx3PMeWrMS6Fda5l3hDwOx6aIivdYFzXG+7CGIo2CxSjW
g7xdaHqAmxFcffKeeeoqTgVDHByDMPy4dv51SkQKaIfg30lplcKhI9xzu+JyZF8TTUBftTftYB25
hnakL52S47kskcTcZBLad0lz1cw35ifx0rO0YMnAgbs9qU13ANkuN9X08A6NfA6cF7kB0K+Ruiso
KorocSkYZLb1BsEOd283CqVvBm2zmTujZOiTI3GSiG1P/QoQ8LF8cN4hXJERYAPDEpfs3PkcRfpY
O87bU2gk9xKqmflCzkG18I+JEDGXTpSUyMNqQdKquqS/TNDNusIqzywz1xQsrMzaSdbU4eG0to3C
l8Q1nJtcV5D3jiPHYRVOigVcLKLqrKHnLtZrAlkF4bdmqoiIaIv3vrc6rIVvGbBTXyN4ZH0fTO+/
jl9oNMv8IGLFI5NOnURier5Kt9EfJkfldKzqc5sgKBFE0WPjDjdmpd/esjImAyMvQKvgA3qywT3I
ufHDLxYjUW9fGC3+CDzfZRF/TgsNxTcxxnlfcvKqBmoWYC/YtYoOshTuLF+x/9DaJCBcqZciKdAo
up2uwaCPTjpGMh9kSp4pmK4Y+L7aYtWV/r1f6uQbL+1DBZth/YIKnHyc0DVEj5ebhAi5zKIKFNCe
PkSeWi8U/Ovy81rEhH6L4R6oTrY066mvWdVeaUo1JQfHGHC+WinnEexWlAm0Qa5vHK0ODKVf4EQM
p7f0V2e+BXtOfREnuTLlEv6a4k9CWDiQfrSYUwvgJVYwRNQg5fsrt3+KnQeilHGH3BWDzF5S6zAh
QDhd+xzVD8FSeKqifKaqaxg8KMRzK16xgBTiKiQ4fVr4Ng9cq32SNGjZPQjPEAvTH0TwNAFbKQEq
9NwLjTpdIQigrUzLs815nToZuXrl68VtuxzzRQ7HAkkdo56yeE5eX7siSeCbMzLKlDd18e4ofpsR
Ofq9rfweJA3iDxAhM5gQPlWIR+3P+Qp3SqgiM6MvrEKCBfOy8y5D8FtIdnwYFXOg+CTnyjp9bJEc
FCusaYwSwMbFvrbQUlgGFjeiHuS3VBeG8tKAmn//XOc+en17HlFEaedGsYyGT+wUnAO7B0bDoLEu
WFz5j9CSUvwiPHPYDPob6mWEg3OBLqKG5+Cb2p7Wxd0Mqgk55x7wgHnw+p+qDMDGcCglDpJ32OOv
6vwBBdayuGVXWJ/L7GSOnG4fy1LWKOjfLj+Gr/RnlTWsPnLXxEP9zDXZd2OwlkBVxA7sPQv3r+WK
M1UzhIC7SlT2aNU6wEo7P358hLyvqVfOrPP80BRZS0FZHEuGscEQSBlhywBdubCxZzyFgOlK/u0q
u/VYRwk1FJDKAaMsmPRvZFfJHAHuiYwoBPh7XpTcroiXatw2R28qvZ/CPYaU1C4BhF24yhCCY6RU
mvx5m8wryhOZta1XQ9UVAd1EwiOkp2lNg3vD2kPYFX23Urlgak6+geAtKAfckKa4NtP6fhjhN8wk
75MCGOjtcVLL5MWyQcQs3a2+Z5/yv67VNRAbhwT7R9gYbWfAm7Q3Gnlqo5niTGh+C818jdrU/SBG
42XzJmRn4Lp5x0t834JSSyFsPMO1MeP++apJHTfr1jDBJ4Y2Dkf0AvnXwtamI6MDiE0QL1VhwfjV
twydlfXgJsjMtIZWL1Y0jyq1aEsNG6+PZ+OGiw5rx33rtKbhCL1E5Kfdi7Zix9bIJikHFoLU8bZS
jZki7dMDEhijPg04VyRKtf49tewQcJRaMiSrJuALes+F0SAJzIj5QPkk2ifuWOMc/zpCYHl5XdGM
SkczM34eBeBAI1MiSvpeUKzRPSTGKak7P7EPJZprS4zloT2MjYPuYpE6vp1rPMKRwpmLyUUZUkNp
RJKgJY/hQPCFyPNk9Acn7EPjcHe2NdmJ04GgGDzOnOI50+NCn9GJRA2YSJdo61TL+u7E9eJGKC99
aZ/Oxl2fbcG3YYorzXi2NaihoxyDVLz5lmmk/VhAkpp4RK1j20vXrkxZ8GAVafxwYVS0LUIqaJay
qwrlvo5I7yTQom3PEwFe9BJu97vMoVoDzs9ZW82QK5l/7uZ+D81zkabDslNwrHz+EsHrAwZHcK+8
yWKsMvgb+oVVeHoLKNktk1/9wXJxoEzGn5z+uHg3hD4l0l7lyKiPWHwmE2CfyWe/Nw1jTupxHSfr
j1nTknyeQeENHHDQU2JyAdfABzhubkequTUoRaJ8rNpWGjTuO37b+2VF0YBec+I6uc7DHxCKrFoV
inyW7r9cD78QsEjAI4YwCmHK5R9NagIR3I18AcymzZH2oSuBJbf9TaQgmHV0akUrKXXhcpi9f9eJ
j8MzbYnQU1wxb2ZvsGNVNFSMQrEJaRpea4sLPpof+vCprrofGCMWaVOSJ+8NhtkY8jLyKDyQzDFv
SQ3Zhqql5TMl8UtOdj9TxJvn01Tv57lEPAJjPdi5eW83H0s0VXzWml017b3Axa16B6/tt5BDvOdy
wgD6IUxZbHYh9mm2GA3dCRx4Ayx1aJN619ob8yU196oTPUS8F/0WGkO172UIh2Jr1aQAiqxC2iy3
Q3OR6yyEcnhh+Jzjbd7Am1i3giVtxsytnDbI/tZY2TDzSlpD4eAbAU1fccQIpuYV66zBEqO4Qpmi
opbiwRjZ0j6izgRz6rO6Wb2L34g4HTDNqNQec8uh+1iU3W3r3N1ri+WuK3xZO2Aqu8bgRc6XI1ng
JHBy7hCtzr+Y8S4joTvvPJmYZgZQkGsgvRm8kG5vq4zeL48Nk5vlx8VZI06Q/8Y6g583XO1JW8yv
K4GtX4kGXHVLPpbPz7jNA0KouNc4XTOn9eOKfEPkXnt9eKPGPFt4Dj2jmRyG98G4MaAjoLQ35ZVU
uZbns4se/Z98irhWD2jLb5VvayCjREtuYkruVEOQmpxJPP7+MYm/m6aQ7YHoGV2p415QdK8/s1lu
HSKZGLsdz40C+I7Go2RLP9ahU47Rpr2ymyRYWp7mTDVlfdCsCTFNG5TnNTv67TfAmn2YbXjoqLoh
fRnOsSg7Bid3UYHZSAoGcfjWcMAVnpgD1divnW3VfvxNQu570dCQcBMg9kZT3NqGeAyAcV+4z09K
5YQdAgjQW7iv0lqkvYVtRjOtuVkVAe6S7zErP8hnwBEHUMz10qvbHByfXI603qLiH0OygJ1kyO9z
D745F2898sO5LLjK1FtADIyXCdGXAgzSSmsxi0+vM8vTvEXHZCU+6tIls8PPKjNiMZQI9FXAgEwH
RxZ27hwsFpZJAK8sFQpoqty+owalWEUVtEdOv2B0+JtOCAXQg93AJyu1QlMR9Xz2AWhzU3SCcylt
O8GTJcBu6/PL+UbBkvjVbxyLTdjd56O5ZwVzneX9dMID5n2tFmdhtboT10D5kDf3VPnKQXQFFJMV
1STEid/aKpIii9czTFeucM3sT0Yh2pcZ/R9mdV9pzRpNa7DeSG3HVBKDWnAa3dKj5HANuIv7gOxi
FQfRlW8/95jGjHoGXLzSOl+gU/2X+nxprbXp+dVP+x8vFMeLY1RvsF9ugsrFhnTnAkiUDB5/eYx+
/ZvUTjwoWmYS5SO/uLlfBftNDQA/jclLg/BDPBk/W/OO20OYJh+QJpzpFW3s9PS+lBL6yn1+zdaR
QT+nZSO3sEcosKtxFflEyUDg2/BRk92+pPkIO4OqsqNFgOb9X6TdYc1GaWhGsVIb4BBVpjI/aKdg
+Rs1+/we5UKAnVe8/Q5iJiWTsaZPrvkvQZsWOzaDfNbxohlBEzGcryRMblFsgcfKG+vl55lEQ2/w
e0f5EzgY0nMu2gsE96Utfxp++u9LazU3AWjV4d0WIGe2bdbo3aoc4hHiijwloxGK56We2tlQ/FrY
d1VGMpmUETmK1cT5Zzf9a9oUWHP24kWjaZ0620imCcoFweZ4G4ILZc4IzitarbTu7ZRfLY10CxpJ
lgh622KqkDpET6HqOgLl2uqWEifN85rr047Z+GhPEz/Fn081KV5aYKEy8uUs8TxX80hI4zfXEHgm
px5pgdjqnz0OvAJ9UtJrG+F5NTSATznAA0wKuPzdZKofB9BsdU+PFdQOaICPkl1IpTpKGHXC3Ibt
NLFlhXFG2BO4J/tCz7cvu6AgFpYTpAFrTMSiiQ1JHsoMlT5p+pUOSehnNgt5dfYCUzywJIxxp5oY
hT6EeNs7LV/US+mS7gMYJ8RukCrHEEbOje5eRCU1MWYI3RXcWK0ZC4uQDiAK+r1ojBoxBbCtnvBG
iFrrUyzf0Hp9SzlWBAQ9EgOaQHQDhia7prau55gxMcdHoH7N4EP8i7e1ShhyVpWten8R4Kgowmbl
Z1zmNd7xF7u3XOPsHRpFY+N5PcszCBeqQBb++QSMu/To5cZl3MpkaJZtFq+qYWEiMaNDlG5Y/zNK
jWgfAGtp0UyuPphq8CC1lByrGhsQ6nq6b7RQvZs0eFMgnU24oAhjXyotsbQjrWRdDtwtNeJvPFZu
W4WSBABGa5nRJzWagcis8Ar7FrBrgkbWQ0UV+LFBv0SEnWDLbnoY587hXMcpSvpqPvrvBBiOYj1Z
8k0+s4eOxwDxujbjX/kvesqbC7JYJei5M3cxRrSmoZCTCtvWtCFRNksrr4jsFIMDicox8KykrW2w
5KA4y+Lr7z+OJHiZLOuTmw8CDPqx0Q35ZSkFLWXAG8S/nh4ziZEJ733e/XmecD2vm4tRwyUPY3bD
6MnfnJ6NRgaeZN7ed8CrKSM6lVa2hD/0Uk6VPzlAxEFj/NhPqo10yOlpSV+njXnLtXSmTEVhMetF
N4BjtDhqgKtvkyoUdek11yPIvILMyqUVruwkgqQ69hnx3enGzUcK+LqS4nRfcSG446052G9lqRL1
B4o/e1XHLHgGve9f5YxcMA/FaJyhzTm64fB999d+reXrsABhNurCuKhXmrCBx3mIfni9telV+k/h
9Vg+uyTvUaDhwCGDirIrgnGdU30iFyBVXoVeDA7BdcgpekpJGT596OVF7XVBIWzmuizVu2hcopn0
LEdY0aYgIfRA+nSEtsINWmLuiMtvsiarqJXVZjvfN6/2cH6JQsxW4Ae5uq1b50juYrt9MhYhugiL
nOim/PhWqVWdnG92Pv5MG+DWVLflvfHerOAuXOLUD6Bt9RNXMZLUNxZVGIh3rhwKaSTmKdnukH02
T7Aeu6P9KBy4CZTH5k8rphu/s9w3N9aUEw0pGaiRBkZAmNxiB1q+/Z2etgzmVeiPzrj5ToSRATsI
JTp8Ki+RHNIBajtQHWj11vyqlmNTcoB1VkIcsOXjhMhjj/lt9/AN5Tb2K+frFSBiZtQ2wFryXS6r
OBeKG5Zp38AK8byJQsumZtv7NrhO1ENu7ehLYDl4//JzKsH395Msk/6cPX3wL9RjSPeoYWsXOACj
wv1c8rWQWPgUx0ZJ1BPAvy9uMDxeSnF+j/8Ayg2GdSkhs1vwBpxYHH7sqSg8umwO9beb5TWckBy4
n1K8icvVXKlcUywdFwUrJ75GtTmrf7/IsC9rJ8CEy6hExIrla5RMH9zTkwEhHi1UlBvNubyOIR1t
fMsul+niIEy2tGWKZT93ECW5w2tgCtDg1D+orz42bYvhrYm5rFjxpeAPIy5LzdmSVyG8yi71hiqa
JeeelRK6CE9dA/Rn6A39W/8EvwrEH7zWilWfI40MC1kE2kDz/lppzcMW/MATnpwCziejgIqPU0zu
yTClwn9weJZmwDGl8oVZPnJwbjCcL2XcaJ5oA7PlWgWpO7nP6niOU2DYnlyI0bkPusp4P8j3F3F2
hAk5O30kYPFQN7TvEgSovvMl0D815vw9x1V2iUNxYjdix+SGvEpnZfE7gjcRG+aR6M6VjepzWXM1
qct0gogVdsCbuy8ZDOTvJQDcROSvsNCs6fAz5uozXnXlFMpUayjFiuzK8iOMudEhD+iZ3FVgdxi0
fDNIlSxMaUxSMmeaRqTrd7s3J9eMw3whiChrEcXcM2RCum2oMn9JlQSdGp01KcHrdJ+OWxWQOqwT
gyCMF/TwrQNQ9uS25mxmwguK/WAdaAodi0vPIoZkK+zPI6qNFu+6wDPM5SQOGVN+tvc6O2Twk56J
ffwhOGU33xVtuZRo3zbPPjTSlNn/UyltjtnwzRhhdH7aw4SbrRrZfjHldib2c9bSZPi7tG9ZYwUr
ldnCZY+zMTfIcSz3yQh3PA9kPNmMTN+gE4dwNwfz5fPdHlYOtcwg0WT++M/uGkcAKeZPIjt40fPv
A8zrx38sr2wWmF5NpwfhIlpgSZU5wMyH2s4rJECKviqkYvokF8cv6oaGRsfIvuRBqGdkjrZIVJ0P
xjCGhYK7VgM1bBNCz/bcnBb6tUGRX+M21ROGvMv6kN3hWsrOufbL1676HpDUhBYtVrT0nnwVns/W
BUKcEjiABHgw9uwIoHJPajPfe+ZEJ2fjjcNp0F1sGTHXIW2FunWJP9kBdwuaeWuGRW3wA1dffs/A
UAG48wha0yCEZQ8H+aNcuxC2LHJ8+IovmP3e09mwSBYVVcTcUrdWSHnFKOtFxB2l1cRaNH2U/cS9
tC+QySAgh0UfB6PmVji6FRolCBbdG/UCSi+KhcqIU/GDTZUYHs5mng9ReeEnGG2DaowLMiwaW3Ql
FwblO2ma6cU+95XecUTXMudKCYGO6SnC1eoFi7vPapb0UTXN6FFX6WVzdUtZOtf/bkU7JAvxqF+o
vhsP6DaPK/1MiM9ECUmPTI/zDhQ1BvtzWo+HhR56rkHfxV8pL22c8QxK0Z+0Ey7BFmFxczS8MD3o
L3e3OTyUDdMBCeHM6tE/KxA6urWIIZxPNaBxI1U4PncxEhw/j4/EeFvnx/iOj877HMkmff8Bx4mh
9KrEVh8oUHf1fKjx5QmactsbPB9k0v0vXK9Ll4onQReC1AvghKVbBGBYyOWD4PD6smM1kHPD8n5H
4v3CpWWAenp9ewDbKtraiOL2ScwFXWQVefGf9Cr7i/goOAh3CE7BEnFYTbBiWznIKO6sPLdht6Vv
QkduypWGs4vWU5YLRGGMVzgfxSMHd5Bu+3bQeMvhMNkzlPCYXf5zFgsN4O20tpmI+STYTLtVq16b
iEXiRtCAhi6kxjbAMddPzSR370IgRKUDMOt9AMGmUo8e4yOvWmD1NgtAhEns6Vm/IbiRmrsOYyLB
FcHVDECkCfdcvSjmZsANpt0oREQwJ0bQvHJmo58ggm/gXagKaOVVbvi9cqCE/e++YAered+Ly4Xi
hFbWDbmTqd/7btGKULIDMGB0zVy7sri4ZMgUcUaYd+T7bHNmtnFGzWEuwM3RGIlZMCvwrF+TrG9E
BVQMFAL+vZ6ZgtUyjE3V4sPYPFfbJkaGI/XKBclR/yCtGTOOMnzaDmH4mvY5+ClogcBq8SK9wjz8
qpjzWkxrPzzRvajXUsGhn2zPe+GeiwkABWQBUFfWfu2pZ2pvRBshj+2DpltrxDSyO5lcv7sZUco9
+4xFDXiW+YB/kqq2cJ0LVbivTXsOMPwtvViNP6il6/mnkL2qUBo9mlIGh8U5Co9/65RDTAxl9AP/
SayKAQkZL1OFRAhtx9sPuFGxhev0+o6ZdRwJBiB2rQdF6xHQT69aij+2DZ1sPeR/yZihRLQeXaiH
XAlb+bo4P4+4tgcqYQZTFyfF5PWGHvRDi9UOuW51xXhvCVjZvEbIFYcNV6+KDJ7tHNVPm1mihb7U
b4ll5Fpl+MsmJA/abywNXXLou4HcJxl+FxC5id9V/U61kDfAT2HTq8X+XB7K88BimMg/RH3nX9XV
WhPHEuRAuMw0BVn004R277eXjmGRoeT0ENQLFAHQ7+zg05a8RC9jKcd/zMiaoyiKciqIZtAWpKAR
cEOkzSBaSuI+2ugewMkOPv9T1UwTSUEeU1/8PdGpnbYf6j96ud3XpS2EYDzA0IDZe8HKo2e5Lc6J
o3os4oMg8KwASr9Qag5ynbSBwFEDZQPBce1GHjhd++uuGXYiGwbW6I1Q+izh03xslGI22OstnrL9
f+qMZLMoAz3cYmWGt5But9RQOtZyEcf2btZoyW6joDXgKZqVW/KmuNBQtYxBUQmhejKhnfPyaR+Q
ZwbUs+WcvUN2DIsjSyf9v7CimdsiBMh0U0ybuZ1vP4G0AhBUn0SFpHXhuH+mfMUXjCq7oeGLESDl
XssCOhzKkFsqPmAIBMih9eGkJ1rLIlU3hog7iseji98tW6Dz2H5wb70VOLz5Ok/lgqo9b/nGlvi+
oG/ESFUcn+IFyKumW9/FA9pQIbCksIcHfwVca6xaD8+yJIKC/XjmcMz7u5MsdpURUgSB7ZUD7N+v
KqUw/1pA0LfBPkOqWHJzzIoS7w4JM71rq6H1jFAtkmAz75uZYn/ENlYE17ywGN/t7vLC7KM16f4S
LV+58AiOSnRM+l/6RrdUw51ldf9d9PbBsM3nXCV58YvNWNYkmctDL9yyLKDh5Vs1YgToc213ugJ3
/OMWugCRbbWBi9qAmeCiSmtjRKcaoO00PcMwjf/6dKTCUJ/HPr7D57GWIPMuCNStStPNXtSaIPF6
OFYH4S2JC7KoFgiUBHa8JcODlh0ypCkU/kG6RKsvIln7IMlHzzIgGapIfYpjQbM+98Agda8sZ3J7
SLEHoc3ZU7DDRbB3F9YEDBbDokdYxMFHbsfqcBjVyV50LD5AeMwpgAHZAYoz2xU3kPN/fijeeHj9
AWwARkko6peXelpnDOTm4/a09HV58divt+KVJgJaA9tB3QC7KKj9PPjn2QWJtYOju0KtzjCGmwWR
NPS/IbrFuXZSh2MSd+Ic2prLvvM6/QHJY3OyPaZ2mUtI/ecfIkHo2hQRirD8BkVq3+isDMQVYavP
dsRDIDThiyzxtqTuVxQYjpLCJioCHOmXpgivLu02qUipZyBIIqQM1kiN+v0MFOeetDVdfG3ml2i9
TmXMTqhJErEsJNQBT8Ro/knDjgm8/JqlW2KWmgiRkK/9YcPkLx90IBQ5IJu4nd+cs0cjWoXgqmNB
dDFvBp9irbfcGZKfn0I92MkFL5OnU56MFOa38fjuW+lbk3Gte/2kk0oRiTujmpRoCZRaVZ7UI5WU
KgpAUOahYhDoU3ulNdPWOuOuMpU8U5h1FRiL56YLB/MDF2QeekEbuNNI5c7NmXSeusEX/epj7KJf
k+O5v0dSaPV1X3BtPFSgidBbCof3kA06mjd4NSYo4g5YogYWajSXHP8UxF1kc6E2byhKfAf+taln
oL18m8uQOURz7VpUgWOu4zMXSGiLbixn560wyCxnrbKhvcYBXwVSHFrD2o7cTlDq+s7y7aO+qRT6
l6FOS8ygaqaYc+I2J5L9QSRxS88jl+gLNvx/JkqGo9+3aFEg9HWEXWa2FR8EoL2W3Nlnv3owyK9m
/COPlBr2QqzP8wjgy5/VfLJWgsayMcwRZlJAFn0K6zg9/V8Spk6Wa/6h8e9m9rwdm9aK2XKrrXuy
bI6Qa2UHowk2YlvCr7XF5fcPv5Wlw+eXjDOtu8wboKMuqqWAC3NEzVa2MfyCxyD8oE7IwtcQXe6b
m3IUlLgRhRQjMghl2izsiNuQGw+Ilh+lJlt2kU4ZJQbghXplLPWoD6oQEKbn0f80/wzWDuo58F1q
qjskzxqXc3R+75c9uzuQrUm0FnuRfqXx7bI9zPjAzJPM8zOvvQMyKcPxcl5Zxn03p0NicD9Qaz2t
aU4uZ+AgzSIHt5+0MyRvwMiSNXr/kQ1IruWOjAYupptgViW1v/GcmnXIp9yNZky587sOY4XonxeB
xgszvw2vbyzlg0c7H8HWv8QghiqtSeAwM1pXk482Mlj/QDW3+IGa9pjjM8PR15Qd3yMKkIdM6WnE
naZF6HZS7xODpvlArbEp4mplv1/BAWa1ZT6ApL1TQmCWNHpsu4+U1HxChOkYgv2K+/nl+ODsfaY2
77tNbr6/5h1z3rtNYzS0O0+jCbgSZmIUK5yJCElcWUb9n5/xRbLNwQ9gU06VQZ6/fksF+inuQM8I
/RghAvjeh3PDkVsQu47IP20HNB9kmS/Vdc29cZiMMQaEE1j5FJlRbX/QUVjnBSQjl16vqRzpNUCg
cWHDvaamCy+TJhmE+tEADw6ibp0d6JwggNbDqYZwBUbM8M2cowRr9vf+UFjTpFTcwRW//BWhl0oS
2/U3bNUk6Q+Ru1guzGUmyCgeHxpA6GJGiTOpuJYD+CjfQdycuLzfHneuOwtcB/CQNOTcCG95cfIQ
ncZxEvAcvir6kXlaztAzL6Wd6Igl0KOb/gUZpFtz4w3ir5GUqv4Q96OZAacLGsjKABVHWZldkFUQ
E5qIzZeIcHDn/r7EXGpxy9G9ChyupN2m+4Uoin5w5H4xmLp24meyR61n57oNcweE+RRyLs4vuQOD
hgUDEYcFhS8UAHdTqWEyI/clJ05weE4ngKOB0BT5ItaAuwwCBjj4vddfDmUv4LAexSk5HcWl6uD0
UAsEmdavqEff25g6KC+BShg+Y4fcYrkkUd2srDC1aRpOz7ck88oUehVruigp/j9y/hYhvyFPNooa
pOUNAqHl9+AfseCAs4awhmw3J/yBesHMBLAEjdSqlbzXUg5t+oeSNfS8zW0VyUp/TjowtR84EAJO
YN45iNbJv1KgMnDFAeZvSRMmVTsqFo45uC4cX0+NYSpHdhIoVDeEtYinYphTH/0OUDa8dbejbCfF
2q1dQm/A5aybBWXuidZeDrCw6nYX32qdif/i7JPVd+mZIr5+9RMxns76uZu4cVpB3Sai8BKgDMKZ
huxenLIretVocGS/fdxxgTNRo0foxMxS0dWpMRY8zq74o4weyxsALizyvYGHhCYB27TX4lzueeJY
wAfS1DXZcQdxojkIS91mZIe2IRCsTVMhfetBFHOJBRZUTIOyOhr4YSNy4EkwvQ1H0y/VQwW555T8
z+zEevtxt99WkQMpUEj9GpyN+eGHbFUgZeje2TuF8VJ3OIz2G/187Yx3RmhErGdVQo3jOFMRExSS
Xvz3a1gnbmc5CLOWst7HLdyOezJD3Fjxr7hVdl5HHPyE66P7rN8f15Pz+Y2ShNi50qfZ0MMEUgZK
rnbNzB81twDZWpXgGLq5K5QfzGD+MxMtVMkywf/SG4knxvBL8IHkVIkK3V8f55qvc2KQYw9XvTBD
c18sfFTuryr6TxiwOgB1GfAwHd1LfcIx2l5dxudplKTM2Dgcp2R0vvdjtCo4GfgRWEvrEZnU+kpq
CKiXifkoY6r/2M+BAkhCGEsGfVcFpcb1I7QG7YlYJ+uK9igLvsoB/GkbbXTyuo0OuRv5VLGexFff
B8J9KY0tf8cwpM8axonH20QIsHbD669LW4eGHEkjEoN9B3qdIh+2N5ioF+8T8DPLQxW+HCAwiBPR
i/eqzGQJVtnlGpI6FCM9ubKtlE6e73gRoMUirmzWNkKr9MewN5h6S5YSF/z40KLOvwPX9vvCe74t
Lmp/sy68z5PkDnuaOowzpu98Ol8QLqXGE8RqpRp4OGSo0r7BIQgfEAve4CnnU4l77ylQ9hgoC5Wr
BUzAGiTYSNkO0veNVa4fQ/+tje0JHPcUBLoGlFa9Phn7JQNIdx2HLjd7I1qlb9uF6MY3r3RyfQYV
cpGvHLJKSUrGYjIN0dJmLgD4UnXgFgj/khYSEIsDkveK3aEp97GcNFOJgqsJkfXQLRlg80LG+nRy
lg7VZ5/P6AAyy798uf0/Wvc5nKFCI7SPhqdQoo1XWvXV5lD5StPWZ1fIV39MyxPtIfTuXJ4ac3ms
wQwY9/n3gAwGXN1vvqrTnOBbCtBsq55Yc72QHNYTseA9mF/fJyVmURrQ/aUpkwRz2BFZ+laXj1nD
vRWILMPGUQPAQnlbNZo6Ie3GIp7hJ8m1FJQnMLGukEqmoVR8HGJgmBEr6z4PdlCsgXnb2/GYaUdq
NxBeZQoaAtulL8QW+h38q9fJcGbQ2+gJAJYbKcdj1C4msVaEMTHu1pz2ChQ4RLPoUluT1x7/S/Ag
nPWZ4ixL5Hh0qEGQKlrzgewkrIdY8K+ruHKYY0GATFd6rJjskS1cJLorJA6785prQ6q8YLDL47Nl
GxgKohd7+p9Y4/gJmb259fcDcko/yPtM0W2M9FQnWNxaIT44vmxPrjQcHmKEOdbpyXfRic0Rjrxe
0VDHXKy6e9/YOTPgvWIm1ZnPxtF7Q52sG4bJCPK3mDlo62thBC+HM4c3EbgL+PinP/UaLhWEskDE
Z9CJzx3XkMwZLPgBlR1BfNO+wOcXN+oQylkwdXYP5NhcuJceup26lwJqhwXTqR6oeirH6GrLYzED
G9BTOa30Tmo9zZgHUL+LjBDzqiu+FExO6Iff5LcC2xLYTK+jXIQKycivya/jeUwquVfKMLBJDDeX
U/bYTrx6MUDREJ12VEsy51Tz3quRal2+fCLQg79Smle1J388GHR7xPbLMK9bxezoXOgbNfyjplkV
Vb9Dd94bnNgoW9fRH2OHDtr/gtjCs63Az2p8RoLo83bgm/kDPznem3g0RkfbdmV3d+bMRamw0Jp6
elMpJDY4ajC3lt/XtmVbTlkk6FCAvLDM6yN64pRiwAt5VRFgcdvtjOCeSkaQ+fbcwC9+bdR8IZME
sGga4Kh7DdYIwzqofijxbrtNjgyOe/gXGzTD/ztArMKN9V0zEZefSr4t5yAG7oCCaZSA2dp8qO9Y
ZQsNBISv3GdMV1tZTdPeSdLh4zMG9HC+0NiKrwjY+FV4VY/l3a/6QpQCubmVwCerL1wkqL9FCbOj
ZgapLErinefq6AbZ0DbX3BxjpJaGjL78V+Z7vZCAzQbXhpDUO5XozdHvpODJeTOXjyyUDBsYTmyM
3WLbEheLvwUTiTazSKFhEvOPXceyrYvdXCPpJbJGQqwHshYRxwVDHnqOQvP9OHj37Zqq06TJK4d1
gew+R3o9+eaobzZxFhK3ulvDxKfw9jt7xzGMZrpUV1KvsqUf90rxBYZ7hEi3bcUmLTylHSneStgc
wEaZvkosAJoGSzWcmb+WaPNPAbnJ/qUyXIC4DlBpfxqNAyKpPyVuGG74QGb5K5jQ/cBtc9BNxgQF
WnAFBS6fgDnDsh20Vasj0v2mxaMYAMCjFVSztnAVQQzpIKNRpW2dQAGcITULz4c9LHsD4XHCJLn8
kS0DL+s40yQ29vHa717t6Iy8perRBXc48pNrCNmP9LkX+h8LcpX/I2/LIdZplquQMHzbwo/UIhCx
n4/8NH8qPs1f7Kip+c7ygI8ERsdUJEf8RQoi+NGAg8VqvBlRIpMMMevXhvDP1b03k7nQjRPKqi3P
VN7ThyNynBufim6mboinx2u8676pqYBens6pZIUVKQXBdPamPLZQVX4EXboJ2GkCY5UWrwphD9zr
LXurdvMtrA4yKlo12A4DYeD37bScMBkoW6sIQ9Yda1IfzvUJEjOrPm4GbBETBGaXvDKPNGBYs34Y
Mul1Ryi9pvHkr4Z0CzSe4c1hwe5yhQ7ccUPgjxP3UqasEXkCKvZqYv6SxLf3XPIT/BV07I+5sHu3
hJ6yVq79lG3BuzMvmB44PnDkagStdaJBRkXOo+uKkHadwGVE2veRl9jkJrc5MJU9cPsH9goe0vVI
O/m9k/LjY5CpekG4keEf0/su8iV/gfcST5TWpPLeWKRDKkX1PfdN4syZ0TKOj6yyLjtQ7f23gN4Z
DnANCqg6zPN8bTb7Busxn/iaJV0InPn7xpKrb2LPMz3EI3D7xFIHdPJpwxdd0+1LjPUdPWfRaZnh
MR1/nBLs3shVB0AhRBJqsXBMA/AFoHmn2ag3KRFmgLyNE3k01+oAj2mjXIi0V5CO0CzbHvBvXurg
Ax6bmvvgs7jY/KRbSkbqDnkOWnG61l1v8t5yvcBiWgw1dny9Kanq3kWvi+OjVuSF/TvmQnIYPKtX
LXCHZ+426Yw/g0R0L6z0Pwce5H2VnpJZusHPcXtrR/67/StNT3EM7j1HgbhJxqsYwi7gkI6Ib508
ZO62dGWNuTo7uxUdn84Ppp8XwFa0jpsV+GIOD9ztRbalvv8nizS+Z3Z6pijsvrb5Yo+EgC4f/ewL
wah2xhr9tZiCsPzPMSl6tYOY6Ewm1IUF6Dw85yeWe3knyoXv9yZ94NRjvBZQgqUzfxO85CwiOg9i
C5SxpEbvUQ2VC452ErINovOv9zsWIaVac1/Wia7D+xzMEnsrPDz33cNkPeSrZ4KMecnxRwDLDaA1
ljAwjHowFEszYqRvERqupwTWiOKvVE+USRBCzdzeXtxERT4Gre5iQuOaIFDGZL28Q7kbw2p918Bc
J0jUAfGaIGV1N42HTKGXKReRYQG1Bkx2wUHxfTcM8ncPvzDiWcZ/xMenIc8jH+BvsM1AA/54c+vo
Mp1ijabOLi0NKi7CPADzeZDNIDEyPrvGeJZ0xaHJRdWpTR3e9Jbmzz4r0fYo++TayjpNP9QAEN5z
2jcRFQXC/W8udK/RPQwm6QFCOzuNa33nD8w1AoosACaXu2UjdbGmR55dWZIODvIL+EmhXWIKj5Iy
e1YOCra4UspzedV/Q6n88kmIwAvCxzmKWS8EpfuYYLfgqNu4iZCKcXdcQgN5MXzzV3N1UJSYnbLc
PLsqCqp2xPwU8AaLhhwJ8X94nXtbVxP8PhB79Kwwx9Higtsge4Sinayh3E8QjqweOjj1qDaGYd6j
Vrdvol2gUvD3FAr6J75wbpsQzsRo7XB9v/vis+Kqz9KTm8zPryvRZf/qaqEql6O4s2+lijAiPkNh
dyZvghpOCkWBPofIhN4rd+3BgwExdB2bz/6/Y/mSsiNx9k6oanyv/8z2I4BsgZMS+sUk7w9iBgXv
L4Nc5+p65W/gzuKphfTo/a+G3OGVG0KpRzqa7e9rbBoypVRCyXAiT4ICpsNDYIL78rP/kPydLF+i
d/hyqoDzwXpcZvBVaZzciBoQRxoYDb1rbjGSxVjOBG9jr3qUy4vsoZUGJhgCFOyvF8Yism16jbXS
E64qzy9DEBMIr/geZAAvA7fB4bJunMMLUwmU2Je3ov8QFa4eHMcXMLY4NlCZZivy1kDxA4j/LAml
vV0gnzo7uE11eoCKcog6KISt+ymWCy/iafx2LZD7zgQptty6SC8FLmJk7Yh4ZrTe2NrDYb1Fm37I
sCyg0YTW0K0aaxChzaLLDlWerLq7H+OxSGevtquHl5ktVbpePX35PDJvWH57BIOtDELGzWXd6RlD
N90dmzxhsSy8oJknRlzlsZ4vnQp0RLT97jWU2FuOERcKgtgaraovg+R7noghUvxkOn09N8GL/DmF
jaFmNKMzhAsIbZOsn9a1HweIDWZrwNKCO0NZvu2c/g2HNcFD+Nf5z3cNI61aJSIUzedvJJLWayJk
/zdv/uqF8e0MKoCBxWW+oFl6MjvDC33HVTDeYVi0xBWqz7A6pidludygQqer3aXvcjG+V0LVuZ5j
nYVCdh/3251nRgwFExsszeJP7aKdTun1vBBumTQzC4z3TZLZh8/yhF1txXtQTHgvcEZafu9q3mox
NEuRj2Qy4vdHIYlH+5/qTa4Pv/MQW85NjCDN8KZFMwETsSPuDCEti5QUWjs1xLlNP7eD+BCRCgLk
HwKyviaIuZ//ylTqDrkLJJ6f360LI8GSYiQiYGyaw0czwkkin14SuU14uHOFdZawz+KPyS7Giol0
+ZaXO3ke6QeiJRjzLtFzhvyvwkn07ZMGdTYi8xvsnP68Pi9yc/EwSz8tQuQIpkUy1NBbMNeoRwm5
RazpioWjDKEW7q6REuLxbB/CKQMVuGcr+1Y5lgvMCQZm5yn9DlBE1nPR5uej6bd8M35TGyXNwgBO
2rO8knQ+gth4KOSQXfHWfx2bxYYpUSMdROKIYb0DPL563LQGrBwX/yj85ePhM1G5WPjZfayJiep+
fJYC9kyrutsW3WvZetEXEw3gaHZ35LRScicOo2l40ZCndHCZqIGJvV43nzbLswWulpFPzC0vxvoq
IZhc6zJ8Xu7V6gEvpo4rKyFLUlNhOHaBK0yV3DXGI+nWamtjiT4W/+MvOxG7/XSaZd2oqNVzuh4i
qOo9zeaatOqaPXbUwZJkhzicvDYc5mi8JWzvfVgsb4sJVwBpNuGyW00PxkZLyvnkIvoE79KKotut
5LYYw5E4h3hC23MYLqzX2LxCBIlCd8smqVKJvNsiBkwcky2eQPR1EmJyY7TXScUzL8N30tCVNsMY
3S/wxgKDxwsvfSBtInojJga12LLvIFVZjqRRNckF6YeKUuBz4oe0lMUSgAVfkr6qw5iNawwyREYX
zwKlM7/ou1T05csUxNDwqYVdaGMNAssJvOEXmGoIZFxWpAxHltfykBLyB40U0ZV3wdxHFZ2C0gPf
w/UHHbWpEQVI5iGfocgMrSi238tSEwMeM9Rm64QlBhxrrpfukX59tNpEsi/i1bsd1K3ChgShMd+f
2pqbcejq8j5XvUJWI1ScwOjukIz/2xqgfhX1yEv1oHF2MoSqUuvujLbB+C/VJb6tNymuvfw0YyEl
Az5mAbcb9eoiskZV67hB1LkxJrJiwIQ6g80aj0/fq88W4EsVAehh4+YOOIdF08HaZRfI0M1xcQ8p
1IDfj3ZBkaX/XedE0gLHOicihqvBCIeMREp2gzpEa3rcqWncE1vZp87PPDoraPSEMgKc6lvS0zTS
HxbHdiHbXgTUauaR+B2iRTasAb8tMqPbMhP9j1altE/M1IBglpXOYP6WRNJTaG7pkGxiJWIiAu+H
cqhvvf5ob1hYw/ELKTxA+kseF4JIxfB+EMSCLoYsb4Dm2keigj78CBAbAuyXZ5alc0hCM9TAhd1Q
B4jxtTZ7b/p9iigE/KsnqIt1QgdNRKVAPqxjPPNiMm2mFLZKjPPGHVbjdNB79ttfi5idxUmqS4HC
7Pmly2h2jOnfv1VVJkawKv3MovH3IJzefYpDKTgcpLia11t+DTqtWHvL+TNGf1Cs+tXAEZVFN/YC
1hRVKsAZx72+VScFy28HuU3td2TyVyG+hQVIOoNgf30HZ3bu6TuNh0kIMKNefQwCob23xg23oWis
wK7y7hJLB5h6yvNLaNv6oJKAB1yMINfLSbiQMwbbB6RpvdRg9WnC2rxw8eUyrM5YmzQDqRzyJ6th
zDANyXMF6kS6C8fmnBimuNQYD3tby7hYx7idat4qLQcdM1kTlhRU5CU0yYnvDFiKOkisGF8juK4a
VwwQQ/TylOZM7OTpv6N2zsleK0fVFPRi7o3AZLurvvsX0VgCQgpdOYBL4E0yP9bkYbsKop1ngETR
BsB+n/EmjWFcSN34IZTIZP79jpBWvcVFPHQQOr76+UVEEaW4D7pX4mNurG7LrUS1YTbhZ7+QTZib
uVwhQrCFgT3UUpfWVFnomCfdCt7Kf71/O9muXg1xepBj12QBsbxTyQPbrc8iHOi/faXS6SHLYrsI
e6ux0cvnK8KvGPc6SrHI7/KqAwuprapfRucmo7k7ZI9nFMWr+M7tT6i7aTFUz+mjt0mWxvX4O3+8
MAYYqK8gRY0nYFzO3fMFn40yYXQb1ZwlAWoFKjpBdQzSgDyAyn7D+sYOeq7WgBZ6nKVBn0OxiagK
hrhkWEla2/NMdqBQvzjKFa+WSE1UnkFkUJcu3aAKSrDrumHOXECBTAtCcR1l/JscztzGI/kRUme2
007j+Xydbfq/YkV3tS1fbcPcyEd0zfRc7reFu73r+tPaek9va9sXeN3nJjn2AKgQMKr1Z/DDtl1U
34C2MJXl0vrTPRyX2kgw9AknHBDQqcNuI8bJmvj2M0eQqsqeg4GFJM1ENvmhVKu6QZ+6O046+hYO
LYh04fZPVJkKE5bIOT8bZUm0eErztgcP3o2I89YgiZqjVMjqFQhCeEFKT7kal2+L18KwHvS3lzB1
q4wK2BQVORsWG5PV7oj5NwFKOHc7CmoEc6G+tci4A7A29BxdrzPfYctgFZ4aHExo95PFtg7FcJO3
cRbf43Y1Ry9ogOE/B5QsQhI8AdSZAXP/0FU6dsH2WCFOmlKESVgT5d2Ootcktx1DrkVmCXEJi/hw
KZApGDI35KPP1ZJj9I9o6h8cCBqplybIrN3Se04Vvcr0RCffFuK02co+A+80cunwH1+YPgBQ9pjh
1p8a+uQ6ky5V9Wb9DzZ92sA3zoFHjTL8czmy/BsAGtknBURf1YtvJEMWfmBQEHAWHBJyxFXZAsTj
wV0iUS59mPv/Wewlg6JzQaLCfsRss3p/aH1DFI+iJd6r3WOvezcAPMan6m6kbPdo1VrAWbrVSF1T
JHLPU3YlYOOyhQgU2GPmApYsvKbB5kpBBNQ04dH2DD3ASan/temtBQFK3s6EbWqk/ee2igDcgfl9
OlK4hAYevGN2gNVQk0fOVcZxX4PgnqPJL9JDdgs9Z7jqM9Pjsv3COSlnYy+cU62GJFwmJ1H1tX3A
+SlMD8602h8FeGY6ymFZqMZpMkJy7n7uMKSFVbXYC3CS3AxIjljzL5fqH6o0yb07KuRIzHPTRz8F
BiZlmcwAERj0zT7wnmIm62BxZiXHtGqWVSHKse+UyjKIJKHefJXwV9vfXNJrwSla3/La2j21vEss
9lq6RhQi0RNKWNY/n1eVnR5t06wndbts8QC5WauS8KCImxETP/Hxdp4UCyJ2kSKejISRsif88FnE
H1tW0b71WXE8LJP+Ph22lSPiTidFp4qhV+AH7f54dhY+HNRQCyAwh42u0S+AOkBbgOSOYoAWiJD/
4gJFq6PieLCaV97US8ahijK7gvj3/lq19clP/mWnudnsvqljRUm/Ie2qrasy9fjuAQfONLewt8l9
B7ckYrW12VjEaRou63Uy6KVPI7YMAE1Osrj0yIbrUB+uXoeobzh9J786l7o36XoFuoh0KJT/53Ga
Qg0npFmIcjV047pbyzir3dT40hsElKW8QsY9hBhlvY+1wTsv9nFOg85KiQYs1TDgydNdEvouyqU2
o6+yciSbn4zp9WJ6qOB08RMNTSoXc4ewHHtCVd0HSFZcPm617fmMM7dHoxVrGYBA0l92+udtVzV+
FYkNVLUEkCfGJ1S1ev66KcZtrWRH5H33JueDuBnZH+JmV8t13D3NXiBA+ydghiqkcJN2uAB886SN
a1nxiahouL0d414NP+A9r2a2gAXncjIwBXIvjhdlBrTDdsCyUBKncJqAzcEPUJVo/jZG4EwBj36r
MJVNKZML03Bkd3BpzFE4vlwP0NZELu1Y3WNgikSbtrTVYXAXZCbfwRXtlIKgLokmteOkHvZOAVTN
UyXe1g1tpl69pZIklvw4PE5ohX46pZdPff2hANeus5WuBkZQUMJ2iMjojqAXhGmedGqNNHuN+cmA
3MuO+8MJfqs9JqMTU/1c5Ntp9Py2+V1ePunF0ypKGqZ3s9ZUwkceZWQfUng3jaio8u860KbETnT4
b4kQkqRchKRl37WGpGB57f27wsXrJrjNiG6MXaAY74239+3pxLYHGOjaHa6YtIzLItV/PXvIrsz5
36s7CVHHziRDkfDWzU9c2n5Z3fDeMyae4ifPsLWSCQWXt2HuYPWb+9MaBR5a7qBM+Mhwpa41TTF6
560kJjdFgNdYKR6FE/BIxmPyac5ok/j5XNwZasty/9Bdc+NOwYu8Gi9aoO5yYv9t6GCvVu5A2Xpm
u3BzjTn0as5NysZGBZYucjyMieMYCi+7IFx497wHWD5q6H3ZXcgQB+hSA16VFD4qHBishFDTzMSB
FrIgGbAiqSfL7nD6PW/tUgSQp5AuILr403CrgmtKpxkVT789j9zKIiYnlk+c91CeL+6DR4mLWB04
C/qrrQyam/zXdtL+Vl9GBOZT0JfwFuqzOD0qGzMX6JH8nBhs2Q0SOxdwzEQimlr4HbNRuAR7gHl4
ydvHiRXqOoMYSVFwaiFNDfcfTAy0f4bRy6a+WTAtGmSw0lCcLMNITmWTYB1zlu6KfyYg9H0c2y7k
y7/FvepIJECRW/5ruUJUXOn6i3ESqBeMYS8AQvjQFaUYwQBa0CiJHl4ulKAhqtQn+0E9sdef1OGp
rYbBLgp2IY3AaeP5Tjtmf33LDCVvbdxzi9LCrKU8+FGiDdtbBf6VZSrDWwgJ2tHNk0aIItBxaFYF
Ehif9QLSu+DSDXlzRfEVnHgTD/WeXmtlHvBhVzuI37CyJ3YvuWC1S/EvdWyXy9Dp1sbLTi4j/Xs3
iS2xS9FliGZecK/5IwPElijwERuZMO4x8ySYh6LDRlLSlCUba8PLQmn6ozUwGZie8rYkx+UBCGJO
q5uSXaWuTfLNsWkMBi9gzkhYDbIEsXBOF1LJOuP+YROVdAPGhyltpuE1qhRaJ9Z4OXqljOkNKAZx
P2qhilOU6dVbxklXZz9rzN1ZkcFh6ej7z1bXUofpknEAgfRzichjdk/6QBwcFoswLt0TCQEgpDh0
Q/597tngzMgAL7WQBnsdzvfU9zcZhOjJTNhG5Rc1/Lxcra0p/SYbfGxkLcEotyes6wfleMzIa/1f
qkae8VNY0Xi/Y+W2m1J6aCzkZMTAd8mHMOWBblKw+9BUtTvmMT3ToODTl4e8cczbW6HoqczguieE
ammRwZpxW/q4iON3b5jkedh2Xaeb1tv0oqOeysyDevNLf+jf2jliEAXMQA6DkM0DYizhDRHJuRG5
MumTUiZgB3PMbON2UqmIOsyQbupIyTl78SxgAhWioDsvhpctIxAaRmkLcrKoZ0wd+ZcMZ2TNHTn5
33xGBwn7f+SZhLyXH5o+JqPGwKCwe8Zr5Wn9ArLM/uWxqhK7B36px/ARUC4kuaYkWJf5fYNjJjr8
QzdN58SJrayOUGwtViicEYBlJnHRxrCSTUPw1xusogYVFloVN8yyZ9waFwHc9bgENM1/Xs40vvgU
HanvB8mwTRQOHoNujzajTNYu+m2BP+2oYV8LJeTYUPWmc150IQNwnlli89KRFs7T7EolYA757Af3
adcFvmXPjlxuEJMJNmia8ENzJtnudXMSpYGp8il3riKGy0MnCpwgXhgaGvxAjG+x+ZMzu8xbNmjA
jTdfQHXVPGjLarM4oWs1ynxhvl0K1KS4EsYOdIog073uy/swbyMgGlgX48lygH6wn5qqmPYJfxax
MFM630KMvVYjqylgLuEuLPogwDgCNwduYV3NFHcNvjY3T6xOlO8WbLjDi9LYqZJgURJbHg6HRT+h
d1hb1cJlFN6wMUPcg5wNr8PNQdNpxhf5lbEJ9bLir0er2UuJ/GRrTL73Qj1fFZdowvJ/MMoRPTsO
W5vRHgBxeZ5mE9YTw04XL1Bn7fhS7MJ9NmcDVptGWzEPxo8Cq5SkL7e5Pi2wNCE6fzPmmt745jXU
wIf257C0utyxVGZrD+BH/bZgC/nCNkhlSjA9xZBHWA/n36HkAxKDnhEirJ0ubxsBF5udkCZAihgt
awDHmrFP/cOHcYvslBu2KMBSMaNPBtH8iTvYoK/bMYJ5wFiCgX1Gxg0yeeeXniOP4wUpPNIgbc4y
pbnZ3oCpuYmpiUSSc/8npNM/F6iVUxQBI1PCqPMqb1vYQY96m6lbzMeqARNML2OHOkgi1Fvgk7/U
Dny8QGzUKtJ0uawhK+mJ9VoWkw6JlJMk15mKetivyWB8EUvl3EpAkhpvd/gL4ITIJdVqL4f4f2pm
I4Zv6DRYc3TIYViYs3LTc/+oc4mCeCq2vmz98xerixPP2/u05evb+qXsk9h8DmFpRIsTaPpp/X8D
6a/fewScqua/zLpex0Aq9NqIOsUptcF6zk3LiMxmqodk5NTB1Zxy7igPYebmrpwbBMx2sZFo7ish
j0DOMSmeueg5FT1QMDY+XQxGtc1E/zexGKdBKK6kod32L0X639dmZEmBjrx9zz1akQV77vMyYp58
fPm9pqVC5ucmVX/UWMRSHOr01A/aUd0tYMsJM4wvqJohSet6rTLOC5KGZxVqqtK5/GYgJxCHw1uQ
M3L5he6kINljemQjtGFy2laHJOBS2L4kh/oF3NNsy12+4xL5YrdnpSwowJciHhJRYrcGuleGg9H1
P04czsMzG83t512gxReIk8xgHRO3zOXUxJM816gFTZZLfLSwZbZsfhHI4OnQLuIPcv4DwpvRcQ61
D6duTQ5vIbnwnNC8r2JU4Q/t1D5lIMF6/OJsP/jd6035B7yzkD+HAzpB61sjHQLv3cd3isPsNkI9
eiPMGMXqKwgoJH4hPjStj1Oeq3K6aNZSn+vt3cVS2VpHUn/P9hTxEBp7cGGpGwsOi6T9v/KrKpSi
jTQXeWl1xAk2DGapdyMNt9TjYqflK8m93o+xFBUK+a0K8ncZQeKFPqJP2NxrCOHt0F3Kb08IZaHt
gKyqxE9/LyceSVuWyHKhRzhJflnx+1Dm5Edo/VzbtCPFeqlb/7QVtPEgbNo4dH+nOeFeGnSHQq/8
eAnuxJlbM1DA7Z1dKU/NbkEkjgGc2D3fnb+tEKt0bIUd2tZSgStcrcbrL4miWT4A+glS6E9CGgos
GMciJafpR7M0P7uhNPC/AZB/Q1VP6yEBUbFa8HZUXXMA2jibowv1IWu0ZenupoUT9uf5nQsJDWnL
nOsT1TrwI99k8BiHhsJOK9mqoRsb8g/t1tLDAFIY7bcaTKpi33U9YPLTp4yqjG9D/MxLsJjTmJkA
EwKC7GQfXcux785EzZ5Hh2lwP0hp5xiAAOmqy44/mANwMqXUGwJz1BSDzkD0E4sKFgQVjQrfXzTZ
wvLqwYZK2igYu9gHiWNIL77VheDKSwjQh2K+U0TPK5R8RNIng5nCDI0eIVxjZA48AfQMZMmrCeL1
+rI19xwKaJyTb65lkjS5HiNrZ3dhIpTfvp8hCqL+Q989+IVo6GSVAfFPaGp4j9bbKp2/u8g2guTI
g6eI6FGR2778TgQUMts2ULVCKkYX0ZpwjOyCFSKvSB274kfuQEC7arzN8t7N5/MuOibtVAZ2GDcJ
yKBSwcz0jB8SBosMj9xOG/l4dvMT55oHQImFTmSQQXFioHWFUUJpG5ku1mwBqniJzBARs2Jt3S6O
r2DGSSop+NspFwwr6wu67Pwy3dZlQ4PYDtrmTjXY/zk14JqNeVqLslKtfvFScJCS2q1BEjRJgJbZ
W3U3evJqC+YaJbGEBVXRnPoYd/xgYW79Z/tywqMRG6+BgXI3WHZ7mPaxrBxq0xoleYJnw/kkhSso
imwDsQfQnyZBDYgiJRcUKssAcYEKBtDAqLdrUtqIuDAK00ZSOa8kFk2GajN6Qhfv/s/5/4QdB1ir
KZg3dKnbeYVpj+yhszofPcR7DwohJXjz6xImClwkrsQ8ckgW2guLAmtDNFx7NuZXq13hDa/Szq4g
nRcFZshYepxRJWy4//8hJkQdGxtx2cp/4ojMOGdA8oDrMLjs8SmMSeYoFivroZPdwAQlxFUNHV6T
O3cpkNZ0GucFfmujK0U+xpxwprmWGu+XTRDsbn1lidEuTpZFCspDHZdLnvDoHO5a/2YxOaLtdXlM
9ILcfz6E8g02D7J2WjKsWWhQYD2OCB5oCCEaB6k91QE+iWKYr/FMLAm1zGgmfXOXBbvA1bMAIMZ+
aQ2dHHPO98A6IuZgmlqmJlqJa849yv3msNIE2suxdcInOvL8+9LoaUwyQF491U/5ZdbjOy/otAaI
ly0WdqjzJ1LRlg8O7yM8Rm81ltY1Qa6mFUAB0cz/8eOcHYklMHF/P/l7kdc+DhHm3A1ZtPFO+80J
G0tgCBHVW7zrFWgV+tOQUfDhbFyXKpkBfzpqr2N4Kcspylfr+TzuVwBL5RemH1rob4YSDhaIKK3I
iRfQAmmJElak3b9TjfinQSoQa4/N2ZtXcclT76h7lS5LHEmoXlvNxgnmbu7+A7467aEoJ0/Ec9vh
W4XUXn8nmdea1W4ew8JByeUvXsQzdfaR+OQZnzr4btfXJC+MJd1skwcpyDs4cMNkcDKwNXDmJ3i+
+/9g4rLQCJgnfCBYmn3bxq5Don6PgbGPz0ork8q/KsEsiXSKczM3K1hlQ9EWglfrhDzPhbdb5DjK
lhb5Xo4NpBsKvqtsZFS5An3rDrS8ij+DwrrWBBjJzUmUEN68fN+QRUcV49YXK68hUYRXGnrjlDfh
x8xiwI4CpiZoT+ZiQ7f4MiRfR80HKpzCtrX2j9J2xqYVsJrn23ddeLM/oE8E6NjqbR5iGLx+Sfgv
VfWWGC2e2tVSrGaU6woDSS0XIzJ/yJjH2YBG7jX30p27M/l2fIYIoS+NFQzqwG/Posn20Dk4+SeX
rHVPQ1SFPukQtCFyn33P0H9W6ciWr5GvGdysf8qZqcaZxlxAAvcDnEJz9GCvREY0uLpiC3CN1UFK
M1XPWZROkuwDirgNdNoCpWoAwe75L1g7UaRdrM/EM50uchdYXD6nS7txeinLKOGMYbxXF07M5ZS/
Orpivojaslu08ukGZ1J4nfdZ2NCOekrDl5OodY1oGr9clrFTcNxW54qyUkxUw3IYJdHMLnZHu1tM
OvOGQCP+yD9fEqiWaijaJZpRucxUj+HOrYkdBIZyEv+oJDOz+2M/lQrGcuErBGbiwCoHKfDQEWGu
Xisrbtf8NXbSKKzxpXB4a+juGl0yufSag83XvXz0AeQ+d0jGDt7BQxsRi0NAAHYjkGaGNUSVVCmB
tzownJx8havRpGwhuOzWyM64BogLXQS1Vzs94Xq/Svfwt7BMZvwiWw7YwVBG0XREeEhB8XrmLfgT
yh9wigZemU7Avz4iu7E1e5P7Ncfkuc7eIdhLG8L7zm6LgoxzAWYwGesSwG6bVzwDJr8VXN8jPmLJ
8d0AH0MngJLWwlzuI3pfLaobQqgz87RJ4t0ZvdhFYNcGv7QPf1G1UD6l41OIku0hE0pEIRlOTM1W
V39vauIAeciP7lWJJ65oqubpw/wTNVZX3cHEjaJNwvX4y6+cvR37rzjjAndmp5YCp9lsds2/eb1S
eHeGDjbYStrkYiv1xBj49eCYYnhcUzyVPKuGn+x73GLNcahiqDV4aoCsHHYKceIuUVaMzumvFJvT
sE1FmYXQ0ri4gRg8wstbQT3K04V8p423iwvgCKAfIcm+/gY4Oi5Js4tp5BZ5VsrNVpPyUjfTaLi8
V+tpvenZHWbkPcAw6DckLznDTuZP9mB4C78lsLhWWgUbzsopMvXdS3rHV+Xwr2rwk6hlJ5HxiQvw
pjnEm3OzL7S0bYt+XnckAS0TJjHSFE1to3CiRdlmJ04J92T5aDC3zxWgqXkNJAB+bCKKOoBewY8R
oRgsbZbGbKpkW6hzr0lJWySKr3elSf6eU1sVoitfzFmAS/Isjc49tbEOuuOSmef8ttixUg0Q7GhN
rvio1xw+L0xR/qCt5T668Jwp/5e/9IpNGx/ue88TUnSXYuuldM6iArtRUzJt8D8uqY6qvwrxfMZN
184Vih/VUBHmpE6aq8humAjxm3VdDfsiLe235tNK/Sp76vsjMzsL/RUrfewJ4MAgf/4xYcMFV0AT
pVdHIz9ymFUgMvfD2gSgi3oMKSGuiZJkD6dbskkaIkBh5FigkqOZ9qk/RK0zx7NfSLlBE95r+e7U
7ib/UfSlDfqby1lf0+0HjCMt4YbgADyBHKvnrgBkeYL9UqJ68OO6YG6ztObDGEbn9mdsmZYkWWmP
yFcrIdSC+iivx7mw9D8+U0K51eszyBRbEjUCo8xOn6YCyWI/sPyXqZjSZC5L9MiaU/eNyRnvheuB
Y8Sr2lAu/MKIwBJN8uNYaq31Qv7HYebsZo1kcg9+2JEXqVGhgdau4fGb8ElIcjwP/E5UaCisiaTV
n95otfFe/zcdJvDN2E7kEuJRNuiGrTwGdrZi7FDQIv4gLTMagOd3bkGXUuyY3hsKkhpuzXVTG2Fy
vMXSf9GokBxemnE+0MfmdiuQZdBznEayAc+SOLoMKl/4oacl9xaXRYJeP+ahPgXmsvGt1ynpOQ3L
WwDkD6n+5lVHH5viIde5v7s6gXS0GZXy7okns54RrstwaKMtn5qfA8ynVU5JA2d9aTv7QaQQJVvd
2oNhMy8vSk7p3VbukZy3hM79ucS2UUvKxmIKCiRd5fVK/oo7Yiyx0ajqKdr5QbZM7NeNRIA9BP/R
ujUSzF7q8lg57qzDGjqeIIDAMAaW0o7yf2nVr/u1Y8YpGL2k0k+9wnshtpGFuKc/Rn1SU3Uem/An
jtX5XKf0aPOEK88tsE2xjErmf1tH3z0Gu6PjqOrPe/SusnUIc20jNxFx6FAztcAGh0EQYp8096Dq
KMtkFfVtVbaJxg8M/pYmVwmegGDke5q6XY21958J8OEamgJHrygi9wiLfZd19tjD6xwwsL9GGy6i
ah6Qm8ls34GS+pxWDssQ8GpIgvEhRx4Ss0VY29/pHzW6mACod2xUAYCNP4j6heOEjvtIO7OUzFTI
vZJPkNp1VWEup7rHvXrnT8E27GZAK0upmeRd++W739YKTHt7sW2VB74OfoM8MDIETaAf3fTZERkZ
vZZL0IHjCIXjwf8TFiIyFiTl3J8eCc22wPQrhkxkcz8PAlE5ev5WZlUIUqvWKfnW/V5rm9Mi2LMx
bHD4K01+monxvDnobe+R3N5zUM2tIDA4XtGa52wsIkMwm1Dq9xV4LGi7lcNtrkPWTpEwj1TLeS/g
m527JAbdGVBH1no4ykgeTpXsPKCoO9sgxYkt4KmIA/keWooh4n+oYH15v9GOElHSbEb44ZJK9fp2
2/OOSwcqcx4Qo5ilayRuWVlw8HNUmBFxcnm6xFa2y+Wtljw7wmCIW+xn0/YwfVJmEfg20LkVUQse
bCGwRKaMH1nztlhb671vPCRc4F1SlrWhoZ3asc/U1wzhXuVO92/OdoOuXhvrr2ggenjXEbyvifT0
e/RMrnXqH3tHGqZhybAThO0zc8Cd/ZK9h9YwvYsGjSgMRfAP4rCMfcGJDdIdauBSTDArDogZpPGy
gBJR6BEoPSNW7Mra7EysFzYaf+mLBvnXInGfdAadN7vXd+fBlsm7p+qs/Cwojg8f7w1J2+3LFZlV
m/av1BqtEY4orG9UVCpHzjGMO8S+UChOK391/UICQaI+zf1ExZK6DEsg5UG4njIXYQumezXPXQcf
PO/0lgpgsQVnBwogFzWKu74E+CGAxv3wFKVK7yY+/UFFMypOtbWfv9ECiV/0SyMkDPY1rai88lNV
6eDDIychOsdcSxxM106P19WyMaBohCXEN26BJjFet11J07ZdAuBiOaTU0sDCL/ptB+UJ8Z+nXYwP
qW9gId9wwavy6Qxrx7OKvnef5DdD6kYVBKKPrSyzsPqwjZuDuFnKPsg+0ubwvYqbFHCwbhY+ekl4
OXSkwrk0J7PdXB++U6BljFNsu8fbpY940HNyOp2/Imh51dQINobbYOb5h9nhpZVF4TiSwd7+so7S
8btikWhvCrfj/fW1wz6yYWa44FnEQV7OCtPPTa9FGJ9t+U9HdDDkuBS+kxH5oQLe+HrEVy3XFTsw
I1/Uoi8ASTczoGJmI7t2w5se4QEPdONCyNSrsdyr6+NT0gew+WhjaCADEWnQZhBhTBCyRtQ7XsoX
6UEAbtQXnBvuk823qfF732LdDz0A68l60ETSHIJ2gHH87nhcLOiN2Uo4iptnj/ub62eo58d2/IJ8
hHb+Eo6rHCGE6cXtZilcd8tilxBxGuu+3Ls9fih/j2BSz+yQoGmwrCHCCGZGP8frMtN3hMAx0gF9
a6D0T1QonHid2F+FgJVtI99pxyvLqz1ImLaqXsXK6oUcOdaNhM+pYI506qw7NRvluqiuZyto5zjP
gQpMvisGOHyyPmwoa/WD+8O7/XWg7hRYQoTwJsnRgP/VJW/2o+eeZpBTulQlqz+0z9O8PFJsglwM
vSfMCr3hXLSzFsUxvZxRr0pjCJ7mekk4bKmQOeMKGsTHreLjl3+qgXqvm7ovF/PwStbnQ2vAmN1c
yI6qcK81NANGbmVB+g1hnY5RqE4ERdDuESZJhZuRHN0geipcP7iR2F514eUM7jOWouBe5ZRzR2gX
a0bqom7mMGQLEVcrqfXicun/3OUDQGz68eZNon96kzLwei/bqJGmHY9wMlTUR+3+vuxCC7yEx2Wf
RjiH+/t3uo2q94DJEQkF8gJ7GgN5bgc8m2kzqoMx2r3SpNI6x/HHoNUT7XOsKoPvOEzn4uOf2GQJ
dR+o8Ti7OJUwSkVNq8t/9xZHsy75ztwKDKu5wj7EnkUTev3fCGbK3yw8QHXO+dviuzyT6ZmvFRY2
p1EX8Yd5ZYyCxRxPAyDdkikoDKAlV/IbJ/DVvnGKsxl3chETx7Tl/MTx3M9a9xsiH3eaRChNoVix
pwSDnuGJ6lVlZb+OD+HUVm3qI8+fIm8iNHy/U2FYyGyA0khchhsfEdsBl+0jotcRELAfE8b0xv0w
ex4q926HKIlVPngN+LCBt/s0G99oycnRMppoIuXsswf2sMFyfcoeOBdGLVis0GWYlToUAlHvZufy
gcWjZntCcuYKVi+IheBXM/72ZiKc2e+Tq21uA+FI76mOjg181q7UR/Cs3kHN8sg/pSXsiisRVsjQ
XigzuRJCU/GCKJdIbZYT5EGXla52XxsP8ycltgYz8d7fXGvKSOLxp/CHuITfoKcX0KTVoO594kgC
mYzm20vpu73ieDyRA+x/32DtD8HCU8J55+0F5EpTAbt8XSnXymZkwKSdd/ld53JCrBbtPDLpjB6X
LFXkHLuTGS7k8Byt0c4t2r4ycG8XJL83+Kk+79LDiT2Z9aaG1dSxv1BBxertnPoqhpFx2qNRpUZ7
XReeWB27dwmCRBwWLxQLzzrccOlDsawa6NUSjlK+CzFCCdAo/L2xw4E+7KNm1cU4U1l0xTrbg9if
iMa6fnU8VkgGP+Q+h4Ebtd34ZdgpRmALwii2vdGiivzy+xc94tNAPAQYCjdMOFgVj726uTCYOJAV
KUkvi24GLmXtz7ZmWuIIPMdpInYLsC4tO+/r7h0cXtVI8eWLa8bSu+t9iw320Qhj8nefVDF8hp8M
CEOURRg09wbDZIDwxOoe9VpABrdoQHkpsY9Oct0MILl865Wznf98dCMH6k4bC/MV5b4F3+zqdl6f
XpT/+V6h2Je4a/0ylJjyZH9ifdteNtv2GANQyzX++Y5r2A67jLjnU29RJowPKbuIpr4oHrlbvHgj
YYgFqieMR8KLYW09j9tF7lqy6S8uToxZ9fpopUH92wmPh26OsYjaqlAX02I9GW5X/RRwYKzB0s0C
8miuWH6RCKuuQNAR93C2nnkPTjleCVex2nuRpdbXba6oxLNlveWYJdZMxASSLlj2ihCxCrsoAJ6O
b27xVeahgaQw/D7scO0DSzx9EmFkeZQGIMGX/k+QhbjGwK869T29mKITxsHPP1dQg5iaekCfkYC9
NuGKomk4DPRnASDAxCU+U6lgKZSZHYstIr3kFghA3IMglsU+rvqhXwRnhRR/v2onbctbwnWxgsZw
RI4rIVUBFBknMGUGkexDzqQhEdKRmNnivK9YxFsnt3Oy9WnzTeZHxXFsKUc7jVwQ00M6S7tAaKqd
rsFbUbnhshzF/omYnoGInjgqmfz/s8S5CNqwPoEWmrgwX7F9Lrgi9sYh8fStKjt1ED8WFk/Ea/Fs
lJDykfWLGyVsQjVThPkWKRX0wv2l6PATOUE3OoZvfNAkJnI88oTdrVWeVzBqSrM3/HKtmSevXDgC
WiutM0B6bnK/UB1ivenQrq7uhAIbARnDEtj+OOU32SBHxeL5Qs/3SQL6GTHGfFzZaoAlGXuFPmro
S04ebkJc7K5SMxGmAvkNJNX/iuyXZk0GQp4uPr4B+Kh6uNc93Qynlh8G6hZax5+iqE7DzUmsxtBF
QVK5V22G6oGubqtUnkjVhmk7tRilqmZThNzb6FV7n8wH59Y2TZaO7I6zxXNdkqf6RB7mGKLoFC9r
mpoqHHb8cUX4KOGXxdEaJaqBCo5h3qzXoECBrAqWXC/ln4s2gWpS0A04futZ0r8r6JAB3213NyH/
Cswv+CUj+jNtXjKV00N8b/rn989wsgAZdm15G6HjcsMd8AWo+HAJEOfofA6qkX48V7hmXfk1cqo8
GfPwMhCuG6Nc0ec5JsKhz0gtMxG0tlGS/y3BkLmgEsAmaF3/XQWa8e6sJ1+uJJ9Syq7Q17PvtkQk
IOg37cXkOSpHkSWyJrVcFznRfKBTukydLTG+l8gWB10VqbUj8cEbzlfhmmQjZj5uyTwc33SWup+5
NILijEVWtFhTYpKeqi5yh56/gRggdPoRnXMWoy78K3GnVpZZTN48ugicR7zsw7Purul6a9eM65dH
jiqtonK+iCGnWIDYLZLCKwq0/G/M6WSJew+1REd6+NLZn+pJZ1K1H0Bp67kFjPushGZShdGjkm5g
zuvxoVVO6rwYf2z6kPbdqXz2++eS4gs8It8frSY8L3HQdrx7P+RMOO6CzCvl5nH0e/eFV23tZMUR
wiphwb60+EcMM1Eu26KQK8TE44SZwtGOAxaAS4sv+XZ5jUAgz4qdmHxmdjo358MGaGSSWNuqNI7k
IOcctD7eEekTY0Xy4Cmkx+7mLJqP6Z7LH1ifLK4P4rBmKKOB+Qclgt7iOa3bOSxGwZLWMGgBF2wP
mlcv8xm2KLwpFPxlV6jyMfA+imiG0edBWrTKSp9PjbX+OTWQTzkOKUzh57jc3WhRqEyGXLGD9eSR
rUaYLWM40YtlbCBB1pi4vIl/xgnJ6Zt3r3C5NMmdNtNr9mJT6XU/aU+Iy4wA8Au+kuRtnjqZ3vYm
YdDSIjJ9XomAu30t5ot1N2yGlEa4X+2cVWJ5v9cRbet3jF6xSXXJXWkRd6Qq95mQ794cVr+ZVVHk
LrvbWc/B3MAKB2N4RYL5DOiq1Kp7DloxRMUMVgdmIu7+cxL3zSn/uM79xR72k1yO4gi6uhxC3xvV
PxYLRsbTXZerRdFDlNlOxsNPsoKZ+JDH90UQ+exyAMrLIxPljCUC23/F2wzZ5oQsvQw6uv0OYj9x
dnXYaKKMy6fu9VOu8dFxHINrFKqwsS3Ga0aBwkSm1GRO3yhlELux9UpyLvrzfPnp5Ef5Prnvwnvo
/l5fldOeUI0Nt4YVQzfbuTL2MrBkQxgW9IqkUHYkkRDUION8xtfks4t93cHWqR97zKYlvCXPG8Nu
RilpdH2++MVkyjA07sl6i2tBZAI7fXPIZLmQkqlpHKoR1TYgZDlKU9ygQrPUsy4wXLPpQiy4qGOh
8s4H2M1gs7R73Tj+86ciyTbUpnCi/VtrTCikDUlX6Btx0yin+ZbC5z8ZdwVI+aLuOtYL21eUTGp+
Ye19F38gjpnTTMKJg8JcvQr198tKZtq1IuEHDwrsbpyW31LJ0yUXJQ77fAgvZwCbE4+3ekb1Mg2Q
jw2IaamjCX+gMf/1t0Qj6EAD/JXDn0qXKLKDJ/+WKde7egyNshDSl4E/IkwZGXtmuQIla5q4Lomo
w36YGzffL1/m8u61cfg2Rjq3SkvRHenE/QjOcgFuXjFf51tPjHB9p4y5rx8gBxZWU9yxVtDGQCU3
fXDePIcKaB6aSrTc3X0AjxoAHcJghYaMVFNUwDDHoePcasPOjPOgDxUJiVB11kZuoJ7QN7Q3NHeA
YKWcGw7bH+Bnk7/HlUAm/lfsvehN9ZC8D7kdn9bo/rSz/NOKfBvuJ9kOWyJhB8R7Og4f2Fu3DCY6
34IqVaEvFqRF3+d+eLHGwWbyyde76Ken/axnaMM2LcgaK0qk0uFtYU7RYsUYUOpA0+OMlS6N4BFG
UsNVGdQXl6IpuB+AU37077CnaGvcWsSVWbCCGwpYEBIpcfLjMOg0Z6gFj628BFDFEfU/0hDN+b9M
91G7kLOGnRrOjHBzvYXFMxSfvLrueitBSvrM1NCAKn2dL4zrrdcyy7Txlr10llHDLDxHyetnr+nw
dq/p3px4uXl1PU838WoYY9L7CNLpKnlaq/rJ3UB4/Xt8hPhIN3A7ExELnygRDOMN61gUSwTPNPOn
geIlRHaCDX2xl1x6Hq2CYKtaSVU6W2XtOnyihrXeLN0edjIREA82wqpk6w5qbL70Mbf9zDfVsMjg
Zf3HqUiNZKO3z7nveSY8Kos1AFQwP8xJH54ZUevzg9AmlSi6kArmeEBcS4PYog2XkxEtmMPNB1cl
zJvchBEBl4yW8jx+J1Bd+I3hQsnHI3SkdaKCpjPLxLoTgFtRo+jGUJTcXKZCAIYFjefv6TtVD+Nd
eit/oHebJrZrGh+Yot7AX/YYV3dcj++p0kOp/QUs60j1sMELB/lvMP2eBp/clhF9y/XwxE4Jia6Z
Lv6bgu3xCoOorfSuj2l7Uc/26kJmOQt2TdDLmqFopAmso+rKue7AhuQG2OBld/4heQrjLlkWiTXe
XIOMbh/kRChB7Arv5OW/HVFEuYy3UL4kdr6Wc1G/VTJlHQViAsC3MYt5SYXKIcMslThdqhrKdubd
KDkepr/6k6hWI2Q4qA79YVY0WyPiSGvUOD2UoK7CbiVR8lptl89Ht2SAcTgiJpgK0eXDSQGYWkmv
tk3RN5YYMqzeG2OJvDo4ekOT4TiLXB9rfuJXEa7sms5uoPQ09pXYUR46OkJJZpoAU8l26cz8RMjR
E7GlKkzmK5kLdMSyS/w5wKOVAAR9nCXtcdfK256jRSlqm9m1PXdEh5HLIuektnCkyXrHBlqCExsI
yc1GX+jGNfwbkBf/dwKgZPoLkZzBXcxBNIEMOPKB8lGJ1wsBm1IJpktj9baCp1+cCTE8VDMlsBaP
E/NUz5eXFr9U5v14Cks1dypBKwgXtLIH5gZ0srctu/3HS/sY3K5QidKXDaoM82UylA66REHoCrkJ
keXSkEsdiDdtK3t7O1wn5bHEzDWJDqUK9JACYUU72RrzTPR2YUNfH+a2c3qyCKJDi6IHLtGWmpLq
JsDYpF/b+sn+25dkQSlWGNfrjcIUvI6MGA7xbkGM9xGYMaa5hC4dV6U9MMjPNmposseL6B8rmwsu
dipHiDulb/3pLpOGRJYzUxr9l6Vd6H+UbsWvRjd/+cFxA/4HfDgTDxWsaCjOGpotrv54s2/8RiJf
zJDA+yE9ndvPK/l7TTWSyFc82L8LLPCmpOlNhSO/jzdXFmHN0AX/RujpFYYYHDXHTh/XMJBAxpZC
Ue3ShBUhjW3x9XKk4ORarm65uHX13zH1wYKwcvEl1J3fZdl7wCVKFXixnTr5XOF4w9IniicGH//o
eImL/6rOmNFeJL5KyQNWNdeewT9mTHRg/K6xpTJJ+5yZ3Hr7A5N+otVzd1czXEInkHfuGLzsyqWD
tZ2zqydigYNRR5AtURjHJzFmtlGDQD2T3qd87VzL3KVL9pUyjMuuSlm433HXNqE8t/sQHWP5P1a2
VADK5uRVSAbcdv03BrC97sl3q00gdbklYTeTsx1AdXq2o6aF28m6VeeFQ5p5hG41GXi5/IsZtIQn
SmUO8TDQnS2j4fNR2PGfTC9UrUvOzDkPALMMibjV4BC8Cg1cP39j2BYfWwAoxt1pQiDH91/28pcX
krGaGa2uzgI+c9+7gCEWxwmQ9miN/9BJ/zj56C01muI+bTG8odpqaUr7QKcYvkKXHwOtceJV7KZK
99jSCgRumtzWyP/LGa8idcwEV9kfZICLEWhCQjw7zuEt3h89Sf7rzpiPwpuQdZz4dmR2VT4M0/YZ
fsbukNN6YUHkQGenAKRepEfNLl5rSY2/2uEbmirprQoSnc4omxlN9hzcKsOKfPc8AFKj5Cifze7Z
xKmHSaqdlrPgU6mvms9A0gtnx4OyLl0I+4QtlHqoNCiJ3Xp68wGRlyKwxSMnGG7IHXxSSDH2ZyPV
qmzxu0G//1o/+5gWc2yv49DLlPpdgWKp+bjLX4VT3jhfRMMciEprWK86H6zG9hzIjT9jb2PlCYP/
gN7pX9qaKQvJD577dJnQrmbMNilyoIpaB0URad9jQ+tXw6MVX3jdAzlgBjwi2KF7VKGa7uwWBg9N
1WrI75YHezaLKwWVKt8Mh8i5G3QQoaZharYIqEx4ZdhdxouJYKRhAByD7sW7Z3zinuUGatv3oyri
B6i77a73kJ9YWFBaL+J22VZwWwljmADIlsn5LTQiUVEaJVXUAVrys6tUOy1jJSE+XLLtDMwzZjEe
zLGLE5UJ3VdFeal29uhVoS8UbrwPz5DoKutgudl9S/va6I4Tu1B8HeSKKP3byRws+P8A0dO8VVYO
ZnqGoiZMIJ+c2/OGZFzRPvPUGf4CP/3qQs7KvZErMiT9OGe36C3kkjmO1pZIDtOi506ozu7/QaK5
CwzZD8a+BXwJwsXUTbyzrMGUfAH4VkeKTuHvtXdhGg7dzVMsY5TN7EzSl0ZLnu3ST/E5MhOfB4Tg
bQvegrztV3t74+VpwF57XgkHmURiA0VqQ3pn1y9zrDj70gmEXoA88ggorYY+quimHkyj8T24n+Kt
HaMeSHMB70xjMkxDrKl8Tyku3NVwAjAoFiOjap+zVTT6My/xijD4ie7Rk3UsNEfN0JHAS5dZTfne
zdQppfal/nfrVoPTOVim/0B1DwQIi17Ofyrnl+XMA70oDZ+caFEFeGSdZY7r3vXInKGo7SRb3HUZ
ecXG74Vc5M1nZLliHX79DfkD8aEBFnAbdDqv5ADARFmDQPtYxh6w8ey+/NbTt99Pg7HoAlNlsX9B
XpPeFUuUe4Yy6laZisw0mBAJ97VRqnqq7NaeQ8N0VqrMtbzCKfXIf83ct8fjNOWnLp66mi4a5O+R
K6U+mU7PcDHMaNMEusaWW/3D0ahO0/36yo/MTAe7ZGxuNF+liHzc2JSQ4IqfaRFiIKmuWEFVV64U
o8yeZpzxLJVlt6HIdqVUx/hnIxj+lclHaTNKb9RA+VrJOVJ9zFck2Hp/FshNhSzJ1tEplVrPSaAH
z7zbWl5sdk8okcANKle84cWgdqoj6pSAh95lW0/hBKho9i7v7vQ0KbW15iOG6NdQabS+dsS/+0p/
n9NQb090wdmu8mC4uH6rMM3cYPewpgK2qk20/yb2HYbO6Wr3Vtj0sTyFoQ7xBlSYiuZntv+lkBTb
m4YLQBJ0K+Zt18i2BW4AXcxtLrxuORM8C3gpEqHuLqZdBivJMXdll8iP3Zj0QoO6j3vnzvzrxB4G
hmSZV9jA2WO8Qaks9shPdCDG/+dK8SRjL7H841jCVrApg/jBFxRqTTeIM2kn/T9jkug5tX8jb3vi
an6yBGIpf5XQxmuOgFHfjYhWEKOsEmNjnR9JjBAuY65ILlAN59oae4bfWPIlBXvZoPaxFoiHP7G4
8Cok0l95QioLFX58NhG1ac+4dcEFxYtscwe3io3HP8+stx3nASF2fRIhoTeJ4i65KxXNtQLZ+T09
20Y5Qs1DfV8ia1z7cCBE5ESkZpA/p1MhkNZhRTbZPf6w3CnwNOxvnG7A8P4fOA6gui/tHf1lzCAD
AB2XX6Xhmt61BAbRm8JdHfjM9Mkm8cRt/QquUOImk0uS8WcYWEbkUB2h3QNjRXlbYvm8G3i0sFvE
XVfGMSRviY0y/yvNAu4UehXikf/tAY4kydMqb7tbGi1xdEDckMJL8MvzfksreeuuxrMTnykojema
cGirFw9W5AAEcMiIYG3JYxeLwSv/ipvl9XfK5F0Vf8RNUXtKIB68uzPrk/rCwQ5UlrhiHZYkQDIt
wqJyJsT1o2/cdjnV2dNEQ0B8Mp/H2Ci6cXh3w1U8asPU2Vn9emkHMInZ8w2m+PVL5LMTIMtVMWvp
YqVuwOqyHfGF3WqPCkcWYu1dVQjpLDQX+ywoBH7Ka+LYXQyMncaumcCqrFkuxOIclsP9Ao2TvcyA
jI2faukd7sO7amEQEgIb1TVemMIFzb4uSZcHDphHvgDbABrEwWhmvpI46T1TLBU6sflIWszfjw3E
gBq7kz4BZh4xlGJtKq1RorIm8I8lU6en9RZLykIAjZ2+QEX7ZF7jfS/bF1m212CD5ftOryhysP6Y
sw5T0ydfrozFwDck3XBLtEaxAvqNRL5NYoVtvFBLTCIdnBka8B5Vy/XWSj3SssNmFtvrAEj1hiyq
WBLftXtcsxmGbfLWlLNMBs087YddED3hKVhMtKEDhYm173prwP6wtvu7amCPVxbJYt/bD4DPVB7A
fYH5fJ5sH6oYC0Lyc8QJvM/AUexQipeg65686Q+mlxtLSWrbKrvz3V/wsEQJ1y/2YR+x8E2oN+NN
dI9ykncTNohQs7xC8+TqZbAmHJ9bwDAF5YOX414sSG0kHZWJgqCKJQc6E+cDdUuSQd/aBkzGMAoO
RosvCExNNayYMfvxFaloahf5v4kIdBrLvppRftCMfbaOMVa+lPi/8q+5NZsxPQZg97RDjNGHFLyM
acEwaIRbqfWBBXrK3upp6tV3YeDbuDlOFXp8EcsiI4XeLCevNcWZd5XzMDiR71z6AcgtIe3YqzzF
EKietagvyI/5RopfaMwZRg5c4swfkfljYhMVgRaAkVJxIAMo+xe88o89S3mNTzmxik4bW3rRgKtx
c8qQ48kNuZIXH7lE5lvgauBv+k/IEsGYO+OWZxwAXnVZkHk/JB0/Y5jbNHjqEwfJjpalF5s8NIcZ
nVyaF9NHKkMomXtOnVjVOkLWYqFkJtAwV3ippfGBiFqdUR/k9ci4zUnlT0eD0GWXfowCmrWolHDy
0cj+uYKgW09l30Wge2SVBiw8UVuvSPw9R23Zs8YzvTdCQ9aSCTk0wd6XO+z4TCOf/Eb3jLsYWcBB
yjexlMgg4ArPSKwZHTw1UyOL5RHhOGvtRBUVkKiQRn5TEqRvWroXdlyayPAW9vRvydLrG5yoOytC
8Od90h5hkfOWUaLgUJnth7R8C1bHrnzPp4Uw/56Exb5ES2cj2uTAoDbd51OMtDAn1r7niLomzfk1
nsnwBif5iGwzWxKcxAFOCaCIJOpMXJpr3kHxlKAF9Axc94bAncCMqKd3Pj9vG4gCcCsBTMYVQpdt
hah65WhNbI/8z84rUlFheVXtjArxoMsLUwtTWimEQF5yTv1zkP+4N5yc5gECl7dQlGn6ArQIqqE+
8lK5/mEYiRV4T6sKBBAFMVuJwPvo3mn/fdIdMaSmDWTS0Xf/uLOpYic4EaE3T2IrXeTBvW3zqa2O
XojaQuE0lhPQGV6vr6GXWiso+5UhKDzlRulhjVmGpQLMMvYnJQJBZse4yDQGmPH73COZiOQWLe6g
pnT/8RxyUtHVvJGQUhUzoQIyU2GBuqZpCVfCYvfaGGi5WMmlWpmVE5UYF5HMa6Mg6NJbx/TI39Pg
nZt4drmOl/QOQKl976Tkax5yeO9GJ9s6BZKJqqYnPFfXotH3ZZx24+yWQLJNvW7B4hPGfHJPltdT
U+qNh/MI98+QlrPTV/AMHp3rlZpnZ/lFC70lesxMv+ZRL4Y7Iodpg9v7vLKX5LyO1I7yrate7/A9
PAs0Pt0MyAWrQuzaPXGBf9lRu1wzCRIo9M5ORP1irMuebzmfAWQpJ+cF/5Bi/o3eA3hJK3eNGzKe
NopJYFtzdDnpRUI3s6rVYDthtZbAu9QN6OD6KQDaSqY4DZhiKE8s7Q43Vj9mwMuOVVodgsfQe7Rg
71+Jo5xtTAcrPssRLQW6AC7XUrSdH0EOJ6YdUkdYOkG6yFsH9xVBi+RS88q1nGRaCAOYyF3iP3YP
kZRBXK2TvF54jnU5+eTmohRE+PkySrUSQAxflzescX1opD3kHS5mAzBjDiKrzQOpy0qT0ISlTfa4
L9pP1BwH7FivO/CfM9JrO85+o9YEo9YjdtG9g4De7yKp9WoxZOM7FCbT2fH2Jazk89hQ0sqCPGhU
5VkGBdXpVF8Zij+Bnp43HEnONNDVAIuXMFHLOjVIM0LAseRamYoiWk3ykOAbKN/x+d6Eb2ZAOKgC
zmhVEa88vtIAPSji+bblNjyVRKtXPx59paRao+2hfOjoL4liMYSQVtYlnTDsjmAp0pq4rWcZ6yx3
kw2u21eXZ6a2miLsrcybDB4QC4N9j+hpN7xITKX2kkFMQDIByCFAg+sABSe8es0NN3Ohm7Fav8NU
cBLjIFUi9TzukCpsayA7vk3I7DYEuiY8POHsMyLkGCc14hp0qglXsdGP5SujNKSB9N2smrfr9QPs
Jp9QggKJ7Xitu6NCaMh5rqAYnfX7xKxxCrFOsTPT2WMkqhr/ZO4y6heOkQeSy5kQPruDjJRgxJJS
3OgbGi4fMpwSr9uPfWX9qcI54pj2xRA4OcRswyHXdySdlff6ESE13LQBHf+sbaTJgt0NRQql0Wfi
ABJhBoghw3X8tG2LH7HSkVkI6s9ABaG875ZjsGO2YqriRMBlZ99puPauWsRKLGKkkbaTH3S7QEhX
+oFt0lOl5k6KL9WoUhPdGsdxN+WXI7tuYaoI99sNi3PFDU4LGIzC0Xw1qwzzuULB/9vw2PRsNGvK
fBWoFmQXG/ue4oA8SWL9bWXnN6dm/JiYQMDiv37la9O4ovEX0eaLeZGgplhHb4bSZZUKDna3SGwc
4HvkmSEZA3H2IB0E0wuw/By39qAAzFaaNwr6mGi3KikUgU4nYP2UewIMhw10skuBMT9f4d/el1Ub
6ykUofmX+ikfg3MwI04gjWZRAQlSn6qeJMCyIGyyEVGBMFRNOah03QsAQ97X5EKlJwxVLgtJQ3yO
xw83bmig11xyh0aUMpZ2IKqyV6+NA9rJmUG1pXin1OtcF3xxpFPYH5klyerruJTfFMlK1Md27cvq
1p3dMXgchx3eNU2iZui0B1DDlYRAWN7MwB4aMfNfiU7SHhI7tUssKLGm+m7PqfaZCXj2E0iM+s7K
/VNBYX4IaZM6EO8TYOt1OYBbkkgmSPIy7IqE0LEL/GhCtJS5Zyk/npvFxGAAGOgO/rHD7OWzz4y1
KYGeS5+iCzmXP7moY8i3zHgBmpPKNOGczLIf+/NA1abD4slPeYForaBcBLgm7CGCJPfnzFxhlBdf
HoSOd2apd8+b71ZGL8dWjoU0he86Adur3J4nDg6NeXUp0XYuIMBHN3Krl8kdSHkzXlB7DZ71ceLG
ahXslCNpU7fhFshUInuBbaJbByswwbqxBLaWAo1EafPD6EHA5cWhYKeDzPgpEhXfOi1GXeFYZHNT
1wDWLT+OwEU4zt+bTzB0UJaJ8dsdaOXfSlbznfIPzKTkjI7lfe86QnIE/NaFVEfBymtyIfFHqSYA
Z1bpgMxCRpI5PWgdO0pW/H0R4EHdCwpCPV6ENLOuDqJqEjejBhnOWnFB2D33BN5qF28gukdvq7Dt
8ZfqeXkG7wT7vAbfOHzrXXl0Kk6qiSVJk/tGz42hj7CHOZ2yuo7F4eEdxpdP+2vXdsNDawjBXMLX
Oc/qPXRhOvdxcMwRoLq5id46N+/IaHVgjZ55gLHBH3mZ0mSKgjk0lCVvJ/DrT+CWIPdy8GJR+nCG
3Pj0fHcOtvDvrEz6TzI4V+lODwWoovsbTENrYwSPNqdCXIcLwUM22Xii6EDw5HxQlujUPN05ZFj7
RkR8fdkRMlDirCIalqmNchggCSQPVthPsR0uoAsba9WsXNcd01IUZuZJqUnG/HZf3K9bDxQASnbQ
u/dba/it8f0fwbrnFC+HJf44nO6DqtVJ1eFQjARzG8JpMCDF7DcvcuZ8TM0Dd90MEv6fG3UuFd/9
bMPQi65AXAKZEIR7pROEsTe+qmS4HPAD3RZXbwEEKnJVjWNsVmg5Zi3hGjpa8yJ3dbTUAn01T452
4JdJgzfBLiYe+6XfAmkbzFVcUlMrgnZrHpONvopUi0G/hj+5W4Pp4c6UToZsgBJ8/qE/hH6jJceW
H8teYUSRUUlwu48nYPscNJWRR9608D5T2Ibg7l3VMFrkttl2zGcoAGk13mDHJf3NYC5EV+fTl5mW
thi569q2I/EIOg/KJn09B5pmBclHQI3pMgVvodsKDaA2VFEnTWro6A02XPZ7rrode1mqKVGi5rlU
axCkRyYuOjBh53SmbkiJDKoUMBWcBwH9xG+VzWAgspcJFKuOpjMdJ706vsEOna+0n3Z8kVO4FDWc
pwzZ/Kmu4T1dIarOD4LxYZDt3CJbWh9/8FymynWy9RjgFxe8024NZvICU4KL1vy5snUTpFQ13CL4
/lkn9f80ialf8KZch60lwiGk8DUHbUKWcwZ3pxZhxrmqS3qzRWgcJ2tZ4M0d7KVc3QZVlV816BKf
lMGHdeKkjaXTsweko5fs9UKJXb6a36th9HmrK4lJLupi+pcFiJpkNZadNQ2kDhbxaYNuanDiLhlQ
OamVRmiGAXWwH+gSgm2RGpCnDY4N+9UCpCWIiT2CPPZVGCkcl3oj2jvrIrGVlQMAPmAxx8otd8DG
7kNQCX/F2DrIrKI2+0olYqXmwxeD1gHxvpkKyGjkgzJfF77bkV99LNKjxYNRJTFJL5js/hTExMQW
p4PnEcUYt3V5WbZJ6uayqr/tqjOccwnwfHSV4iA+VtcBXZ2jGwgeiZg19jJG9O+0ndEGgxYgP/Zd
eLV4gB8hfbo7v7PlMmiA5kuhzO3D/S+hUobQJFyUptXdsvjaHd8EUjV4UvoDARrVkURZgJapnbUw
M4VqSacn8aF0gUBXM86wrLUIhuWjSJRBILaxea6Taxlhw3TNhQTFaHQIUayiRMFbEn87Cq03LqGM
46OqXF0wcnd7F0byP5qRYiFDt6Djz6cZkfOoc2QlLRN2m/Ogm1QKvDc6ZX299OpbcAzQtR3pPydu
NjYaMWksoecFiTIoHviX14HbhA+umLI1mSASEOsbuEHSzfIyv2I1on/MvdoLsFlkcDgrWrdheLTJ
PXVKnPw9OdYSN7XE9ldMYeAPYbedxrbraMcf56AjQBc5iUDeT+6iQ6AmjHFpsuWnzidQKmbFEUEI
IW23PP6pm+fdu54AL4vjfTbArNhzbLgYa7wyPI0ZSD5HLsKgsBS+YyDSGP7xlUhURCijH/0FjsXD
c1qxwCDQufQ+IkAGfZqrbJqhUuTC0ji/x0f3ViAw7y7rFzphTKDS9ybboV8zO6kecr1xNw1TErUr
fdw+J3n3kFxVugwbn6ebXAkTz53iFAwXeq3l55rrRNiPn48BhVZxLv/L6EXoy8RmO46Me6CrJrnc
CuPPwFsI1HZDf+tvXjh0PAt8TrBXSbYBzTqDuNkCDPRxo09Qlzz9VXIi4lPZWxYxlcd/xvXBl4iZ
KYWfnPqx6zHiNGAVG82cSPPMbtpDdkq0ue4mx/HEddNY6KhtUXA6ZbizWR4bJvPyvIgzuiNSe9Q2
uEaZQNBsM7vbOfQNLPT7OxdiSS/3pjaWgg37TfgCgDY7zadP9W8jdnQeZs7TiIRrbjNBykhv9Ifg
HXyOltXN3kU8ShlEauae67saH6Ig9eI0q5vO8DwxloPyq4tDzU7NZHNNqPAJCeEN7e/KU0NeC9zP
sKpwL2oLtCpkIPNqXNzOTK12KidUugbmr9XIJ4pYLOSaKvBGkKxQPSn9FGqVihMPN/SGWHOxcP/+
6wkcvspA067+709EU+hZ+rM+uJBcHroJ8CMQfY9mJjcOsUVDEX+c9g85CS5u3dcE9u4m/oQLGSoy
QqMh6uaS0xxh1bg27+K+32XeU0go5uHvLMl1r56l/pGYf1S2xDSkPsMngYS2czmGLLe1qTjwOUbJ
pV583uUhAubg7khY5PAFsq022mhwtFQXRm3pXKv/LPB3pKiHRD2ZPI+Qz+jA6tM+8pA2MoAFYtE/
2m4ppcPLXp8Bgila3zDCemaXtzMV7EZ2NRcuqB/DWNwrD8FDM6iubQK7KK16gQKaaxXtdmpN+xzz
yw924tIvZro0GKeVfQZBM6dWNEGRXMyLU/91+O36JeW+1dpoRKUMLm1OA+XPCgq3tAvTDpfOpQrf
VblW+gDZDOxHoO/Nwe6X4q0hDHhKFkNRYG/d/sEkXqHcKZtz8KFQ5pvDQSK88lb1IwpDbDZIfobX
MXbyFsAF2s8W+dl5GbrU7VAFN08P9+H6zQE3cP08bd1DN0BkmMOaUADc58UkSCBuFkjYQhLPAT02
Mb4+7Zu59kVScxeVZgAXE/z5EINx1x1/sfqYx/PQ+0TISJNgtGeRyvHgT0w2PT9s6MFJQ+H2C+yy
CcqENs+JeXDGkiLMzSJR0pfgHGbHaZV1/6Gz0hGBXIiTA9KF2LJ1HNXadajlHSxmFYd6c2lClNw5
Tnh58EYA3nKg9VcCdfhhYev/t8s/P+r3D9mlVGc5faO8gqD6eGnZyJUqUYIGZaiTFIHpk8kuYHSj
c/wvODnWmWY44KX8+HV8bd67pNknp8un3KAUZvtWjz86TvpxD4TWGbaWTtRQ53QBUTdvpcdlGToM
G89wUqKg10ABHYoT3U5ayu1yIXCpNkjypcwbA5HtLJp9FHa5W5RvxeWZmPGv9dMLMzqMExBfbOe1
HTdwI+wummVxgDFBOS7T8wIaXRSQPZKcdUmHVYMCO1Exc0bOkUMXKjiAbMYLJiXZq8zSC0Mn/DG1
bz2bOVLuG61k8YZAWSi54P70NYAS5cVVklE0zkAaT4i6nFoiZr/yIcLmHYFreMucCJCINcMQ2oxb
UNfx6oNIIH6Y/3Qg+Cv7w42pR12EO/+W8z1XpcM920AXPuyPcE8OLQhZ7pUZCFQKA3a3mcJTAJCx
uCnKUKPt4dW68eP30bVtyDo5KAWpNFuS2QwHJT7b1QmvUd2CymgBGg8bErAvgb5GzYf1VCi+V+ge
CWs93bpcCnU+PMoyYLOCKDNnY1LfzQ2KpJrWmQXdlb5qOhjJUyxXVHoW0DHTML8jLLiOGr8NMLVx
gbpBdwT+9BIl1AJRRBxnXNUvKtiv0DkjdObK55dUEj/w7PSt8Yrqy5Mcsr449ZDXSG6F5xNkjwwc
o0o9hFVc68YK3eCZryrz4HWOZp4ZdVj5lKZepJVlXqLnT8YCpfX0IOEW9ZonSgEf2+Vj1e8dRENX
6N3Kfua0xITmalBy0kVb1O4nWtIgWoi3MpspUpboBh4odOLsg+YaFwrhrszKicKAuSeZCHkLLn0X
Adw+PbfG+TVtQdMMqIPO1626YadhQUoslGBZDxjvQ8BdAGSal7U9Rff+ZhDLwoVk9Kaj2yvwvhkH
GOLitm6wmtuu74JtS104RPVu6jYuYGn2v7WmHrsTPuv304Wty4PKwrnVO/HDMHPOqucj98VSceSQ
+FRP5V5fqWDE/gxBcHXTFL0iOO7TfkNMCepyWwrPQiTFcS4HEG5UywxAVeMkcVRYGijdoILrnHvV
Ujx6GEsn9AlSQDrBamr8BlrKFstUml6WOgyJBaTYzqEzHRnX+QQTqsjtAKGwwBNmzwdNitvpo+ai
cs6HHgzXxKO7TpbVhjQBXMam1WlU9KvDS/VHZa3wIyVcbB0dl/9Cp6kM8oGln22z5ySQhIJa5RMY
AQ0b3LftL9AIySdV4PdKIEid5+FJqqpaGRYm782wy6cV7WEpQCoQ2+C9mnhlAPlPgStEXEp6GT0T
rPCaJoJYssYpaCN9+sg2Hyje8Sd2vvCpQlTyMJJKoGPiPOsOneZd8JqpVhizmNZwzEnmTwHsIG5Q
c7GXVGNhUbGRgYgf5QkTFUEw0hamtSYLNqwTjEEaYTewhSIZwMSLTVmHUQQ7rmBPnYaPwghDoCAm
x9TeUCSJ/fyPCVfLf8zkXdHg5ItMHmaOfPnFh4dnJyc2wgENnr49oY9tdt46xdXGSSvzgKdXh4XA
mfIOBkRYKOKaANhOQ826rxkdJNK35vpUT1KkR3gRsYJGcQmjaA9wRYlwutR+TmjxgS8TxsrK2KAL
IptVRKKg+IRwqVF5gEkIZDr7cepYCxgJgG/1QIkLxYkarF7w/rd8rP1Npy4ewQ9imUUwZmgvWwty
BT+vdGZp9iT/guzTERaT8aSP7OEkbpGjug+YUdNaYXspvXi39vhHZH3kMJjHK0KPV6Lj/E3V6kq2
eZKiGWSdt2/CY3rj3KRDdnxCWXXr8wIVEMZUKsdNTdJaQK7SCaT2PpoUDXuRs2mog42o1vZL1VJL
72J8VAexL57hCu8TeI6LX5hKJCNOB1SedUO+wjj81hdqvV3ZItBhKftqhnLdDrqKUvWJPP+5IslK
7Kxqpu7YtPBuHMM/pHQW221PPeqhV1VzlIHe1WuEFX2xWeIhjNx1iPXmoxYwMCdY8ovLtnFowNg1
6mNfia4rKPZUzl14G2IUhkB3dTmfAbUaL8+X9ifUZItrIgG0zTWEeAYPyP/TVosmpwxo9yJiAAww
UMmNwZvKYKEmV4gzSa+DGOpePELEFfUUNzNrlU2CQbdDBjg0Wm0+vGs9adfzDwKG1jAsLRZQB8iY
InlvH2aqxedC5tvXZgMFHo/BCAwszZTHPENBi25bFHRgS+Va1j9cWKkuVKAEEg7rCg61SuY0THS6
VN88iDMN0wZUXetGv7LX9On/FirjB8ki8i/flc/A2IYPD0BkOGGwibQCvy8I4/l0MQiwQvOLSkre
POd5AwWwX0Y2gH58VohJdpjTWCVnYBhnA/ramSshUzh0WEfNcBFeJLblcEsy371mrtIz3i4r7cvG
Q/3lZ+1ShCBKjTZbuHFv53i0tbkBgLpAYHtfXzAFs2ixjh18ydT8f3gtsGJuuNZru9/ssl1PWASF
pqXSKFNi8o5KhY6bGRp2tEskt8+I9IBHLy48Eq4otyTj5oXBvrw+9PvR4e01fMQ5mSyqHjz5rPWH
LKJjrKBgXIfBWt8KOHihceQDwPGLoHlY1zE0Jfiq9YjSZAN0HEEgLTXh/QONPmh7r4vIuonMs/m8
h/VSaC4rZXLCFuWolYRZzu2fTc3aNUTnXTP7WbT9aGP1g9qSt7/mkc9SX7UhuIXs63Q0AKcXz9iK
nH7XR6hOZSiQM6wAqzdFAznODKAuSZrVg2PjHonZQRWYeha8axIxfb9Qqr7wnkAQ0tfQI9wvisBt
9cmSFnlcj5Oeog6tKP4Q4Jft3E4jo3E4YsWWz4iSKPhtuRADRhbLhtAw1bamg3z8XbZ0edt4v4+R
UNhxzdh0M2l8qOFInyw31etFrU11ZSq3VPNhrLydoyhx0E/zVJ8RM4UjTw34czvRiSQvooqeg3SK
YE1knSxR9icLOdhSBpDgXeL0Wm3oK8iVIKabeixg4FTTfhDv1jinmXV7tAWSnnwXu61bsBzGZ9CV
2vDb8rf+ebJei2wU1lF7CMI4gpUB+CVbcfhh/EKFWfPlQ8ReQQ9wRmFGtuMsv8/audXNC0kx/Ev4
PClfcus0qN5MRpLcoDr749yzM7odLB2p5vLknjxuwZHRQze71bLl50jERy9p8o36c62EeO2+8SJ5
YtXPVxGCl0bba+cL/m97WY1BNOZOgrWNLG1PBPNDVz2fbZTYXqmVtsxZgPx3lWQmC1wgjCFt1MgV
p3wqWgv+KqvhLe3LvoISZw5gClahGqzkWOhDCj1zS2eFpV7rwtUjANphoG9BiVPFp4oGiZkEHC3E
28Kl6nOlJbf4v3eFoN7ATsMP9XT4rf2YGIKvXT5wbo2YHDXIFdbrtdGZkdQ2/y/lFwniHdyfFNv1
2ALWVg2/u8VKU6mEiccM4ChNzyQJvKX+Im0KnKRFHS93j8H8lns93qcXPixwveBdeCHkiNQbdLkF
Zp1O4nofMiwbT/S5wH0e3XP/FhzPg9CKac2pdXv5Pu7cC3ltOE1VtKPK7nFR9iyE22w4YCDo5PeR
wPr/c7V44/SZJbG5esUOnycALyia38ibZFX8umJ1xESmlYNQsi1oulaZJaX6X/ST/RyWEsCbL+yV
5lHDT8BnZAadZpuWN8dlpf6DYwW5R/g2VKgPVjKMqnnIjkq/7zWT/A5Rop7NinH8JhVA0wOqA8BA
YX5/f8Wtux1STJftQs8xYoRHS55ogakuRgLZmLP0gbrF0hXocPd6natZjvy7guNlaBCtXfnMJlST
5iBhtX9OF+08iQjKXIwktE+uEbX8hlX6seRtn59Vmo4KeDwJ7dQWdCMZbOW67Q0t9qhlOj3kQO8r
50JKGltGNbNV2zcAznfy2xiobV8JxV0MM1ZoPf9OAD8Btnag99RVQLkmTf5uYYx81ZNFg3y0PPO7
DPZ9/yUsWj+/JRp/W9rlEc43OJomYkASX88JGzECzD+YaixaIjrw+ZqUJ0zOKvSdxh32fGTonqid
FOHoytYjuGEH6g69De8F3tQEXfvzbjXY5YthD5+6Sg2jjaUQXICN2iumdQphJl1k81bb2WJ+db20
dA9Z9zgxBLRPjiSbkdw04VHtLB7SxP54FSggioZJr0JEuvUqA0SrZlMZpq6aqsL64CwmizH/bWdl
9U3xrFIbZ3Odnzj8Ves/180t71hqU/YNFAqS8qIDr2zmuFWUWxQs48S6klfHpue7UPQ/uROH9EVu
xFevC3ANy6/5GWIuvXwgnyoirBcqdKB9kh8Z6d3SjSxV8NrIWSWlLWMRboLXRfzXHrcyunC8OusD
rRqhGLCoqDrSraf/tCTveQXHrf0QZnjrKeNb4DCfKNww5CLgbKbsONLtuHk/EU4gh4COMIll5o4e
ycakaNgKLwFA6LXYhqDaxDZKR0gOcYOd1vesUOg8SbjNvPTCpC0JtVMJcOzxVprwEPaKXPj5For2
7D1V2D9bc1AtwzOhIlrPc+8CiXGKfOE1PT/ukf3W9/Wh0cJdz2r5B0IgNIfBjLRn/4d833N3BXEC
SnA8SIpiB++IWgwFEGX/P8Lj7aQuQDPd/YcQidNgRgoXHAkw3iyT8V7PeSSiD00Dl0ypWoQDynmK
8WLmyLXh7OUcyDOo1m8uQ+I4MhypVtjTFZKnw0hLaOFiJO2lAVSUzr/1sRvP+xQtHrVh4JLXPFtb
e/5n40zXh9ej445szxzyjIYqfuGtu+SxUR3DiwGzHJZFjKVTKaFoJ0wG8MLfpV31r9FGgG6I2LA1
tLyDISXfnwuL2WVB0nnFbQKnUeWBnjqvG9S1WpHJmrJKZ58p9dCPjb/B2PNNGfTH2t/67wekVqkq
OrZkShIpO4jT+tcM+nAm6POkBVEDX219k0nbneCuGV0TysABkyR2GgXbExswjg7wfA9nFAuG1eAp
OlSM+HFmm+006sERWZ/JkGsbUnl9PGR1s9WDWaWVbxFjJ9XZwJ8SRzdSjxI6mqg0CXx1NX4JRem6
u7FEltQs9fohFB+TQk+GS4L/60gCttxnBLMvGjQ8AYVNsZ67YAaUtTFb0v6DH/c/WGQ50M8DVU2X
4Y8pCHIwNpxoq1uBgI0eKEAsbnBXC1DcqGMGuAzq2GQ1gjrp2hs+g9zSzwEQEDoJd5Jk+OxKniDp
35YGflugRBD+MZnHXL8RdyHUz9gRVns/KMYFm1RH18MIFITmYVgUgt3FLqRk+jFFT8nuXEH2l+Na
FyTy+/OBNYz5LT1Mtt9SQfCRzF5m9k8CpbBJgpnAIS8xF+C4GvXU4FRNq+gkHjtHi5ucD+JI++yx
VQtI1cVaT8cM9YcorUZR4vCygdeiKO31lMaumdiBocVXpTMnno3VNXYfxpifjiRNe6KAjXgaDSbv
5+ABPdn9E7P+i9sVw4ZRZB379PU2Texh5kK+jRFOIzOU80Wp6IJNVZOhJ7aqobi117DnhXvxJVtv
2GQ/ZBwZYG2S3eFyxLfowQyiwclvBRHFrWvTWvJ/gtKAKm1ZVrBE3QrynhVM//CLLgZ267wisDtJ
b2eDSkQEOmmv27tk1ftOITa5C2C5NnLw3MB9D6QH8E8GMF69UkqkHD08hANOZmQ5Bs5fDSXcYn+1
EGyKFJzDFNbSsTaTiQSeXSiNLo7KDwH9KXsp0QrRiCLnS7h6D/eKWZQniYnhnKGaJeMK7538hKQe
XcOeEuzJZ6zPHmkl7qre3BWlAoLYnRNmPqs3Elb+sLzgByRs/HfXH5KtRoWN5uP9P1B6jXHJ5HSe
sh/6FGutPqqh0Y7VhekZlRfBd7I0jbmCyrTIZlJ4kWJInlpCBEV+Oj546IDa+yXiskKDf7KGL/JH
Yvd+vEOCM1bQfQ6PLNf8+BmCQXHseGboOlSPqFchUjKU7bZgO6LmSV9vvDRWDNxSGG4sY1H25Daw
dnOsWi3YjiBKVUkBi22bCEHrMbOKEQ5Owran6Jz+g6XvSAMu6mN2x3+9zrXNpXOvkgqAUYZbOfvB
PWIi+jeUmScIyM5uYkG7b9aeA9hLSNTj1CanVqE6+PmJeWBLAg9AFGsd7OI6fEFxmUBGq2POUpDg
zeZUpF9Ce9IOrWlVgQU/Mwkxw91YgZIKkW6Pd1/gqWc6vQlQGV8fPo0kFnC8Bqq0+ZF2Ij5e0vtS
itxuQamVxGsJISRZ3w265WTQdVLwAw9tvFqCTvTyRo0dbB5kKFlgUblJYyXC2erVYWht79v+vCTS
y1z2+tX+WJGFZ9yqJAeOPFYINfd3gXi9sTKHwiykmjygPJXHbir7s1vJhEJGAeOUrPRcK7sehDPg
lRWIqai+NaUMsDSRLpuDyjg0DgnmcBF/dCc86tTZenAjJlNmLH6GlfP29zEQ1mplITCuwxbmafJe
F8QktdWkldKhHi6QuE1inIyRtX5Ugzu/u1FNamoJcBJkqDUbX+pUsQHTsXZlrGvtEPTwvS5+obYM
ZXVVmgXe6/PX9io3JQBQ+a7fXJFa0bumvSfRiMgDJ5bCtZ1meGaK2QZ/1mOw5F5Xi9qBD19oFvL0
RFy6sRMBajhJ5+KbLd4gmosYv5laor0tG0YyhatZehDCGR9k4jOgy8d/Zk7FvmateeFhiIE75cZe
rwrJaQyvYYSztLZb1RIkj2IzlQfNcjDbrrRQXY9XFh1AGkHKjbhYvFWZyvDIE/v7fuJLMOghwN4p
jL3o1tiBs0L2UrVjNniBH1KtlwTbtoVPPygKoanYEgafD8fPMAMWt8lNw1DW0OTcKPVsgsFl4tb3
VjCnvEy0EBoNW5hFEs7Td1w3IU2A+er2zHeKKojYwjYo+zcrEWI72JhT+/TYKTFxmqeVYfTyxfrl
JWqzAahZF9fpP5HFfpROtoKd6OZC6yW7mhPsi+/hoC7ktMfQ1H/pBNO2IYFKuxXlqlurWwmTspfJ
mnnW05ngvd8RKWYGtARMVe46whKfxtn+Mi4W09D/jRipFsdg3pFxqCTzzvxuyKuZU3oSOOeF4zwW
fOVO17E0koQq0/5NI6Co9yFw19kiNwDsG9ohVsIFIU9Be8Y8PCa9YKf9ldH1pVg9mWLzHWF85Xzw
M4d04Be/ZWRPbxwwqdrwj58GzDQQN5kb/N1wjJqLkEFKtsJB/+9pQb/epXO0rwAXGlh88YZcXGzj
IBaWRIx5fsleleSqDJno8KPLHD/LSq2yHWcy27WL65lp7Xi8WV8mAEdVhYSEzadWQE4HPyXKLoGV
IF8AjQQ3owdm1CVFw/Tt47P3wJYioajVTwB9Ruljt+38tMpnH3LqCI4Q+xHwjAfMpHSK9IISDTGf
9WDj8iNL9BHnrk/L2EPKCUGhrGt72Of/neK9MAO5my9ZuIfm/DVozYxClUp6x2HXZpPt54w1RH/Z
X1v/Fj//pE8c+qdp+Uq3gtX81togRPR6aYZ0xB+YV9/Uvg+Dn7xWw0y1zHAk4bzc1pXQskbcvBuY
EwYjCxCBz0RQuZ04UbYRKCQc4hu5gTz2OgjckLRa176ydzgZTppPUbp2gt4Tmq+oTUbgd16Arp+8
9JCO1tuPqUWbvHB7vyq3j5R7HPQcaxESzXY0zubV7nFbMwbLdg1ujyMA24IVUQ8p5Djkc6vAXRE+
BLUj/Y5ImVMVu+NqO+cT1vebAEevDp3yRcImNEyi4JlY16Y/R/UJk1Yqkp1ZCfqBa0n41VJqw1q0
EhkpJpANliEpm7ATuI0FaZwoGZyFuvQA0ZT890aWk3CdDQVb3TRGlhjdUpZ5WUMrgM22GsG3iVaY
BK9MEMz6uDkWcJUHncR2KwMez5TKnjkYFzc8yFGgpKWwyhPcthDhXvQBRy30Fg75EgHjXg48bdTM
+tphWMylLsbFcul8NgGtzln1TMhZbobSInm3mkbgm5T43ore/gi5DH3uuVLkM4t8PNQj5WfWFWCX
jvJRpFY661QPjZtA79GkRrBEIJvEHM68owOvYNrASnS20SDdpHjXze+koZN/aaC0Q9NseDkeny/d
2sLbIFM3kFHTCpnA2+EAzZ8FNyr/RkBb7EN/24aUnaaw1OuaOwhtwmEEJEvcZa8Ep3w/o0mNXqX6
wfjFCGj/NLDE9F3C+SRLCs6UtaSsUv4GSWqQVxeUuXwsA6JSb1Jv9rup8aB6+TLxBO2MCyoNxW7Y
bTopTNbNYZaJjEHNuqh6nATkf1AEQrBptZbiZW0m5oz/3hqXvkOuerfZFGWKLcDGIMw1N6ikWh/R
b0lmZXZ5P6pLG19BPO2JkJCOtsmzfYBw+uOac4oT+jV0q7d2LUw+eP6fb2Foda6BKqWrNhCr06qO
9t5NYHFFgbWnbfiVPdsUNA17GPUo8e/hG0xKzwiBue12UBDZ9f0M46jWTcVEf+jiVX9li/uB3CNF
+ZtzcJYESsIdY290r/gEITRPHgnCwjKaNdlw7ckT0M/Zu3NyxAqljlaPfPYPSE7MueDH3ibtlYt9
q95rdP9OZTSq4oK0BgK+GaQ4wpzGus+ioUkLThKdlaV24pGzjXxB7ZJ1176VAWzfq5R2TS0LOphr
WRWAwmxGsNNR+PFDzUksSinOBVV+1tjrTEJKbF0SY6Rb2R4omm7MFP4hg6j1hn4qot+VeWSc8mcE
XAel8TPxJxq8B+HiEmU+YFUWokkRUioy60ctGJNKbKPhvyaXb5qDE/oeaTeuSU2uuNpdKfetP7IN
AmbnoKL4/7+evBJ1zJT5eTGZ3C6Psz+0gSoGPQgxPDxTi59cR1A+rRfIl7xP0x4vH0zdti0pylCn
bWuh/S11nm1WRFVyB/Uf8fPv+PrWdEs2GruteaDPHQCFs+FVggob9/6z5tr3RiPnC2mO1olZ1781
4e15dzZu5/ktQ0CmVZHUo+yR1fPSMlx+B05BWuRa3lfMuzYmfm4pPDCw6+rpqvMI3sKrgH7VfdFc
burKTgH2xkiPUnhrTotv3S+BnJf18mH//JSy9Kl5/5gK5YJIaTtbz5xRc5dPOrHjKC4hp3fLb6GH
ZXNrlIFaJ4QNbzhmbUwUeSbOftXySz6j49eODDH4GkHo5+cz6i1Tu4GyXyYp2uraJmpfjhokQxyH
A3/zJuPRtPmxzXm8yNEO5v1Qslm7N2UcVoOclU/YBOWIJKwjtDCoCzrgwofWu2hmYVXpRAKwVPaA
WMYTrReCnomxN4hmtimw+pM5ijYLHP45IVhLjxifLWeP+iHmsmVkqjD+1WtJeZF0txreUNOg9aO/
pw0NEEC/MNc1nfCCRvguAZNcE+kaLBrqlWSzooxyAWCktonpZvUmS6mQfLGPg4eMQA+iJXAF+dG1
WGEOpgK6txDCXwzouZaRwr3zXK1D1+/mYupjkrW+qnuBp/cNSGGH1TlTe+eWM2CR0qpbYaAofv1u
+i8JvjUq3FHZ+wixdwi/LiWtukdFYcblWYMppzmtKZp1S0jhNo4OOa5Wdk8L4gs4aneDoOCtkJ8f
XUCKg6fFyol7C5PmWl+liVEMWtF/Z/CmISlK4GqCRObDejBszIeDwCJghSMp67H/dhdtdYzRC5E+
vrZgNg+3qXCSY3s5D4GdRrEnK8SdKkCnT47s8QyLIJCM1j16Hy90NBhO5oJjfy2hpVX9tA5obA4N
3PWPbZVrZNO5TLhQAMw98I+3XrkFF9esmqt34yppL6Gnw0buA9W5wzJn5eKhpl4KQoOffd3COa2K
ge8wF8zqm3e3viNKGlvZBeiolgVtKYaYBGb8fnhXblSCOwkmrh4Q0FvyeqO9F8BEICUrllA/34WW
qvDvNqRR9ubkKyQaFwVvUUONGoDCcB9IdO5Gf2ASP4xzfvMdoJcPX4Bn+xWU7C0nl8O0E8wB1iPb
cOebBM2fe56DitW1vm083EHlELhEXKjN6dnoPFvz5D6ELCa5yqafVOX1HfWayEWW90CVUOLD3JSz
pIdPeFdY8xHUumTe2yRpCqCyV6AF7SJv9vvFbHX8c2A9MskoXaGdYOm/OnhR5b4cXDBuJowqu76J
uR6EsGBu6iQ7tXkkyFM4wntUr54aitZy+5jEosbncAof2NGdNXrTKE/tODL535lV08EFvB6iTnVD
U/ZxAG72jI4lYbiKi3H0EH8Y4KF256rEj5i3S60eSBXIcaXd0n+VE8b8kUl3nhHkZS+7faQDENjH
Exb8lJ92sQZGvpsJY13T2nIILhtq8NVbnPxasBM6e8lFLplmHIXsvWIpgo9hFq9VKJk1BKQNgtL8
dFRLpuPgSIYJRUuG044rjWQrcY5Bkh/mdcmvCc+srY447NWBEuDmNbocOv/4RhH3g/Y/3ohPRwgF
XwFUx3m134V0ONgu//Y8umvP4sNkmM7JKA/3iqUZ/7o1U2iaE8S54YkZ/bSjR7qkE2yW4WRCdviH
Gv4aIxvYAL0FC6jmehCJdYApOEiOospuynzIkpManvTCP+u8zZyFQASwsv9L/2xA8Tvz9htbY4Mg
wVnmK+I438EKug9f+Z3BONZGn8EtykuwDGRR8xIyYkpDISinB6UT/zRJwlQYJL2OH16DLziJSA2G
UZNQIlliWKrW5/FLPte5vOgwNwW53LVRbtFYLzWYuuv8cxY5z1FFIE3GVt7ORMIUMFd5O+mqq1W7
nQ0iqGomeMSeT6nlccYzBLPUc8Df3XIbBHvzC1Yc4BDE2c5oM7TnSVwM5Wd8qhtt584ZqVgZ5pcG
du6nOomfWUMX/3JrjyHHRW6tQ01ulDukE9Ncv4h6CbQiq1HqMEvQ0R4aaszRFOBQf2EpMS3Vuw5o
QTack5+1G/nHWNYjXKovhmNSw3WZTKXqovQIu15OjViP8w2CsloIGpcZjY6uLFGEMocpqw5Q1kUf
i6UnVuDE56e+fzojxgUDTsbt+4n8RKAfhSULWhcUwz0hfLFeLk+qlXahQGdN7Jt1/kJGKIaBbBvj
7vOofMS+WdHaoW0lmLj4RIZB67qG2y/wjy3uHa8jnaZM9p/P5hNrqwCX1uTPrl8MmfSWqm9NYZkk
bC7UecnUTTdq5JRox8e5kIZRx9jLQAe765PFPfD10AfDIuuoOqPW3+ZeWSxNCdRELu0AoRe2cZhL
1VSEPFwP6GyQB24FYjz8EB/Q4i+y0yZZBDDWoSkX4/uuqb39Q1yCZBEaxv4RwrU52kLNHILZ+DZv
8abG2dHSvhnB2QPmLTAE5alsfBv90dO2mhzsL8aZNfY5DXsb9KsY1NQ49SLaWwyHfcCH2UvXfooY
tMEZxGPHT4KdBW5lJiWVaRSNJ/wqmTYLEIkW3I7bc0gdZ4gWlwZT1vqCZdZ+zMWjNpLR2wyHiicv
3S1SRAg57GHgStIdbhXupCjmnIGzoH1vc5zsZnMhcpDUY59rqCm2BNuelm+Shrw6c6YhLAMsCL+p
T0INA+bd3JAebG6KuRxOO6hKuyAmSnNuJjXF3e3Px87WZwDg1XLRU/5HTl9CjA2S1VLM4CnG3xwf
FLPcuVu1ja4xI5gwbBvCbRMIjM+mdG+FyylcQ2aAAAknL89lomeJ2q7nj2MBgajiv949TghPS8h9
rmvciCl07HHVn4itQ9ZRYlBxUMdhAlfMs1pW1vwy9ZZF6t88pwD5em7AZU/Bc7yfBVUwRAIgxB0N
UF96K9URrHk28tCj2RObif5spEq8VMgBMXwNnMncpGx3rr1DwwlF7zOIqVSGp8ZJLP5dyOBukP2Y
Y9aabCfaC59UCH9rgpp7fC66A97OrXTcFSb4bZhIdGQhlqabyjtX94oVstmF82/Qo7iUi+1FusHr
AJFPeK4xOPgN7xw9ZBSA35H/Q2R5+FiygfOX7lIU5kTthAMhs9YtBfUB5tv8kjGnrUsd4BIV1svP
DGr5Z+C6QLAk8mVsjvAm3VTCI6B+dBhXpOe+tuzc9CBLdmr/AYfuJvljw7JXT06O0cftfxrbqMFn
G7QtCUSQ4L4TS+e7IaX0GWmiRwlBHlObL8td4okxxIxhJUzxyEZrFmiAZ3LRE3yucXU4c2yWuLcD
DtmIh3Nwf5kfB3mbpxkDVifA/ccafQes3LmA9z2PqQV8R++E7ErQmc5rKlynsBbhHck4mWGzBO1L
dK6LWDswK4D2alceT/PpZ71TDam3ExgzvDs3QpnCGC3BwC28mmdAA2zXRJttcIDfNrqxUBZ8W4U0
/JK1QxRY3eWLFJwiuemlBc38Bkma30Vo58QosxlTIAiYnT6x2exT7L/pX2GmL50VS/eBvrBR5Ezd
4GK4lyU8cq5Ul/9Aj+sIABCYdGbTqKynnx1RhtpTWHvMIaUBne9YP813B4BBdOcQllxAnQ/llZjp
wJX2Czr5MtI0Dx75Ib6ycC11G4SIk4JyEZZyeZBBI0cnZ2OxwjJWba01MSFH38fylFoprPJuv/Ul
VguBDuSQMMoM5/V6uiMTlJvFvGuueUkgesnewhB8qByg3mXnev2aPT2p8Z8w41coIS8o1i8Erx4W
bfUgut4ZMHPilgDsq3NuGU/Yw8fY5tLP32OUYr3O7lE8Esj2uuBgit1tHBDLkIuxVZc3JNHDZV99
2I1Ug0ZIv1BhgyT2afIrXzHgFGbuo/RqAm1m6VGnvgazKKbt1Rsc1gZWxI0fJC/xRuA5Nr0+OuUS
CXue3tXHG4V6W079Ar8QJ8vjE0UQaSPLiZ8b18u2pC/uVgFqT6PZEOyaXvsOVHauVz56vQlEseER
VFI4q2ZuztdUoun2fEPuB87SA05okollDKtjqp4jb/Nbbgs8Pw8fuc/G7LOuzagjlUyfFL4VQ3pV
drAtCzZFi50T/yDZyBMOuI1iVel419kqHlOYOUb2fA/Wn8bMhLFRZA8iKjmzRqz7rI2+1fsjZ3BR
I0+O7j8E4EptZqMZ2F3K6NSvxkp4KvR6TmKFnjQ0UOuNaK5HqOjGUVOcs9rNucs3l2YXRBM5Z2lk
KWXmK/5BZNJ/u4GjPJBd8JfU0TsmqcZdVCvIQYYZOnDVCJzg3/6AAHvS45KvJoEcCS+6mveUaTdB
MZwiBG06oakbrC2MWLiSi6pOcorX4zcBPCpuw+FxrVbgPs7B2wXn9ozePZ3dXlCKhTR4b4939E9E
5GOH+1I7k6yf246LBDQyMBE0+3Z+Qo8Ow+IkIc1rLH/Y8pyj+RXfdzU3Bfh2uensOJFhoDaqbnge
gRxbwnx5rI8hcQdW+Xei3euUMJmyJhOioTBMjRBXpBmzlRQXTZ7qdFoj9ixv+4V6RMnewPb3cZ8e
7HwXsSRIRGjhBFN0Z1PWOyf2wJQ0h3OcH8NFWGWv67FswC1ebnbnWs8XSP1DOWUwUa6Wdkfq2oy0
8hI8FPdj99F04dLqp5Gze3JRh3ydgQ0rkltJsf4HEUvpNEN4iTh+HCr413QUT8MSPZqATbu58qEV
Tl9mTbB1+xBeuopbyGcU3V9Qz07BETrrsyD3CYEoABb+5gYtD31IwapPklr/mVoxGoKijuVYS3je
H4SeaOl8bpouZmlS88p/nobmHnJRKe3tQsAOLNfTs+N6GLyZDtr8AE6yqkWvKCTN65ElJhNE32Qs
yiRKvvIgW3z4Dx4EfI9Mk8fjSSVsIEPfoXEqvd4TbzSRi2+d+z0hykqATaDc5eZWaFRqkK5xfUpC
WhKxIwBj8dJz6S78oI7ypMYUe8KWA9BggiiCTzfIp56hQ8o2Q6YYemffrQsTSGOLI0kj+GZzdwmg
7T07N6XGwOeE1bItgMHvD4WabBzJSbdOOz3ErwK1X1HmqVhNHIWulQcLJJ3Lv1oslgFwXM53KAgy
OEPNQtFmKS3uBOI5iiGt2FSwOVUWvBaqkQTaoliMqMFI+Hg6+5sNPBi48i2FEElmvOFW77qs8iua
qPgVWe8ngoAu9pGCS/nzNSo8DX+VQVNONE+QhLShYEmagv9LHB2JTwSdtm5/be0NdU8e8SEDz0hm
+R6H4IyBNShWm0YgQI9Qf2jmf8ibImfpu6jgieZohPXV/DiR3bUwWc5cjs7UFY2dGuhkOCthm+Uh
UvTE74WxcMW6uZKOsK79WVwZdk0rHpe87BsNZ8PyuFjFYg/7g1vUX0AOnaUQSLYggS1+mk7d19wW
DH5X8y3pvPBuxKPJ6rZwClgrufsuibRscCKfeutZz2eJRFW5Uqp4e5SKEtbi4j0g+nx3Z9a9vuOD
juwR9w58DEyAi6v+90TRcUFI8kqKrUSaXPytxwaIho0Dp544pE4fF1IaiU619XXH9fcR5oT9axtQ
rpHGq8h/z0hyuIR2WGltAqNtzL8XcYA4Hv9Rk9SSitcdlr8WcVGIkb5bM7Z1Qdm3Q6f1Ft/c+uOD
Kn82+W0FJ3y6tzeAXTqZ7122azIRt0L6V8pLe+YtlQcS545yoauk1plXhXUBfAWtzTN65VtWaJLB
6GRyukYALDWhThnRqxmPdkiJqHeXezr9DFBDnsJd6RjVZ7DBsNcSbj+rJXLRz9Y4Uy/J+Dy6CDSd
R/wGWnK/ZoqgmEd60IWq+0pgm7vgESft13njLTl6zii3vD7Jtc+Jk6eiNwJR0FxHlXYGwU+pRUGw
HsugGEDxqt7c5Yi9VbC3cwyzFrb71jS6v0tE3FFXbryYqqxiR06eqTkI3CXbX7A9j19t/RaeqpGd
u5rFgOcm8WTCDjTgZb3foIvh/Sj637KUqSkDpEwMUuDbbjJBC2rWhoekika8GAM+xFIQ9Wk8QEhb
8Gw7paR4W/1T6OPFALwN16BXa7O31y+ZHkI15YZvDIr16aUYxrrWZ5A2kaHG22IBLLNtubWciCHv
DXn39uJuOEReh+xafThv0eB60G9fCjb1Tn5KPyMePDG8wQXbrvMGAVCzHnrBioWmDKKQzCt/GtI7
cNeP9MnRG08DMJvkoagrkNhLH8KtUFHAdh7oreZCFIwpWVHSWfg8E4XGYdwq0DUeozit7G+w4An2
1fjoP1JAgbBRTaEM8giplYRaZ09d8WP6lAtoHK2F5I/8Lx9iePTTS76zyp1PYOEGGJae2OSFZXkk
acRa0LjgKdCGkjqOohqTmEAk6l7TdOYeoDqoJSIKM7dGRL0F+aqZKm4Fj1KEcHxH1DPpofY6ZZ2N
zjW6tHzFqSehNgtjmq5+gjaxfibSZUd1DWfAsPOmHRJ1SM8TireyiK+WZ3cqsOvFheIa7KG53oHW
DMgDHdMAmsEL0zwwFApKAo67RKv4yJv5CJZPP0lIwj5Fs5/Fj1HnMtvUe/Wc2ORLP5NzzRXC++ND
LbZWg7FeZ1NGGpRZhdl8AyeoNX2AEABsawSjCgC4cqeQmWWxWnlb7yJrVQ4W4wy9eOT2PMOrJxOA
FkaQVVQjiiUu9xsH1LpWmjXV1WQzMkQZGw25kG2LRwQ8T3SCwzVZmHye2NIqmWKq7dR2VSJkEOc+
orWSSVgZ2vkbpntoTlH806TKeSu9tRCcqmj53/0i5gT3zMr/SISjKLM9RC+hlXPUNzCojAXfQNvX
GYsJhOSy7IvZnCOLuaEvQ25yWFwP16cutAlkibTgjAZJAhuJScLomoi1qonUmzIKO+U3FpGDhDWI
eyb9frq4Ykp6VPY3sV1GJO9wl2ypgFmlrFS8s3zKo++jVjsJpaLt5RS94iWWEscR6NbJsPexkJGe
tbq7bv8oasdXIVQAq3kStD4/snudkcdZwhWFatgm9v0Fv0WGvGDWrrV4gfh45di8XlOoLzEhyfzS
1q/K4TWgIzHv6V4ViR1ekyQ4/cKSx6/0dpsYzYu7wvyxGXXFgOgpZcHep8HpHVelCSmPP8ngLNn5
/wz8VUq0tGt22QlhK1Q1jaXVIoq3UzIZiyJRqEMOSYW6bkePQeFBtoc5Wgw3AhPvcbvxyA34h9oN
Ux2ZmG7lLqtJFpmhSDDbyZD34c+x21deAOA7WJE0hh2lsupFvP+wkPsh14HsFbRQbIQSE8kai2tt
m/kwOrPcvGnyswvm8kCu3m8Mf28FQxmKsPJYNl/+4c30Pqe6R4LeoQhzzph5kBz8KxbGwRReT4OO
TT5erCw5c1IHNEjYLf2Uy+gFesAIaRB3vpwax5/MQTksQ2zRFPBnhPqcltjDgQxOISu8MFsSyOKr
bR3PXmutzic/OvqkNFJvk6AJI9PTcFe9zArJ4IjqS0uGmOtL+WYLaf3VVoma3XJ9HdiEEr42hnPY
8B0Dh5RsjiHRxxEaIAUNFzU5Inl8dKv4u5YTpVnWRzba7xMs7HlSVDnN1b+Q12o+xkvfbqfnQErE
7IsGKVFLwtolXQoMYf/hQw3xfQPgE627JScYIejD7tYrWgUUoGSl1x3PWt1P5nelv3w+3nyDqDgg
LPApjTxmwCsaANyZMU5OHxBasYLB34QgAqJv1uszVJRX6L2nNQyHfHHtm3h7YBdkMVv7i9RMZdaO
EsgBnT4QxiCmQjfNCL5VvR4qxgvuULVeD+VivKsnQX5XgV/GmDcVDXqAlMJp4N7Bvp8z+oDbyzom
kJ0G/LOzFzsqyx2hTXmbtizpb8SByu0sRWTvU3vL0D1clCKmKBnZFIib5ewLi5Ei7vcBV0h0aGa0
tp5IFA2ivugI5eeZLmR/QUNx3i0nV8wbmhZu8rGMKSCtiSpfVLVq8sYVQkJIRjshLklTQi0JmL56
RPzVTmUY/ugVN5bFR1QSZLZwGlRQSautcmglgDI/Ytqsah+0GLHwVu72aafroTBpxaJ7puVCAHX4
N/c+HhCICC4ltwd+oDdxjqG+D74FZb5ElyLev7Ly/5Rx4ceOephH7vWXuqfsXJiuAiXToNr9x8iG
jYXHUc1npg4mJBZgP/Eqp39/FVy9n5usDqVNRcgQRmZSTu4p9dKNmwV4vXVHZ2Ix2ipVNrTXcPQQ
QdBesoOFzxRfIKbzYBA/lkfOpobX0kPMcTfElo8aJ41vdHz5DR83YtFjpnTNoo4ygTtaXX3rF1Sc
7SH87BtP96YX7qks1mBwrM1Vh91HCVt61L3u1h22j259UGXxNxH+zGQcdsXN31B2uParYIhu/KOc
bYAGg83+3HHc6zFsuPhfsnMLGsLgWtEpVqb2sk/grE6hz/xe2gL62tCVp8LgDfgbXaKdoG8MfS8o
I7k2WQ6Bgod4yxKfuK9SvmmwWfd7XOEdZ4AIF2SBCnASg4vb9yJVqneyq1LN5B89htRdAlIq4VeP
mWDLLKckdlasBMy6MflBE3dxucAXbBEjp6gGlOMwUZFLR0Ks3ukTcK+rPeVDYhZiej38y6weVTNk
GhHV/RbWRl9U4DFxGiYV5X6HRZfLy3+g0sAh8uCg8GrT8WQ5TrswHEmp0geXCsz9kSioynbNKb8s
mldVnM1iJvaU8rsN2bNZsN99e6X8CFR/plgLEh/TJWPPmL/U3kINVUcTwQ//sEWjcSXS5A62L+zm
B8MPaQuaetBN/l604jMNwDLvE2TGd2+bChwaj0yEFfttsDv/3B3lax2wtU1ufyrzDLXNIFnxT56h
AjL6AJo5GtFQ6Ovo7pTKUztJstQcSYd4AksjV+lPRQEpl2TfimJY4XXUZqyPQyaEr7ffbTsCXSSq
IfDHXqS1GZf6yiGhznklG6CE0hFGqyE7poE0BLO9Atc5+d80ym4GkxEjVKVr2t35DrhZImd+EAzX
Q93Zzvrgx6MqF1UjkOj8OfnqGeZ9t2k0yguc/eZQH1xI9Q1NmpGtuEYtg+40c8YbWrhRvQH+hpE7
U8DHq3ZJCHvT+6oEDq61S5gvD8bEv7gvJ4fVGSdMBXnYjzK1fDMSPKNDo7MreKpnnisgX3hwV0ud
3wPA/fSRHADhbcLCAuqkLWyluNX2djtrjoJnzA0/zOTAiHeWb0PioJLYRNJn1tMX+ASLFPUType8
nTnqO3/OqtPx88uWFuh76vxRydJ58bjZqR5510tURh+XLtohopYPI18Pz+7dHwGeXXuihNBGC7Nk
XGfPlqw7YZujQwTib9npHvIGY36rQQ7irCefoFIn8qllAkdzT/YgbpFStuDK1EfWE9q9GlgXqIU5
KhB+u5JlSwYia7Uelfv8wzGw3pX7aQ7KLOftaZtH2bPM3iKxVN3zcmcZPL4Of1r9Mze1p1cCxNKY
rWd856qoEkjbHyI4JJS9XUWyINTHf93r6NRuAU+6Qc5KhxqhapigKGT0L8wlB7v6ZsaUv9fEfuV2
8+U5+zoSqEcVOdf+KEsXrLfk+7jarcfVfSiyZ8lXkYssUpxUyKEveCLa976ozMI9JY0SzfDwIYPo
tO12jZQ9eVVojuoL7Pb7FvB4NKgKzgqTULTFgmPof5kkFkf1iIEAAhMNUm35uThvOcrCec0GAvpZ
sfiod6xmcD4CMYy0s/3IO0Qta+2uSBzx8InOf5d4F75PJ4YtcQy8xoYU5u5n06hBJBF6+d7Gu0Ib
+drBuQM0JhdIxjDAfB1TTpcCqbKv1CekkCOE4FvagsrOsyrgL1epiFOyCdIsC9X/tUiFGoGtPVs/
VM5eZIrNs/6BWkdBFHHjKgiTwfQApveqjta9gY8Bzp9q4C82tMDchcK3k8L9jY7yyYIahh0eAOyB
TUg0S0lhJZz4A5Qr9b22spf8kqlVmdES4tGiB0UibhRVzTYFfuZGlFjmDYJIqAcG1imrWRmnyiIZ
JOupDKOhNKWqXaEut8wN/bB1RWCGOmPnyo3rEi0pHT3B5DCnjLs00uymPTBSdPHaJWK6gC5E59Ak
fGTsM6JZ3Vgh7nCl/Us+qJ0NkKWyGOudzSYIl+X5g9YNF1DHsl/CojcnDtCp0AL4NgE9Dip2KuK6
N4FgKKQTjBIswn0LhRGRF6BZCLpa8GN3Cs9rOxUSksZmvA6XPn9LXYfQRpqoIbxI3fshu3k0UnOQ
nJc78iOMKrlLMpP3RIASHyjKZltMjUr34yUGQb0adOg349bY5X+tp2slom7F1cInBrLM0tqN0/QK
PObIbumhvKXV0mUilzm2UO77B2/4lxXv41o6ixNXYw1by5gu6y8i8OFgGHXrF8oKQDHswDkDecq+
ARt1hp3tzoS5LLxk84yZolLH7g6zDe/MhMsGMQe2JbRxKGRBGbW3jV0oxI234bE4wf/4T+knLK2G
fGjq/MCxbm13WdkHU/6B89QMzBwMD4Zo6hEo+ImOZsnvv4/J4LYJzRclMdSvpGCv7xPVbkGHNouZ
Qs2XfSscLdhWjVFsr3RuHquAjHY0tMasIqE8uDiqaSil0CRro571MDqWApms750/GhFK9OZxGBrB
C6/YnZmULjGVxiZnaOha2AIrQ/R4Pp51L8GULINvJWsFBKo9dZ2SDT+fdwDRgQaBkVWSQ+tj+H7p
HI31vvLIpiCq0bkM4S+M6YWaqQkPgHQ60DkWYkPcXYNOXTpsnK/g8uxazCr4QjF+C4i2YCLs44me
pBIWD3p36onTHnwbyIWY9z6uBagttIQwaF7smLWOspg82qJd2nv+49UR4CCmnVGOdW0jZN2GShbz
yi3+TQjHXdjlfexIEYDOFd8ovMH/Uf2N+5lezRh+/MA3KpAT3/GB13RkmwVkiv6gTskFL7/XMKyL
XLGId3JBxPOWIVmFhwCD3IbQ2dtRzf8MNMRA6ZY/m6+qdpUFVurF2tDdSK5R8PtZ4euxKIlCyRng
8PJW73tcYnRAKwfvRWl/t+eaDtoAUDnXB0xi2OUEBOza3CekLi+s3beIVvYYk0w6Jc7a9ftz+QKZ
tfiVbfVjqMLadgCfatxlt18wYM2O5VsKES9zMsjP3f0pWHtDiMhsVGVYrx+brn/hiRBTLSomQAfV
hKpZp64+D7aU31uwrnp6nLWjxHPVtmK+f8OD8l+X8h4D8osqaQoN0Dud34RnKbzPBpdCXvW+qTf1
beuqHE7C7Xd5GNexG/1AVay05VzrB5fDKge2wjKfzvibR5+JeyGfELNL+dA8TZGCqW67MW+N7RD5
2J6LklIukNie0EMDkSDoQKmwbq5uOh9BrGIqA84/3PyTxLX3IgiV3FHAPE43vn0BUWGGILs0cLS2
fxvjGeMt++S71UWGDil1sovpQH/JOjEmxvoM4DJzpuU7dxKvtA5CvNYIbY42L7t2kzrXOBoT9wqM
MJtuYjAN+qv8EmZGPaTgLVLpOSl36Tyw0HEkvbjFZFZRIZ8TWfXFo/O5yfOk3SZsqzzBp5EG1zSo
IO6jGPwHYsar/ol5gpfEBC77k6m501XeK9wq8hjSLuvqUyyBcyR9t3y4hxzoCzmddCkNhtNSeeDN
hT/bR+rTLn6OoB4u5ESmrIqclQ96DN8/S79xhp25/33VuIwhCx7uML+LzA3trhvKyB+kURt7BtgC
hmoLHun0EOuzcozVVXF0uv6qKzvmYKt1MMrzGkypTbciY2PAt/lQw6V0nsF//Rr6z6vhXF9rBFjm
7MNhCCM3p0c5LsPQB0oT8ZnxrdpcuxVqbBNslohAdejf596LqA8GZBLM8yDySvq0+vBRZupdEVW9
qp3IiuOUFrqyYOUz5daNSHq6PfaD1Np+WiEwge2oeq0kGSRd5P1Nseq+IYHtyQMCIDQX88r1d1g4
EbfEiARuWjtd1exSrxEDJL/feEQlG+q9t2aUDy7+JYQiY9Nfy+tdDesZvBR47ZFgywufFRdrE2Bg
3MW5L9YLNpeD60sBVPyOaVyXJGZgXa28GVu10LQ+YsWCuVW7R8DDV4S6LsOieyy766WPk03T6+Fg
xdzC7duoNEIM90UwHk6oHx4Jk8FGcbE68nR+iGMFBfI3iyqfo2boFYS4qar7NSu4Z5PFVMR+Z8ta
PGVBzc+B8ZCD9M7+pzTvDMZzsUvDRtNTUpkjIzgImxaqx9caPhMZcIzyRjGah0znYf7HWWzCxAZP
dkU44p/3ffMs+d/Gln2iCsi8X04VutXkI8lLalmEbOBW6zAYjEaS+Hod2R/c4Eu4tHDUY/YgErLB
ZPx+XXrevvTClfKokQhuE42KrlYjMTB/deTem2Dpd3M/9CNOUXX1J2DUhxIWQzKrJMM+XB/CsO4s
GkBKCuQM2cWraUUgomsaZPoct4W3X3RSIBfxq7uPcYwxibRXy7rsvSQSWEngjzSj4cdQsBonazEZ
Cl7DQdFxFSod4rErKhhZoE4XTnwVQ4z6zbYXoBaOgI7BKpVx4xRJ6kFOz7UbAJqb+mWJTsxl2DpX
rBSBuNPIFhR2O0DzMI75SkKmA4Fm+f8dQ6/iXZNEstG/paN9x3Sx5L4BG1xMsjC0B5QORaRQSwFM
8K4km5PC8C/8PWyoQcW0OHJIHrpuhhs6ZgxFHK90hVquxzz6q5ZdYFvvqiyaiNrhvXwQJmzPYXna
MS9II+f2/zzWCOS4uIjNRF3K8De5Ia4pC1hfqSzsn3YLnwSeyL3AB9fXXXTxqi12NW4EWQ2EFOUM
3VNqAs74uc/V/auSg+zCXDB2DE/WDn7Xwf2BZ41ytoxsksMO/aAaKovygdb13ka1Uat1uFZh/9iN
nARj+3n55VrVy8LeT/VsYF1P2+dS59I1lyAX/m/o5uji546tNRAcIpzeJApPeQuaavnZ1ilS2DMo
QVwABTtRvvbIu+oU72+JRtAFgnZsbMJWcg9Kxibshu1yKFGBfZGXeEuVadUG8i0clJFpe6msNe/e
XzqgvfyWqXK9h1pmrQXZTDFzM4tvHpHgMQVYw0OhLpfGsrSnxBnjSoB71StQfTV5honAcqeAFKdA
gcfXaQH2XyzTAdEaK5oO4joiYoHXXM7kaMpAH/HWAe7KrfwD2hwjwH0NW3TcLCqzRUyffWvXQOBz
Bfl48ta7gRh6lXLIH26bTyXfFUqcdIhE+dcN4FVkqywhJQJQX3rQNDNCspDhBSFzt+OIVwoIkSgh
4jEzZC2L91XFNNsndwseDTgTqB44Il5uLzkUGGJLBIJYaraGYtELnxtSJMWjp7Q2YYVQNo4cY8vJ
2nEkcd8TWbP7oL8DUbmPhM3DpW0E7/hzIdCNds/CW32rNkahwpmuhTwK8h7h35kRYkGQQWLdbevb
F8TRNIDAikaQ06mm8KsZ6UKqRDgExlOGggOUVvnln/kVY1B1zyC2CQnXXuyvHq3NkOPXg/vBMRyw
53oFKrnQT8/NDWnPqt+wW7LczGoJf0s9nBsguTsEuyhrj0ExByNQa8otPk40CmtBjb4ELjyvcqf6
Qi7PwC4zf8QDfaZ7mwzFkV9yEVIYyg9KQrRBBd+FokDtZx16kGtT6FEMee3+wSPeYP7m3zTSzlMR
QF2MWqIuIEFcdWU8tE9q8p1gOS8LdrJuUYmSNfITxnTtu0DjdSlDZwNuTntTkEQvYJbap/oMlR7g
KSJ1534n37TOkRnoZ2RXbEkVHdxy4bg9DVumD8pRhz5sBZ2MS+f+AUAun4vOl99agYpVoozmptSR
HJE8t2VVhjbCwyJ2vlw054m2Pypi2VCP+A5S9R3/4EfSCiiSkhHh7JIXjTvkun7aFwlay/BdHX+p
2t0EfJj/34h8qUzIx2P4TIgKZM+dz7SjXFDH5E+0Ww83Bx4bNI4J4EHj+OqxDVMaZcKE1bYBiT9F
8stBNZ5T5EdQT298nMj9q5BXhRgoFwIjB4JZ3F4CkPPsrQF5i7JP8Y4pmA1HXmXpsfMYZ00UIySd
oJn1r9M45sOH3Fr+GbMCkXI2IoEk1dEVO7urYVevxyS1CIPhh2Vu2j6pMJz/nHdHgQB22WdUkTZo
YOOXjsK1ovaBxLAqKOFld4aEpx1mTb/O51gHOHl+AJbFiG3B5Gs82VGuQBvWNOG2/AV2YbmEysQb
zsHJGJKvvThzCVpCLJhdJPgvC2YQsHSn9zQapcA6A5i6/iE2Ix1riNCho1ARqVxT3dFTSZUMuHx/
jH9s0dYYJvbXnd0axiwdR2PI/Vpy77rRRMEILoZiGog64MkDgUsP8jIWHTNjyI29PIfHsx7Uylrl
n7AJMYX4Q2MkLF7t8vgiZy0C2sUwtvADIjoY5jnMXZ0lSF15zsctJvQkWh1WRrJ1eIdk/TxDc6dq
jPPcCZC0lGz4ZXpZ7Ea1VBBN30beczQl61LOhOU787mXTA39YecVyHI9tYeFiK9s1YzWN+D5Ikwz
/icbggKhbe/VcXprynla0YH77NpJzzl1lfo+rlylajM6mgVFz/B49HElEFPgsTVNIqAmWnxFd8fA
HrTDUfhklyVBvkrJG5rpKS5ju4gOLT6oBtXYV1Rw9PDEE2TfEeJomtSGRE5aoiKqYW8NMmho97wc
t61vZLtQLnVYAfMxCwR+CUAc/RA18TfMG+e5cj34+hXM6V6eBBHfJ5456FqSXHxGlSMKFj4TY4Do
pMd5LbHTlPVNMu+uyXnPqIzCeI4ULWSc8KL0YTknXtln34WMJPEfSP1bL1kGIiZeOgY1Trys/7Qr
wUII6KdrmkKoeR/liPJYTTTVXcbHZ9QD0+pzTh20+LVUtUnCaVI82B0SDn29VK/5tpqa01EHR3KW
rMALtX+X3YUxSfnJGhG+ETlpoaRcHl/+ukI2Luvx09luHmhmAk4987abMZBxOU7AXSPhNnyOEy8E
AZJoZ0r5UxXRRZ2iS7YkdQDGf1jAQjX5gSLrdCEH8v8dFIFgGtRbz9CLbFMcIww2bz8MYfp36+mE
nZxWZLcDoBkBD4G+Z6tSpLGIyDPtzuq6KB5dQNvbMT9a/+UMxjw0K/Hqio/bvrUfZoesi6r1Qz1Q
1jPRM/e+atLjY+UdqOiId+odB4HWEG+mcEYdnseVyJ/6yHhA3VFZnf/3FkjH+9gR4fYwl/Wv8dow
8guzIKQ+izd71WnP9RD+DHZLyxjMy7sIUwfunc90gzWDkDHltkDvrUVP8pJY86kL8gstXCsLuxPv
7bdbRBNiFonmUIc5t0cg0A42xyT7BXRMyp2fYiQqKx/ae3EyIOyLzexZRgRwNTmtq7xvoq5DJzRg
or47c9ZiVSKcdvENO0Vy5zgH9/QLU6uO7k4xjs3c+FSQDvXvVVw8d3XqOJXuzkqlDa9oW9fAdKI7
RTBldh/wi2OB/HgtFLdyP09mBfK8IWueAmsaA9BNg+HQ70mzoUqN7WyOgdIUtmT4OMy3lpfxLboq
oF7ioXwvTw+H9JuYxKAWs5kYFMDPNGwgW1yMa4FpHX2T0sl1GypiYQ7hfxWo7WedhD374YGKQQS+
joDdfstBDtNKDz6G1oHXaPsuNtE4vswa9HKsoud4vRMkTbRrM/Nesbp/0JHndEZjDQWzFV0+rC1K
2+0XQWnn3IE/NKaQQsRckTI4lM5N7c10TDyI/tQZ9fZbHU447MTEEsgl5YveMt/C3oShrpj/zFfG
iWfX2PQBZhc3z+btlTmgw2Vxvr69XM+bIBC7TskQZS8dIkgJa9D/94qepKLA6JqGGP5KoGATjWKE
ssGU+DFQRj05YfZmP9GT8U9oDDf9jRMYJGYqCQzEV0Oo/v8BaCqwZ3qzgqr1eB6ZLzWGPl66/Fcj
/X4Y67YsN79ivhXn/Nl3lhSs54gGrNtyY5M8cOdvwyICWS03/GVGstMSDdTbij2pfWwhqB+Hv5B+
vfVNgwT0b4k/S16r2/IS/0XsUbxmu687iy4STxOYEdeyUexLNkF5MezHx//ZO6Js8jrmzNDwya3v
ei44eDFRfSuojxjV6mSDNQKbbVLcwpJfue3gQPVqE4xtdEHOjr9+Pn1V0sa50FMrapYWJBfXj81n
VD9kPwxxQccoVMFVo3DABbvBwnbtvvFJEgTwe77swgZn1o50u+9JBfMRNY5hoAZpSGICAPCWseda
8YdxnTxm1oiDrynM4gst0h6aTTx1sgnbGSi2s+ztjm3EfGSS8kUOAbtxZzJsz+xPX9Wcoxwl5Imt
4TwQDGDwO45tc3agPUABE0mrgTKW8ohUDwfJbd7O3gfA4oGCYRnCiQZkalQk3I4r4+AAYMT4LEY1
DxYbYlRpmBVcwS1Zc7y3FUZyl5gRXVA7y2FdaYH12UoZZ8TbWJuBXaMKp2kz+0l9XbkXYclnDnMg
pLG3ruFPV/MhGR6kVXvUDg2WtLvqRxrN76rYWk1UjtHQN4+DMgIimpu9vzF6CzBDR+cFY1BYkJMg
6375X+eyABIlFlUSTXXZRzDXWaXNyN7iOeXG8AYp+dCD7G+48b9wH6h8Q+IXnYNcWkK6sBh35In1
lkpTnQJ1C3X+tWtd5dEobVrqTmyC1MxQp9l0g81y3vRAbwOLPXMhHOjSjx2Tjf+EO4u17xbmHDKe
8YI9CcVWz8CellvM1j9ZGOe1nvxQpPzzOICNT1O7zWJI35F3fxRJb3Osw003jEXA9W5wHuNATTwl
aO17q4+Ho6P4w1xnVdPeQjj3crZu8zpGHeEcq9FXKi/iskkX/Q+KmIb4tD7AaxJ1EFuz2FKKVaEv
ROm2li3DeabLF5R51PSVGcly5zR8x4k6VDRUGRx4/SBQwzJVvCdyE5jXBgev+hbSciAMJuzV5Ll9
nfR6tmKQ5uWE82Uoy1XBP+egpEdDBZ0+Rp8oaxCa9XanXkCuorp2OoZPrz6K2h1Iec5SJx1NgYhb
iWDBQRjBoEGm98qRFR8ctipenYfY9YSDvnoPPxryCbkgTrANQoVmHy53EfXrcUL9DnHwcL1zpGSI
ccbiwxkIkIcLYxM0jtLl48tiUlluFF0BswG6WOYOjEAvuJePQtVNowpTS+sU1IDMnKn96pskQ6FC
I4anarxhSM/USOosrwbc9q+2/KrgMJqIHwmqQFB1R+dTwk2g9B6u5ssECooIsl7krRGpfPuYgnla
sM9G0Ktvn1+AYq4oy7LB9vmeb1znpBX+CAl/nN1Gjc4YGWi0j8OBDDUjsuwJUvE7xVXsT2H6LFJv
I7uIW154bfNKYkRt5gNUPSc7Izvk9Wd+DaAvHcR9DsRq/zBs7s5c/ji6BWEqEb11ID5YD1EXudcP
r5KCcBPvg5zVtgKOzyyqfQlJI/VhxTc9xIYExr15ds1vr2tVZi6cytUTuDwTUQSG4wtE6fwSP6/3
7ygEqS7WjGSpHpTlBSjcM+BA/C9oVgkCr26raNVoFaH/XLJARxYFJ3cvJH4zexLYhg5SytDCbjPX
2EZPT8BmUViqjcdDQcXD/2m3ZskHA3AGmDHUxgYIiyiYwmY0rTBWmMBl0EaobzZLSJ7HPF3fM7Mv
Es4z3k8jHu/r2h9f8DhAPkkpvGpKle/8HRpZlvDybFtx2wqotFj9XF+AOamQA1nmmt/+4zyos/KI
d3MEIkKpOdQqahZIncV5ykmhrM/4dVY47pLyYWXzUWkQLRowURLW/J0QB7kp2k8NSANVDuG+mCNU
/S8Kr+JyoUrHaGVXiPgBTwbyfETuQ9YVrISYdZjWMJhJ+KIYZeqYxpqA81wPstMvF7TUmoMhMBHV
XjCnyhi/ejl5xeMbremK3JuUGKmHCddBtesOe9iI4ZSr4dWlAxBiUSLqPwpy+QXIxO1iAL3E/WhD
EMJ5H1r/Gq9wZtEx3tw8ja6wkbloHW0XIO0VhRzwIDuMHImcsYF/cuFEErgDRBD4hoL6tE8Nmrgp
gEDZ2jnUVFuQCcy3+deL0GSJ8+M2KWIrhYI0Q3L46Grl1ETK5KhTIQ2FgA2CoUWVXw82GnMPbXc+
DYgugJd0cpO+zM/5rgaL2NWOxrCAN8RZ35dEtuPNhbCn124Oj3WjIj85eHONHl0cNRTXWtPd/szD
Vz2VBC2nh5wO09wsbNRhUdts2/JU4sENwYWx1mbkUe/QpvEmeQw6Q5Rq7tt2YfFUZ/m43GuU+/+r
823mrME7YPBeBJcLQFXtQPjL8XD+yLOPKCtZ99P4ADORw6pi0E9jFkbT+1Nw+MSu+HGW/FMD5fo9
TmOGHwQXBWaXRrZgZV4djxuyMFFkgT7GBZ9NDeSUMD8S2A69m86WlmdSOYfg0mgGccncPSf7/uFJ
IEz/4A029gg1bstl7tVLcz7XDa1bnA7Z8O4f3vBS7xO2XyLqBXb+U024CauvMp0Lt/ICnQmHOOs7
sydJkj8K+BlcyyUMbb0avDFt3T6kdSvwaQ9V9rq1yaMh9eH1dOk7RRqsr1cL1kJ8/YrFngHP+9Hz
TRuwjRQocoYkqLlaSEC+/C7SVLww0rCxTiVenAvj4rvG3OCxHYyrXae3zB3kMHGOVfmE1YK2lWIq
KwGRjMPMVWrxvZT2Lw233/7wUjVyA6V0zqoE/YynnesJwSkeLl4vvzuh4hfYxqa2ZMi9ZEMBNsp0
71kqOvlmRMYpFZAlKgh78bNTae63oJG+HKRQjJnyqwaLWl9NL3uNxbiWo3L00IPfchSgcBfcQxvH
lPyi2MXBMvDAdwQVDKZ0gzPP7Oa6ic92bciYZJsSGhVeLs+6F2KPW5LW2zxAQAaoLXsfvZBP+A6S
Afq1Ey0E5T4uodDdKQkP484yJ2qz7Ccu6Nr1MW4W7vm6Vq9s7un8wNGl4CD/Ef+E0WchtH2DekqD
umPEPfmTSQeXKa3eAHb/RaG/OhevCYAkEBj9U23YQCOEvFn2VSb4APegn59cv7HSo3GeWHCsOc+9
KHQ3o6/DWTSrEeLOrkW987xmkstKhGpLvWtKkcm3QBGugGlERPuvXsFPO93ZvKCQah8pAiqfMBcN
pSR8cTbDtT+FCGjTYOw4K+Sy64y/thsovCMOywGuKvDTH71IhDRNvAOJAKmbMpm74mv2o5oPbvbe
DLIhU6vAD1bIVPIW5zTsPRvWV1SSQamJwVAmMe6szXv/1dVG9BwGp2POpRiceiMhUXzUHrQYy/Kf
B8ZZUCa+hV2OD1KAiP7IAwfq7aJaB8u+u8HNiexmtNGV9LkXAqO+j3ui+aYGqnXxMxZuB3TMnYxD
m/KnOgbibXML0EGwj1A3/Vs4SFmK7+Fo595bUijMUZ7IzuhOo71Iwr5rkUjcG1WOOzNH3uzaA1gJ
dPDxxncryi97fm5TuCG3Tkn3mDXSbhXLH5YAvpndXKTrfw2eGJAmvGqXMujMWPVyjS5lJvgPteUT
EoiTrNKIAvk82kg2JxPgbVVSgzVxpvshc4DsiPW+V+sJ/cVMnCEYg/Qk4wAi5iCa+VSSE6m5CmiC
V41I6xgPxfev/xxxWTNY1EGYkEFVkMR+oOnJIuEcqVF4BWjA81WHFg5d0wuqAvZUzVPrllQutN5k
tN7F8p/zpr/jA8wrdvEKoufuI8/kTzmqkQ30UhCj2zIufDmh14RWN552bNbotXmmFrRH3Gl6OLWk
tBjJ1AjV503rLn3jGpp//jU9XBvez532UzSudtgAKEuwi9t6T6toG/SpsjHBRM+/dwX3MDAj3YTI
IX8V3/4/hhL72ZEx8AiK/jW+fXAkoCKjNp5x1gb7pVm0fGxT0//kP1Gv1h0pzTMBIOEepGQ6Mgbj
yVSsmLUxZcnAxqvKJJFvk7xIcF8Q8kq8eKEW/wADNNuMGrUkivptLsq9DofvY2FQVCL/ghJNxNhw
pssl6mBajGD3vIQhnbob79KKI3fM9Edl0jHoBhUKomr/Ttc3iNyyqu6K3A0e3vVmOULFiwgX3aZc
LavoEt6ycoRP+TkyjGk29+/Uw0YqGgAs7gdcuzoj8j5gg98d/yNVIecT3vZkCrfYHWfW/LOWjGZp
vIpj+dk62pwzTMKwxtAqIxQhlTQ+ShHiO6TofMNT/oUg0y9KPCn6oJAjxnzWDQ/ynj/yMT64hjqM
bmtRTHrIXmlGlm70QyTsAsujsehGAPffq/v/KKHdkjrWnuVKk0LI0ERRy6zq84q9BCVixH1Et2VK
TqMBy25PIVkFlJjM0nfraQ449sbZWndUrO6COxRHhX69GZleLgGzVIbJzmz/fN88vagAjB3ZGiC0
nB9Ci295Hbsh2KIcaUfsbhtdih6i1kQGn7Cw7kf0+RsK1PddPZTkJg6IuPPTbnJv6ex7NTZjwztQ
RivMyU5bh4lzkH3qDhS4pZEG7yUsOElnovPKvkCv5/SoJxtZ8tUtHV6w+oKardIPJ+di0rpmWsBn
LOjKLNSy8e1nnfvHqR/20XaJ6mytyKe7YlB08TMGUuZj8UXP0iFGSKDcEqobPLfZ48qUfcxeRkA9
/uLsdyvq6RVoGfsy0m64HCqwZymPLp5Aq/U93q9zen85v/wcYhzx12q9whgzMlMcJa29evXjBOQA
L0wmFeY4quMwrIm3zSKKy9CtEUrzIRo+JKFqdhDBNdlLZXpO7zawsgRs7TEQ5AabICY4C0LJniJR
hIVYEnztDVahaJLlFSBbTslPeR+LuqbmhRQ/8Mw/IrWU4ev7B5bIACWCNVIJa44dje4LKwzs/yXA
N3SLyaEodRpIrTzpXU2kkH2fEvLIVW9RJSFxmPXtzM8MLQytjuHrrVnn2PnzJGoOrdWfvm1d8ozQ
Z58mq3GV1wDsQukSuDxARQdDisHHASWr98HcUSPdEDq+1TZUqb4aWtFjRZOxpqNlKKb3EYMyIe+H
duql70hHbl6Wr0QNFhIGNq6nczWLAaUsciatKwSD5rGiG6kDuu8tIf9U6sEalAcK+z26BCir6Fq5
pfKsziCkRLCTnABDwU88xInMTUne+S5SooFHghktSwBeLgcxjXZ/94+mFSZbaJe1DeOZlOpRCT8Q
LLi7rNGJOxdqMKHuB0Ga63XyCZuDjSJbkHRY+5OIOlmO3UhsvGglNaLXteS4nQrpWxIB5zNU+OtB
9GunmjYJV+w8w21k1PuC6GpybfYPRliVyyVoKOMdGAWvjxk0OVztlQgWv/oH69acx9AIKjKNgM5Y
5VpAb14Ywh18H3zZZ9Evm45STVEtlgwlPFxCaMZwWhtNdbHYIvocVENb/v1VhK+Zd8WO84H08G4Z
qpitFlE/0X+aGqXi5H66RK3mhpi2l65WuJmEYHMZW7T7o6OiNB0PRfgBYz/J2TCs9belfzZmzSiU
8BJ/1EurnULJLfzWOUCh92ZjPJv0x2uUoitIT21GR0wFGS0AMlaOV8QJqDyVASu8xDAw+j1ByspG
xi5wvKOrrT6KmYp4UebXDAWLFjhsTkCoWrR9bjLKVjpYPuZNqwcuHW+/MrZdYdI48yHJz/nbAmJa
vE+rudapqFXjQy6iceF1brz/ALvp4jhQ+aPC9LtHKFWBQVDTcmByWe8BaVxgHqd56+xth2QZGFXz
K3E4b+091EZy4L/auK5yHM+b1GxJF7JoyoBYQlG45xuE+popNdqQAZHvXKNXwnWuzkLgovnr6xB8
M6tIx8nDjNxZZKw7Gu0Enu/0ocw7dCq1jPv+jSCqVQZ0rXFC+RY2HgXd2x5Xb2adAWXZDs8TXjGo
HY7Ch5U5kPIHPEzpdr8GLcqlqyAQxbya8dFJ5EKrL6Tya3xgTi4cqaOd+cdPERWCGtmMwpuUqf+s
OPwsftxGq8S9mf+eKAwDkswrobDK72c2t8kwpPfW1sD4gvJb62xXU7ihWWpwLEh153nYriJNZ1Ew
SqD7yxcDEhWvJCaCBY7MgYAWiNrYK4wNOd/MZnh2rYI6/rAdSv1IyBPcW7UAMNiUdkqHIz4oyhS7
wD0yBpEa8zRhTHT1D+xSILR+ZZ23TQkzjwri3fAXdW0E7nGssD+xAdDHrJTLSbt/lxbrzMfX4H7f
WSpoW49qoejd198nT4LpgU207qVSS1F7N+srYrkQes/Yz5PpPdhCRAaGrgVHh8wpHVClLGb2G9gp
sBQ7qYZvJ9WZpyMVAzQvHPQ6AcGZYF160QT4QeX4aV5TQrEt/dIOG1/NIM5OdCWHWDLBxYfD3F3v
oLJ7RuMctBsvexVnZxwK+4J5PkhGcpukPjfFpUlrWjbxhAdOzQkNGmrssQk8rjqNK+KzOpIGvGWj
2f/p2KpcZXXGZCJ+dcFdjaFTB7j8xoelx92z8lNM3qAnkl9dATulcMZgqIHTLhojvHmXRub6iLBD
eZBNpIQVtN1m0U2C3mjyN3bF/8u8RwqT4Iwdvpxodm9EIElg+45BsDmy6BdYurof9aj4TjmIQtwc
0qGqIC4ofTp1EyXs8MfBg4n4R+VQyrKQfa88LtHB/kNhgls9tESttbPTsLoCvJ1RfyQtelgdJONf
RVraHxuN4KERLTy1dxzQSrWZbOAGl98BVwtrcee0nvJn7k+g1zFPSKDAyCH0m6f+x2ThOsZ0xX7B
z/Zz3xJNvtFMdk0mcDvaOYLpWlQdFI/le4r/VGsLpw308yNJfQwrQjvMtOoYTxKsWY/Lsw2UyPxm
7zU1cOqZYjn3UW1578mxUyS1YNlbb8yKjGA4UMyhXd/Oh36qAIUMejkxJ0Rt3PdD+EQCq1P+5kf1
3PnFkOA8fZeRFjrMhQq9wT8/hH6MuSbbI41EvVYfvsKC971o9hWjcV2bCEMJ5APvINGhdtds80mm
uadKTCbi+T3kR1sfvJOM6aWqo8deQoAKJsBRRiTEm0j/Nk/P6PXpNdQL275W4oN/6IySwkhUC33l
8AWtMY7jpArJAiPFLyY8wKNt2uQWgb8H6EqI00Cr+mvZr1Dz9dKnDRoEWcfU80B/mM/br5Futovk
zCWsxdHYGJpc7+rblrZy0rDaJlOrFPiAezlGYwpSILxxsta70UeazVJ0f667OBlog4j8JsosxT5V
BUuEJKc7mUD1q7dQ2fCx+L4isTBSWwGUKkl8GUw++1xlgqr1Kwb6pV92xG/P4wt+rWceZjYfPUim
lMcBFFc0fZ0AHy+F1PNJxWMjuhfhgfRr6rrznWH7QON8wJQSFfsSWE1qelv5Pf2ySuu4XkX6faSu
z2JJM2QJcFdFD0DBBFBD7uLlRB2OSTG2zm183SY2FJ9i7BRnrdYP1CRSqckKqSf2/EbfK33qsRx0
yd2mjEu5YOQPKg+7jSuNccpyV7mQmgcFkUmnCjyAcpa36ju2biL4OAm8Ru6wW3GBd/7TGsnR2uTT
LxBYCNbKjkR53+rbHeCgWImtwdM3guMP1qT0uSalKi3n6QeOzVKiwfmRhU0mTEgq8FtCN9AXMNTG
L+fCDVgflsAaEBFU+zGVDgETkjMZf69TLxhYSVF+NxxjSRoWrGRejSS3LpKt6zJzkTgf4I1btWKi
NVrIKoYS5RakK4Ft108oldEaVC7ACMzsocw8xAMTax3cm4nCasz1X2j6Yt+juGYXqLUmEN8aCGR3
tWnBd3aD4RIJp2YQoBvPAZI4nLg2KirCKLoM0KHfKLpd10m+Id23qIjBXBSjfAPsxAyRVkfnM+WS
wGhzBjMKWnB04IjMHOnEA2fmaCXM8JqdJBsk/p9S5+HkR/ZYn+xo8d3KeZ67RIpWXMjOnoufVEaB
EA0GydPf3tRfy7XIzeJqSWk49Jaq3VwUaeQ/JMkQ2H7RCeQyVRKgbrb3V0K3Hy5V0K5vfRQrnpPp
6hC99leX6AP4KC6w4MQ2w0HDacfJ3H2FS8W8IMxztV3UNAxOqNJzNBitvu2a/XxWbWqqjpJtLf3z
7ivf+abkHB5gJg3446JMOaU9sNkL9IW+InU1AE2C8hMOfyLBURssnR0zcsnqs9NNJS/R9rO2LDj0
4uRpJWh4hnLqSOpVE7cCrNZn9ExUFPF0StNFN8VhcfnKwDUcDElzByuCEFiXDT2uPs2A4w0YzTg1
22H5HnYPNBy7mejPLRCqz6nxI7znDcNXrnmcVteoa3YV9Ta2+QP26oBHe6C4xMm4ExAhzUMuf2c4
alV5xmznLifOhLO5RXVx9MXkKcqsjxbBnx+fmxQUBg3Nv58PKrrsa8ADBvcKAJ3QK9OvXd6QJlfy
v4xayY3Y27WfX8XSVJ2ls7aneImbRzEMC/cGuoQTpr8dL7O2U/QguuTsCXfsmXd/gmXftIbqcx1c
VyJyr0bEJJBjRbnyLX+r2xn8ZmJJudkj+VP+ev/eqWGh7bGLlriUwIYM0UEjsq53oOK++HZ6Hmp6
lkPOnYlFiF1Wv3iyOyOo/z7VzWCQV6hg8ZTacP+H9OPuwe4JM9D3bsmAK05yNNE4tQplLqv0fui+
ENyS7XMmQt1htygNEZO2RAi/2hx5vGOz4bauACLulJ7qkey2f+HjXtp43xanXwGVt4IczZxs+1tW
Z09kBeX15as//IURu0jXhbYoOp1ExS9t3aXJAw7LKTF37IekWXxlrrjhRASGTPb9HpusCx75Zdoz
04P89Yu44wh9MF2UU1ujwCplc3Y6gjmaUDHMScVw61SD+G3VtJmBuQVrlQXZlOUJR7Exw0uwO6M9
WzqfWZY0SaL8ZEAB9VuCiDgLzwdBjeVbeXhNSsO0RfWZk3B6YKyAJyvsSoQIkc4SGTc3L4f5yc2S
VTQ+T7HIv0teBf3XunTZ7mpu/5ZJAUa287KdzQTXKNP4Ru8Nw7/bTkmV4f+/6vEFyxO3mAQWjoL6
fT7zQ41OXai7u6mHEI9GVFY/VeAkyK3T6GnBv7GCbzKPNXhAbPgSX8nocqObsg2hwKd4MiExU/XE
94dLDLuEEql1x2i2T+vw0hHIqkvVFpVdghAyJqcFJYsGF9OnWRxxIRPDzpW6jG8A3brjtxpuulB7
VCLKsYwJBSSPczjUVBBF9lBRhhhaK8hHv0znfAGe7G49SxHm9107K77i/qtr0y5+ptn9ggQD1+NL
luehX5w5ABZQgy92RR1JyL7y50DYqdPTKHsiBwv48GfQLEo4/imidMNXURq11cP5TvpGAyxlm6aO
5V6P4ZPKT0sw8yacG1wcdmVq0t3CGA8DVEtuk7l4btNDZqI5S/6zbeQKZp5ZoMUjt9QT/8Bqgwdz
WICr7q4w+Lvs+JJ8oNoFH7AkaEcUGGe7Q5q7fTfXJbIb49LBZNaModQ0328pxGlgzoCKoWWTWJo0
anPoJbaFjWWC8u8Fp3BvPNx4AHmP5Ri5QtWquwrSTXEJYI+xmYAoRFOnVhsvmvBSDsUtMc7mH/nN
HJKdKpWdBy8KpGZp2O/brnekLuBCQTD6Luf1vVunq71rLDvPBogeaN7JMTbFkKg4VcAc0xwsxeZj
DP3Hi8w0Yx72HG8x/iu3xitbTfWPnn4N+va+blGZadkZupf7BolsTld/2b4HBiyD80iBJHZJZ48u
c5CsurrTaTxtcwNNGhjVlo43cQ6pCVAIQUmdj3fdNb7F0A3too7eTluu3df/Gk1Xc0bQm4dpUGbx
bXWUeHkbllM+ZRdamT1X/hqmSwzPcxX8w3wJQeK+iDt35awvP+iJtlzkjkvlV+ArYlTIHGtbdE0L
ZdSk44pOwSe5CipaZpseKfkcg2wMJaw3JxyrfjUDd00FESYDY21qWkwBDCjB6TnSLETU0enE6uKU
E14ZNkXbsgZsSLYmKeFr4vNzb0dqXqQpPkK0UDFMFqqxHHYjZTG7t+kip3b88qeIa2PLgeI+RkeZ
MyiZBeRwjvc6EAUZR19ix0B4e8iPJJkdhhWLh6cUJ0eHQwLejmL9FjhTKqQmyam37UL3YuF/Mws2
e8bcFXRdgq2T/P7BG6RIK/eb69/6m2MMxjbvm95dHNux/JpotxT7ZM7kohTkQVuynstS4QSGOzTL
9Dkm6gBVSr6v3mle7gO8V9zv9C0JxVWW0D7JwlNiX5p7Hd0BdaiD/iHiM4rjqB7Fg6dZaOzCVEic
Cb0hOK0qs4qzMQ0CBdk46+qlKP7gHZdrNw9mbqa6W+E4xmMyEJ66ISrKgsTQ7Jt4kqg72IsvfmWP
XSXm9KIR/Y6N/MkcTOCJVSwXHDuJz5cplUhF/UfHg4db5mMwju8SR2QzNAaIN81l1+cMePFUkjR6
WUa8LSkYOULpgH0O6Q/flSb7rg8gT+0gtmmAmr/PClWquefRweGQO5OJP8hamdZAwVyijeJKUruy
4gpBoOFIST5wZb6VAevMiaB/qXoALHvWyeuNIP1f9KhRjm0YU48YDcxErCKEIVrame6AqwOh16F2
jFAKdHP2vkd88ceGlPmsYOxY8iXEDGSDgKMRSW8YB/1NjamhupY8gExEL0Yhn0TlW+wY828Oh+TZ
TmT5xfFhMLdIMfNwA+OuKCkvYtQ6wTMFHLJsTgdU5lTNbHRjXGgx2/7Ayxhv2N4nYFX+zr0CyZ/0
k3o9bJAAeXUMRGa5Xz+1dItzOrx2uyT7Rgh78wlUWX6iP8Et6zROSKTFT+Y8bfX5x3A6W+gwBLgn
0gsz7LDvdmriHJuxHChB2SPQ0boOjrCtpD95zXu13r5IiJ49CYHPj+hW2v5e2ywjxftr0kCLDiJX
q0A/aVN3SgX+TFeSQmp3DyRD++gQUPpaFpO7AngbEoZX/bnKHyrLe5uiJ2hsckWzL8JxkvDxBu02
8NLAps74StpxH4EBVxdhFZZlwY1zv/NZk4lhBoZb+whSYd9WNdEAcYWLuPP8z+3O/zasQ32hbSGu
bfYRH/q/z8M4kq4BYNe3xgNgT2Wvy7MTVnRnYyTts9LcgiNJJ4YWAOleKRVVPbxDyFXd26RY5kuN
/8LwxRA/8sraT+gaTN4/m33X4J/hgP2l3J3VFlMZ7t7w36eLvRg58AHrVVqpMeU3N73aqv1gbDUj
M5UT2n3XA1frZC+KA9+JVFdu0PbSaMk4Oa0TcNIT8am88N4VSVjvBzJHaQKOmvLjXtkUu44Tf0uV
Pdl0VV4swSJJem7EABT+oJ7ZGrkZRBwCf0LzaoltQJCXfu9LqLyBhotiVHQHJOLQs+dg1KgPeR5n
Z3BCfqrw+tBFtrl3gU41clrbPyPhGfrFmPtQBXpesEFHf8iwbnmlqBghDhE5Uy1CdXb+kw3KL1X0
f2MWyLiCIoGz5ZiOlpyVf/YVLg2KIuL+fJpIC/d2QGpaBFxNo0/vI4G3fqR2kDiq+fgk+DtW9RoP
NrylkI9cLQN5R9Yo+6B3TXS/DVV1Z96OP8nmgKvVvEFLTWwJQZ+hwp8p3JlIAYTUft0p3j1Txhyx
skiu0Lcr7x1J7PW1JNENYb1UD71QhUWb6WtvUfIQsMz015Hsx3mbYoACxRuwus/qRFkrZCImfpf+
pcHaqd9VvfyW5sdQ15F6PXewb/ZxeHDnvcAAw4lb8ymwf9CrrW2aIGQNCiBf9Mg8BeHsesCVyfja
O6foIlh3hV9/m+6DvWvUTs+qIGbpQtxn1U5Sm0VoA6qq2IcLDykGJBVmDJv0IGdMmZEFbJ2rloMC
m0Qke3ZWvACeK4yJHYjX4aJD9s5izVuKBeOFdznvQ+JHBD7tO6KUx9RQKe1rlahlBrkBBY1yOiSr
aGpwNPWjunH2dmYIPUGGKX5/z1wy1cHW351K1qFLSxV1qTC91HLGcCQTg1VGPDOHuvgAM9tjBZ7T
7zQ1ut3eqiIAzb9jzD9UlsLtNsKzjlYzorTwnXyu+DhNbGoP7McuQHqHli6RAbHEWK/YLx6kj9f1
a2VZTm6WCTpN8fGzJm11IU6uTXZ0akln5GXuQJV+Wf3vxOlZW+hz5AFsjrnYaJm4OxdS8lZFeps9
/Voaay1O9b7LImb20x1bk997LN3AsZVjay0kEABmjxKGyWEifSXL6e/E6IuWyRMFilRf5hc+YOvn
3NiiR415YwGr/5VYncILsGn8zShnEkujGr6N1iBINtTrEZStdgYUMs6AUCkhw8bjVYTVSCr6MYF+
9x7FFJbB9fJx69IrZp4URid6CpkigSlfv+tXWnF2e4oFz5p6QfulDGbSPTpL714IEm1GL2oM15XV
9xhI3hB2E2WUUSj1PngpSbqoAwtAbl1qOG0HEecx2bUYOv39Ai8QqpxlJGCL+RjJAiKwna5gBPNU
k/Hpywz55rK3ydn/fcEoMsttyX5VlJeDcZrpl49B1A8ckztN+Cts5GP7LVUjYaUlPxrQwsJNr12b
aCkShFpyzZcdhZ0RhQtcTmc0PlaLy8kZ68BR0kL2uDE5NJMfOSinHSO8RYPSumeKrbl5QPMiMJee
jpoZVNNzL6szWXVXQeOpD79VUnDMIhqSeo3IpRo+S4/MrEXWUWY+iyxSWUgAk1w5Iy6IDvOCJuWo
YIRLDlaRL3+K1ZDHz6n0Z3NYquZk6ZkyXuFNK2nA2/GGZ9e8RiR0/v+LrSYOJ8vThkPasmQUEVv0
BoTnYjCW1RR2HUIYz/BUNPbyvCMqRpZ0mrRK2TVMFiF3vcE9Z0kzNyaicDInM2vr1UXtmyTRv9MG
JsWw7cdm26mG93S5kEQHoi7b6P6V0hkphVEJ1DfDRijoyOcRGKH5gxpGe+nZYlBABv7KLxpCytuV
Wsp3lBC32T8/oZ/okBMlHoZQq1yn/5R1d+v+UFh4Qg6wzF3tLFqBFojZpMtxgWcdoJHrfffr950w
Pt8B0McJWTrMWhcvXBR0BXdfCQ9Q2e7g76eQRY3JRV59xgKaNDgNn9+snnk4f/tRoQn6/FjWrj/v
xyD4Yio69DXBUpbEs5eGNx8SuYOqacUPiDxIPUhpLDuZKRGmCbee8VRPXJxh+MRKYQrpew6gtFEt
j7pb+zp/6JoX59U81YPui74WQdrAsrDTUT3fdIbMMfbn8k81i0o7KD4cPVLDJsG9P46JcbR0Lblz
J7Y1SJBW+OalFkLEAZkp0plsReBaUZgl3blLD3JZdT2ivfKQQHydgNj8htM3snaOH57bhn/wFAic
6SbzcTnhqWHvuMZ5UvHqhDLyWGiiMSZJeY5zb83T69qK3s8n4HyiPuakcrQKGiRiSlxOHe0xiS3a
ZNSTZin5S0WYBcRMNQEajIhJXpxRoR0faXm95y01BCGL3AtUj3yaAOVKtJJcbdsPRw+sX1Ef2YmP
AthACnz7AuLHqWHhkxjhxFoSY1Ll89pOFY205pX3pV4BN4Qs6DeFWiWw2mFNh1/y/dCVK37x5TpB
CqlNd6toCQk6hQ4Wys+kJODdSWXmp63XRU4AXbxuNxfm/NY8RIplPmbSUi5NHwGA128TrzL82uBV
KVagjr9/a5eszH5zQreaUkv4Z6aJuVZcPh7+pPoAoo2Qx0esy9OMPPwBKcDtn8YnFOFi4xj6hOX9
NromoTBkR/BhNh99eC0OgYh4IArSOn78dSX6jvNWT2sUZHp/JsStopLunmW4Wr3MTDvwAol6lHUG
boaUQTQt3kmVMONEcmfJF3SbLtVNN8deQ6IFok90Xb9nQQBCF8tADctNuKII1gaVB8NLBxQMjGS3
S57I57uV99xB3Oso/FXtUxoHeioBR4P+NIq8+cS5QkDuV1gTYNf3Z94Lv7tcXf2TD3YmDkuUTbdZ
glduTE8QubB+jXD5ST5ftNbZvncqZQ2i+dMagDJltVzZg6Jl8hRj0FrHfjDn43Y5NFf2Ojdl0iG3
YOtVE5LSyTtpx7rxpfnXdnQXFQJUkNJusGAWaBvZufcq1vaWmsRN7ZrTygXB+IB7Fufl5ib9YfqX
57+9KJhaskW3j+G9fUb7HQd2+I2D1M6FIVsJT6eh3KCamJWxLtRpCLcEIVqg5+rHmbDh97icunZH
mPzKCXBl80x2HAzFfMD+88VS6/jP73TP1FRKk0xB1mf6FDiHLMyR/TWSuoPi9DdwFPEBnSBHg/ns
UgCk3LFpy6aAXEfcgS9PjLxWEW2EoI3YmsF77MoYrL8S7hm8fwKmcdDv6q1M0sSmlMwkSv7WU4S2
ZXrOSTuzlU3e7yFv9w2+ru29+yQT5KUvm26HJupC8upV/DhofLukcm9SCwvQ/ZmRvF/r3vUMkerD
zbEPcGSqzYAIFlU55ZpFdEglQy8Qz3qHcuAUuVPRI1b8FlzUOimkfOJZ1UYzMS4cfNtL+RfRPTmM
5sOHlmNoYuiWVTgzVXnALH+mrmhuAfTInGgtGp2pvJ2/b8e/K2HVkwoDmqBZsblqoun4I3zUVnYe
HsilkEMTtJ1zgkdJxFN3GxHdWG8pQRnlJpO3LBHk27oXRaRCsBY/dl3lStXNpgMFITym0tHdmZq7
FcezNzkVJnGFJwtZ5BYApG9QUAq7Bjb27sh4b4v0E9T8WpU/9h7TzBp6t4QanQAt2qBY22ESKWaQ
eehp24DJhhdlJPVi+2S8OorrLWzshr8XF84fSASjih5SOklMsDQWsX5heV8z43SHgKE6QIhYGZRh
uaFsbirE/p54Vjfea90rRxlP3vfHeIUdjnU4tDFKWZ5i6ghJ7baN1C19LvqtwYw3LtKlQTovi6m8
chTavtcnrplBvbqkZl0w8+J3K2Hdu0lyiYSpM5pGnKdJCqkF3CIXjKTKfOA7BDh9ciiO/5uv/n+O
8KTqCr8CPDaE75be7n4Tk0lCLoPGPanhA/gb/SK7M8BkVWDqAOJdSQvd1NVBo8DgoIhakL8ERhAh
+I8hpDsXcwKmaRHlF3YiDLrY55D60A4iL4Vf9sPwYNkyCNEdAYZhph4J1+VcF2OtMDKBrcd3khNI
heogBv+LkadaBIyXTifnH+rvF2fQ4haGgSMji830GckST0FfHW60NLy4XGy+yL3MAbgXUtYj+QnB
OPSBi3yRB2riQXSD4V+OQG67bTQRcSuCZtfKlU9UZjaunAogEiXcbnuOsRp6R35DndpL6CJsKvdO
PLbZ6U20WFNVHXx01YZW2NjGSKmxU6gcvvrAqtZoVd6Iub7815lInYsjoIsU3gpMVIPsaGNfSYNI
o8FW4iHKXgt9bL8yG17ur6Aey0G54dbUshzGcOqYVgPsoyt9jxhHHllO1CzGeESKfWewpo5hDQZ6
vwPEAGVdxq7A4NUVsVrnPcHsDuvSXVxzzFgO0jIqoLHbjQxjQ5blkY4cCRX/gEObGXjFNFK1OQlX
zLQst3RJe+1JRcno+EhVzJJdDdnRQq+eCelyAwsQgSmz8a32Db63sdl3hOEn4p0fvxcEoNN4qfky
1CyO9buoO5M/JG/+vXbD6H1RNlnf9vzMrPmKV/892oL480al7tuno2XPRcbjQ1iY7mADWf2mcW5F
pQpT4hfYsr8w2h2gds7n9BOz2HXy4a7mcnTfvT4vFmKkHDB+vrTByV3LnSugCiDplx1cBgjy1JcI
mik+Q0Aic795SR8+SN0Yw5OdSaULZBOEugewOAXQbOtNrbcw/r1b0iRnNbaU8fVO7eJnwThzwN0t
Si6DQ4ZGuVG2oZQsLXa5Jjtcw9kOIAHaMXGUJ33on5bKrLDrcGtqTMT6A+5hyZRfIpg/81k/RFEv
a2njaGAvlrV4WKYBFt7Ldy1mCH7RukA/wE0JPHm7EOcu1G6sPT6Xk6PozK7PKxsh9f8UjLiTIxz/
ZeZdPSjUg6VTvqaqziokVnutxc4BSxjkRu93tnBPCNzBPo952GYmd0cGdKLssNLdqPRJWvTI5Iwa
Blwd9FfvYlXaSP68qi/yfPCpnjFEiv3eoFNTjY+1YjaO9VLCzrIdvCQyaBypLnUlaJ7Mk6lirK2k
/0GSlcwfGiHOABEz6E6091eu46IZrN0W5s1i+EVDdxfUdmQaH8o6mkpjcVBTqVYdyvqdXxmxc5Yx
of3aROI4MNmsREAUfBAmJI6d6qTaBSUnb3AJQsQ8TKsRolvqi6wDOv73+CV+iWC1uNyCqfqxscjl
HVS4dwgq8mDqxtVEOg/IyjS6wv1jPMx5sXOB8C7Uzw2xBBFWQxBHVGoMelcJkFwf98KZZlCjsCe5
QaXz1XWPZ/gf4Go0YoJJ/NhfbUCHKVzaucyrSE3GENqUTD0FDZB3yV4PzbcRdr6UPjfImu95RToK
EDCDNNscmU8K2nIkInGb8DpqBTty7Km6Xmn+qkrBVGut9/ygZbgS2A14vaukXrnzdJxYCP4GwviW
B0ToH17TEQnCtNwfX+GXOAlJoDP98IeuWNgTr1LJkpCgKP23Caa1KwvX9F3haEdf+YiK/7T5HTM9
UhzoZJO2ChY4pgs4UXL0eAcwiHZQrjGyhWb9MMKO5pYCfyBM4fKY6mwOv1lklb/JRm7HeRkKGIpr
GNmxBkR7002e+9mCKcNwVX6pcx9InMG2aBaCys18C4t3hskilwFQ5le+mtiw7SRksq4oI/UUu3/x
AN7J0vpabE6vmem8Yt8l+4U4Ao1mql2ls8X1Np9279iExyPRgk0xN5tHHgYO6xpZv2yzQPDKSMYn
cNYAhW/4wW7bsf5z40jTKh9qStQxPguP2JmQVlbOmeqiTc1de2lptPwa/NZToASgaz7CZi0XAQvi
sXPPXdRUHoh4Zgk921qzc4s/CusJKg3+1CsXq0y0ChXsv8DT+FRybhbEAWnvOx+hZVtvlkhLZRT0
PYJ3HTytWvVPUjd5wPaX8b67ZFUCtGVHTVH4MNrxkKVOx+8xhPnMN1pB2Zoz+HpCPEacQtL6fraV
J3EcrAyEdDtLm3sC1MH1NozUCc3KUGPz0EjOP9iY09xd0md6W8ODdMdIzNacq319zML65VdEE9Hf
ivcvwMY1GtFaVsr8Cj6MR0ESv4+CsESrM53HmoBvbHxsp6IRvY4bjEyKHNTPxitmkkiY4uV1RYPJ
M9ymM3nh5YRsUKV6sk6/KRUjLUoMm/z0Gh2WYtxiRvPa+pE75TCuPBM6vZZTAeZz/u6qTGGikc4w
fgJE7YAiN+HmO/BDsyOEZHnwAEp7aGSQYvLwHu+OMr1brUqK0VYODA8pJHRa6VbugfJq5/6Bfr2F
ZRwjdYKiMa2RolNV+U8jgE6zy6Ngb1W6wOgmpLj3aWRMnWMxwIn/Nx9J/OG0heqgAGiAxS4GmVkb
xfjL68uyjhUvwuw/XKGB6lRRiCcdKuYEGw61DHMOokVTGLa3n+7c6f7z4F5RK0jfmfJONqxuin6G
g9FQRbke/7fSDKT1kErCFOa0Qb0gtPbHn2VKI9kgra0CZOdaXti78Yc2EnGyJDfSa4PBvbwp0Sjh
ha+AfZ3wGXFl6aed0qzR/h2NEljQkQUMb1QzffxTcMqkLPkV8BNAfFZoInsnt+ABb9p/s9Q/7Zv5
MjzlmTYesz8xtUc+Gf+jeaZxBBujlGJMh/0QSxcQFPAKHgBWDZKmb2RYOmXhrA+Qz0tl5bmpWEZw
swF2ekmw0xDOp3v6DNTfvaSWPDiuwQ8bUZ0PlUdIznzzeia/j7jlB62NcaQ2YvPLDUKIt4n15H7U
FEpCg3ej9WmAEpPuqAVetgiSa/kwt9cCfdBRAmVYXJdEv0n4sN9ClWXub2rplzu3KwgBnGX3o7Ud
NsrnyGsQ4H01FS/fbCHzmdw1Y0eTDCaY/9HZbyTh/UDODroLaCAbAgtLWHkIf2Ovpy3BhNRyOQik
Inoxlolm9DN8HlQAlrEh5wz/IxEPQVxl9xZUvclNAQo9BIp66ETIEivpiYXWYlXQA7ryYma/8p+o
ySPUzNv6A+8JMM2ZPKHDmg9oFRjl5qvi2WggMpOHLd71bMUBmy9yKekRNPI/YWfx8d1mzaDN17S2
u0vgN0G5OAOx+euxuBon69gtjCA3tM8ZypmUwYfVzA7sEPwJNT1e0eGJ+scebwAAlDqG7iPjJU38
3nH3qbEwFV0NVj+KMVTiljUFfPolQODj1nqiKCMCHV/uCwaDXmI+uyNADbMCD96IpF29+Io2rOo0
OHJDU4VJk9ZM7Q6aMqQceayigSThwygK1XJrHuk0V5pRjS94W1YJQVLKahJAH/IKfFkPu4TrTs6x
kM0Nz99RKpABdVUUrBEryc38IBiqv8n4hSxX3ZR/7l0Aigwx/9vRLYISdNxZSpSuF3OTxCRb6yvD
dQXhMP52kiPhpZzGKUPNKF9JRAznNldgW9BTRw6wl03fQjCWQ7SIFOzw2hf10XKR9gGbT32xUuIB
kNIvnk4Q2+RminK8Nzzwo5+wqA66DfChf19Ke/Z7m71WuRDfwPBdG75NprhgE75ycM3DCp6kCsek
UkhQrhhii49Mxb6b2/7LIWO8WYiBNWoE7+ACK3QYlowpA5ZSODyto6DuqFpBDKMciVmpKrXyll3I
GGOHpE9o6QR3nZWtmSOSWJfNiBwMBslavO6qao22b5u4Ua3swPZtr9ivTvZ9NojpQnatVbWNfWMu
OzNE0dJ/+eu5zzqYzUj459JkR3Y1HQ/tfpWL+yT1YY9ZwYBsOsakN84ndXmLI0ZTTkSCeasqjxrG
PocnNDMSi0rzw6L3GUZpvRoP3050DGyC7Ri5V63+yW9wcWnqo+Iz2q5cCMkbOrksAw/FR4pP6yu6
lywasNcA5l4CDHpvJVfkZZ3nefbLlKKsqrsPLBDLIpxyKwZ4VZ+7zF1jCLkRoltJg3+Nq3GLtgHb
Fm3qL85c9IAZoltLblP70dBbSBTZET5xBoHbS6vISdyOHLVhAEz1Qg1NCf0dnGugcYZdsljXpsLx
7bT/TL61Ks23Az01UkD7XxgplT/vgveX05UDJHiIlhkhw9qJ1GU1Tjc0uXeuOv9WKkXZNtKJmqma
OLhYS0cQRq74F53ESZBhBYbMqI5tgOrT31VnLjwdP0mUhnzp/OQzWYrxaO1RxC7NSM08pzpY6EX/
VnNipUQ7MBE1ZFpYpQPFUCv3x397361ygwE5n0exLUetf6ZHET5AEy7d7yWY2e/j7pwDz5DtNvpJ
0xrHQ7nf8aL3vj0kJ7/7nKaptmKMy25kjlxpswY1eWfxQWHfLOnHHeP6Rw7fYplmQnlPRPOqe0Wy
Vjjw7fgUEK+ptocVcQzPS5es8aKSHPAIUWAvO33k6pnSRrlppKqlzQVNOb/K6oRwl8YoQBvD/Txi
B2cLsT0UZSp3T0HPUPG3YrJPIawv5f9wbjBNrtPH1V8bOhEW9vp/L4+3MhzA1d9j8jdKDXEO2b97
8+e6Iv9Rn8l2kZ/kZKmPshiy0NbsVoAPcJA8ZJT1nvO6Vj9OnpCubusl3vFfIwbohaFDGaqECuNa
+Y3Nxp7548xg/8mr9SidCe+RowGX4oToJOfgOC+tQS5Lv6VAqJTocV4f3Fs1fCJRKhULcyVZgyxa
2YJtU9UWpk++vA/uePnkdTdvD/9aEl/K37HfktGc3Wjt6lGU8peSdTdJvh0A8IveDd/22HPkyW9h
123dwqj+TAm7iBbccz3fsgJ0pvghztwsAeFqcAXbmqG/tK5qZ1JJErFuMWltwWbqwcc40Ksvhd9m
CQMcgK8yeDIeELBCAFBZgbwrEkxMXxIeg8V4mekRHJHeTJCaNMCSMByb3XO5weGhsKv73nneC1jU
aCjseWVDtdx09EFWRdj/fp2acCjfo5NZX+tOA/C1ZzH8Yb2kHGD78T6qEuQ2Mb+h/QFXzzNR2wnm
FqZnSXxVPdWy5B8S4FpuNB/saEOfuSYZtxKe6c2zbNime8p2pCWoN1pJImGXpQ/BGnmhE7nLB8Ya
RtosJzcAJ2DVlw1d+kua8UjtCBHXIQzBN0Mi9hI3wcvtU6GppsMGrRrI3PIYHFnLK+rPFe/icUo9
NTuuATeW9gASTMI7Rs1IUv3JdyBGHDom972aE6BrKhI43/vZR8fxWdXZ3mpAIvSkKdnTsYUkv1BU
cx3jXcAA0ONvJ7GvEDQEBoX0wbflqobEpeAqp5UhQ4l2xIxFzg3kXyAZ6mP5plUnM/QLR8qWmMcS
mzIUn2/OWRp+9n8EglXHGQjVUxFuSGcg3HyTmGIFZ2zT7qk5eyrskMHU1cTm5SqiVy7nSgJrM5Ed
GIghyDs+baCuxJMJr1ODoUoAL86B9CPn3yRgk6NYXllxmCz2Euq1XHHt+bUDGNZxlHAy9IWow7D3
0hoPzBjx3k2bnQEYgr4LWp6lGJZPzmrg4MEH5ijIbKztafU57cOpS3QYDxKFkXN+KLwYh8DgICl/
qDz28zKcF9QBYU8DlxrGL71o2JkAOjWbVSL1hQJ2RL5jQkKRjORC5JIuroi5rOXCHuyzziYpknPX
q/cfduy+emMJ3xFSCYPYCM+V4kKbEOFxnjyBVR3QAj0j+L+KrhamE0s4msaQjUlMZhTZRoVSeq13
8HKmF18NefUiHffRi+K0x4AiLzY5TtNFTFK45fBw9+6oPQlGSHYbNz4/SZPjQp4Fd02sddByGcxm
evFy8ycjXEqJWTUwk2AIm7+iuAs4HQMTVYH2p4bnedbsio02T2KJCZV/nvMZLDc4aBYSis66UlBJ
D5iuGudxUp5ywnZBqxyLYHEJ0xuRFAH8uZV/CK5AXYmYU3D82nYIlv0/FPsV3j/3HJegSxestvC1
B/uL59FuLuY5DdHjuCHlJe5WGgzekopaDhQsXYNgR5JmCiOk3v4ZC85SEU5ld276yhFY0bsIGAei
zJWIrSnmOML67xXKvjWQow+vGzEPRrh6ALCiuPV6HtyJA+zbaxBfoEvYc3DxUM+Y/+7A/TMIUTNg
UgrQVqDfmqLMZwr/8C6FgZsE3T8NlKUWRbwrZT+0yF0NxWpmEq0N461Suh3KEA+vsvVM2VBqfxLC
1/p5A3G+4Qfxx/tMJx1Nxg7UWweSxKgatBVIGbXy6Jv6ULhnFx1g3wBhDgHPojjeTod6VSDQec+r
Au7N5wAq7l0a+HTGR+f2R0AAi43rnBXmi+tWKhVJi9rOd5yAPCzRIr2aCSzX2Nsc2WVkSDAGIjVn
zkCZl11PbW9N6VqQOEGhXwphIsRXCcpH1imIpBpqTPenAWaPl9T2qB6ZSk9CTd/m8yofFBSU0qvF
dFoxf86X1Wy7+JcvqM8lFvGmGM+jjosU0AuxwdhqeW4oynG9ITVwkvqPZpGzx1N3y8w3p9/ElcGY
ZhuLQFGCX9nmA+aLthqEhxTKGT5gHxmv5Yh8Pm5g70MjhY3MkppJA5RTUi7zoeYOMSTQXUW7Tzo2
AbEPJyo+hAu08NdQnjAGthjYu7NVZG0I/G9oG1w813H3Nh6lnf5q+M/EuNtzaYDJ9SWvW7W+tYCg
USC9xsUYQ+THTHSKk+i3KjhU+LSIuE+yXsppdtG1H/RAYuDeL4CDQAvjPMAs2cE7eiziUlug1wqR
jHOYJJZQJLvN/PUYe8UC4Mwt4WE3tQxoyJ+XhVt/wNZjoZs2mh8piidM91a/HpWcOGYrnp2vVQbd
EfdSl7FJ8KF5p2+f8nL3KL2AyRJHwpcRRsDlNEXn55reSqxVJCD5726cxgYmCZkNiQBdZbJ5Egvc
7jaZIpqkpHSQtMcvZC3zH1JESj/M7id6TBdUmY/RRKmdenj6OMrjb6bEffhjBSB8JUyziDeolOtB
2NV8i/myI2HfZElYeL3U+/mvG9STRDx0p/veiZ7aT8fgmBJnhN+tmUzWrusfZnFZI3qYLe5nAWzM
14HlE/ADsouuNeVpzCVvrJNtocnm7Cj46a/jUCLy+CrRItgncOfrcohaVKH1MjfqUcPkEwc/A02A
dxVUKiD4cx3RU0ZTtfQ6rBW3yIyvXBEtZ+4B9pVlwJubhx+GO5HuPf9BILQiGFkczmsthLsetVWB
C14hduB1ezpryS4rQ7XXGIwdPThrHEVYrSnwAwVZm+rzg5QCQ3obrGH3wxSeLg8KB11Aga2MuW7a
lSYxrKNcONPpdKGdVxcHqqeCiKELpTUjgHS0NNY1aLaB0rfSHcQoUV6s8SL5g8LFMVgsG/kzGHT+
V/4j6acXgXWb5dpSMOYS6n0zJp1epX41T1ik8fKX+vspF0hwAA7DWKBg518IdrlVjyOKFI3fKp82
L09OXCaxCHX6MW98Mt6exEaXiUPCXD7o3ljR5XVAvlmoyCEXQKDtIYCljtE5OB7taJKP+tVrzemp
FXGlhoBQTAX63aO0yr237sahDJLCtOEttCGNpUQZv6Yj1fz843TB6QcbHz2IPlC9t1daqDJ3hyFk
Af1nzXCtLgqK4p4e1tlWWy7B/RcGdjEznIdmBePp7oAJs8U7F0ylIvG5Q4Gj9uxAMu/Gw5vYX/97
AX4tg4W9hFg34XMcWxQUuwSUbLahgTljPHrnj3Bq6r3m6/JJUkqqdKdm54WDO+6zcLuMpRqkHEvT
eWgYi1j4coPzgdWPc2liVlfNyedKKKlRKSDMl1R18V/wQ4ceaFMYfKcldwkPPhvwOqAG1nTIUjG1
GLfjJisH6qrlDLLmyuUwmlYgIc3/BvtRxIGOGG3BJTYdiABLJqfwP/G+nOYnVqW4iOF0qCg4Kom7
Mp0oU3w5n/DFkIQM5lvRwQ4Vdr6AFth9a99aUO3TAQwq43SNR0OfKG3LBwMtsj+Bw2Wzk/p27PvH
lMQzq44ZngeneLJh5FMkLJzdWBnTX8S6vN0mmcC8QXvX+F/5ML+h5bmb/yQbC/97ejnEyLfvW7t0
baCfSG6THeF4N431BDpPjHml9d4fQb+zq9qs5kcQhySNr/OwzeNne7pqO7pEYEibMNZRkXJ3KpG+
hsYgJmpbkLPymo97rMzmXw85C515LD7lfu/5kImBfzYEeKHB127emfdFxJ3hxGLpiEyPtOUW3ebx
a/D3JfJ4IuoBX8DiXniirzVo5qeIIJffuYXNbI3WuC6dNetx7moS3NxHz0Ui/7twrvS/Iiywm5zl
gI4jn/XFeNROpvmIzAgLJfGKbNmC5mg+Jreg+mXFlAmDk9sxmM0Mt/Qy79FaGxWTMUJ2RyEACWB1
/RQJmKaJY4BAMU9jZNpnYCqfe5H/SV4S52yryBOuuLviqdsmnD77beiSStlIOGYlnkEbJU5e9IyP
o90RG+Km1+c3xfYy0ewH9e8KqBLIwwhJvBrqgXgIfplapmO0OofuYGxjdGWJf3ocCc098WsZgaTf
TY5AQFnkRv43G/KXHblIil2iHe1FPjU2QUk++YLH+HcXrjW9dNGAPyy+HTtKVxPzGcEY5Mq5/8J+
bh5H9Ki+7s+f1AYT4pb/FsKRD9MR0pPqJqfUXKWrOq3f96sxC7MLRtBl8gMQ/sxHYXdgb3y2Vsw7
BDAdwVl/rWpLp4M4dOrpsYtNlX1O81Qkex1XfH1fjDClBY6SDiJxtogDe20hNLo0jrgyCSw7PpJY
IlXxZwurz6hI56PEj9BY3lIGBkurwnZp+bqWtP0ZQJPLouKpYQY4thqnY8PmGwXqNHxeHsRvANDO
hlkpb2hoco0UrWDeHY8hZQwgN2uwzG1pW8X1gTjCKg5TVxjsaM7VQODG9KnWsztFvSvzLVkCmLQE
Y8Er8KhWk5emfS0z/cs+9IzmNXuPQOAUGQbM+3qa7SYpeEv3KQXz5UJOTGwsLrALuXgepEaQzP55
hy1RdwpzeFpI+e5UsuTBPuOSSjivQ6N2HAU7gnEXZSI4+vz1f40Fd0vZzuHfpqRD9PM3LirAYKUg
3KzhYTrrwrUjSlmp2K5lsQpL9EQraMtCT98dgfY23p8PpEj/21ddju63bK6ZkCbm+P7wtiftnO3a
Nt9aubU1DPlnHSEYQxOQyckzekMi0M84JEIn0l98ZtbXDmt0Y1Hzb24M9GbW51M+jp1jqt56vOpI
txcO1MqUlG3DRmCU84CakkAEH/r6Hwge9wEmJ7T/s0QSyWhyNY4ewlEkjwUegBx1qDSe8t1fPQA3
FjXgWLWmEwpH7uk0hz3AO8LxxXa+DzLgalhnrFmgmiwnG7K7kPcZxWdTi/HGHCcFYH15x/+bPyUe
zQuFBDz6S7/jxrei0+xtY/CDmerKdWfLBNCo0Aa1ResDrp7n3RtqDIPjZxlaaNl9pkugRiNOcGMt
XyTkRbsXncbik0mSj8Fn7w5O8NCP/69AcoKjmg00A3DF6hJe1x/XVCM8QzuNRWDK5uVwTRSX6rpl
3Nf+fDgOnq/R0bWJ6sEdpi8X0nubVJCkZijCzTxnuCAfMEuUjR13ceegQAh2RArlenIh3T9ll4E3
Zy0XBjsTe96DMO4Qp1vhf50FiELVhczclc8FglIJsORdojPQTRP0KEB8TK1FT8YTRAU8UXomAYQ4
aU0B7bLSfjpPOioYW09l4mbO3a7LqA7FnkIyy/vnKTm2+dIb52XzGNfAuTYmgVIyeNjAzOzHrLGb
DxlYfnnhxtP3skDJ/UJ3vpxAbqe2g2VY6PJ88u5otfnpbbrFb6i0FLG0qCh2pZ7zAPK+Fi5b4Gdd
MyKx73xkqsirl+EDfZq8rJInL5poEnCSqgWCCEiIyR98z8qRpZJlSVcZfG0ULJGMBYp6JboQXZuG
bAmgqbLAgNvQ5kG0u2BUyTC/yhCvQhiK/yYCWwo/uZAt/r7HNmGf33RP8boW7/Di/8zRMMAYnJyH
HIVw83NxwuEEpeJ54ansm6MqZWETum2Oa/jHwBVQTF4gCN99jc+IDD8OPIXniKPbyhGGh5Z78hkp
JAd0pIjm9M7eSdZVS5YK0d9m962l74WJiy0C7wn/fV1VpZVD4uciYBRvzSKFGz9TicuXk6AVKpR4
byLu/TgSy2wGOHQL3Cv65cZbXrTnkJy9d/6RFGmbbFyrfIfE69oagqXVn3MrOQNXgpzOjmTyoBAr
ln1wsGBgcjpcESXfS+s85D7VEvOZBvK/hHcUSqGzcJas5iDKaTkZ4RmRi6XCyicDDwT8Lr5XDKVV
dVwxJFr0T+JCL1jThASxQPwpGL1s0I6x8a2UoLX+QydeZIBIsG6XfaeFrQykNvc+GDJrEg2Eqefm
60kb1KVTKMQVDKsS5rRAlfMRjATjFN/Vnght+HcF8VRJrfHevDX5sdHpaC1MiZW0A8JjIMPLhgWm
DrGoLppR7REFKK+hzoJg4EqyH6A9U1FDUL6+jlhACzRnK/8etbyKrOW+b78z0g7ZjS4ivgVyRvMh
TjIVGms1edt2pCVXMtdIAo0LvRCtt25+jjKMUDyZ6dBcuLSS0D+n33CnF8NkYN71OyNQ7w17De4D
AyUFCrLzNuf5yOipzitC4YPgMSXwYIZBfxHAAeivG8SzsWYRqw8j4xjRTgNcNfJwHLBattDvy8Nz
Bc5ZYmbk2b8Jb+5q7Fk7c4UUmip+6bLF8zUxmY6yLq29cTzKK5Gb1k8IWVhFKaG1ETQIUAseOmcx
gzmdm8Xg722Cb7TKg6vNcGDljQHpuNA/677gE0Z4BIjT0woURiSQ/vo0yEtdciLhr7UWbAvMm8Fs
gRzhY7tD2gS0oxoMTSyYrSgG4b7LKz7EmCmnlo2sTziIi2daLChxZS8IIi41DwArTqrQ0qXhMBQ3
GnVq4Rct/rnbtVtf+O1kZn/CHqgVLIYb0dUiwFOmGGqsLvvhMyXGkou6B6+KXQ7icm6C0EwrYIWJ
GxAmUi02uPbaq6l/EA6xfya+HJLowfG1S3iZXZ34yiSjdTEZZWXn57YTiSDl1uLSdpEpsjuoMr5F
uC9lwNDZr6hpbJjW5i2Ag7POqMgSs/OrwaUQ/vzwQ0qnLgXrrHHnfhXJrOF2LOK8+868/EmpN6rq
+Z+mkfyoHadM7QiUyyWnzVVeW8Go9G3LFumT/dzX2cssoWNo9t1oQTuTU9EBjcZGwfrxNP7Wm0HV
AGSQ0R9ZBIvD4duMnhy0J/bcO8K9kHfrkbmJa+NDILP0iVfq2w+UqPbIXUkT2lxX/jwKsDDXg/YD
W8KNBFcs7OGPBsjnZks8vrhGZBYaLlPLK80JUqLtTNLvECwmbE7+oqeA8hhxSyHFjM7ETRTonNf1
+LQMfGWUQa4cRADJjhvOM+trhxUbGgKnhbdK+h81pYHMz8DpGU89wq/QsTU/XkwMCtaT+u/pVz6+
XnMKvmQxf4yAbZeBuDZNO4NKHSH7hSclfGN3+Hd7sWsMH2k7L9lEdugfLfwCMvP83LMy+3v4Fq1U
aq9HYPOjeuF6YxqWdWsIVgU74ocvnRLBN9XLszhSrSGN9CZR25uKfXsoVLtc+P2didfD4AUhX+8j
wbvj63ikhm6twaCW6f9JfXCQKMrRjXuWofWo2c0epJUn+6pc4YC1o+vwaxwh8cfGld7e1FuBd8N+
tmAHndTapFYO/5u5klKdHjhmiO0f2moO+X1wpzxJ3QB/lRh6BTPIkr98JQIreQ2XwdcdvrRLZOaF
Ku4VVE83hMFz9r+otTUsDqULkJynEdCYBpXYYA4T86xWyRZxfPD9J5DaUh1jAltf9dcM4JI0a0fJ
luzbLRxnHBbnWHLrocEfriV2Je+J+cxfXh815KFhJGdOXhARuOAstQOKmSOhhhyLeoUBm3AHoYrD
oQ+xGxX0ShzShiXWXvzbtPRdIdXzeMjjBQBVLYZMJDhW0AZjBkx3pOWzlyLzhygSw0ZWo6mOW3Sz
qcJ30b2KKVOd42KoaY1qtkfMnnHigi/Ji+4PAMLhsemS/U13Om/WDRv5k/8zOe9QpffqtRTlwr9O
1TwhrM67aW3SchxPMpdWdz2SGrZknaWyUX66usAD/ZAPxKpuHtjkLHVlp0XFiBdn3cVjTygh8BP2
aiIcIZM10KDtbvrBlGX+E3IDEWESx784Jf/LWotV152v+VE0ABsPab7PUZau0SKuGCmP8grLyvPx
+XswHdLVYcEW51MyfMbotUFg23XB+Kn3jHgsz+5ipeCzo9DL1Pq108/vG6xGWb+9rKA93PzYcrL+
rEaD9zldY2d9RoDxtwawuu/EZVu4nZmByqHYElr9Tvl8UCU3rpnRpk3Vi41uohUcJnkMR/KkuIc7
UKg9znCRGuldNk5bK6EEZ9xfl/FuTEYQoQS/Kk6iJGymz3T2PMXz+1fuGrssle4Ew+g808+O3Op+
xuoKc2YdAJAOQsxAmalIfuOSL2bOE2SRW4iamCjVVIAo8TwjBU7qUaAJCw3ldes7zrkU6xhFs+7v
HVrHmZC6SOzAhJXV4rSnYQZ6C5fD/wII+SU4RtmyPYkXIvsFXYTvm79+3LIcM3PaiBfHtFcVyTxy
oI6mOZDdzk5tPVF635wDJ382eqK2Vz7HldhsLwr6pv8Sw7PoHE722KxjngLGcQoyGT+nMVGO7ECG
RKN5X0qIHzeXPq2qQhYGaZYKTmVrcCTC43GOQFrwAiWGnqgtdEkK6j7flv02T7rSIfbeqqoXBS0E
LFUcRcRgU5RHuAUYcHEs+whQyx40I3JNQIqqvzmvELwHJjepJDp2NRwWE3UYT71TMH7rEBa5fZ3G
LB6gyfAhfDsatACpIbMGmX8qHYaCSSwvsJxGoP+G5KKlnNBjEgw+x9HH9113eGi4Ez+w8I+orP6u
UyAONMcVveVbiLdUyYOC+CB4g+JtLKHt90my9I9u5unVtEJjvFAUPIAcRKOi7m6HeV9zK16W3Q5b
m67L4cg/G/egh1VQHBE0MaqYXhRHdF3X+5ZtMEansR7t4lJRxZn5jfofuCEWvCxBuGwymI757/oM
WFfCdDhHZZRa3NoarCh2tFJhDvR75nYXLK5mV1a8vu6qiLZrPMqNBeAW9Zm1fpbGBvFRKurm4vzN
9iAPywiFYhc9ML0vA0JuWnjXuImxqpsoh9J7yTWrHHJOk83flnXBmoZ0FCS8N9v7pHyqkFmNoMqP
6TY6jm/GvMTtupdlk7Ns16Nrq0UvszsgjIahbbWikwNBEmvjbpaShDGBUTsyCb7xWWR7phyxcWRq
/RZEF9t1IAyUIzGj5VA8I3a3XVvr8y3khO5QSloruLy4kAQebo7VLamFYBYrf8E4SFZGO4lf1p5U
ZzsYfiz0MJb4RbrkUCY3/r8WXx8R8Lct+l2CriLDir0ImwdmOWiONj6BfOMZiyQTmHSHsoGutguD
T1fHhWGwBxhJHwVnQ11PRcqY2ovsM/I+Q5TiDK/9nJXNaLs/B0BDruXuuWHzA5zJPBqAqHbjiHfp
NOrpAwCCG3h8gzOMD/w523XMbLtsjO+DqUdzNtftg1uvQglYIsLcFGgu/wCdnZBR3V4moKsl/7LM
+8XNz4FEtgrmHZHkvynhQ8Hr1fiCdAqLiSTysQrKqr6XkRp8Kx28kYsvZp0d0/Mzm+bfzXtLMT8j
iAf6Z8xoccUoqB08tdMvXFTuU1OEtt8+beXZo27Fh/fR0bKMdxZPVEknWcmVCCCHbkN9QxYpaDQi
FD8UM+tHk0y4mq77h/n6uxscl+Awk/6LTSzJqwgmlszFAV0YffwXekQOyWmh/yHdF/eP8Q7WkYTA
qee83XgwxddFstez2sctTuTVLcNZPG/MhL4cMNS8LQ31KbSaSgtUsgHLS+I7NZSdDHAIuoZjiG19
wxYFoVcpvZzhmsMJ9YSvICHg5O59IyXv1fuiXAQk1mlpExhqtqp80dvdnRqtODn6bWfwWSLEn6GK
I7IUzRioCM+g4hMcP3/Lzdmhm12KivXRKvOu/1rRr9zjq4afulXV2Mu6Gfi3jvQPl8F8ndPwQvFA
Oe/ean2WQObrwVEY6YWQqN7SZYhon/2hKqsr72FYKeVOn+ib7V+6njuoD/11+Fvn7FrVMG+HO4qc
nt6UGzHCpLkSwVjcqzGbUJqdB40QyTYz3vRJJTaE/zQKD3jZ7Z31drb4pjsB+3jJMaq9Wp2D7KZj
h7xWInPvWgOi7xXIQxxmAJg5Sw+QyiLFIDAHk4pFVMzSPSlCRQK74d4Lqx33cfb39UI/jlRZrR2A
rxei4sbFhsorqfVzu2e9rh3mfizSUIxV+1hNFy5qHmVc4T7FCi2YFOC6Dbhm6OpKJ2pTzj6qg7Gd
Ng8OhUhfbXeRC0R2tohNiFZEEgMdhvjDtqZlJY8weLyc9e0Y0KO+oPwqdp3bXrlKAeKeLgr0Pddd
zg3y9FSIT4ni1/vDdtu5+3mNVz2Ac4eLrQaPA3elqBCGxHc5+kyVT6Dhcoi5racjxR1CKeue6Jut
m/sNLqxeAJeOrT9WhAc/0XI9KY9R0ouVuu1PGhkySnCap6+AiEt9zMBo9DdsP0TbbY1q4lynWBsD
NSjHqqRevr7q2an5G4iNgOisN7qFCgKCKRAi2nnVNxZHWw8F6WrqHw4//xd9N+MHOjTkZ4bTlnx3
nZLmzRrzk1ShR8ygFAn1qxbvgoIv2VS1kUhlevW7XibutkhqdUa6IieQi5N0zvtbSDzZdcCdAYYD
LJAdeoEOPx17lv3507nf9xNTSxv4uogYTfP3PN08kOC9K3mHet6h8XK8/mjxlzzydag9PpvQ/7Jf
BbKzsG9RpxXUZgH5GUIvcXboB+2rqNFddYBgS+P2H5Ax8tSdX393siKAm0rhNH+7Jz40xOMS9Ppf
NYfGJQFT80CBFBTg+BbkL3ohhIMff8BZX+TIgIZASThUPdyqvKeg7D1oY77emmo1QaIzDzobYEMy
PwLpgDlIVX4NLtd4EBGFFKo8YUwsHJ410fUINsPALGleCmiYmOfgBGAKBfK2gUCSxxhBgfR70O/i
9ej/03v7BrCvqBUW4l2pUiq3sV0kVRdFqSFfHvkTodrXatdciBfJuAjWEB+l/uyKRr29NUVSpn9e
k0C+Hgir9RTyNCIUO31vtqkVnE83u8ub1mBLj0Rt2iNnuyWQCyhh0lmHxwiBcZUlJ2u4LXJB41kk
5tLkpqwQnEjz64fphmStHBEPW6XLxVSXPWSpTPmrF4lFgu3Rb6rdq3PzYzMSlUbsg3EJjfJJPrqL
k7BRyTZpH96IMgd7MZQk+yABgdVnh/FJEfhgksxXMHFhuwJ7zpZuET4wybtDSkGxNLhILgiemlnl
eCMo5q6hvrXaSTXZ5hiMSO5wfJtP2Tg1hKCpciVx7lvgSkePgygaFnIlNq9nq87UcdfzlL9Q0KrZ
a4ajPS/U8Ug+b3PZmnaPp0u8KQcLznMlD4Q9IkK6BO91lEfmm9KF5/5T++fCfcDM3hradozrFTQJ
ahc5oIIZDcOfuS0fQj0YeqbtQjB1I8pLqQQ5bk0I+MTKUspqUqcy4VLEdd7bTFFCc6JksmkMi7/L
F8WklFO5S3PiKolV++S1KRJjw9wLGXr7nm9mraomI3uTvzWwqmsrlPjlTGrtNafyn0VNg43uEpPq
RWmsdbu+W5rYJURPmlZD/Q9iwrp/elgt8FHYD3G7WAJWGyTG+pLyOxA71qFqVwS6et7oq3+Ondnc
Tcp9DfTTnLvXCxqoGWp2+FhD/JeoxNQMSdzVi3XYT6xGbdhSqzOmt5sn4xW0V5+4CUPUEhFU8FEd
lfxfip1oahUGXCovhk1wQ6k0T7helVa556+aQFGGRyQ5vncIUeOyDW8RFGK7VUflw+6MEV0YPtgV
x4urC8uMwqpyNTuMQm0IjAK6g1Fkw4WIZ25qlu5duur2GkPgL/yG+ipCXmfJjjwkZ+uOdiWIYZSj
AQBIb9R6LUsRNZrupiUKIW24sBZfbHkxsD1++oWrhbUwSDc4bpUJhGbsZ/UFdDeO3mF00NzX4ySG
lR7Jixo3xh+RkZUW6+eRbToLfxHUW2PxpjevVBVdmIcoDz5Gye88XwH5fhJ6eBMmphpWxQmMBz2E
hwV85rAzTbN0SMjQCO5UUxtdz5b8uXLwEjzbhL+F0LUi05J5OMvU3V5Y7+K1s4js9u6+yPeeJn9W
LG7b/kYEKo08L79VPffshSINB8UOQKhtskVN+FsbmaUZshUqGyRRPF8B/I0QklxETIplL4T8pWNp
5y2sWAs8S+7dNQc8mw20YSJsDfRV1GIvdgXIc1PME9MhYMDMrCEYyZwm9P/it7t5itL4EfqB4GYZ
lJctx6dr4BD77L5ESh3McbTH9jHZebUi1pYpmvB7yzWuRo6qnyHlfqDJ+mQR9RJJRV5kGCqpFb0q
7cneCSjy/Zo0wabJfC/fnfBSd2gNqlci9pMnOFKz77PMu61Gnq5qYz7OQ8YObPXigY3/QfPi32AS
vjL4LepK+n4e7sxYEcfOGZXgFXrS3MzdnWriISsTZBzm2s3UaWbXchYO4xLoaqUYJDmDP29IBNxk
uehW2P0OHQkOF5HXoKv9B6B80UhkxiffUpJHwmIzZKSh2QSV0JyqMuzwe/V2JFQAhii0f3VBXnm6
S3EPH5Q4sBDUV8EozL63Yt+mbn1XF0GPXM/jYlPh3YBXlA2eErN2yM7Whfe4KfW8L9hZXgHHBkhP
BJPKLVFOkylNir+iPqNwjYoA5xrEtMfU7koYhHmKsxSLszHt3lpsTVGmcPqtdgHzGYaiKTAEjsSA
lfNSikPnEUjDXl2cTDCWnSJyiSyOzji7jHLVXXcNfR2qh1GMY5jLRMTglkXJ7wljGZfIZtfxlo/a
Wemvrb1iMGjFhkZH6DCOc9abwWudlfjZsNuynrcxnoCr6NJ1UXf3o6OQss/7Y+ArhuEBixD1kEXX
dcb6Vhy0V5auI7AgVDi8pJcJ0v2WxLyuuHJm3sk5o1oONVo7ocVI2mvUu3NJCngyvY0IK9H4fcpz
9wjG2BwTf7aFusHLLPT3uwklwzWCUMSC1msUEBXi77WYuEpG0lpDgYwF7dDMtCO8UDp1PkDnItJy
Kl4UWlUzitjr2ZRTxZEDhjPdeADu4Rbr33HfHsSEjqPabIsGcby8jU/0a4svb2jFCT8d63pN22qF
EXjokLDv3ABT8LxC6eBqygnFeQmTdXV+5wpgEVhzwZJfW+kfbFeec8Yf0fHk4eQStEIgDHKJ0Z6j
GAgCmHrw2pkAQNlYF0N10MMTb34ZVZ3nfBSbF7sZFCnC9mpmaSkVs6fxcHmz++eK/+RGAGsuntdD
D5ETtr31hI1aO9vhIAYPZjKNgiUjQ9exxUw2iWi37XXmoYIprAqkjHzD039iEX92ox//+QxTKRXH
jhImX7HSCsHHpiDCXvtQFPezTcOFzPoJbttivIFNkEdaWbkK89DvRDKgqpZpf+zo18XwhMu4qOtX
8ZseK42nyUTuHJ1MbpWXDTF2h5KmB7UftJkyYjqHkq0zkLpXNEFJtf5rpzqAIIXm7vEzUu5dHcZT
uE7+CK3MMsSABkgBbm/DeKyZ+YUjSo8dzjdOqgskXvdPX3X43D/8ATJI7iyfpbT48+tEa7wYcM14
vR6CcNwRHE/kVQjsFntKw36+Fla1fsegrFjtpyOFpCZb6NcVdaM+NK1FNVdC1sBPoHn8tLEqw9Ka
51znneN0YfzatQjW7ojRR23D9u7M36M51EhQKO0C+0G5/meArRzDXaSZ66RXUYKIsI3tGDnAwDSV
bmo+0JxNmBg3K5wiA0BOdM0P/7A3suka1yT4PQmqfReSxVzhCn9IJcQ1BFnvthKHQWpTSjEnbM4l
qYKKQ9AbuD6SKFu7WrXDcnSe55tlOfRk6bZTCUvN/Xs7qBVJkiThOkuvaQzocRRBXYkm248+Q49D
cH8wpMkPeW+FH/d0/EUhlx3fzKJIwNJIRgyoL+eFvy5dghALu802mlcAUwYeeFBC/PLeKFLC+drU
tGfTlDgURpWGxVBBKileuLLxCSWuiq2MOO6H+ikfvWVPar3llNcdlQnThSUAu5S+R1ghl9+Dq9cJ
NUmi5WC8q5Su9qTTIDmghEdbJqgrud6dcR0Tda5fxS1YMkONhEOcf4liF/VJoRjNyWRxwtdMoPBT
sVdlVh14PdyZAagykvNc3H4/YtB9NzRrwTj1UQPZb0GsDchGFNo4v1u4g7HedDzdSVTGdoqqwSWX
ELp9abgwlEaz3n0mrj+hBQx0Wq255300yOuxdZlHJKQTOpmu34jql8uYAzpTDTChzqTHCScrNuXG
QSnuAEWxKJOiTTcTpXD7HsIWaaAPyHiud/r6+Rvv1Kz677uVT4tlRJ8gbG+oUOMsPdjfPmedcCdh
lqz/vsYRrPLol4dNmBoVhJIU2yhOxrHM+W1/4ncIa13euJgjB5oLxgjC3IwXSbQiJKMBt9lFYAR8
0++pLtqPPqPOp1koMfxYwinnK9isIlPE6Grs7HM2105jypS90G7D5Isw/7I5S559W1h/1GNHcEC3
Bd1ClAae9DbG49BNTQAhxFQ3cAFjcEKJtLZMobYEcWG+mMvXjYZ8tv3IBVQD1wNwhXTdNRbVQhrH
+jcPdCPTiXlZsiku6ZyVE54GwX215VlaCR9BUb1+i4XuqLmCfgi+ktAjQ29dUtlKEHmbgjRaPNGp
O4RoCTQRLOWB2piNAARWPIsAB34lPeecfSpF8KYUC9DC9PcYSrP95vev50v6PHrA+srjMVw4TcvT
mLsKJeHImj+7spyg2uRUJhaytl5Zq3APv7q/qK5CXWOPV2NZPGD5cV5JhyczT3hXs1RzYXBsUOIw
764iCFQNtnI7nHvDrkgROEXziB/GafdWQv+eKhX1xKOemnHLvl19QzrIjMcaAxVbnar/NaYSNuwK
rYOH3nR1n8gTeCcTmWYomVc73YilSp1R14cSJRB5jFOs64Avhf4qw5L3O53w4wmw/2+L1eY/EhM5
OuBURV6tHiOwr0wXq8ojsE7Y8Jib7D1FQel2/hwi2wdxGwo36m11BobUuBW7A/+g4WNaND9TINSa
fvrbClr4wo0tvrOHHb1fOZnVbbeY3WAMDxm675PwD7u7wNfNPQSZqO45lZigfoGXK/kNI+U/Pq27
Q59Vbb+8AiSxnZl2m7AJa/4i72E9LePs0SVMOEYampmYXZrCZRcDifgWmJUBSKdHX6uh19bVpRot
yng4qRIsVNXz78Ft8x/PotAI8A49b110y4iSHfSzrCf7v3gyPyWZ15a0taoDRAnDCqCBWg4E+xqf
1s8IblvsLbtfAf0qncNRWfGQiKt0GNPIGlI3qCTREUDIQMHOt8lLGSeyN6ovxBlC/BEv3ZhXYGeR
nlZ63tPh2J4QykXGzxAjFe/KeiE1esKAP1JXAklpyfAglDdPZ15GbIfFHdK5gBamvBb2Ld/phxks
X3B/INpBwJbhmGRffub92DEIkBfDe9E7K1acH2LP7hvQUfNKXMs5epzombbehk127koVWAlBu2J+
7SBNtfs+DezVU+lEuKN4h2o999znR+qHk1bUwDaJJbr2OtyCnnZhSoDitvPtaECi/4x6OJGY2h0y
P3hVhW9YeoryictLMSHWagHbQlCo7yl8z+EXNIqTUMUK+xhvgKI/OQLqrdUckkRWYm6ROf7Mbnxy
nW9vGPQIo/mlJM/fJbKcaJvvtvegnEmqZfVVuD8GG+0Rz8WVZ+NkjUNaM6Nj3ofDFdt9drJUx3Z2
sdNBZO+dGYLeT2eQ9jTeMwjwU08QNFrJnZv37ag0bJSAaF3JHy4iQlW/WT1Qkjtd9oIgl5g2kykt
szCRs/Os10kqVbOfB5u3pCnhL93gTNMRjUZwpyBWE+T1DChrbDFrjJbHLs5Onr6FOZwF2lgh5TZ8
Cdwhq+khiV49d5FgDKC63hwdhRpXtC+VUnCz536zmIxD3lIPA+K/oJL+CvdawC/UfEMHf7IJDZjm
jVK8SdiFGT8lzO1F0/DnbBhHoJKnC9C055ewnUSo9wM5KG/cAiMJGWJoGp6fGyfLswkzd0pTthjF
YQl+V6Tran35ypKI/2NAxy3VwWYTwc3zUxUVHde/Sifz4qgAQ/uHyT6s4FYwMaH26XAoQlzjzQkI
5sGFwgcb77i9stMH5P+1FeZ5JoOFK4xkxqzaHGHMXhpCdF8U7DKrnLAZ8o9C9Bk0q9r9RjhzafCy
o7/1ivM7O6Aj6J55zlRwztA7cEApasc53rBUtTSq2YkgxqBXMmDBA0I10uHqQSmOG/yzXn0j9GHR
zTZ+UuTJh0E+1qYD2kvHVishikD5JW7yzGb+o/lHXDKogYCHOUk0r84lQ+Bsuh5cPd+w5T4mBKnQ
BU8Rr5L5Zu3tzNTmTHPpjWhy3Pytlhj42WObYIQusa8qqyDPM3JC6OCeIi8ZwTSy0ibI6Nsxt0om
6TGVYwM2zFr/2SBBZ3jTC3KX1UAo+AuF1878nDrx2roS57fMZnQwjBSukvjBRBqQmHpBNCg5Tg1u
xEpwTLYqBLfU7cOF4OW1eFKp5wZpxwVmKBKfM5GLtNOy/2eVvvsczPtuFCsuY9WexwroEz5PQas3
DPgSqL74m2ae1WIqaiaVJcez/x5DSytaetfCZ8Efz47A10Kb29PMu8q+yb4Jpzpj5Sy1uqx7y8Rq
OULhwadUwcj7W9Wr8l1cwffV04Ajwg1jzAFwg15nFGzv3kYSDprEUkE9mFDKupJii+/yn7LaQ5S3
A3W7evZzSFBCJwoJy95WRweJP9xN4P+WDD1yXPM+02eJZ4mkryRESBzszI7V3+P2oyXzUrUjZ0eb
pGrg5sa7YFKOwuzvzR4eISYohi7ejHWOKA1gMBsGkvNUsSXYwV0dk1IiYWffpiyT9yKNvqzzbo/7
aJTPyN523rDRUTdZn6vbusEFGhR4h9vQp33D2ZtsXJmjIdNMAWu3Rr9/wT+X1ulIIxKid0V7vW2C
OvFvqA3Y75ld8yN8s2wMJGdkAF/jzArjG/T45uNTVwiSc5lUxdegBmOVSvEZY79UYJGMmkoGrssg
jGX41F6XKqqQrvqSFJHbDWodfE15Yz2aJjzo91b0aDy2pgzfN9bwdD6CjdBYG7gfiJLljYzjcT3H
ZdwlmE+kqGlARU32cLUZ9IXJCVcRAeK4w4dmySZCL3mW6Z402juqtEfFKEUm2QyLteHYCJraYlG4
DZ7CfzjgaR1xEDas1rM9pMkgNxobECtejDqRB/6bPEXAHjzSxv+yMMd93tp8F8IsiPkePpDAeVCR
bPnLxKRmeW3WhV2KNAlloQqUvYmkLfPPHyLRV7WMIQhi8qbgNLR9LzQiDJ/xTrzpXku1K/qRJ1Ie
RB2PNwWAFCN312r91iMrgEKz2zJMuGK3TYMewsVkPvEPbOIUJnzbxtqzPrjfYCtG+4/320uI5sNG
vGbF+vuO3umNZ6XUYZFi8WY0Ul7Ue9bqdVVDDBS0f2U/Uv1RAMeXdnHaVHAG5Awth4R1F/L0KZWn
iXk4NBz044yq7DrzHgVmjRs+UFq3NXtEH1FLsMVgw1PWU9odHVvbnS0FmOBrrNnqSp91Xt2dn3Nq
VYfvX2dYGdYVHczWiVxBekX0Oh7IdGVr0o+fhfKKLrP7gwLP3wr1xbLVW0Wk1yqOyzcFdU5PWGlK
Ym6E8zuMrboK/PKjfArRPvQJbUUl8H9vMDtpnbJThpUW8Ms9i1+mSgrqF8qYmYUSehuDSxzJUWDw
Rd8ST/2MOYskY+750ABq4PuE5Y2+Rk9GstPT22Dwl6TdEEL4gnsMcGRHYRlShDnsM/zgGJVRtaJJ
AJu2L2LyR0T40NP9HB8G/vkUq79W2OToI8SNregPYuz+Q8MPNlUM3AOjSpgXOoGBtmhfGsFFsaxq
tybtDoabz814RsRCjwAOj5jhvA8/z886T6S746Thbn/tM1EOMpEyz3dYaWmlKnvtSm71qs7o283d
LBKRs1mRyTYPI3mAVB8itI2Hh8vtf3NNDG6x+OV5vJTivabPUd1sS6ROgFgQGDfA7XraqpNB69BU
YWolkI1H1o4KmN82mvdGHJsg7kyag3XPOG3laruXGWay82Vz+fTx3jo7zEYzkcevWgVuBrdVIMuE
ant0f10GQIVYMUb4VZJEMbdIEPakoGQrhU+P1RT20G3bx8FGEy2T1/Tvx8vu+GTD4ElnNDnq1Hka
7q5J+Iz0vHSTVh/nv1QwjIgc8E+WQGc+q3lR2x9cxueM+gyn/D9xwCFIP9k0fjY0/Hsl6xJueJtE
Q+uW8CvbTLzXHiTushKIBUW6HnAsdsR4teZ8hUKDopGEAAsCLlKVizBUMvKQ/8YUp1IjMulC4H3T
FKu7uBbZY8X+83Ur+SwQuKCqAzeC399A+GWJBsSuggLmoVYermc7DoWhSUlUQIhoUc9qKHGWYO9m
8CGvAushHDqTIRssbdyZ4M724RX6wiIVn1s6mWCuRR/iC+Wff+V+/3QcF6w82ef5M/lAPMrwLlMc
cmj5pRHF85TRTbWf898ephg+A8g6WMuhimiNxhxYeb3fWaZI3+6GC6MR07SGBSKDZNW4BdIa6Ijv
v+SZXiNQ1xnY7T3nfIKUNpes2wJKciFYAg1FNR8qvhYbhxwOSpgLfy/iVBofdj+YqG//QaNljQ0M
79tmnXL0N0KYUMLb3hRxsYHWbkBZwoobPJT9+IeBc/4SmJk+JsVFmUEJEcRKRWmksBw2Je+LOFXi
8CNtLvoZQ6Rxhs2ec6DYWc9ylHuguPzziE+coOpDORffpCUVdYH+RNzScltvp1YOsUrNhoESdXlU
TepCSiq+wdnChihXllaMx7PjdwdKVxM8/WNoJPZPBO2NPSt4SQAZPQCxHTcftN3TFjwwBWOQEW7p
h3U5/6shuuZ7e6oEudKkbOrMpKwJEszQGz3ZhbJC2Tn3XeL/MtBz9FdkfKv8LwwtsAhCn3hKcXgz
ijVQ0p5eYr6op2QpErCOgOaYk88aAJpLdzQhpQ5xzpL//+2GGOJeXRHE1mxeTE8rd6VI3Zc2XgM0
PO/F66ORsumcxW5fSyFl9oiYAt8GT9Svhlu8LhUnWC/kZKEftm1/P5jm3J5RK9LTSREgmMrbD0OV
a4tTpgE0GzzRZUfq5xsJEUHIypxOXB7vK1a3GblmECBWSr3mqX4IdirE4sWZQc/+QTzRHwaorZGH
7H6rtG3Oe1zactzsyFDA9AyuMaUAZUme/840WuTrWFluxFxHbn5Rxyv7uzTd0RHvwZ3vjdwO3613
4aOWKk9CEcMaeg7EnNcdhvAUkYokrkEGGA4HqV+Om0d7xn9JIKNxHoY1djFxR0V0Q0aj+VaoDa18
wYMxndndIlohTw0dosz1EIXCGjC8BB2OA5dPnVmzhsr6K8A9F4sppJgbbCJby9MmIGrtts9aewN4
sMERq21GD9pjxfAElbDFMqdBSetlPRq7k1vjqH+KWoa08gBf42ZQOm0mMKHVYoxn13jq1KIAeCiL
XkdhJEdgbUP/7yGk8opYZ3lgItrNLvSrjrfEVp+pLumuoAyk2ECf07ngn8LvCeCJvfLeHYwCWBsK
PDuL+5UYRe0RD6O5gagtwAvjXfvvVJ5Cq67utrEi3oDwAfEGY8m0xzcTTyNuWGOzi2fEsBDkJ2u8
e0A/i9DyzZxyeQfEbRw2ZYHTQsdHWV2wG2Wfso0dClSRBOjOJJMyxSBryqAVpehD2G5HW91mJ4Vz
Bkqe6LsiH4ypBpT+jGv6MSgOqfGCJYxefwKtPnxu4vydjxQT+VPLCoBh3sPr42GphlupjGL1Swye
zmWzvjdvAxwfV1CN97CaT5ovd7KggTmwlwFOiM/LwXvcUT+byE4x4exxH6oFxD7RflJJ7uCIzzEQ
EHA+Cu7GCD91E1yAYujk2XNS9OoISmhvzOdefUdGTQo8yQ6MvgidUGVVqJWy+Kq0TlrT+YZ23MH+
Ey5+UU5B1YhyyfXVp7z/aQFZYZn539vh5Psn/AvwXTiaLS4D/C2o0xthsBjVYSrHZ4QuRWtIPz3A
dqHhPCzU/qoGkcCtgZfVRu7cXvlgPPtP8FXjP+dMJ+GQa8X4dP2TW3dPUi9ZM1l1cbn0mabvZSN8
/4eGKCqJVYuXeL0NejHQF5kCYsXyxJO0rKQbbnA6+kI93vO4J47PbD+bOmTQVym922wcc7DbIjo+
4xhA67J1AwFlX8PzIeG/4YxjPIiHbYSVLF5khMzGuT+jRVqo2ukZH6RSWJLsEuzrbvr/iQcsMQz8
N3TkeVsYs+vP+bSX8Ka+Ru0Zjn+YqJMgYLltf9zy5NCOuPObEH+aadOrvmVPdAqOKUtIap7voCIE
A8yicIqQU+auXpZY5xN7bQz3/DW1fvgDwSG+VBT0lRkCaRc3mrmmrg63tgapD1yWWOtitIkwgzJl
rqM7sxZ+CoHVOqk18lYgOtH94MuiEJXjrd6d0303ATXf4rwCIH7mqKZt04r8XmV224Na36VZWdQq
fgJ3U4H7NJoIvxTizIoW4ZjfELAxYFaR2hMrieRk37cFymPGf/dVYIK70W8wxy+n56Xq1ldzx0ky
jrX/1OsWASISofeiWVinpkePI5uwRxngxVfOmhHd7NcTGqLt1j2Q2jGoiMuMD2oqwfZhT+bgwvQt
ZN7QOrJRGawRV1hVRLhvY2ewLSGmjpQgh+WeXrMavwHQDBPGZrepwTBJ5oJFs5qzRk+6iJz3g6qi
yGZEiUSyKRG8TFP5mdDkNMq/172iNwtWcOQC0VUOtzO1vDrhayRN6gr4Q7CP9tfi2W+AY1/aYwfi
HBp15/1t8FDrPhwdGmU6ycYxIGsJZhhN07XaoMc+5iCfQZPSfw0akWghroL4bEHDZWpMf5mw9O2H
X0EnTm5+Stj/64fcv0FvK0VpBvFxuvyWFn29UEwfQPYMOFlO0GoZ3LN3m4l2GmhtgMHtXfM4v/Zv
Z2eyEHU7rk4x3uNixG3eS0Wxq1x7CQtjBMqjLHIKYOkee/4IsyUmzD5LSZBH/BXJfKgBt78J5IUk
idDVlqlauiXOUI/tH95uPU4LIjSePnGmZJUBTLWSwpiqVqp3flCvj9tSYeDKx8LceMQNTbd0A1Qd
STKa5p9OKfMTaZp3Np2dz1qvR3r6Pd+ygRfgrddZ/hHBsuJMDnaIxhJoQIz6LctuuyJuaylk9ZJh
jOcTcV7Gx2PuB+SmgY7arldOgwbbwaM4PBlqjgRPgVl+Ca/bDAOEgz6R9jT+ix3IUjSfoZ/pJEu+
hi8iyrYJQs81Tw58heCi95XIoWABPM0s92bPbfkeg7bZkrXO7VfVMX7U+J/ZV4fbYLmniJ+zrHzo
0oOUyzphUKr6lOIf0jvW70IwRkSA7kpEQKBGMjlWYIBB89ZLwi2g/e1CUgJgYnElpqxPJ9rhO76h
Y6q1Sj8fwlI4guDDvJfL3F5qN1Od+688Isbq4zCMZfA+7iphPCXxBCO8wDZbDlb86FQaYDT5dW3X
LuSTKtEwCOSG32SpELc/nOuw3PUn96CyY14BECYszFL1RGIVOi2FYFis6dOSFxhPZyY7Wcy0v+hM
mTIcJbd0+db6EIsAWzllmQIoKHKTIT6bzD9TDRYICRGrLrkbIGagI7RCVwV+0SwZib9/wEcG1HKb
OQvzGMLUPvRBXE3BRZx31Scr9gREzmVdOkj3ITWARpZXnCpHbaM7HlGTJP8pdmj+72EAvAL6v+4q
pACOQZ9zxQWKLujlpFPWySAjOVLkbwUOTfXvpi7uDVCLE43IqyNwP8fCbUxE59fO3Be46Lo3Sepj
UhOtcI4uLrnjAiT/SX1vmfo0lVUZ2b8v1Q6I0XOwiDa8GZwHTW6ggSeHkl5XhgSt2Qu4tHjY4UiG
gVfqoDBV6fKt/bQA6aw8Jyf530kqmYCMT33+W+4Dtm9KUlQCt/mpc2FyvQmhhtwXHHiVH6ZGEN1s
CWOVCG2dIel64LIXDqRB64xZ6yYOrdh9S0b38wPLq5votFI7H/qYyFGh+PyM0eIS+S67NWj6RTxN
DZr10mXlgq+mHtIME9JAzSt1ISZcbddJX28rklzdLlAyJeqz0ynE8OdnoiG55f4OGuuVwLFKNwfN
AdUzmK3oh6qLJmoR6KT0a7A/i3qfgXW16lphH2w3sjxPYiIAIp85lHSETHXVxkeloPPK6HL68TTF
MAmr7xU5E2REUdYS5uBUacdagO2LzA7omvgh7rsDw4aYqLp9zwNio/+FQomCbW3uoxmoKAAQVOe3
OHWDr221PD/bqKe+opXvtpB50E54ze+NU5hcEGS2KF/OLi90zWqOtYjw9kM2cdPSjFZ/LWVG2r6z
Dm5WrS/pKa/kqjtH2gk0UzI1YQUbFNhV8KY/pYCX6t5Szb11pKWReduiO3879JqZEJW14YICe+ft
Z8znQOj4Cog4BV1QuzKiqt7tGLd+poyw0yHck0kf8Zd2FxxGYp3L/5cpnK8Ue5274e9W6vIVmhiV
o2gO/m8p3yqtiVC0Tm43fLxD2//FqfsXoBCAhdQKcBXIuTtNSLdhHOnoZ20GeF5HZZIKbrTY9FmF
dULLp0GWtyD2/pfWcEmffgsR0pdgxMfvu1h+7Cb2m6M1sEiK/QFbFoHccMu6rNMhh+45cBDhmJPK
IJrEM4L4F3WssI1gGkOw2cB77vgSJdHJfDSa0T5Jpm98X9w9FXEmwM6MDdDhPL7s2kcjVHBkvz15
uR22PSRE3//fSC3B80Di1oA+48cYRwCfYeBoe/ATYuSSVgEkEWuO1GoIDApdt7PvZaNWdKh13WLC
DhzHdbL+05hnU492BwqEn93bG13Wo8pwROy5NHYiz0twYJ+ZSa9NEGqcd60fyfkiMrUCayCB9pVf
DbZRh9plt45avIsFDJIYLFebWFFPpC1JnHqyIq3oeL4jzThN2p7N5Gk+p4jueORFUOhsOFk1ITqt
f8p6epf7vLLB0mfKrDimOSvZY8XkUBSlmFZ1hfurugCmfjLWWh8K7/vknXRgu6x9007LufeEOMS4
m2fJuaLV1QMbabTKqIKJmK6K4AvnsLdXAChFH7GKJi2gX4O0WTDDu4nYMXaMbpCFY8RFf/pKy7cd
Cdd/5iwk98QimimNfskFPbIG55CBl9GCFkbxhEBqRr3+bP8jR1A6hr/+VXXNrnCG9cDxXmn/38/0
vNoPK6rNTSvFtxxSChvchaWzUY+mlfByFibg9IMbpvn1h3Kpulx6d6wzi1SrGq/+qCZ4UX1x6n6H
TRWuGab9tRl5IesULkaremvS3bt1mCOpz2rCrxmwTCxr4fCQprB2mPuOUXwHZ2ldUTRv8gLbEHN/
SrGnp8hWc87E9uOndq8okRMkDm6Mqw4ZceCBDNHuw+9keXD2aDSpQOFQ09k9mDk+E4G8CGwam27X
2iTYz26qevia3uwNYKd1VpPc74rdTPnoCmzR8985+hs9ztX5E8CwIOsVP3yZlX6bKf+fSUB/xCAI
IWdLbSREvPfIYbIHlQ644oavVXA0uO/Zi+GimLeoDOutla9iYQn1rga/a+5DIAK7+quyf2umum2R
T/G8kkDLk37j1slfubGkQA4NciaSYPtmDdG6Cbt9gierbdgbUBCS3sNkYF3U1RP5aP3fwkux2X59
biLStuJmnWgj1O2U35W+xVCEmEbwrM0pL7wa40o7v92sTwIyk8Zb+vPHt+7+ezsrqChNR/bF0i3Z
ix3/dbzN2juuSIm1Gvs/IUbOp5jcI7SYtPemQDU4VDS0lxgRGceyHbgPgdwiJ+9npBhfpGHbu6dj
vovqhVhQyaK8ld0oK979URZ+4j2ycp3xfHpMMI8zMKJJyYWa3oYYTACDoNv1MkLHdGWVk30IqYnd
xNVxUZIRIPXsvGC+7Fg+Rn9/c2djiWC4fYKSQpfPWdr6dGGYTQ71CeUi6tGVGOLvOv2TEqTyKlJX
GGugvB+9TZYOOkyrBXiSZLdQm+Di/jB8FQWE8gOvyIPPG8FHNQkYRe6saIr7BdFqtFLkOyMM11Jc
J+Io1WWVE3orpPUXFOAZ5SZpDBjbahanPOolff/PBue5ESFY6LJuS4eaWJ3GPzusyjh+SIPwJgxw
ISvLtesKxl5cShI7nTTDxdsogOUFAXIWXHWHwFYtj8rJid2vatc+PDZTHMLHhfGntiZ48JwOsKGR
Ofpd1WgqEy7bzbUH3ayGXKwesHFsxXKQx4sUPly8mRNKDftEurWLfsVcFMTnoV5Paru3ZqwY9JyH
ytbe/1hxgheVwzfT5R/ci5wbafhceKUl1VYNSM3cSXAmiNaAyEhebwN70+PE0ssIUEnpDYBHAPaU
xL91o4hDpFcIr/p2udt1LeTzyAJ49pu8WO08i50KN3SSA/YPGc5subqtQISrtRe3fjkKB8FzI+L/
d2d+a9/BZhwAYBo8G2hdxTINU/Obz+Bg3ednEdy7M7zC8FWAjT/Ar+I7BEtF1fpY/YuDaPdcKJIn
7BVw3cB4ptquUfszLvPmEw3kq1yQdvlvDN7gD4Gs8pPPXz9apHVWJUu/m+D6+rAL4Pve5vGmltCd
B1x0ebSta37seJ7nAIiCUrwwt/ZsEVD3XnPYvqiHv2jmkJ5wcee/oX4n1kdf7/jk7Eut/withgap
17hvKaLXoPM3q4kQZ+89KYXBKAvsg5gy0J0LbbFKQKBm2gbBplA17s27Uh+6tvBMA3i5bDty1hzz
yk4ICHVegcHTTLh5pKf0RQKorjRm+svwRw/zgpGVvKyS7faUgWjuW4acmoV64pKsFEMXsuwiDffT
ZLmYx+cZRCI8BGPHucl+PM4OLP6OVeJznHU7nPlz4nPNEy0jL3De/sNGP6ZwD9IQxymUrz4z34fj
UxReLxB+pQ8J8BjuDY7sNflb2TbfucJuaWDLbZY+tiKWoRb+wpAf/8XB6bVOz1esH5Bu+zbwka9m
tOOY+0Bf8Li7sYDDXhW4x97HCi3wpnLExjKQQh99Cg6yl6CJi05cP656+E0SnsN3wPsd30E2bziA
C6INXYIzxFEjL8ute7krSHYOKc6o6k+w6PaqVQuOEQR/w+pe83uuIIq/wPGkfJzoab2+mvWkaJkn
xrSW6FKBEjU/FA7MTqW9Y98wssNqPiAO6znNT/HRkhbXNpf8YQxAUA00ya0iUZPVagxwJgMaAMgU
ensU9XvMpVvofjZ0/eQBC35sMjZiaKIG/zTk+edOymJ52EQgg+DK5nDy5+YjDFRQt5voXM3Pt6c4
DHw0m4JagYjwcfYK4jVByFIfk0pUVrt4YKHcy3wDEMJQqzLKoA5NRiT2HZovhefZzas4eNkNVa6T
n2NgUTntRTxCwvcX5GIh7sUTNYcFOoz8jl7UojWeqhcUz99BuNLjpROQHhBTrqkeSb3o1fAtL8wk
d9yvrIU9kFaG9h94lu7t7z3h0d0BElnUUAt76fznybfTrvzgAEJYdryFPTWxjhZVKOXHhcncFb36
jLb508FJxlqub8yAp5CrxHlIfLgiw1TGL8hjuZG8l4XKU7ecj5kKEFQ8rvk+zW0JyZrq+ZIiO8jP
U2GCPwAaX2DIpFQ5lTbrTXL2jIBYXOBv3VJ24z/sIN46JJFMemfYgP6CF84Iy/7nHHsa6MDiNTUE
fPgQmtcGA9yUsdiV92RWP3C5sRQ3iiIYA8xNwm4qnNUAqfj9I6mVVaRMJVGmqCUMcWKWV0RMA1Fc
2eRXMt9ZNIPSiFrE51Za1AWfz8ElevTAsxC1n9PPU23LpFRcLnXy5bMGTMdzDT0GizUFUCPl3CC9
tdj30lcA9UGHl6Iynf21Li9d6ZddPtpAEkxj31L/cBMeUqWxdzIM5pt/l59QavVmpIsIRQTC+KOA
+lZ/CxHAD0Q6waiHS27OlSPp/MPKODl6SioRKgoQBN0ysUei8hzZe2hI4A9Si78SSRvvQOSUMgsa
EBE9bR1rNgvvXotphIUTLiglnOS2MSFIkWyV+VzetAo4+wOUUF5qOe92AR60o4Nd2P+wu87w56i6
JAbTDrX8+UBQVeERRJiSoI/qMd3i+EyZ6KcCx0gPG36KBYL1F/szCO7PjiQRFCwhAuRozt1Ia3FC
kTmjV0B3p8a7ydy/fVcXYaUh7QHKMN4+UsbB6H3rmQvmjmoYufXUbW/hQFZmVtBpuo779SiWVkLR
DaYK1lIHVyFyCq/dr9H6fBgl+P8eMPHrVzzDVIB86HJELFWNOb9ZKBNEZynaoxE/EJtQb00b+OzK
jeSLvYmI3WEk8ZSJ7MUXsnbqQ0SzkQu50GHpynICUbVqzMNxuBOJGlWIKC+NgSvjw0MtKKfpiUuQ
hZXgIM9FqceHs3u0xIXzpvSQlJE2AphX+nh9dyRP3wbao5b+INw+iw0GMbKK5ECCrspbAQnB/aq9
W5k/oUeFKE9XdenYgqTplfL3CbgmjNEJqr4ehtbnJ4YV3gfNdF7lgDO3nn0n9PS+/g4U1GuGbDRJ
mRF9ux8RXEKNt7uGDyDVeA5qHseP2xVTfPUtyoh446J4CS6E3r6esag/bf/UREQO7ck+sil/E1Ix
OOCucxMmAfDtFakxtsILEnI9VLt7fkOCXZYgRD4tR+3LgiPUH0GARpdPTxeBM1815dSBMwW/aX5M
6cz/LHTz2rUrKdDCbGvLDKT0Ww6r6Fwvwn4MIPn93X4xDJUT2Y171e9t6wkzYH5MQLahNjLWa8QQ
SK0SWiFscLOocS814SLcWU8Ib6V5wymP1wj4uHX0qwvxkv1lE7XlY6vRCAoV2bSk1g52GxlUmqRv
vkm9Uj8G8XjWtKaWz2jil9Y6p/dSwOkX0x8zGa6cprLaDKmt7Wji105UKV647KNkR5kesdyPjzkb
H7EQ+XzSEXlzBlZFzHNUWSROKd4dLHnn3VidQbq5zIy0zfIcA0zPqV9U8ZclIWVRPnhNFC/CsyG2
40x6MU/iR86qJmJjXwsGlmJ8p6K+32/HpbarBLRsXelPlDTJk8hl72b+fk3Tszkvg+iRwMOiUG32
A8tfWSGEu2V+LGxK6ZO0jzEMxeOE8bpPxgvDCZEZALGsJyU0W0q0mo3ikk6zsVCLMMkw/aXRKIcN
ExZ7SJc8ZBhNMgqEESLSZ2dSdVE/XXQ8WHCXhyYDlwuyKmnF4oAwDlTGskAHgj1Uj5q8RgHeOTfP
owhFGIx1P2o9ZxXEKCOeqyynMtIK+7je+SUd10UOSwG+r9of0NNHqhq9DRCs08DaVpEC4v2Yrzbk
qCVEWzJCuCRBgHVzPYskTWBz5y4SYGtdD7mY8BbLO7kuCw+/Z1jr3PdeGGWU/tZku2nuF4cqFpRH
eiJKGjPQALYq/F6ACE+8s/cEe+O79fiJazliH3ES9yB0crnvdxzpGcJq3fNSJ7UVZegps5fl9OFP
q93mj64c3rFeIeJRWCMJ2t65txjnqEE8bQWuHaNcELJXUQJwA3N5stuosDox2lWiw2K9qYT+DOLR
nj1qqCFAL/aw8HxW9CZw2Ldv5MDWS9WHIFwd2xiQgzeeBQUZGXA8dq53FSibDtV5wbf5T79pAkCD
z+HhWHBdRHWcsksYTbWs0KX+VS97M2X8RjoiqJmxlMc4zJNta99j8ulnmquLou/0mZFbFq/2h4GL
SiZzUJIN6NoHv0wezjGqtkW+wfo9NnqbnnAEdZKea0bYIbwWBUk/k44U8+MCRrCOL7ODGZiwD+Xm
arOJZ7WzA7toVNn9ZeuMDKBR1kyy3/jedNYqyBMfyIrMVESo+wV9KWVEYkCoDqy3iwYmpbTr1UoG
Jeftp5Ilp022rDAG40eOMrg0mZFcbGKzkeBQHEkzaraYRYDAmk2Ot07u9xHGBUnmHALLV2ACGvy1
S3AYaeKUfDNw6dmt2nYm4PBQJxDcrE/FIEcpVsHSqozI5+W+scK8z6JiTX7HumXny3lWvIroSJpL
TQ78N4JEC8SFRB/V9kMAoSuf9vwJqv1vdSZ19pferPTpsgirYi26WgaDON9D1J9uw/xeuMUR1Guu
uYFNkIYFDWt1tEVZWzbI0AwoG7QRazbDGLBkHt7zo+2AR5Xh9c3NCjZizuDd3HVBYwAL1bSwxpHk
NAhKOzlixOU0GUYp40zUBP8utujCxyvMs4yRBfU9m18PoZb8JBqXe8pE/BI1DBXzroc5bvNSqR64
e8XJO7u5GuJ+BqJ0iiZcRQqFev7EojMBQSJwburFNRxFf18kh5Mxo7F+uoQPvkMOjdRr/ETDrnlf
1CLWUEN5oAC+h+Z6jxH6ynnF9xat9zz21X4+suBkDcmcNsnq6vHqII/Hgcj6Hn+vM66z7FeXINdZ
b2aE+gclel8z5WB/uAsjvh+qjDwEENEBjabeyeMMOL/qeUSiuU9XI7D0NqvF5W+YyA4Hpi27WMeH
szlXWVzPPeD2zQ5EK2rGkPfLvueiZoZxpj3sU1Pv/GhKhHlG9lDxZk7fgt5RQwX2MAxfbT05Pi/g
BapmRqFgK15qHi5wcyrnz/VL1HNsSZ7RmKHY3j6yPHysZ/LBAscO7wTTiMqCXHNXy+F3WLvB+lMd
Ot4erci03oTFQdBK9/2smfEQBoE8+66Tk2s+4mtKzEIRPFWK+SxcXBRDKCGnyStYPiw/HU9nNZ16
RvLC0vhbxqJFBof6POIiTWSky8sVTK2cLU641lOGuZY3T4Zjodzf0+yBPdp46Kcabd8seOIq4ONI
/JMi6YMhR4ZFH+omsVbnG5+Uhs1MYS4QSGr1Gprcqb5eUSNfYb0bKuwfhvq/hn/Xvr9yhU3ZyLgk
m5LntdCNRTL+pNuOLyB8fYmqm+po0L3iwz0wmU4EmcVwIJZKhtgnF4Piyt1FvzqSYZCUNevhaYg2
+Cn0jgtm69Q6i689trX4+akIzVdpqlpAP7hU5zFKfz/QYPqVCWLOxgSlD37uOnx8ExMw6J5RL+f7
2wSilBvKm0iJUHJAjFTGguAQb/ij+hN+FBtoeD9msnfEKR1joICH3QNzxSA8MBZG334X9Ym1t4fD
ildkAxn2OwzDARUzSzoM20N7G4XafGVfBKU3FblNIQzwTiIgjg7raFTtAaHBFPvCcHvno+n5uJay
LOEXap+C5SaobvpyKNc8z19RE/uLpGoiXSmjfiYAOtcgxLcfr1uKjjA8UR3UOnbcloLeX3GNWJZB
OQcfL03UVHRg3CBOFDSqvnTwKfh4RIh8ka9d1x1k6M/BGAurT2lzk8E3Z2IZkcY0hVysZiPoLRl5
GcFR+WJSLr2UNb0xpe2AMEgsHp6HfBvESOU1oXHbrH3DVP6tmJYTV3EqZF5+swGMWlHDCGbcSlui
0nZny1ZR5qyknQWFlna1V79I4+olitz2NSmrIz/4NJpYav0nASjjOVfozHdO7UqE096RBtD6DgbL
aDNhquOeDCndIokMIphgR398Bor98Knwi0abHYdUsK0t3BzfkhXnzKQH0cx0dNGWJG2TiF718L8x
fotcT0/3YQ8Qzq5EsIGLKXu8xgSzSayo6fJ/kg+d+sHC6EaczKUEOUSko1cAIYWiT5RysCqEx/u6
Ktgq8FEuW0CV5MMROlmrwu4V+ThPmhy98IGxPVSgDJgpey+yVXl0cgw1R6bheyAJFQKDskxIwZLd
+BG9ypY20bgi0HU2mnQvgAeMjx5WsyT39xf/WT02nVyCKmlX6aDh9WFsjEdekkunbxpvGAroDiuo
QcXyktG5pEL6DbQ9m2/pG0qEVyYAtNA+N1mkZrq30C+Ycx8/s2YNAaWdjM9rhmUbu0NU9lc83gw/
K/cMHJ5Uv0kQW/UNiykxJZYC1ait/bFdqqFnuciVC8Xk2lGH/sGMyh/ROEhaQ8mTu3xdazVV2ov9
P3vAPh88+ALF2H21UaWPHz+ZrShrxcowQ+Y2aXiQIKSRTe0O8AdGKx9yIPuj7gW6dDh9trSiEsPK
Aw3bBhy3SQgyamrLmdM7XIWeULXG3D779dcbckObRz/nGJEKJmr5uqB22KrvFYeFhsJdq93vHR3x
VotAKkH2mizqqtBHmlAzHzvvAUT2Y2qu2S5hDVrjq9cXSbYMOcRWOIOiv44JnZWRruORBhSSoQcQ
Hbvoc+sOJyT7TOqgNrPr8AaX9KNCTpOIoeAZXYFVaVxzlevohnWyKegi3v0m7jWcytYFwD56unCo
a6EOw5o5aPKD15MnxZgTSSU4Gf6yVmPEpNmSMTpu5oieXLaEXOgsJy3SgFARSBEV61oMtoj0grKZ
OCj5nxS4ZS29jc9zgJooACeWhep0fo6GCfDj1BPqrC3quup8iRRTSoiNIaPimuarE5/A4lee8Eeu
OmTXXFWMKi9ImPBSI0aSSqcJjtFJYR42Bq02WaoT3vXDlmbAPy1xB15JngJHtnvPJteTy86tLwbC
K92UH80p03/yfaQ8gecEKLh4R7pyE7mHD27Z0mmbaqJ3Eb9XGJ+uuDooNKZ47y/b/Q8szcs9M2ky
eniiKZ6G8U/ywhcuAcznDtg/eFwqBIqg1mVrV0m4nN5UULUtteh4zdqroJJqSGPDqf7OT/U3krPj
YnT4l9/73yEkgUi/OOE+WGHWySQSONLpFGRjPVd0I4rz27rDXMufFTDcfzE8G9YmQglXcl8IpaID
4xjBCKb1tEf6zgbCax/lSFy0jKqJ1gTkY1POnxAYP9zSfjHRrylhiVFLanCG7SnhrkIlApH1YvAZ
ZFaF4Zbw2OzH3fNBIFlqFX0Jfgs90d6HWnG6x+l+EnjYQwnAQtTycOZbv0uGG06Od4k5n6gDJwhM
DNt1Uf+XDBKsvFQUc9kHrRofsOqs1lkG/35XXT3oPVjyquHq8jsHJNCg4KlorE7bJt65lZXOO69t
hn1EjiR0js6cEJDGZ07GgpWzrbISu4M+KT0Tiyl37NoU3cVUVxZshrn4xTg6VCh0OLFlwdG7oQ0X
dnD2ZepV4zJmGGEqHf1m4Y2tGPBs8KCpNe2MNECMGvYdLqOCanWS18PIEQp/JhWKXEJ3AnaY++lp
ErnxnDSraIqdNICqzOuDxuQpoUL4KcUE2le/X0L3K4oaiMEHmC3t+NnqoCTB/Eh0PPV+S//wig9/
W37Za6/CNcNzgsR1jxeE8XlDxXOAWSHYrRZ+YlBHFyyaOFH5XkG84H8fDaYAnELdewAOcb7UkSj8
mGYHJg0crWDKhRt37wwY41rFEbTiibpyKVvnE9qc5b6fhUlou1VN5c3i3gyc3OwzlRXTzAZ1//Jo
gDp/MIFDRK+tzxoZoK59KPOBibUXUd7ktQXl+VYqD73GIM9Cqk/jQPr2RuccSgkZVcVBXrscYxQa
pbvE2uin9e54e840j7Lmx8KEp3x35MPl5Gygj8Ncl3OrS6QIq94Xfct53dGAAKI4+qJiOq8R710b
UiZvLxQw/JZr+ntfUFoNal9FVueDFZQ861IzLPGyvcvMfpcf4liOzSjW95DcYZk75aX2LRa/XlJQ
q7AZBgwJ9gAa+oGjspw2OXTVHo8uaCw9dPmiE0HDla0YdYW4RNGUykaz3Ti69E14YUhDrLBJ8zNG
IDGIw2cnm2/1fqRdLeVUT6zcKCtn0FB8qhu722sUCfZURNwQnffWdFfAquBIM6pnjQXYuVMIvkMI
Q1IZg0ym5N1XB7PvthQj3a8tFnTqhbGaPDNTCSTVJBngQNVW4nUkgG/EjCt27WllMI5wl7RjVWde
64FlYKqW2nqewXffHknwH8+mrPjpLboXBMFibBcOsHmyyyak83V6RA/Pf8AyK769/cEZwKpoba++
a7+d8RhyGFgrmu5WJW93fdD9u2GY0Al17KLJsdzHTF5SF/b41IKHDuaBJsl4PRaPvKmJ33n05Gfr
/YlsjhDsDi2hk4q9jhK5kgMf6ZBkxpTm8LlCru+6xWobe1vrEYyIn0kftv+8iRRFwuW/4etQEvJd
xnWlyToMTVjjsYI7XOZwE5twX/yIXhJijbpFkQXPlYVSEKZbnTEg+Api0FDfSTA8z76U5UEkqb+Q
Sva60qM7QYjMgskYMxpCY2jnB3q3UbxW3vRQSwJuXIVJ96sgMiWiliJCTvXl9xF4YM+tMvBCCofp
8dvqyCPMdpZQUBh2UuY2TEENz+PI4d0HPGda/W1Vd5u4RcoJQOgVQ1HTbXUCYGwMGQp4ddnC//AM
sZ5m4HNDOSEZ0k2VH1LDlbQUNxVwGPcQ1xjhxwktztyYoSOeRafNY1Gry0u/TtSWwWVOEa0aPc76
CovfjJb72IcTw10FtePPouAyAYBRrKDGMCsCHYq1K+SCs2VEZYbMVsddjImum3djbdslYrR8n4vm
GtPFQ4QjNNEf4kZIV/2clmYhmgbrwyy0rI5cB22da3Zc0gfR4/89vvsqraGXdkmSAKC9yZsW7i3c
m89BU3SwQkZ7atcR0AezNTisxYhtcwaCFwkWoZzLEIcOSVXxcPSH5eD5eKwV/8bMDCrMp5W+X1SN
+ssp/AYVmyNRsavMmm7UWAYxq2H9Z2shjcgzc6bSfctLza/qLSlzgYeMrrb4Q40O/f81uLG+FF7w
g2Hw40EFoEayZDmUK2PKWSYZpQ+fIbTuzKYWk9ooSEUROQuSG2WCpMFBkT1K+QLuHgFy0NZmKrt6
v5tX/1aPcJUAkiwwSzizPl4cuedtOtcHzCHbRzPsoxceYd+CdjgX4RuIZ9PsNo0AcYO4pTsHoGm1
+96gDKCmES7qpiZWQlcA3irhyEYp+XjKjUlRkNB0ChxM+ui/rT4ZOAeE7voUl0VTxVaGWDLWLPHe
O2Wb9gaag/M51xIKcpqgm87lxYHjvTMWYBjEyF7OCw1IsLaipSxtTJl0OAQf9LMQbkCdxN1QA4iG
FnJUnhNZPhBY5wBXnxA11rxRih88WB1mPqYA6ZqCJUftle9QNOWMDZ6dEkxgj7BylM85g+tPGiTS
Y3qzzxicf9mPQxjzJgQ8ZMqPCdZdQP78shT0N1UcHdcROiXNQJTKxv9rkcesDY1EnOtaTiAr+MeX
f3fMJCjTBtiNOhJ3MbNAvMQ78K+dMIL2KxeZ9voKmzbgX2kAJdfkCtNKhyZwWhlWkY87939am+tQ
88Xybg1+gtxtdevfbq/ErJnJirLnmM4/iwtDjoEsXVrOAeojXzmIUIOqHp/DPcL5aiUs2Y1JWu4H
pKB/0TgqKiLOiCYa4FFIODe4hAJLMiAEPf1RZtJfJzItRyMYnYzNjaPo8VinWsOibm706E5O3S8W
NVnMdq57edGR2WFmG4hUe/x/bYEtIOfWrPrWJb8FwZEl9ltybladPWE+0WT9Jn2rj4PnHGbK39Rf
8bcrlUKC2GlCKR04DmEEkYlpvCMnxHZSSuQMqj6QjXXQSHAdVjfvlMVuiCLwM359R2SrXoKxoJaU
DDDXWcz1aJoMWuO614sLb8PXhtMX+jVgBGBEpgb7qXOzLnKPvCaSBaMCM3l3/keN0wAjv5PHVITt
VgLB/QeWtNcIHRM2OwA36uqVRgM252BQoJqq5cQPW7lr6kn/+sRpHggLgCjrUMU+ZCwnBH/Rr/Q+
wnkE2t/JDRQReNBN2mznozz+HskgXJiqDU3u5T+ptRGcXUp1QxIlAe5Btx9X/GxHTSfB52fB4E5n
Q1MahQ67tn5plBbwPw2VHpBGj3tXiLil328tnF6vz606vGW++Y3kT3cwOng6FFNfaqWHZBGo+veI
TtLLbceqFPkMuGBtJ7ADAhzbLd50ILzRnUcBb8GIiqhAMQ1lqZjYx5NEPOVGMz4G5oJsceaoODeM
OTC6hq5uae3uwk09nUEsABupehaDPr9dQzDtS+vwqh5ZMcrD33xL+QOdaSSDQxwrhghEzByhYRYJ
Re1wZiJi5ITWL+rIXc2inby08DFogEyaTihQjXCKcVl1N8PT3t+vsb+7562psx8peL9Sg25QjdL3
v7swy9/gbBk2ATKUJnfrQWI04KdWSmNeuqJ4HbcZ6v0aVv/cR+1f8xJLWEv5BPxToV0Mcju+sSsw
0tHg6PBNTqxsoe6tnESL31Z5VhcJa5GcU6ZQMMmKhHExx8qB0IdJLmxy8wOxvTs4TMPEG+IDzpoz
d9yrWphCLuaWVxRdy/4BC9byZisOWSahBOSOwkFCLr6rF5f6jNJTZkgSi+ol46wh2I9vi3/Y129V
q2Nl7BFd9DDKRMa1jkT36OFWTm5Uo83TfBRo3euIsPBAyt990WAIHPAU9KmiLR7INrq55lsP4MIf
KaF08Zk0LzbTucetmtHGBu20rvHEBizaFC/stM5wFBUrSzKmojOPqoKLGIpKJaO9yJIj0skv+lkK
HNbYvjOZ+LmYcuQR9jmr3hhtWyzb7Qh+UuDc3lL9YaIrQSg6ntz9K+Lu2Sr0Z3Nojd6ckDFirP3H
JAAIMQSDxzhHxSvxkwOR0nXlbGvf7jd92/jF9Qe24l1wvRAhttbNrcKVJo+VGDJg/dYbDWOTPote
3BaPC+1jSTwpSwz2fh3VKpt6Lj/ygLYNdgfXCas66BAIVKkTRA2ACusrVPZyT/4/EJshbgpf+Ys9
D2WJAdgFy/w+p01acJHhJOx1wP1FWJx60lRz88ZwGa3V5hRwSgkt33PVbGV+t6oOrc4AZjXxvEW1
Y2PwrSBS+XZDtGjX1Zq8A6wYbQxAMIDh07NhDc7bUmuWiatbDwm0IoJgXq6ribLVhE3h0tvW0jpH
0mq60IE/MyIy4TpBNOqbEKDZB/rDwZu5xnVorwggciXjhnjSn1uH4NNCVbHVb3Dp7/p4Cx342w+H
BCdA5bs8JBnuSSblhA44TdC3qRp7PMU6zIHchG962XxLAdY2xZ/UCteubbgOgkPfbDRUX6Q7BEUl
3Hq/CoX7jPgpTemhRKoVcZsN4sojJjr66MK7taQfl3awT8Q1kbW3V5hiXD78Jx9ywnVlreFYtp+a
nGVxhORyHSscfedm/RNN6tDrDOVDoSZmYqmVXB7mNorkC/TBIgsWnYH3dJBQ2awfDsGGzjvdaJ9a
EQ7sXIizkCP2w5yzahoGpM0pPt5NIYj2HM0S+94OMnH1sdhXFYAiq5zpxITrk8MYBWvLLbKdpiYO
jg2hYfyYNiXOHywVzurnYLVdJ0JVfGnRYI63O7yiW0mMkxS1GAdi+vo3UFycKPBtTZaucRFI8oze
G0fMOJ2qCXqHBlM6erQV2+41vhoFrX263gmkW3l+HoFJnJC7D545Q/ozPbVk2lzWUVDnrovuTLfw
feyWUcdlvwL80AJRB+n1AFhCVgmB62A/tQr13lOvXUtUeeb9pal9YL9HLceF4HI/57W049x7A74w
sZ1GfNStM/xdx0qZp/HhJDH6gtIPNyhMo0aKLrw05p1BeQq2pQ73tt3ZbNKO7ILcLi62W+c5FnPO
h7Xq2AoSY56IYGnWENelOxpF9bFLYFto5L+ZEL3mRuWGoreHdgZ3Ee1izSmNeUN5Pd6PzQY32sO5
F0zkPPQyz+EjvdxAiKWpcSK3up9wx9fP5RzFCyl0/zeoclL3nbQScqBBsMZGxz6kd5w+H5oM4MAk
l+UnRSSx3vy9Kn/k48g5F7FM9O5YrePNtNj84Hf9Rb4hhSpaGw2dh1Mj4NbLA8Sx5glFq1CPoxVa
KzyjB2HnYaHMzeyJPtggxYUINaq6E7mVP2AkE6PE16QzGSnNnMRh9cBmSzQIOOS5oF7Rs8ZyLCQx
BkPv2yxUvhwL/qNqYWd5+mpPBCKB2ZWyOUzmh52utP9vX5ic/vD2MVKOZnWBoJcX+PRMw3Z+sv6R
LTM+JTDLr07le6aoleekZ0Uw8AAxXMt5akZDWhMASDMhJh2jrIHIiqsA8tZMRTUlf+j2hMYEakS4
8RgBwlZ0BgBbGksBLDxmIEbQ9/0LgBA97FNvYlnKDGPSWaDNtwxIqLpp2SZOo7vAMG4sygEcVJyL
XuvwNtsbqLg+NTPSMAPIIlsErjUNZ6QGeOQCel2pwCSiQDbFS7RDajfWnCybQr/w35Y3h3P/r77S
aIDUR0rpNVahP1ZHc9/UtktFYNG/T3y0FBe1pqZ82GBwl9rc7F1pCpvcXOdtT9KtYo198vzyxi5V
BfPyGYfSkfv0lRKT8D+Z+Ul6OEXp5Otc0WWifl/cwkC9TpodHm7Lrr8X9ZhqSWSp13P3C82d7zqH
YGeHHzB/oEaQGSqHzAoQ4Y8nQPizN4BMcANp0iP6JGTrgzSCutqsnUDz+fYKyEJanvQE51d1fv5S
uxso1ybYmciDhxg10gqhMZElIGo0p8CJJdwotlt/rTbXR1acFQVrqa1KIj4f2MXMOgLe8iBFOY4e
ysyNxdPHTACCwgMFEzvNbgpNSFj1sHDxNKPjxkXqPradxueaC4fCHa9Fs961xmhKEVXuiKGbiH+4
Nk3hBHj/EQPrIlSQNLtIMK4yfH6kCc68r9tTuVYlp/N4wti7yVdOuL8nub0gwEL5ofqNwDE7nZ5c
x/vXhoiFH90HzDmbJYEQ4mUps9lJKDx43pcLiRLlA0gKkFJ2guiTRzzh5aOwSfcb1HX9T9lUC6Ry
1TycbOcywdcfBbD3LCbHmzBRmKg+AZ4twQtGrLb7FlMi+6hfgLW7/QWpE2XJyUoi/ZhW96fuvLgn
Nmp6bC8owqKR9OF2nSPg0s1WCv7ZakM/AU9TPqH2xfyYjA/KIBbgp1uT9BqvMzlB4H1FGvSSq0Tu
X/XAL6PUG3JWBIss6jxornpc2h9lUgOTF3huEe3jVLzUcJb8snacYlmVbQA+LiS5Xkmv4HGBQRO6
UT6VUL+D0Zyyq2RWz8X49PZHoLmSupuEsqeXA340cJhYAwv9DpE096Ct3Hk4MLUa0WiOV+QZez6Z
rvRWF/QQbbh5z307sAk5QANIEpYZMybbdOQyt+6TF9FJNh6m7JX5cd+taak3jVV7ejPFNABXEkSu
ZsNteyThoxUPs5v69ks83gtuHtbRQrdBuVBoaYpvPKwS/w7haJ/gugke9PEs56DOJy5E+aGTnbUb
qLHULij3NGpFin+Orblmj2tPVhG1Z5W+po81AwjXDdxwJMrxbEDU6z1YNxwQvJNgellTGZ2FZY3i
Ksc8+GYFwGWSLvsAi7kLrn+E81L1zI9ifnGl84KWxsjDWJiof296HgM1klACXNOewL/QwtQDjasu
KqGB7sERxRejAl0VBCwAY3BipSllzuNTv8GVmJZahus2ogzLBaEVpgksG3k5aik83DPYcTcpIej0
++em4euCvFz/MNUpt/lUFFcHvBD7wbmwrAz+i1RyS7CSYH9mpPR7srO4pQlvNoE25JtApF2Gpomh
TijqRZDYsu4PG7E9bxbNGQvxLkDcjpgnz6+TTV7DhcDtdCa6LHVAPlH7CWOIwsBVTxryMrztLNh+
q7ygtsTC+EyRYz+6u3A0SH0pxQOb3qrWulHdlVBJNfgtLiuYxRy7LG0Po9cRcRgro6YovM45GaFF
Z8frykoMZog6av9awisUAKmwMYEBwHr793LVw4pg+16238YYWomV61Qdd1zYm9fm3xcchKFreJlz
l4Es+KMPAEPmzM1GqQ8P7OnuI6oFEu8Ntt3zZg71KemJ0ewUcQBR17YIA4b/H/Cy6aGSf0yFr1D6
OJf6ThjgD9LGbs5IMhZ4++GAiffbkWIIquVhjz6IgkVkihSphVr9o2OJ8kglPig4P4t3OCkjk/b7
+jjcy6RMsZ97OvWXAzPFoi/rfPKAvpfuejNJgq/+0Zo/wSQneQSBrycI6zC+AO05JsUEQHFxn5Ct
LdPuERoL2+Mca+U3AVvFlMdKSgYnjKgZwzAijrk3M5ATZ+PPqDkVo1/XNqce8QkAuLh4Lfkc3Pg+
rnFsQS+daqVdnuSStUNMXYgLvUzZbjmMXSLI/H6lFAQ59xUUlXWXXWIxu+nUIAegGH4Hvtj2ZOsS
Ovy7MzvnEaf/pDGhzwZtw1qH209y3dpHqYeywmf6BT9NmXv0mKlOo00B4MKkPtoJH2i+gVyV7qzj
XBEHVWDzHF8P/vSWrjA/5+bOwzb1D37yRk+I1sUTbIsplMUwvM33qPPYEmVZGdlJzuRESRhmsx20
TLFLKuzSoJ8ue0nRULcUf8DcxiU3X94kCb/h/DPG4cePapmppqjHUT9f7TgrLEeDFz8FFQ/Ktb8h
yvo/Kab0gOrdsByhZ97E9qKq9PdStd+GrmNGUCf8S4gLtB4TuC7y/eGoihcFnd7ZoSMwOFn+adn4
EgzbfNlsk8+q7uy1KK6ntv2gEiaUW7Gr/YtvgPqc8vElA5LC9qUw36Kq+ATHCyiOi8RYNBJcYYTI
VUwWhfPUJFYcDBchw2vHasETUxLBbuuoEdndwpOOpdcyQtB5r+ncxqmUkB5wi3Ze5VGuk9vj23Jo
xAB4jFP0BXRTdamG9qDTGML80YKrRN4xz1U7Uu+aHc94BAqTh7/6qQSM16WEzXVPI9L2mYzudUKT
hhIr4yIo+g+LsYE5jdDBaB/x1Tiw16kR7M8jQJF3CXp7J82afesPFSWL15SNW3y+ZvCjmZeGOh2k
Qj0FNwjOGl3Ua+SwiAdSJJ14KKShWJJKvig4iRbNnRTcGuhzyMCWyHeh0eF09dlJTHkOaciBA63P
g59lbHNSi16XnGkUF5jJ19pfsEwy+/OMmRALUclIlEhnj5Fgw3/gxmBzfieEL67VJiNcpzm28gVq
4QbW1br/3hZGxsSlq/VBN++DPpfORPxaMMbrZcOSYEeFu9Ieusv0OoUyTAgOM2dCgBRfhgjRIzTN
vMmCA2XKOsq66kA7wfDsFzvTu7DWBj2ghw8HSmxrLvafqzk3uWIpB2mDQBoFnv/Pc/Iy3ja4m5DB
muH6P1bjqkWJxqpfuv+/ihnVWROrAULDXmpObHBYZMh1tO0z7HjCen5PXnABK06oEImu7KHjenvH
z0M281pt8K+45uyY6YojCOjA/wcD3XoA7bUIAXQ2d4jgKHGT2jz/qZyqm7dtQsrw0tNAIf/bkZVp
7jiQFAbSbfpJSAoegPC5cVhdHqiSobW+ocrkcPqzeGLMDu11vFc/dAciNJo8x+YwoCzVGG1wypev
JNdg8heLo52PTQ9Z9RsgIcEc1/wjbRbTGt4qOugTM8TJxqcJhwoc3BDVH1myktGaRV3QQH0+fOnb
4FPV6JB9/QQc/VMVuY+sngRu7tHGJhW5DOkSluPnzgRdg+22JZr3lbm+X9M/TUVEBxOMyllPmZix
D8u7DcRpMhHzLVppo3yHQ2vuuqv2EIUNNutuYXFpfxYOhwP//lXvqvyaDWIQb6zPCeZV8rnJ2QT7
B/SsAEq4+QLuwM2aJb3YPepse1593IWp8vVCGwKVwjPnO2oFA9/NjyKcOegXE9kj3WwVOkmAVUBP
mPz/yN/38DGS43MGKdacBUlv0crY3vdXJbOtGbJl77QtRIQ3ioeb8L4ZPZr3KT8zTWEoIBNVBwM2
lvdsXcfQvu7MgIBnrLeYETEsflHR5ovhlAIh3PRcZCeMez77oXf1gHmC5boVfCbIHbEpWVUdSq3R
gscETNDBOQYJUwxfIRjjxyvF8XPJV7gLDob6HygjJAINEcY0sJF82HlSV7An8htIwC1MLuHHl5N+
d79OD+53oCUVjWGjMupB7I1ze03NrFVhVdxsVdTLMfNmo1JRKkBQYgtZn4TXaQyzuczs6drkjaUR
2NCWPaudE/ywgtsaLPIARcdBoUptHy6mzFzWmgYJMuMsoZSCCEIsETYISRoFcqzoRLhlifGXT1jY
udbi8Tb93RIytdR49iwKDS93WbNBGOiLOv/GRpUKAo4XZ46y57cgcxEiCjZReS7FCyFwB+79dVzV
TJKzr9ZuC68Mz9ai1nu1QiHQjrOhkebSZDne8SGlfT54GdVQM0I9MDbbuqHrri6BeJAwS0mITK3q
Ffc0lFB4FGg24hcUwy3s5v1rj0488A1x4BgXovsO2i3M9EgbFra6wPyUfsg48dtxQYHvyJiJcsxj
4xq0/BBuEUo2SGwhj4yQD4jUtdmEiqucwm3ckdRKzVO87LakXGSFTfHn+LF+Fa5/uLsZ4cVeGZ3T
GQoXmEPwhjiP74knOHo19mAb8uq/x/4UpOzyZU0MKui1fB06xsLjiuxfKzrDAErVOYYamrByfkIV
hNFpoNCGzbs+lVgWClOWgVUJx9L2M9Eh2ReqqSGbbwGqp8RRSwNaE04uCHlThIKy45nga0yWOcCK
nOXcxURBKDAoJfEAHplW6vNeJtFbJ4URwSMBNwlnqQq7+gunGgN8xY9Kpp9RgU4bWjCeQzuMMoct
kSWNklPhxa2fbXZ9FEIWqpEx2nMxh6XfVv1KxVYfHCjzoZvY6Npv4+OLjTynKBE/o25exz12a8fo
CjV63LbyvxLEoMKNqNaE6zGQvyCXfNXDdsijcukrGVDppQoEG38aJ7Fs1r46RuCvdpUi+N0BVlAT
Zw/7lhTITaG7e6i4tNtEQSk27NaAFsZcxQgRZmh+mtiptu9jJh5q+aA2qFKk6wZuh+nPsp9HrqX7
72AFWnC3YAEv3vhFm58XIGuP43nFjkaqt0Uxcwbbgy83KUFFYEVSHy/tr0x8xaSMtSgrG6YxgaQp
vtJ57r7+LaVNzXRRrACF+SyacNDhRZpWzctVxWzLn+ekl3a/xVZZZ44QUcRj2t3tgnljpGwtF85K
/fUZS5Ctf1riyTuKkhd7B/7bB5iKHbVOfxncwtW2sAGOLzvL1MrHIwmpN7ZuIeJ7E0jpjN0POems
9ialrWRndW59eGwARsOFxZ6JoMIAHC0XtOjal8jakkhklL9K/s1ybis3h9Nn8c8/rF90ujkrlFYr
Dqg9xD2JXbTYX/yZ6ccogPb0BP669Xsd0/zVjLiCQpEdmSyJ/ZMFTdfQd5TjZimppeB8ksv7QGoP
irJMwFY11Lh2IkxweoIxyoNORkMYgGbpD1YP6Zilkzx0PMG9a/Owq1uj2REe0j8ehIiCFUUMsNms
RPm8xAEl3VO4770vrpjlXmZQZOoRND14uMjcK6kdqRxlHj7yJ+rBdrSAan2ZKs8sz+8WR5MYcQ15
Rw87smNuLkuK7DBRjVLh7Vl4MKn++usdD/l/ubKctGtbEweJDjhlq9HbRl1iw0cjYYZsWqZZyN/W
5KdA4C147vyRJ5PiIEK0zQAGQsj3UidPmab+HyXRtGFd1SOZVZ/B9YM5jnIBnuhuTfziJGpG6Io3
/PRKViTIKvZmDdWUyXnrOKSPRS4pndlX7WJQmsNUtwgY7tUlKDQNOAqbmpJEY9AbuCqjf740tKiz
SFhdOxW4hO+k+NaNGkQ2TeRt6d0ODgR2Sglud+qJexYUQatx2YlKZWo3Kc0O8NgBSAOv2+jNq+n/
238MhefLYbgmdjBOEeRGuHwLEY5ZEBQvHPSioZkeRoZ/jmGEm3x8qlidA+bdmcEdlq2yj/idHw/C
+30k0rHoAw7x1iAsOx871FXrVocNhypkY99hwzvx0Ct1ac4GbSln68L3Qd7v0J16nj2CDcDUglrq
29NPXUV6kluc3F9YZqfvtJfd1YR84l6KjFdT27OIEIRqXEUkrzh08T3zjIogEOB3RF9NipmfqYWU
E+1tOuzh1mCGQje/q2eQG9M/cl/sMbRauOKfUO+1GXrqwiTGmt7r6C7vevndiPkwSa7FQCIItiV6
NDd/Qyvpe3bYKsqOtTdIDn5zdlY0FKrfDokHbckhAmv5ENXV90e2KTKFDnsbSKkx8db40a+BC0zG
gaoPapFw/BDZcSAGCL7g6K89LDoV609PmEbaxG7IQyQW/dSrcVESH4pvixKAptXK2xG3xN+n0he0
Wz4wmzQBrWztMZY9iuA2wWmmLybqnRVj2VC5J6mSmJZHVu5CL6cnl0Ia/tT3xXjMqWoojQJ2Z9fT
wRUPugtvm6k1h6v4zBe9TqLplG/LZEzTIrXA+rHwcST7XJOcvU5wzN7h29gPj4iMOTAW2m2S2BGK
RqXeoN+Lqhu6q0lRqM2AQUnKL2zfbbtMU8pMrHwZjcjVfRYp3asbwHn7oFWBIB6dVnRdUgmppYgK
QQJPm2iNgeMy8ht90Rg2mgVXBb+K3Clq+jlMft1IkO2KwKQcSJXGoRwom+ICf3mjT+o49EGjAAuX
o64fRU90x3er3ftjpDO5TJOAeOwDxzWTHCjPLrhSUr9Og7fYHFmTZ2xNgAxM+apVkIULc4eS5rfH
6FdSIgSku9fAdma8mupveWsgiTze+ofw5lxb8wL1jSRmT4juN66xD3scHFYU8Pz7SgmPFevATJVR
8uZhgmqvSCvTAKlmq0Fr7FCZ83nBDUninR6066sHBQCIUq5T8LnCeLa2UEX0LPDVxBkcwiHkkSnN
SpOvd1QTp3p+3k27EXYDX1ywNZ8cW3vGAgyHUi8B2wbl2fDoCU2YEutP38m1zq9oD6KLgrCoDGn8
IccQ2t/Uz5FBRy+iSdYuv0Anww7DBJqx9cvQ3oIBxqlfBXhrCQsvM4V6hF2HqKLLkaFixSVJuzC1
3vHn9vgGy9r0QntyZeRlapJvfzHT1zZnsTlMzSsPWiWqik3C/As5bRz61iWOLRC505FwxITvhxPT
qOVVT/dLG9ZV7S1fs69zYpZN0kbbm+o0mKgpz7eU2IbNlEnjpu/lbr486N9oJcapCll8PDEUuMdh
JaemOqyuZcDMY9+Wfwj/cZbWhiaZ4RiSK+NVcM5SHR3BTeQ10nIL7n2eRiQ05PeExPmFtXZ85EUg
BF3DMLiCcs7WeaC99+Jbf4qKQ0yq7ulAjHLuJvVZx03z3PdV+gmcIR7fFnMMka1UPNJx3LxDcTCQ
5GAHlBM/hV27oJbzA/eDF/q8fsBU6XJ5f5Zp9PBAJCyayZsvaHJQSectwTVWj/JfnMGdVUCxMy2C
xlsy+mlf3gST2jRieUJvanRyxsJxlFAA5NWsEayFr6951PxamDF4363EM/+7owyRl3jiBPm6ot9D
UW0IXPzI3WctBWc0/YY/ofjSg1gPfho5xb6ZMUhvI1eykPgHv3jIIoZ9AM5rHa92f1IPSql5mzgZ
L0OwCUo88W/Tw70tQwMNvkxHKStQ+V222hSKVkObpb/8bmYws9MhirzJocHnp9B2DlyKig9API+z
PMjGXi+LXsXh/+zWzN/sNYg07XOz8M4qKBbwoQtgf2jZGh0N2f2HI3K5sMaRhqL0WwfmPaC8kIxP
asdZlyapN5HQrczr4tsE5Hsr+JqkYygG69A0T+Iwu2PKsg5+W09ch+IjdZskWsMKeHrlLjNfTjh4
aFrwkZUNAZg3pg/zKPZT5SzkgGtP7KWVb/26djPTvYOt6AVv1vZeP3fw+UkJOkBtCJ+sDdIsntlC
CgS/IWgj6tGvI27Y2HF97lR9F5s3AcfluwX8jF/kvpFc81W1XRhVvkjl0Lmk0nB3iR/YSzlg/rvg
tH99XfSXxoaz1Hszk6ULktYmlnNuk8i/r48J+mnAiK/3b6EnA0E++MTeCE3i9HIuRJUP34ngL3LX
fesmTjfArsMlzjTMw2KVSC/JIkHHDwrloo3bYBcqkYZszzXHkOtT5EfkIgmf4O2sH48bSZVDxyz8
i5CrLYoQOKUyyIWJmBukK+bcH+0y2K53lhynJf13Pz/gFkVXXH+n/t9SKbsfKeQ+CcVkih50MtYC
DcNITM8UyqDGteaxXsBVnpGc85bAdyD0INDe8lYc7H+vFl3h5QQExO20xdxoMl9dFC2VITENVIhF
YH38QXCmdHdmJeKPKImXO1KaoHEVW+I6mp/u98xmn7TjqDS7uHDb2MsiqHLWfgaWIXOTS3Lq5CRF
8pmtcbYs15Xrrmiyl8d9LusnN2xvSH8LqWdyZVBWAL3YlQmj4c1EvDXHno+19CJh5aysGFcSqTyZ
EDlColPHlAPFiVIhxFslhw33vS0EbpxcyarRq9+04wAIId/JVmphXjqQaS/JO35y76asu503ODd2
R8/PS92EqmrvfldniJJ0psnbYJcamYPJsvdTw0+kkjDbOsjOBu+DVAZd4yVmbCBtnEc94QXAsyVI
WlRDpDWIgvxJy2bZtbszoec9Uzrgm9wHZVGRYCf6rANFVnrt59NYOGmzUsiIdkArCtMCw7ZUMauq
QKis1IjXBjyHGGm4spegM5UANSHtLd3/NQRPB96GUdqTp8aIJdCrfvcq8/814xiL3aiHWmwiPmoo
4xNhCVEdmHpHImrZ73F2CkfukcB9IlbIfOlCjzVVg7SRTu7MzFVm1fJzRofMSD3/FwHhA7dUv38L
2RNEPKcAR/jJS7K4KdBMqG64Id46Yhrw/f80LzZUNkJMYjFnO/+YhPiLeG+nVu+k8otCRQBg1SZN
635NRgBL/tUA/PnyN+Uz8rsP0uZmJ7FdWRiGIPqxnDXCzACplBfrdvDswK4l4ADgOMNcnsHXm6Fv
bfKPFkTFAza9eIl0JCZDdQacDKjrXmwhaU1t4hQosOzu0NRh17OiP/x1vIWSH3wpN5KP+jRBV5U+
COwisbgbUguVH/O79ehb6q6UDSUHX6cpmwA7J0VeI4L0ccPrgW7XvS9v1nmnD6WoaG8N7Biu3xX7
xdrrqEXCYUP7l+qUcLcMBCR6zfbMK48HxW79LBBs7mur05IyhGlC0OvgQkCSZHAf9ISeXJNi8Lgq
HDa1ySc3F56J1AZxiwzLk6oF4GWKFUPYWoYl0OAFbZ06LTcO/RhXR6nuJGISEg85lYvNlW22+XTx
h4gIyj1BhGVcLT+5E3SMBJkXCJzeBNeduScnepYmu2sJjJOcPT+1gvxKLoVPxHk9rDpYD4rnDpjN
L9pU7Xz9HYBEqHxan+kF9+0wyDbae58ecJIWSuS5i1iKDrGa4p1FNWiRs7QyydDFRlx3Yvr+wz/v
1Pr7LCZJl8+KH8sgc7Os6oUHKk932KbSv9Rf7FtMXyqaPLlpRL1CMVUxKadzEJyzTudkz51fJi1g
ZeBQAapQ8XYUAfGGuBcfyh8cVbRVH0FmJ5twDAaHchLOELvt4JR2Yi5I4G3zNPQXeqNf8ib8Uf6H
IuZChZJr3tgOOn3gOHlX8zfLwSd6xez3YMQt8+8IUBLNSvhZKsggFBNpRvEZBSLtouHGbDIgtpRt
mnfpWxA2iLP7auBbTdDsLuCsw7jEqp+w8WUSOcbr7/UmG8BFu644rhi/BOwFaVJ+pJJqSVAuwQzX
fobanUFaDJ1nLKevv7Zbl4tb1eDE5HprvOUi3gETJ50drnL6hetleGKc+4jlFyLQBEMlHszdAqmN
Ksw3EPQgmLjnQK6jHlxunSt0UuUwG1kB1vByDhWOrcuNiYBt8EfiH0CfL8y2Z7iWL7/eShL3XXkq
0lP+1/6asqAckuncVpkwL0PAG7caHjHbTluiKpTAfIxhSZnge4igxhRM0lOGfBHytBBXhcY/N/Y9
qkj8NWlIU460tbP52RxdyQnInOFUEhnLfGvPB4ij57lsfKjvc/2gy1HiYx7MC+d76A34Cbt9KPuZ
+eU7JAAsVXqewdWzVwLkHMV+cUISMVY1J/2iFapA5fJfecPF51I37Ri9ZAd2aZStvrYzZO0AcTV8
Q5P3fZltkOlTgfPJ34Y7gB5k0hCabbwxNbPyYnGaHQ7OMN24tblhz21TChhGqcWpxnaM/bwam4iK
Z1XhnJL92T23sIm1sCaKzDKvGOvlxlyhnRpcDO602Miw/6o0ojJOptHgzSWbsNHKaRySNc+gmzfF
EIEKIrwisDHjGz+zX++6hGO2eGGcFiKwNMDLGMyy2XdIfd15O7FiJgmqOMX4tFQZYqteTeHNBc/v
DXrl0dmGeeTGj/bOQ0vjwn+NAdpFw5pMB+bvZJiTmt4V12qo50bPqWbv3blqdPNJAIXVpTmwMHog
62Kz88yKW+Rn/2GF40IgRXhXCbN52ep9aGHZHnn3XePxQeb9f0ZdH9ySVNgB42gpA1lkPsMUS3yw
V82T8LD12emBnNbc9IfZ7/X9f5Li0dU6tFdpc+fcjA36imNGpQP7M3XEQi0w7ZkBvEY5antxXiZn
7MrpOADHp+Tlq4LiCgbK5C2nhpaNI6tZ84MdIgP8PtKwYXlR0vtJ0Qy2vYzlAMU4dYvlzuWvDsof
bYecJAB65Nja92XlfikK1v+gdqfRVoscLw0cDOB0QAFBqQz1IdDEo30cRW0o+bpCZ5RH2bOGqido
d2+ZSqh3Xfq26xIPyExCIubrkYaEglz5rJv/0sl9t7RsErs0Vtu7Ek0MdUq2ewIQQBYsVWelnhaa
RGVbedzKCXei2JyUFieQgWFMsCYfGW/CWsx5cnuBD/sohsBSG1qbn0yRWctk/ZejMJMVcGahR73W
kO7QMSv51ol3Errm4KQsNYJNmLKr9NwSM+WbCXuz+d/qypzR0mIHDKH4BWF5pZoIQzWIQIcPzf7R
7Ow50uQx5I0CpEFRciZaH2o8NneldcnPL1wh5zv+AuTXGBMb+gflEzNyPwYnbVk34C6agFehEBCp
KWHfIc1rPwDNGrFyl+SmkQcz7WTqUgXQuvxO+YXgkKGE6/2WAVBKxmaTkVfHlbzeSKjStQji8WQV
vSvsqIq30z5838AXKGmY7TDXNBtAbS7vgU+osWSdeRUZfwGDWKCBaRhOsAGEPhehHdrGZPGZ/HFx
FKZhpM2MHdGO2/YgIHmEkhVyjkN9lU3zaGo4ZGeWPQtL2gVTSSOhISJ+auEfufZx0wSmKQ3q+FgV
iqLakvnPJpiEs/nlBv863CS3kd127h2tc4wwBlymuxmIKNOTVzdJzIRTINFormQmv7aCgmfhBtSI
XD5qRm+BhUZsMtq8nDjjxrvUMxs5Zj6RcKCOZO5yyLt+qJpZAn2avUx2grngLNj0s4WQtPeGPqrB
ZyHXIJeZvzwC7nRq3VuFTYvtPG0CFSWwfF7o5CAb5fzHi/Y1amDrqb/SCU1okzbFV9z5g+ZuQxD/
Qft2TwmC0jZANCoHH+61wZe49FOm+Qhp8iw7+GNHhc1VtRQgb3V0R8lOm7RIt9XoQVyQ05Idy79q
L1+F7fUDYnp3JFLAhAFwUX5OVID6YoqlFKRQOgUlwxSRDpfcObowrldm8rTmeDjGbpd1VlhCJamC
LC85EzvN9EweAJMv7juu93h+mQD+BOy69IZWALTZ3aM1eKHPq8p+0LCNVkLsak/udnxvhGVMl7e0
fCorN/le6bftYsTb4IuJCFfiWDwDSy1FQl8LsKv8bH5f1UvO6xcbT6XtDh5JxCSELk+w4sCpV6RN
wSMyoPkBEMMHl535ZSkYNx3AuH54TCfxMTyNBtAmRkQyNa1JdnwfPWhlYjPvi5pAa18L+VhaONIY
7kBBOW+GOL8j/45e4XAcupbhG5mS3GoKwXDwomS5WI8mEJiPcWnDtYTjD1SPfRxvIisjyiVEILst
r/WmP1LvX6MSsUlG3Jy4AK5tUInDwrRgr8ateREHtUteDChA94Jf1oimArow7vZYyYFLqGkmV0Jn
sHvKL6wYZDro40aHCk/AXvU4WEyugoI3iCVN4gqPXzrDGUK8xvUWGn76hkamQGfEBcVFCHWOIQW3
nngoI0uYF51IXY2Y8OlXYgaASQonVu7y8noGqA8g8HYGHwC11c6OaYjyAMHCBX9GwiU18cuuVLzg
CHueRhNm338N6QidmTF4GZVzyWz7Y4EiDFRZ2PZ4ixSihkJYtAIu07+9wWz0sa26AKXqaM608wmG
rH34ILPraIDRuzyAdQsGCoDy/JXkzVd+DmoIQiQ9Bl3sSiZd761YwarZLk8GzLxVQY9691HnmbGw
cHDqkpzypGBHdPZT7uXuzK5dHtnXJUXJUoScCjzCtL6ta3xPpEv9G9JL8MDLaAwtDIYgx5gpOzFM
vd6dFTGppL2a29l2oxG9GkrePTs8xNSGB5EKs07e3bk+1qFKHczacZRvrSd2vy9XaCeeoSUnY/xh
g/CFBqIY+p3IUc0OO3DRq79ej9yLpReTAW8J5HnYYORwEk3/C9cAtxuDBfqh3zVrf0I8om1o+eNc
D9yxDKy+apby30YZw8YtL4TVVPJtL8p7Vn/CogThwIEnzbJRkxPI8ILxw/uqb53oAg6XsCdkpI4G
73plXsS5gn74mm9nwSP55s7MqwBjeQ2pt98Mx4XX04cUdro2Xu6j48fAGeYhEB/OUsReJVwQE5UI
GBw2jBwneExOYOnDr+oxYDtmwULxNAb838dibZGPVkhHF7z2aje58G8maH+1PRlmmSpD4YkEj779
G40eTJqR/1hLhUhFeuNMsBt+Z7usP0Lclpy/N9DjdQNaTs8FLyAsVH1zNL4pjcGS9g96gOWMde+4
6dZV+FmWNlKKxUqyzkSsP6MCLfxL/hFPpwad2tjxMbtG5GOnM5rOFpWf4brvQ+18KDzaSZfROfa3
GpWY8kIiLOZi3fkOYajfxlbrMpP1lhTzK/qJVrWVs3yrB6O2a82C59v+LHjgVCew2/zm5DIlGSui
pCKwiULRDNejcGfH1/vEgrBGx4ARdbV56ULSNgKVhlEwLMFllDdQI0b+0UVTDt7yKiXZpOcgbsMr
rHlOomSQb4IMZCbhJS2TbjzjJJWy/8Gitamvh6GKMA9J7FXoihqctd2oAL8bdN40jYNbldFq78vP
JCcRXhQKhc6gF3Eu0Rj8Ixq1INY6egIkrw68IMMUP0Y8DYqV7LaUjB3i3BuQIk088EOCkBKcrjKM
Oo+8grYIJWjM4xhL5nsRPJkd2qaTkYoaPWcYkHZc2SyA4n29fiPY3xtHVImUE2FW4rCMq2R7glIE
m+nQQ2AaEfm2uswUuFVsFC1q6h0NHK/NpFSyfuu6ORc5K5VEiGvrc4Z3ytGIQ0FT5ShChTi01vFa
PM+FCG5uR/DIHVaTeSGb820SL7fbk6qaOu6wCGxajyzbnnWylu9lFzV9UWf+Q+iAnMJvG1Rbw4Vt
fnF9NZSA807XtmeVPvh694dV8bCWvscmeznGdmQjxXaCPbK9kNwd0X+PQZQTWvvMyK9pPMl6Jvde
oMhPc8K8YCDMAV02E8iSboLATFodnaKatWorztEsJv4Qlk8/40aJp6vAY2KvS/DyuBBPsMs/o3ey
PWWOW9b5vo+U0JvwB0G1lDCHbHmhofk47MTrtjTgIYLBXghJCsjdp1lGdUMd/UcEZb2v2cHF+Q8N
I3wo5N9ZLQKykvzNR4zdVQ8O23STYdwjod2EqMIuUxeuZL8/g4npTKi5xnxxpEo7sX2h20NF/vLy
RVvOK2ah9LydN4oMP7t791/7DAbk9z4CkkQgFfWbG2xmMH+p+2qLUFThU3J6whYZf6JPZ91P2tuI
aKfCXhO0xbK11v+9P4In8WsYCl4fQUyZpDTkVzMx8tImBlVVZBCF8yFh/qXW0HD1/8R9rCKTh6Da
bSZs6tyKgf5gmlDiYECpKbix+i5vvqk2ThE3gi4c2DHeKRmRRbj93sV/mDcslZkfgFk60tXTvYRK
PZOpEFOVwOWJE62s92UTvi/LRKm+1tkZ7uCQBEGW9TPsEXZAEyxykyexJPBtmtMIRZpkVRzGzhRh
RTfjr3m5wjUxlfhHeurHVP/ImROrOteKX8oKjti7aNxPz15Q04VRHNC7bwdnWZPgYaWpBAVrj1HZ
nBSZ3sZUjDOL2xo9wFuOC0sk3gmJrb4zv0nH+3vDfN/YVl/akclzS1cq3dCGz299hJ5yYEvIlKS5
bYf/y7jGiz9GHo9m06sOku7VzprfOz+bSRd/+OD9x9Ea5Y7D44i5SQbcLSGsoDNSeU+NwVqo3DKZ
k2Ysz33o2eR3UMtYRZ3DsY9PBz93XM3C32euEfTk/YpvtfywU+QxSbWcF3aeEoji7znagoCfoS2x
Ehe+tZ71ALJgEFeSp7OcG4Gv6n3PGhk9eDpucY1DiiizlCos8GwUPLBkmEyrhMpUebIp30jiNGFR
UMoSThD4oI4DpbYWtR4Trk9nI8XlwLR2HFwCcB9DoT3vGsojx7LyCL2N7IGgfGsi+SENFCQCIVgW
PBIbI1h4ip1ObQikVAuEvn/QfvN7bMo85RzSLZnJ5DsH9UAuRu/Qy25rtlYKCNAfw+T7GNqT74sI
hK6fXKm2sJvGQK5CUcbXAGcrbNlBv6knyhCefv+6Au1EpLb9eJUPrHiRNBs22o/jtCk+te2p5747
/RQKCGy3RdtAIp+yuDZvcyVGrbumNA6ivHfCFWRNv1pkomsMX8Ki90PVkG59b9mn6Nvo4eTUFDyO
ghX0iigU38R1+6GzlRjdiqaeG5SS4ZKDx6Deo9O84bBToqd4KK7Fq0dfwl0uFwh7/fQj1Oey2uh9
h1tpcCoKDLxI8KvZd54Aa0AuMJ+n93j0HIzwLflLLXIHfIqlvkpgTx/ZrEYBAhDvbdtkISpKd8jO
Bxwl9RpLZ9HxDx8Dea7bexwxGl7ZTeeH4EGdXs1qk/PGk4IHrJcqpTh2kY+6Ftv3j8aRTWMTiqTE
NLdAaTMooxiD3SpIsvC+Nv/eUJMQnz4jE7rmNQ5W5zyaPCqpFPmrddtlZgXIuQSVTbNftyb19rM1
2J/LgUz+gmSXqjUbPP0nmcYxWmeqWM5XHO68ecZP80cqBP7hMBLgpVd99BM4F5GOUZwqYk83lUpk
EIGd6IdNbHp4iH5Ema+kk+OLa30Wm78dDNHVQjaWE/6AOJFkISqqHX7TL3VkBFAgfN1FGnwzx+6j
6Ia8AET1bo6paVbpJxCncuDHXMkeR59ViW5mMxLO1l9Pb4RgN48iRbgqV4fko2vXHKjzgeMepArB
I9Im954ogO5RF/Z2jglP3E5TLb7U8rTK8dvOEJnNrAt6tw1DGeWSHC2zHL/DURc3/OqhdoeR/W+B
LgLRAsq4G7+Gm1OI3zEnbgnaaT8kXwuJ28/EdZJz5iV7uEx44FK+NCE9Bpuu57qXkpRKkjVyllHs
Czm2cicITIVzdJJB1zMeLI4vSVQOpscp3iYACtY6OEPBn65WU1WXzYnAHoenjjf7iixeIF2yuYcg
3EJ72vsEUwOp32riOYn9952gRU7PqBYDm9/GhenEF44H4geSUPLQ0xnpimZ9fAScRl7QJQs0KmTs
rWukzKUHUvr7hec7kGwiXXMWui9i5Nh8v7ZR3mU06AHjggKsbHqCCw/kexCT+odQmBXKYqPsQGmf
Qrjp0MbagrAKbs1Yy9Gcou6sGRtu980TUTIryg741j+OIcVGHrwrYjS9BtpSfiW6L91iG342c9Nr
KeqbLDs3aXo7ZbLTqjts8XZldc+tPEyAv1nzDHW+yd50X0Ujk3jvqJReZRyfAJrkW1+Vb490pkCu
95sjqXlGV0zO2+EUMjwjVDAeLbwNnCc/W7qrFPwVmuTNroDHfREpiAT7FDENkydx0QutaZ75SzoH
jUl3H4O1GXvUjqFE+JEdfegOY9ah5G0hAfETEiwN6e9j/3zinj+FqUvIAVmqaxZAmnIlte7aVnlU
56EJ7vDHf9vEmLC0c2fVakFD5RkpNgyih/hym1mDJuVrRriPY8tsOnB9u4JNXsdPwGjCPb3FZ6qZ
QiwzwuMwYMMrSbbu887x5yWJghQ/sjMLDp14ADg2AiRTYl8cAbmRYFD/Sh6D+1Pns7KT+6Sd3l9d
9Lp0fUDOq8SwGqWpDJzpXEWpXRZKpnY5PpVps9akQOT3/bHR3cQJLKM8AfI7kw8M0rnipRNnEeck
LCW0Tz9GV0zbRaS0eQfqXhyw72wvHo+LPOO94kePlCidnpSaVWI/AuhY/AVPqUJNSQd1VHhCaDMG
rEG5Wy8elsNqq1XUtotHlBmCNWoKdI2dsGT0HumBuqCjA06yoQTky15Igur5Cj3Vm0jLWibKAEwa
6NL4hivQtjIzwuBCNy3re2wdHQxi6csarTg5X3klXuBzGkRLMQeRLQKSN1Ohonhnkx9tLyzOTWLM
uB2YMhniguHvBShf1ARNe0FFNvqXDyhRn8p0bL52BjtuCzI/IGeCuLeYuAilKiRukJLEhKvCwof6
eX+SB0Xa/65hyS2peIizyRnE0YW5jnxvLlE3iYS3+GM4fCljXV6Q9fXc37fceFuCBN0dNv/hiCJY
C1hh/EhZuDzpbQkrKS7cLPtqjEqKNGnZ/B+aZS7vtQFDbKj/MjXpWEnDEQ9pAYZoaY1hOWhM1Ld2
2ADVySe/aazUgi1heZrkNJuOoXCJrzEC0rP7kzTuBNnAgK+28zNcPnYlI7TL/jO0KZX/ThnDYXBe
qv5kxbPGVL3o43gEnV3ieuUvJo8/LUl6/YNOCIDuGj7279pBAvHyp59u9u5IyqhY/KHT7YrLDtqD
mxF3lUfQe4zoE34aWQL3UNuiaV+UthQWK5fDcBlRtk6FVh5fTb21pcxntGXpf+8zxEZVlfb/a3eg
qKFX7ohPJjMw3GX5Jx1ae7LwuSHmNgv/hjISA8zMbvRBs67AC3oRx2fXEYxTSD3mI7exY/LEIDwS
+GPEnQnxEsLcCC7GGMUD8SHYG/GDfeKLQFCQQfkv6ypHhyy+5XE5IEmbDG20gcBMXQ1w66OYhIZU
H55E/+oUvIpP3CBor4CJzYtL3PzgCBqS3aPU4TMsAfbdU6s4EhHVK2E0BiDcfkEbAMDifXSa067j
lPxelkQZJ70TuPCYWLdaS9hIBYfh2iGSTQsPMaviwDHDDA3dxfjtIijjhMndIWiwwrIBLkT+IlDE
DjLLNinNHBt3LKRt++r5XU6ZoaKnckpgfZFJIpz2kfBo7tfhVLY3Xt292h0v4J1tiHId3TDlKU+i
dRETjV9V/IftXyd6kDXB7s6rtdOipSBE9dfxI45jJrFNEIpybo9bJZ8wYemB7xqObdgCg2Ft8fFM
ZySkCt6+hV+yQQqZnjp3lGl37lNovueS4MBTBdm6sjZEAmxxF61pwQ7NG09wpOTE7vqks/ld6GMO
2iFpwoMzrrUW0Q+TPP8466ANKR5QqjXlJZCXaFegWIipAOwhXlWX+r13GHSP4M4l+uqiaq5X0YZv
9m5y+TnuO9Y015ok7qWB8tNNPInLq0VS2Ar9LK5g+gukh8wCdGI2h4rPdzm6tDKqy0x88v4UMc1h
R8zDZDwzUop2VbgLJ8uTXbu4fp/oP1gGP3mk/1xNYYuRmK2DavqvhrpNSWSo5E4FYhDhlFlNDAVR
MwK6NobGZCVVaJaVqIDlQYOzSui83vH/X02RV/pBkcwWnh+oL+oDBnuZ9p4/eOQbPIlFF+5H+5I+
XZzfV2Osk0SCemJwE7rYS3K63QS2LG+AfNlTbn3/hWLD9ULgqqqwgwmZPrPFtyPnxiqsRySKdpJP
YjvGMKJCgTXZTW2VafyOKRAUhZk1tOTKDU+AA5iZy1qWizOfeu8qTHwLBUxYmfSXXwKuQ0LP3fNC
Bh+niQ9+RxC2iGmljSzlcFx5BTmokGKSCP9qUPCjmMEM6fA3CU0rizjGacK+4LBvqyme1nGaHvBa
nZYu0DNnm3Y/nizMj16XTq/CTrF/3hfGSR6sz6yoA7zueftlvFbSbQk4IPJ2Qsr5YMgHGjSvaWAo
g6aSTDQImGpshzUKEuA7KLLpm9eCDIs6asuxUxJ31qxO3td2QQgS9Kiy0F6B72+clL+mraIAmA41
jodTLC679QKpKiHxz6ocCZ+AGJSaDAvb5rhO4S33BopTd+iV7p6poPxAVYdO8sL64nPfOmTBh1gE
4ELkQvbWf6/bVlDkZZL6HhzEdckuPLXPxGCyMmMgAmYyPZWL4Ndj/lGKJcQ3Yj9CaSTkQBXdj7ab
01Ny7ZT/TmK8Pi63TgsgkS2QEanN9sMNKWs6X0upvguaDmMGLq1HCCqzXkuaHzFfuZrAbGtLxgUI
yRTHHN81irN2y7TlCr+J1PFQKp/BNzqP9l9pQ3o4fr1M0QD0qnhZkuVG27qCX+y/rBKyN1BUDS2o
Igp6RpK7zl1rC2x5RMlLl4urAZljqvNjUcekRM7tjzCVSQSmI46+tPV2CLoNqPEuDzuXh4Ysmt5B
u7kAxmo4XZzHU9d+dcYw9mAnu4Sxpxk4sS0QbyUIr2jjAc56NnmD8cAdj15XSp4To2ysjdoSrRC5
TVSNUcQoHHQJWCpNkN1cuZy2FbJf2aZeDDq7nAOuyAANWrR/dTjB+419wgo6WuDrsnYDJ/3+ey5i
Qk14Pf0FupQDbSSHn22e/OyyveABk3NXPyLUBwGmyzfWttHIwbflZfoB05cVxi3njJwOrMbk0aDv
8eraBUR5vgfjnI65RAIQqs+Q9UOYwUU97Th0mO8OLCkfYZBXFuy3EQGxZLaAPqARnqDgrRutsVtS
gS//jM/p/EbeyHth6FeibDroLTIjfDQVvd44uDAm4NpxsuyRE9H0T8cx06vL7AjewKsXmZMfdiZF
sNtZ9BJTgXCflAPDXbpnu4Eato64FsSWR/uC6Kkia3oMqOatvtVzIR60ahrQGRX7ad4Zjy+hIDa+
1AN/Mk9k+D9n55+55mhd3x6dP2wdxhAlTSuctn99aI40mNVH8NBW28NGqe+fjXW0OKU2jpHOxIpI
n2pNE5xWbYit3CTchu8vGQSys4cpv3awaBcL/CNPNC3o7UFy/IsGKPiflaGqI9BRDuWAQHKwV624
xqhkqILvykA4rQBUqVKqGW9htYA3vZoeq2Let31IRlXQoB88NXc/X90iusWeFvoHzs/QUoYlY0ZU
NGGbSevpF7v8HbQWaRzK+5u5vwXXQIjaq/YRftWPEdjS6IIppB+J8GOnOILCQHCBDrOB6F8YsWeC
JqO6vqryZ9/2v2F50oPrqkNqkhVseeh0p6+pumhUE63aaKZIQakTglgyJh++yuGgLYGtYFA23dO5
Ba9QEclyf/9lzgh2vanTNaaCNgfotrcScIRjPhNPGD85k1Xpv7le1g4PcmTL4eOnIYowHBnZlhXJ
GrVqQhxO4ML9DVNgGFwqzm6Qh1j6PY9UtILolwF4y3qhRd00mLM1B13MvFyh8L6WRJxf4abik2NX
fNx++9LSMebovsDZl+zyRpjlUWMpcw1eyw9yhezrczDhoAytep/3J1L/LA7alp7KLtqV/X9sPjTU
86IEyLMqJ2ey3gCcG6a8q76erSltnGuHb94meDAMdf6DtQKVUEHJ8vG/YRJB4/tgIfOJPFXehLjC
Il6/ml1yL69w9c5Zqdb8mipZph+bydyThaQMOpXbr1RJC4gZHhC4I4dE15KRmemXRDhh87B9Vgx1
LPeXkvHHVsne8t9r5iTixWBR/ProoIj6XBrxcDUvc8PQFXd/E2mQbRaqnKy7xOaz4wFfmZyj69u5
VZzxaHcCrh1z0zAys6xjSpKH5mTAl6lSHXa9uChIMn4OJKQawLfNKuE8PuxucSSzACd1YPYByFSm
xSiVrVvulI49jcScJsyU4zNJc9V7Tl81qZMt7L1SlwolEA9WuBwbUu+l6cUIkBvyjU0T3T2c75By
TFsHlPeDjl2PNi9vmwEsXM6qM4GrNHkJD2Lh+cO6Riqp7tI5VGpQqoTPJt3PKuT96F+EbMgV9rcj
oFlhrzHj2hbZ4gtyIrMvjWdMI0PFKLe/Ogr5iwwb7RBJdVl6e5IXufNRz9cc28TYek4VCFlJLBJ6
xWZTCwZo7/KXbsxs00fGYKq2GUpe+hcngLDs0zw12t5pgJDVtgf9OhFHhUmRongBzp2f5KKzdM8V
aOUmFaD3olVGMQetbhqE75xCmABJ/kvffwJ33omsslX0Aq99AxE2tw2G/qpTWenkIHRzlkJYC9x3
4i80x7vl1C2RpJ3WfSDEl0dbedZqnXoZslihOasK6aNe7LjTnt/AOzW4FOQqp3A2uT4cwVJJZHyf
7Z8Y2LbOygw9QuA/IP+iNLVeiCWG3GiTBCO7WEmY2U4I546iuI+46jVw7vrAd+V49ZXtvzL/OeSb
4qifQ4ihXtdaGLWvdTCCEjR3cjbZLT9hjv2iVkIkDsZy0a5MolFZzvdRJ8Z0P4BLzJp3PMWoLshB
6IBT9fqorvxeDZ7ncFCaTs0iI+IzA8mA7/nuLyBvuChEyt1VBMsCzXWVnHUiwt23jEtk3xhOL8AO
fYSCmbgb+XJorEtWxTkb/9ng4dSH+M9u62wBHnOSxHfyPiBwj2eFeHsMJm0vuQxOgQWOqdERVB9W
MJBnbhlgBGgypRh05DP+oH6ftQelbp0Trfc6ZYW0VYZC4y8jSK7SSPb47DpZygpiBzcPNw7Bydi6
CdShbMDoz7FBhSzB6J3Ea/WF7rJg1Ui8QIHPXJAU7JwV+K1Bdz6YOnNPeAHwD31ipKqviQ4Vpudr
cNjHfZhXJby26zyCtWLhqO0iTOWuVggbD0hOsLMM4nmk8JZtdy1aqe9lxoy+FACigCHCVnf6bNHl
US4X9DG7leax/dZF4A33VClasEpDPhCDh47EhaxGa4ExqDjEfMNSgCPnpppYYmtYLs8kgpwXX2Hn
w3CJu7MUlCGVLfXYNmLra+p0es3H2dM2Uz3pNyo6bL8gceTmROB8jonz1im2sThu8MG6I5Ty7+uq
9k2zWo8Taak/9kjIZDtZ6mJN3MIof4Z6h4JrSYC0UzQTlFepHrgbM5nvsiNw6GZ4ugKsQB+muNLR
2Y4TalL7WUwvjSEEC+zSD3ZR6YqFTTnFOpRuVqIWTKTxyulogVzzA6SPpyF07wwZ6UOzkxToSNXI
T1n/hFZ2sPd4rVn9V9f0fnEUjc7NneI4xfz4DwIBQifDrsqyuDT8pktqO0nLER0GALLshxtYNqnX
cG2S2jYDPfeGktJBqFgomUzT7enc8PzJnGf1BbZ4Ampc7/pLf6J/4bKI/6km9PvE98ke7Dpacq1V
dLBzozqIa/f40i+GY7RA6w7CwRh1iATdVEDeRqdwVwowfvQVrZhj3a65mi6dtrj1nikkah8=
`protect end_protected


-- VHDL global package produced by vc2vhdl from virtual circuit (vc) description 
library ieee;
use ieee.std_logic_1164.all;
package l2_cache_global_package is -- 
  constant default_mem_pool_base_address : std_logic_vector(0 downto 0) := "0";
  component l2_cache is -- 
    port (-- 
      clk : in std_logic;
      reset : in std_logic;
      L2CACHE_TO_MEM_REQUEST_pipe_read_data: out std_logic_vector(109 downto 0);
      L2CACHE_TO_MEM_REQUEST_pipe_read_req : in std_logic_vector(0 downto 0);
      L2CACHE_TO_MEM_REQUEST_pipe_read_ack : out std_logic_vector(0 downto 0);
      L2_RESPONSE_pipe_read_data: out std_logic_vector(64 downto 0);
      L2_RESPONSE_pipe_read_req : in std_logic_vector(0 downto 0);
      L2_RESPONSE_pipe_read_ack : out std_logic_vector(0 downto 0);
      L2_TO_L1_INVALIDATE_pipe_read_data: out std_logic_vector(29 downto 0);
      L2_TO_L1_INVALIDATE_pipe_read_req : in std_logic_vector(0 downto 0);
      L2_TO_L1_INVALIDATE_pipe_read_ack : out std_logic_vector(0 downto 0);
      MEM_TO_L2CACHE_RESPONSE_pipe_write_data: in std_logic_vector(64 downto 0);
      MEM_TO_L2CACHE_RESPONSE_pipe_write_req : in std_logic_vector(0 downto 0);
      MEM_TO_L2CACHE_RESPONSE_pipe_write_ack : out std_logic_vector(0 downto 0);
      NOBLOCK_L2_INVALIDATE_pipe_write_data: in std_logic_vector(30 downto 0);
      NOBLOCK_L2_INVALIDATE_pipe_write_req : in std_logic_vector(0 downto 0);
      NOBLOCK_L2_INVALIDATE_pipe_write_ack : out std_logic_vector(0 downto 0);
      NOBLOCK_L2_REQUEST_pipe_write_data: in std_logic_vector(110 downto 0);
      NOBLOCK_L2_REQUEST_pipe_write_req : in std_logic_vector(0 downto 0);
      NOBLOCK_L2_REQUEST_pipe_write_ack : out std_logic_vector(0 downto 0)); -- 
    -- 
  end component;
  -- 
end package l2_cache_global_package;
-- VHDL produced by vc2vhdl from virtual circuit (vc) description 
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library l2_cache_lib;
use l2_cache_lib.l2_cache_global_package.all;
entity accessL2TagsDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    NOBLOCK_L2_TAGS_REQUEST_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_L2_TAGS_REQUEST_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_L2_TAGS_REQUEST_pipe_read_data : in   std_logic_vector(44 downto 0);
    L2_TAGS_RESPONSE_pipe_write_req : out  std_logic_vector(0 downto 0);
    L2_TAGS_RESPONSE_pipe_write_ack : in   std_logic_vector(0 downto 0);
    L2_TAGS_RESPONSE_pipe_write_data : out  std_logic_vector(33 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity accessL2TagsDaemon;
architecture accessL2TagsDaemon_arch of accessL2TagsDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal accessL2TagsDaemon_CP_2362_start: Boolean;
  signal accessL2TagsDaemon_CP_2362_symbol: Boolean;
  -- volatile/operator module components. 
  -- function library module [accessL2TagMemX4096X8] component not printed.
  component calculateHits_Volatile is -- 
    port ( -- 
      set_valids : in  std_logic_vector(7 downto 0);
      set_dirty_dword_masks : in  std_logic_vector(63 downto 0);
      set_tags : in  std_logic_vector(167 downto 0);
      pa_tag : in  std_logic_vector(20 downto 0);
      replace_index : in  std_logic_vector(2 downto 0);
      is_hit : out  std_logic_vector(0 downto 0);
      dirty_dword_mask : out  std_logic_vector(7 downto 0);
      access_index : out  std_logic_vector(2 downto 0);
      replace_line_is_valid : out  std_logic_vector(0 downto 0);
      replace_pa_tag : out  std_logic_vector(20 downto 0)-- 
    );
    -- 
  end component; 
  component updateDirtyWordMask_Volatile is -- 
    port ( -- 
      invalidate : in  std_logic_vector(0 downto 0);
      read_write_access : in  std_logic_vector(0 downto 0);
      is_hit : in  std_logic_vector(0 downto 0);
      rwbar : in  std_logic_vector(0 downto 0);
      dword_id : in  std_logic_vector(2 downto 0);
      current_dirty_mask : in  std_logic_vector(7 downto 0);
      updated_dirty_mask : out  std_logic_vector(7 downto 0)-- 
    );
    -- 
  end component; 
  component nextFreeIndex_Volatile is -- 
    port ( -- 
      from_index : in  std_logic_vector(2 downto 0);
      set_valids : in  std_logic_vector(7 downto 0);
      next_free_index : out  std_logic_vector(2 downto 0)-- 
    );
    -- 
  end component; 
  component insertIntoSetDirtyDwordMasks_Volatile is -- 
    port ( -- 
      old_set_mask : in  std_logic_vector(63 downto 0);
      index : in  std_logic_vector(2 downto 0);
      ins_mask : in  std_logic_vector(7 downto 0);
      new_set_mask : out  std_logic_vector(63 downto 0)-- 
    );
    -- 
  end component; 
  component updateSetTags_Volatile is -- 
    port ( -- 
      read_write_access : in  std_logic_vector(0 downto 0);
      access_index : in  std_logic_vector(2 downto 0);
      pa_tag : in  std_logic_vector(20 downto 0);
      set_tags : in  std_logic_vector(167 downto 0);
      updated_set_tags : out  std_logic_vector(167 downto 0)-- 
    );
    -- 
  end component; 
  component updateSetValids_Volatile is -- 
    port ( -- 
      invalidate : in  std_logic_vector(0 downto 0);
      read_write_access : in  std_logic_vector(0 downto 0);
      set_valids : in  std_logic_vector(7 downto 0);
      access_index : in  std_logic_vector(2 downto 0);
      updated_set_valids : out  std_logic_vector(7 downto 0)-- 
    );
    -- 
  end component; 
  -- links between control-path and data-path
  signal phi_stmt_2293_ack_0 : boolean;
  signal phi_stmt_2293_req_0 : boolean;
  signal phi_stmt_2310_req_1 : boolean;
  signal phi_stmt_2310_req_0 : boolean;
  signal call_accessL2TagMemX4096X8_expr_2309_inst_req_1 : boolean;
  signal call_accessL2TagMemX4096X8_expr_2309_inst_ack_1 : boolean;
  signal call_accessL2TagMemX4096X8_expr_2309_inst_req_0 : boolean;
  signal call_accessL2TagMemX4096X8_expr_2309_inst_ack_0 : boolean;
  signal phi_stmt_2293_req_1 : boolean;
  signal do_while_stmt_2291_branch_req_0 : boolean;
  signal phi_stmt_2310_ack_0 : boolean;
  signal phi_stmt_2318_ack_0 : boolean;
  signal tag_mem_read_2422_2312_buf_req_0 : boolean;
  signal tag_mem_read_2422_2312_buf_ack_0 : boolean;
  signal tag_mem_read_2422_2312_buf_req_1 : boolean;
  signal tag_mem_read_2422_2312_buf_ack_1 : boolean;
  signal phi_stmt_2314_req_0 : boolean;
  signal phi_stmt_2314_req_1 : boolean;
  signal phi_stmt_2314_ack_0 : boolean;
  signal n_request_d_2331_2316_buf_req_0 : boolean;
  signal n_request_d_2331_2316_buf_ack_0 : boolean;
  signal n_request_d_2331_2316_buf_req_1 : boolean;
  signal n_request_d_2331_2316_buf_ack_1 : boolean;
  signal phi_stmt_2318_req_1 : boolean;
  signal phi_stmt_2318_req_0 : boolean;
  signal RPIPE_NOBLOCK_L2_TAGS_REQUEST_2321_inst_req_0 : boolean;
  signal RPIPE_NOBLOCK_L2_TAGS_REQUEST_2321_inst_ack_0 : boolean;
  signal RPIPE_NOBLOCK_L2_TAGS_REQUEST_2321_inst_req_1 : boolean;
  signal RPIPE_NOBLOCK_L2_TAGS_REQUEST_2321_inst_ack_1 : boolean;
  signal phi_stmt_2322_req_1 : boolean;
  signal phi_stmt_2322_req_0 : boolean;
  signal phi_stmt_2322_ack_0 : boolean;
  signal WPIPE_L2_TAGS_RESPONSE_2482_inst_req_0 : boolean;
  signal WPIPE_L2_TAGS_RESPONSE_2482_inst_ack_0 : boolean;
  signal WPIPE_L2_TAGS_RESPONSE_2482_inst_req_1 : boolean;
  signal WPIPE_L2_TAGS_RESPONSE_2482_inst_ack_1 : boolean;
  signal do_while_stmt_2291_branch_ack_0 : boolean;
  signal do_while_stmt_2291_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "accessL2TagsDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  accessL2TagsDaemon_CP_2362_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "accessL2TagsDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessL2TagsDaemon_CP_2362_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= accessL2TagsDaemon_CP_2362_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessL2TagsDaemon_CP_2362_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  accessL2TagsDaemon_CP_2362: Block -- control-path 
    signal accessL2TagsDaemon_CP_2362_elements: BooleanArray(120 downto 0);
    -- 
  begin -- 
    accessL2TagsDaemon_CP_2362_elements(0) <= accessL2TagsDaemon_CP_2362_start;
    accessL2TagsDaemon_CP_2362_symbol <= accessL2TagsDaemon_CP_2362_elements(1);
    -- CP-element group 0:  transition  place  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0:  members (4) 
      -- CP-element group 0: 	 branch_block_stmt_2290/branch_block_stmt_2290__entry__
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_2290/$entry
      -- CP-element group 0: 	 branch_block_stmt_2290/do_while_stmt_2291__entry__
      -- 
    -- CP-element group 1:  transition  place  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	120 
    -- CP-element group 1: successors 
    -- CP-element group 1:  members (4) 
      -- CP-element group 1: 	 branch_block_stmt_2290/branch_block_stmt_2290__exit__
      -- CP-element group 1: 	 branch_block_stmt_2290/$exit
      -- CP-element group 1: 	 branch_block_stmt_2290/do_while_stmt_2291__exit__
      -- CP-element group 1: 	 $exit
      -- 
    accessL2TagsDaemon_CP_2362_elements(1) <= accessL2TagsDaemon_CP_2362_elements(120);
    -- CP-element group 2:  transition  place  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	8 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 branch_block_stmt_2290/do_while_stmt_2291/$entry
      -- CP-element group 2: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291__entry__
      -- 
    accessL2TagsDaemon_CP_2362_elements(2) <= accessL2TagsDaemon_CP_2362_elements(0);
    -- CP-element group 3:  merge  place  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	120 
    -- CP-element group 3:  members (1) 
      -- CP-element group 3: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291__exit__
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(3) is bound as output of CP function.
    -- CP-element group 4:  merge  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	7 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_2290/do_while_stmt_2291/loop_back
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(4) is bound as output of CP function.
    -- CP-element group 5:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	10 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	118 
    -- CP-element group 5: 	119 
    -- CP-element group 5:  members (3) 
      -- CP-element group 5: 	 branch_block_stmt_2290/do_while_stmt_2291/condition_done
      -- CP-element group 5: 	 branch_block_stmt_2290/do_while_stmt_2291/loop_exit/$entry
      -- CP-element group 5: 	 branch_block_stmt_2290/do_while_stmt_2291/loop_taken/$entry
      -- 
    accessL2TagsDaemon_CP_2362_elements(5) <= accessL2TagsDaemon_CP_2362_elements(10);
    -- CP-element group 6:  branch  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	117 
    -- CP-element group 6: successors 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_2290/do_while_stmt_2291/loop_body_done
      -- 
    accessL2TagsDaemon_CP_2362_elements(6) <= accessL2TagsDaemon_CP_2362_elements(117);
    -- CP-element group 7:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	4 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	20 
    -- CP-element group 7: 	100 
    -- CP-element group 7: 	79 
    -- CP-element group 7: 	60 
    -- CP-element group 7: 	41 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/back_edge_to_loop_body
      -- 
    accessL2TagsDaemon_CP_2362_elements(7) <= accessL2TagsDaemon_CP_2362_elements(4);
    -- CP-element group 8:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	22 
    -- CP-element group 8: 	102 
    -- CP-element group 8: 	81 
    -- CP-element group 8: 	62 
    -- CP-element group 8: 	43 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/first_time_through_loop_body
      -- 
    accessL2TagsDaemon_CP_2362_elements(8) <= accessL2TagsDaemon_CP_2362_elements(2);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	16 
    -- CP-element group 9: 	17 
    -- CP-element group 9: 	55 
    -- CP-element group 9: 	116 
    -- CP-element group 9: 	94 
    -- CP-element group 9: 	95 
    -- CP-element group 9: 	54 
    -- CP-element group 9: 	73 
    -- CP-element group 9: 	74 
    -- CP-element group 9: 	35 
    -- CP-element group 9: 	36 
    -- CP-element group 9:  members (2) 
      -- CP-element group 9: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/$entry
      -- CP-element group 9: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/loop_body_start
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(9) is bound as output of CP function.
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	13 
    -- CP-element group 10: 	15 
    -- CP-element group 10: 	116 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	5 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/condition_evaluated
      -- 
    condition_evaluated_2386_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2386_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessL2TagsDaemon_CP_2362_elements(10), ack => do_while_stmt_2291_branch_req_0); -- 
    accessL2TagsDaemon_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 38) := "accessL2TagsDaemon_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= accessL2TagsDaemon_CP_2362_elements(13) & accessL2TagsDaemon_CP_2362_elements(15) & accessL2TagsDaemon_CP_2362_elements(116);
      gj_accessL2TagsDaemon_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessL2TagsDaemon_CP_2362_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	16 
    -- CP-element group 11: 	94 
    -- CP-element group 11: 	54 
    -- CP-element group 11: 	73 
    -- CP-element group 11: 	35 
    -- CP-element group 11: marked-predecessors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	56 
    -- CP-element group 11: 	96 
    -- CP-element group 11: 	75 
    -- CP-element group 11: 	37 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2293_sample_start__ps
      -- CP-element group 11: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/aggregated_phi_sample_req
      -- 
    accessL2TagsDaemon_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0);
      constant joinName: string(1 to 38) := "accessL2TagsDaemon_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= accessL2TagsDaemon_CP_2362_elements(16) & accessL2TagsDaemon_CP_2362_elements(94) & accessL2TagsDaemon_CP_2362_elements(54) & accessL2TagsDaemon_CP_2362_elements(73) & accessL2TagsDaemon_CP_2362_elements(35) & accessL2TagsDaemon_CP_2362_elements(15);
      gj_accessL2TagsDaemon_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessL2TagsDaemon_CP_2362_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	18 
    -- CP-element group 12: 	57 
    -- CP-element group 12: 	97 
    -- CP-element group 12: 	76 
    -- CP-element group 12: 	38 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	13 
    -- CP-element group 12: 	117 
    -- CP-element group 12: marked-successors 
    -- CP-element group 12: 	16 
    -- CP-element group 12: 	94 
    -- CP-element group 12: 	54 
    -- CP-element group 12: 	73 
    -- CP-element group 12: 	35 
    -- CP-element group 12:  members (6) 
      -- CP-element group 12: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2310_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2293_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/aggregated_phi_sample_ack
      -- CP-element group 12: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2314_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2318_sample_completed_
      -- CP-element group 12: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2322_sample_completed_
      -- 
    accessL2TagsDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "accessL2TagsDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= accessL2TagsDaemon_CP_2362_elements(18) & accessL2TagsDaemon_CP_2362_elements(57) & accessL2TagsDaemon_CP_2362_elements(97) & accessL2TagsDaemon_CP_2362_elements(76) & accessL2TagsDaemon_CP_2362_elements(38);
      gj_accessL2TagsDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessL2TagsDaemon_CP_2362_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	12 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	10 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/aggregated_phi_sample_ack_d
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(13) is a control-delay.
    cp_element_13_delay: control_delay_element  generic map(name => " 13_delay", delay_value => 1)  port map(req => accessL2TagsDaemon_CP_2362_elements(12), ack => accessL2TagsDaemon_CP_2362_elements(13), clk => clk, reset =>reset);
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	17 
    -- CP-element group 14: 	55 
    -- CP-element group 14: 	95 
    -- CP-element group 14: 	74 
    -- CP-element group 14: 	36 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	58 
    -- CP-element group 14: 	98 
    -- CP-element group 14: 	77 
    -- CP-element group 14: 	39 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2293_update_start__ps
      -- CP-element group 14: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/aggregated_phi_update_req
      -- 
    accessL2TagsDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "accessL2TagsDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= accessL2TagsDaemon_CP_2362_elements(17) & accessL2TagsDaemon_CP_2362_elements(55) & accessL2TagsDaemon_CP_2362_elements(95) & accessL2TagsDaemon_CP_2362_elements(74) & accessL2TagsDaemon_CP_2362_elements(36);
      gj_accessL2TagsDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessL2TagsDaemon_CP_2362_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	19 
    -- CP-element group 15: 	99 
    -- CP-element group 15: 	78 
    -- CP-element group 15: 	59 
    -- CP-element group 15: 	40 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	10 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	11 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/aggregated_phi_update_ack
      -- 
    accessL2TagsDaemon_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 38) := "accessL2TagsDaemon_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= accessL2TagsDaemon_CP_2362_elements(19) & accessL2TagsDaemon_CP_2362_elements(99) & accessL2TagsDaemon_CP_2362_elements(78) & accessL2TagsDaemon_CP_2362_elements(59) & accessL2TagsDaemon_CP_2362_elements(40);
      gj_accessL2TagsDaemon_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessL2TagsDaemon_CP_2362_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	9 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	12 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	11 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2293_sample_start_
      -- 
    accessL2TagsDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "accessL2TagsDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessL2TagsDaemon_CP_2362_elements(9) & accessL2TagsDaemon_CP_2362_elements(12);
      gj_accessL2TagsDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessL2TagsDaemon_CP_2362_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	9 
    -- CP-element group 17: marked-predecessors 
    -- CP-element group 17: 	114 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	14 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2293_update_start_
      -- 
    accessL2TagsDaemon_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "accessL2TagsDaemon_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessL2TagsDaemon_CP_2362_elements(9) & accessL2TagsDaemon_CP_2362_elements(114);
      gj_accessL2TagsDaemon_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessL2TagsDaemon_CP_2362_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	12 
    -- CP-element group 18: 	58 
    -- CP-element group 18: 	98 
    -- CP-element group 18: 	77 
    -- CP-element group 18: 	39 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2293_sample_completed__ps
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: 	113 
    -- CP-element group 19:  members (2) 
      -- CP-element group 19: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2293_update_completed_
      -- CP-element group 19: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2293_update_completed__ps
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(19) is bound as output of CP function.
    -- CP-element group 20:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	7 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2293_loopback_trigger
      -- 
    accessL2TagsDaemon_CP_2362_elements(20) <= accessL2TagsDaemon_CP_2362_elements(7);
    -- CP-element group 21:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2293_loopback_sample_req_ps
      -- CP-element group 21: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2293_loopback_sample_req
      -- 
    phi_stmt_2293_loopback_sample_req_2402_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2293_loopback_sample_req_2402_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessL2TagsDaemon_CP_2362_elements(21), ack => phi_stmt_2293_req_1); -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(21) is bound as output of CP function.
    -- CP-element group 22:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	8 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2293_entry_trigger
      -- 
    accessL2TagsDaemon_CP_2362_elements(22) <= accessL2TagsDaemon_CP_2362_elements(8);
    -- CP-element group 23:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2293_entry_sample_req
      -- CP-element group 23: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2293_entry_sample_req_ps
      -- 
    phi_stmt_2293_entry_sample_req_2405_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2293_entry_sample_req_2405_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessL2TagsDaemon_CP_2362_elements(23), ack => phi_stmt_2293_req_0); -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(23) is bound as output of CP function.
    -- CP-element group 24:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2293_phi_mux_ack
      -- CP-element group 24: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2293_phi_mux_ack_ps
      -- 
    phi_stmt_2293_phi_mux_ack_2408_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 24_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2293_ack_0, ack => accessL2TagsDaemon_CP_2362_elements(24)); -- 
    -- CP-element group 25:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/konst_2295_sample_start_
      -- CP-element group 25: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/konst_2295_sample_completed__ps
      -- CP-element group 25: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/konst_2295_sample_start__ps
      -- CP-element group 25: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/konst_2295_sample_completed_
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26: 	28 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/konst_2295_update_start__ps
      -- CP-element group 26: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/konst_2295_update_start_
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	28 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (1) 
      -- CP-element group 27: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/konst_2295_update_completed__ps
      -- 
    accessL2TagsDaemon_CP_2362_elements(27) <= accessL2TagsDaemon_CP_2362_elements(28);
    -- CP-element group 28:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: 	26 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	27 
    -- CP-element group 28:  members (1) 
      -- CP-element group 28: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/konst_2295_update_completed_
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(28) is a control-delay.
    cp_element_28_delay: control_delay_element  generic map(name => " 28_delay", delay_value => 1)  port map(req => accessL2TagsDaemon_CP_2362_elements(26), ack => accessL2TagsDaemon_CP_2362_elements(28), clk => clk, reset =>reset);
    -- CP-element group 29:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/call_accessL2TagMemX4096X8_expr_2309_sample_start__ps
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	32 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/call_accessL2TagMemX4096X8_expr_2309_update_start__ps
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(30) is bound as output of CP function.
    -- CP-element group 31:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: marked-predecessors 
    -- CP-element group 31: 	33 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (3) 
      -- CP-element group 31: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/call_accessL2TagMemX4096X8_expr_2309_Sample/req
      -- CP-element group 31: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/call_accessL2TagMemX4096X8_expr_2309_Sample/$entry
      -- CP-element group 31: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/call_accessL2TagMemX4096X8_expr_2309_sample_start_
      -- 
    req_2429_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2429_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessL2TagsDaemon_CP_2362_elements(31), ack => call_accessL2TagMemX4096X8_expr_2309_inst_req_0); -- 
    accessL2TagsDaemon_cp_element_group_31: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "accessL2TagsDaemon_cp_element_group_31"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessL2TagsDaemon_CP_2362_elements(29) & accessL2TagsDaemon_CP_2362_elements(33);
      gj_accessL2TagsDaemon_cp_element_group_31 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessL2TagsDaemon_CP_2362_elements(31), clk => clk, reset => reset); --
    end block;
    -- CP-element group 32:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	30 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	34 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/call_accessL2TagMemX4096X8_expr_2309_Update/req
      -- CP-element group 32: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/call_accessL2TagMemX4096X8_expr_2309_Update/$entry
      -- CP-element group 32: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/call_accessL2TagMemX4096X8_expr_2309_update_start_
      -- 
    req_2434_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2434_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessL2TagsDaemon_CP_2362_elements(32), ack => call_accessL2TagMemX4096X8_expr_2309_inst_req_1); -- 
    accessL2TagsDaemon_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "accessL2TagsDaemon_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessL2TagsDaemon_CP_2362_elements(30) & accessL2TagsDaemon_CP_2362_elements(34);
      gj_accessL2TagsDaemon_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessL2TagsDaemon_CP_2362_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: successors 
    -- CP-element group 33: marked-successors 
    -- CP-element group 33: 	31 
    -- CP-element group 33:  members (4) 
      -- CP-element group 33: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/call_accessL2TagMemX4096X8_expr_2309_Sample/ack
      -- CP-element group 33: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/call_accessL2TagMemX4096X8_expr_2309_sample_completed__ps
      -- CP-element group 33: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/call_accessL2TagMemX4096X8_expr_2309_sample_completed_
      -- CP-element group 33: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/call_accessL2TagMemX4096X8_expr_2309_Sample/$exit
      -- 
    ack_2430_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 33_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_accessL2TagMemX4096X8_expr_2309_inst_ack_0, ack => accessL2TagsDaemon_CP_2362_elements(33)); -- 
    -- CP-element group 34:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	32 
    -- CP-element group 34:  members (4) 
      -- CP-element group 34: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/call_accessL2TagMemX4096X8_expr_2309_Update/ack
      -- CP-element group 34: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/call_accessL2TagMemX4096X8_expr_2309_Update/$exit
      -- CP-element group 34: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/call_accessL2TagMemX4096X8_expr_2309_update_completed_
      -- CP-element group 34: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/call_accessL2TagMemX4096X8_expr_2309_update_completed__ps
      -- 
    ack_2435_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_accessL2TagMemX4096X8_expr_2309_inst_ack_1, ack => accessL2TagsDaemon_CP_2362_elements(34)); -- 
    -- CP-element group 35:  join  transition  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	9 
    -- CP-element group 35: marked-predecessors 
    -- CP-element group 35: 	12 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	11 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2310_sample_start_
      -- 
    accessL2TagsDaemon_cp_element_group_35: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "accessL2TagsDaemon_cp_element_group_35"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessL2TagsDaemon_CP_2362_elements(9) & accessL2TagsDaemon_CP_2362_elements(12);
      gj_accessL2TagsDaemon_cp_element_group_35 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessL2TagsDaemon_CP_2362_elements(35), clk => clk, reset => reset); --
    end block;
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	9 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	114 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	14 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2310_update_start_
      -- 
    accessL2TagsDaemon_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "accessL2TagsDaemon_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessL2TagsDaemon_CP_2362_elements(9) & accessL2TagsDaemon_CP_2362_elements(114);
      gj_accessL2TagsDaemon_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessL2TagsDaemon_CP_2362_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	11 
    -- CP-element group 37: successors 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2310_sample_start__ps
      -- 
    accessL2TagsDaemon_CP_2362_elements(37) <= accessL2TagsDaemon_CP_2362_elements(11);
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	12 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2310_sample_completed__ps
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(38) is bound as output of CP function.
    -- CP-element group 39:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	14 
    -- CP-element group 39: 	18 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2310_update_start__ps
      -- 
    accessL2TagsDaemon_cp_element_group_39: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "accessL2TagsDaemon_cp_element_group_39"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessL2TagsDaemon_CP_2362_elements(14) & accessL2TagsDaemon_CP_2362_elements(18);
      gj_accessL2TagsDaemon_cp_element_group_39 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessL2TagsDaemon_CP_2362_elements(39), clk => clk, reset => reset); --
    end block;
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	15 
    -- CP-element group 40: 	113 
    -- CP-element group 40:  members (2) 
      -- CP-element group 40: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2310_update_completed_
      -- CP-element group 40: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2310_update_completed__ps
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(40) is bound as output of CP function.
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	7 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2310_loopback_trigger
      -- 
    accessL2TagsDaemon_CP_2362_elements(41) <= accessL2TagsDaemon_CP_2362_elements(7);
    -- CP-element group 42:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2310_loopback_sample_req
      -- CP-element group 42: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2310_loopback_sample_req_ps
      -- 
    phi_stmt_2310_loopback_sample_req_2446_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2310_loopback_sample_req_2446_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessL2TagsDaemon_CP_2362_elements(42), ack => phi_stmt_2310_req_0); -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(42) is bound as output of CP function.
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	8 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2310_entry_trigger
      -- 
    accessL2TagsDaemon_CP_2362_elements(43) <= accessL2TagsDaemon_CP_2362_elements(8);
    -- CP-element group 44:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2310_entry_sample_req
      -- CP-element group 44: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2310_entry_sample_req_ps
      -- 
    phi_stmt_2310_entry_sample_req_2449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2310_entry_sample_req_2449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessL2TagsDaemon_CP_2362_elements(44), ack => phi_stmt_2310_req_1); -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(44) is bound as output of CP function.
    -- CP-element group 45:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2310_phi_mux_ack
      -- CP-element group 45: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2310_phi_mux_ack_ps
      -- 
    phi_stmt_2310_phi_mux_ack_2452_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 45_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2310_ack_0, ack => accessL2TagsDaemon_CP_2362_elements(45)); -- 
    -- CP-element group 46:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46: 	48 
    -- CP-element group 46:  members (4) 
      -- CP-element group 46: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/R_tag_mem_read_2312_sample_start__ps
      -- CP-element group 46: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/R_tag_mem_read_2312_sample_start_
      -- CP-element group 46: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/R_tag_mem_read_2312_Sample/$entry
      -- CP-element group 46: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/R_tag_mem_read_2312_Sample/req
      -- 
    req_2465_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2465_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessL2TagsDaemon_CP_2362_elements(46), ack => tag_mem_read_2422_2312_buf_req_0); -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	49 
    -- CP-element group 47:  members (4) 
      -- CP-element group 47: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/R_tag_mem_read_2312_update_start__ps
      -- CP-element group 47: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/R_tag_mem_read_2312_update_start_
      -- CP-element group 47: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/R_tag_mem_read_2312_Update/$entry
      -- CP-element group 47: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/R_tag_mem_read_2312_Update/req
      -- 
    req_2470_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2470_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessL2TagsDaemon_CP_2362_elements(47), ack => tag_mem_read_2422_2312_buf_req_1); -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	46 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (4) 
      -- CP-element group 48: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/R_tag_mem_read_2312_sample_completed__ps
      -- CP-element group 48: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/R_tag_mem_read_2312_sample_completed_
      -- CP-element group 48: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/R_tag_mem_read_2312_Sample/$exit
      -- CP-element group 48: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/R_tag_mem_read_2312_Sample/ack
      -- 
    ack_2466_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 48_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => tag_mem_read_2422_2312_buf_ack_0, ack => accessL2TagsDaemon_CP_2362_elements(48)); -- 
    -- CP-element group 49:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	47 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (4) 
      -- CP-element group 49: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/R_tag_mem_read_2312_update_completed__ps
      -- CP-element group 49: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/R_tag_mem_read_2312_update_completed_
      -- CP-element group 49: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/R_tag_mem_read_2312_Update/$exit
      -- CP-element group 49: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/R_tag_mem_read_2312_Update/ack
      -- 
    ack_2471_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 49_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => tag_mem_read_2422_2312_buf_ack_1, ack => accessL2TagsDaemon_CP_2362_elements(49)); -- 
    -- CP-element group 50:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (4) 
      -- CP-element group 50: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/konst_2313_sample_start__ps
      -- CP-element group 50: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/konst_2313_sample_completed__ps
      -- CP-element group 50: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/konst_2313_sample_start_
      -- CP-element group 50: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/konst_2313_sample_completed_
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(50) is bound as output of CP function.
    -- CP-element group 51:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (2) 
      -- CP-element group 51: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/konst_2313_update_start__ps
      -- CP-element group 51: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/konst_2313_update_start_
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(51) is bound as output of CP function.
    -- CP-element group 52:  join  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	53 
    -- CP-element group 52: successors 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/konst_2313_update_completed__ps
      -- 
    accessL2TagsDaemon_CP_2362_elements(52) <= accessL2TagsDaemon_CP_2362_elements(53);
    -- CP-element group 53:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	52 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/konst_2313_update_completed_
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(53) is a control-delay.
    cp_element_53_delay: control_delay_element  generic map(name => " 53_delay", delay_value => 1)  port map(req => accessL2TagsDaemon_CP_2362_elements(51), ack => accessL2TagsDaemon_CP_2362_elements(53), clk => clk, reset =>reset);
    -- CP-element group 54:  join  transition  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	9 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	12 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	11 
    -- CP-element group 54:  members (1) 
      -- CP-element group 54: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2314_sample_start_
      -- 
    accessL2TagsDaemon_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "accessL2TagsDaemon_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessL2TagsDaemon_CP_2362_elements(9) & accessL2TagsDaemon_CP_2362_elements(12);
      gj_accessL2TagsDaemon_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessL2TagsDaemon_CP_2362_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  join  transition  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	9 
    -- CP-element group 55: marked-predecessors 
    -- CP-element group 55: 	114 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	14 
    -- CP-element group 55:  members (1) 
      -- CP-element group 55: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2314_update_start_
      -- 
    accessL2TagsDaemon_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "accessL2TagsDaemon_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessL2TagsDaemon_CP_2362_elements(9) & accessL2TagsDaemon_CP_2362_elements(114);
      gj_accessL2TagsDaemon_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessL2TagsDaemon_CP_2362_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	11 
    -- CP-element group 56: successors 
    -- CP-element group 56:  members (1) 
      -- CP-element group 56: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2314_sample_start__ps
      -- 
    accessL2TagsDaemon_CP_2362_elements(56) <= accessL2TagsDaemon_CP_2362_elements(11);
    -- CP-element group 57:  join  transition  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	12 
    -- CP-element group 57:  members (1) 
      -- CP-element group 57: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2314_sample_completed__ps
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(57) is bound as output of CP function.
    -- CP-element group 58:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	14 
    -- CP-element group 58: 	18 
    -- CP-element group 58: successors 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2314_update_start__ps
      -- 
    accessL2TagsDaemon_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "accessL2TagsDaemon_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessL2TagsDaemon_CP_2362_elements(14) & accessL2TagsDaemon_CP_2362_elements(18);
      gj_accessL2TagsDaemon_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessL2TagsDaemon_CP_2362_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	15 
    -- CP-element group 59: 	113 
    -- CP-element group 59:  members (2) 
      -- CP-element group 59: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2314_update_completed_
      -- CP-element group 59: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2314_update_completed__ps
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(59) is bound as output of CP function.
    -- CP-element group 60:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	7 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2314_loopback_trigger
      -- 
    accessL2TagsDaemon_CP_2362_elements(60) <= accessL2TagsDaemon_CP_2362_elements(7);
    -- CP-element group 61:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2314_loopback_sample_req
      -- CP-element group 61: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2314_loopback_sample_req_ps
      -- 
    phi_stmt_2314_loopback_sample_req_2490_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2314_loopback_sample_req_2490_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessL2TagsDaemon_CP_2362_elements(61), ack => phi_stmt_2314_req_0); -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(61) is bound as output of CP function.
    -- CP-element group 62:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	8 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (1) 
      -- CP-element group 62: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2314_entry_trigger
      -- 
    accessL2TagsDaemon_CP_2362_elements(62) <= accessL2TagsDaemon_CP_2362_elements(8);
    -- CP-element group 63:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2314_entry_sample_req
      -- CP-element group 63: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2314_entry_sample_req_ps
      -- 
    phi_stmt_2314_entry_sample_req_2493_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2314_entry_sample_req_2493_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessL2TagsDaemon_CP_2362_elements(63), ack => phi_stmt_2314_req_1); -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(63) is bound as output of CP function.
    -- CP-element group 64:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (2) 
      -- CP-element group 64: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2314_phi_mux_ack
      -- CP-element group 64: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2314_phi_mux_ack_ps
      -- 
    phi_stmt_2314_phi_mux_ack_2496_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2314_ack_0, ack => accessL2TagsDaemon_CP_2362_elements(64)); -- 
    -- CP-element group 65:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (4) 
      -- CP-element group 65: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/R_n_request_d_2316_sample_start__ps
      -- CP-element group 65: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/R_n_request_d_2316_sample_start_
      -- CP-element group 65: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/R_n_request_d_2316_Sample/$entry
      -- CP-element group 65: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/R_n_request_d_2316_Sample/req
      -- 
    req_2509_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2509_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessL2TagsDaemon_CP_2362_elements(65), ack => n_request_d_2331_2316_buf_req_0); -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(65) is bound as output of CP function.
    -- CP-element group 66:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: successors 
    -- CP-element group 66: 	68 
    -- CP-element group 66:  members (4) 
      -- CP-element group 66: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/R_n_request_d_2316_update_start__ps
      -- CP-element group 66: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/R_n_request_d_2316_update_start_
      -- CP-element group 66: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/R_n_request_d_2316_Update/$entry
      -- CP-element group 66: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/R_n_request_d_2316_Update/req
      -- 
    req_2514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessL2TagsDaemon_CP_2362_elements(66), ack => n_request_d_2331_2316_buf_req_1); -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(66) is bound as output of CP function.
    -- CP-element group 67:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (4) 
      -- CP-element group 67: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/R_n_request_d_2316_sample_completed__ps
      -- CP-element group 67: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/R_n_request_d_2316_sample_completed_
      -- CP-element group 67: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/R_n_request_d_2316_Sample/$exit
      -- CP-element group 67: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/R_n_request_d_2316_Sample/ack
      -- 
    ack_2510_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_request_d_2331_2316_buf_ack_0, ack => accessL2TagsDaemon_CP_2362_elements(67)); -- 
    -- CP-element group 68:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	66 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (4) 
      -- CP-element group 68: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/R_n_request_d_2316_update_completed__ps
      -- CP-element group 68: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/R_n_request_d_2316_update_completed_
      -- CP-element group 68: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/R_n_request_d_2316_Update/$exit
      -- CP-element group 68: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/R_n_request_d_2316_Update/ack
      -- 
    ack_2515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_request_d_2331_2316_buf_ack_1, ack => accessL2TagsDaemon_CP_2362_elements(68)); -- 
    -- CP-element group 69:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/konst_2317_sample_start__ps
      -- CP-element group 69: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/konst_2317_sample_completed__ps
      -- CP-element group 69: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/konst_2317_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/konst_2317_sample_completed_
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(69) is bound as output of CP function.
    -- CP-element group 70:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/konst_2317_update_start__ps
      -- CP-element group 70: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/konst_2317_update_start_
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(70) is bound as output of CP function.
    -- CP-element group 71:  join  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	72 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/konst_2317_update_completed__ps
      -- 
    accessL2TagsDaemon_CP_2362_elements(71) <= accessL2TagsDaemon_CP_2362_elements(72);
    -- CP-element group 72:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	71 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/konst_2317_update_completed_
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(72) is a control-delay.
    cp_element_72_delay: control_delay_element  generic map(name => " 72_delay", delay_value => 1)  port map(req => accessL2TagsDaemon_CP_2362_elements(70), ack => accessL2TagsDaemon_CP_2362_elements(72), clk => clk, reset =>reset);
    -- CP-element group 73:  join  transition  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: 	9 
    -- CP-element group 73: marked-predecessors 
    -- CP-element group 73: 	12 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	11 
    -- CP-element group 73:  members (1) 
      -- CP-element group 73: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2318_sample_start_
      -- 
    accessL2TagsDaemon_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "accessL2TagsDaemon_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessL2TagsDaemon_CP_2362_elements(9) & accessL2TagsDaemon_CP_2362_elements(12);
      gj_accessL2TagsDaemon_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessL2TagsDaemon_CP_2362_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  join  transition  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	9 
    -- CP-element group 74: marked-predecessors 
    -- CP-element group 74: 	78 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	14 
    -- CP-element group 74:  members (1) 
      -- CP-element group 74: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2318_update_start_
      -- 
    accessL2TagsDaemon_cp_element_group_74: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "accessL2TagsDaemon_cp_element_group_74"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessL2TagsDaemon_CP_2362_elements(9) & accessL2TagsDaemon_CP_2362_elements(78);
      gj_accessL2TagsDaemon_cp_element_group_74 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessL2TagsDaemon_CP_2362_elements(74), clk => clk, reset => reset); --
    end block;
    -- CP-element group 75:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	11 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (1) 
      -- CP-element group 75: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2318_sample_start__ps
      -- 
    accessL2TagsDaemon_CP_2362_elements(75) <= accessL2TagsDaemon_CP_2362_elements(11);
    -- CP-element group 76:  join  transition  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	12 
    -- CP-element group 76:  members (1) 
      -- CP-element group 76: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2318_sample_completed__ps
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(76) is bound as output of CP function.
    -- CP-element group 77:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	14 
    -- CP-element group 77: 	18 
    -- CP-element group 77: successors 
    -- CP-element group 77:  members (1) 
      -- CP-element group 77: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2318_update_start__ps
      -- 
    accessL2TagsDaemon_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "accessL2TagsDaemon_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessL2TagsDaemon_CP_2362_elements(14) & accessL2TagsDaemon_CP_2362_elements(18);
      gj_accessL2TagsDaemon_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessL2TagsDaemon_CP_2362_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	15 
    -- CP-element group 78: marked-successors 
    -- CP-element group 78: 	74 
    -- CP-element group 78:  members (2) 
      -- CP-element group 78: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2318_update_completed_
      -- CP-element group 78: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2318_update_completed__ps
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(78) is bound as output of CP function.
    -- CP-element group 79:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	7 
    -- CP-element group 79: successors 
    -- CP-element group 79:  members (1) 
      -- CP-element group 79: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2318_loopback_trigger
      -- 
    accessL2TagsDaemon_CP_2362_elements(79) <= accessL2TagsDaemon_CP_2362_elements(7);
    -- CP-element group 80:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: successors 
    -- CP-element group 80:  members (2) 
      -- CP-element group 80: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2318_loopback_sample_req
      -- CP-element group 80: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2318_loopback_sample_req_ps
      -- 
    phi_stmt_2318_loopback_sample_req_2534_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2318_loopback_sample_req_2534_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessL2TagsDaemon_CP_2362_elements(80), ack => phi_stmt_2318_req_1); -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(80) is bound as output of CP function.
    -- CP-element group 81:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	8 
    -- CP-element group 81: successors 
    -- CP-element group 81:  members (1) 
      -- CP-element group 81: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2318_entry_trigger
      -- 
    accessL2TagsDaemon_CP_2362_elements(81) <= accessL2TagsDaemon_CP_2362_elements(8);
    -- CP-element group 82:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: successors 
    -- CP-element group 82:  members (2) 
      -- CP-element group 82: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2318_entry_sample_req
      -- CP-element group 82: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2318_entry_sample_req_ps
      -- 
    phi_stmt_2318_entry_sample_req_2537_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2318_entry_sample_req_2537_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessL2TagsDaemon_CP_2362_elements(82), ack => phi_stmt_2318_req_0); -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(82) is bound as output of CP function.
    -- CP-element group 83:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: successors 
    -- CP-element group 83:  members (2) 
      -- CP-element group 83: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2318_phi_mux_ack
      -- CP-element group 83: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2318_phi_mux_ack_ps
      -- 
    phi_stmt_2318_phi_mux_ack_2540_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2318_ack_0, ack => accessL2TagsDaemon_CP_2362_elements(83)); -- 
    -- CP-element group 84:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: successors 
    -- CP-element group 84:  members (4) 
      -- CP-element group 84: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/konst_2320_sample_start__ps
      -- CP-element group 84: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/konst_2320_sample_completed__ps
      -- CP-element group 84: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/konst_2320_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/konst_2320_sample_completed_
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(84) is bound as output of CP function.
    -- CP-element group 85:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (2) 
      -- CP-element group 85: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/konst_2320_update_start__ps
      -- CP-element group 85: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/konst_2320_update_start_
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(85) is bound as output of CP function.
    -- CP-element group 86:  join  transition  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	87 
    -- CP-element group 86: successors 
    -- CP-element group 86:  members (1) 
      -- CP-element group 86: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/konst_2320_update_completed__ps
      -- 
    accessL2TagsDaemon_CP_2362_elements(86) <= accessL2TagsDaemon_CP_2362_elements(87);
    -- CP-element group 87:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	86 
    -- CP-element group 87:  members (1) 
      -- CP-element group 87: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/konst_2320_update_completed_
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(87) is a control-delay.
    cp_element_87_delay: control_delay_element  generic map(name => " 87_delay", delay_value => 1)  port map(req => accessL2TagsDaemon_CP_2362_elements(85), ack => accessL2TagsDaemon_CP_2362_elements(87), clk => clk, reset =>reset);
    -- CP-element group 88:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (1) 
      -- CP-element group 88: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/RPIPE_NOBLOCK_L2_TAGS_REQUEST_2321_sample_start__ps
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(88) is bound as output of CP function.
    -- CP-element group 89:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (1) 
      -- CP-element group 89: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/RPIPE_NOBLOCK_L2_TAGS_REQUEST_2321_update_start__ps
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(89) is bound as output of CP function.
    -- CP-element group 90:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: marked-predecessors 
    -- CP-element group 90: 	93 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	92 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/RPIPE_NOBLOCK_L2_TAGS_REQUEST_2321_sample_start_
      -- CP-element group 90: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/RPIPE_NOBLOCK_L2_TAGS_REQUEST_2321_Sample/$entry
      -- CP-element group 90: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/RPIPE_NOBLOCK_L2_TAGS_REQUEST_2321_Sample/rr
      -- 
    rr_2561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessL2TagsDaemon_CP_2362_elements(90), ack => RPIPE_NOBLOCK_L2_TAGS_REQUEST_2321_inst_req_0); -- 
    accessL2TagsDaemon_cp_element_group_90: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "accessL2TagsDaemon_cp_element_group_90"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessL2TagsDaemon_CP_2362_elements(88) & accessL2TagsDaemon_CP_2362_elements(93);
      gj_accessL2TagsDaemon_cp_element_group_90 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessL2TagsDaemon_CP_2362_elements(90), clk => clk, reset => reset); --
    end block;
    -- CP-element group 91:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	92 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/RPIPE_NOBLOCK_L2_TAGS_REQUEST_2321_update_start_
      -- CP-element group 91: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/RPIPE_NOBLOCK_L2_TAGS_REQUEST_2321_Update/$entry
      -- CP-element group 91: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/RPIPE_NOBLOCK_L2_TAGS_REQUEST_2321_Update/cr
      -- 
    cr_2566_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2566_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessL2TagsDaemon_CP_2362_elements(91), ack => RPIPE_NOBLOCK_L2_TAGS_REQUEST_2321_inst_req_1); -- 
    accessL2TagsDaemon_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "accessL2TagsDaemon_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessL2TagsDaemon_CP_2362_elements(92) & accessL2TagsDaemon_CP_2362_elements(89);
      gj_accessL2TagsDaemon_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessL2TagsDaemon_CP_2362_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	90 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	91 
    -- CP-element group 92:  members (4) 
      -- CP-element group 92: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/RPIPE_NOBLOCK_L2_TAGS_REQUEST_2321_sample_completed__ps
      -- CP-element group 92: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/RPIPE_NOBLOCK_L2_TAGS_REQUEST_2321_sample_completed_
      -- CP-element group 92: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/RPIPE_NOBLOCK_L2_TAGS_REQUEST_2321_Sample/$exit
      -- CP-element group 92: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/RPIPE_NOBLOCK_L2_TAGS_REQUEST_2321_Sample/ra
      -- 
    ra_2562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 92_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_NOBLOCK_L2_TAGS_REQUEST_2321_inst_ack_0, ack => accessL2TagsDaemon_CP_2362_elements(92)); -- 
    -- CP-element group 93:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: successors 
    -- CP-element group 93: marked-successors 
    -- CP-element group 93: 	90 
    -- CP-element group 93:  members (4) 
      -- CP-element group 93: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/RPIPE_NOBLOCK_L2_TAGS_REQUEST_2321_update_completed__ps
      -- CP-element group 93: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/RPIPE_NOBLOCK_L2_TAGS_REQUEST_2321_update_completed_
      -- CP-element group 93: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/RPIPE_NOBLOCK_L2_TAGS_REQUEST_2321_Update/$exit
      -- CP-element group 93: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/RPIPE_NOBLOCK_L2_TAGS_REQUEST_2321_Update/ca
      -- 
    ca_2567_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_NOBLOCK_L2_TAGS_REQUEST_2321_inst_ack_1, ack => accessL2TagsDaemon_CP_2362_elements(93)); -- 
    -- CP-element group 94:  join  transition  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	9 
    -- CP-element group 94: marked-predecessors 
    -- CP-element group 94: 	12 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	11 
    -- CP-element group 94:  members (1) 
      -- CP-element group 94: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2322_sample_start_
      -- 
    accessL2TagsDaemon_cp_element_group_94: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 38) := "accessL2TagsDaemon_cp_element_group_94"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessL2TagsDaemon_CP_2362_elements(9) & accessL2TagsDaemon_CP_2362_elements(12);
      gj_accessL2TagsDaemon_cp_element_group_94 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessL2TagsDaemon_CP_2362_elements(94), clk => clk, reset => reset); --
    end block;
    -- CP-element group 95:  join  transition  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	9 
    -- CP-element group 95: marked-predecessors 
    -- CP-element group 95: 	99 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	14 
    -- CP-element group 95:  members (1) 
      -- CP-element group 95: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2322_update_start_
      -- 
    accessL2TagsDaemon_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "accessL2TagsDaemon_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessL2TagsDaemon_CP_2362_elements(9) & accessL2TagsDaemon_CP_2362_elements(99);
      gj_accessL2TagsDaemon_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessL2TagsDaemon_CP_2362_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	11 
    -- CP-element group 96: successors 
    -- CP-element group 96:  members (1) 
      -- CP-element group 96: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2322_sample_start__ps
      -- 
    accessL2TagsDaemon_CP_2362_elements(96) <= accessL2TagsDaemon_CP_2362_elements(11);
    -- CP-element group 97:  join  transition  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	12 
    -- CP-element group 97:  members (1) 
      -- CP-element group 97: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2322_sample_completed__ps
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(97) is bound as output of CP function.
    -- CP-element group 98:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	14 
    -- CP-element group 98: 	18 
    -- CP-element group 98: successors 
    -- CP-element group 98:  members (1) 
      -- CP-element group 98: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2322_update_start__ps
      -- 
    accessL2TagsDaemon_cp_element_group_98: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 38) := "accessL2TagsDaemon_cp_element_group_98"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessL2TagsDaemon_CP_2362_elements(14) & accessL2TagsDaemon_CP_2362_elements(18);
      gj_accessL2TagsDaemon_cp_element_group_98 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessL2TagsDaemon_CP_2362_elements(98), clk => clk, reset => reset); --
    end block;
    -- CP-element group 99:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	15 
    -- CP-element group 99: marked-successors 
    -- CP-element group 99: 	95 
    -- CP-element group 99:  members (2) 
      -- CP-element group 99: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2322_update_completed_
      -- CP-element group 99: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2322_update_completed__ps
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(99) is bound as output of CP function.
    -- CP-element group 100:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	7 
    -- CP-element group 100: successors 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2322_loopback_trigger
      -- 
    accessL2TagsDaemon_CP_2362_elements(100) <= accessL2TagsDaemon_CP_2362_elements(7);
    -- CP-element group 101:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: successors 
    -- CP-element group 101:  members (2) 
      -- CP-element group 101: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2322_loopback_sample_req
      -- CP-element group 101: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2322_loopback_sample_req_ps
      -- 
    phi_stmt_2322_loopback_sample_req_2578_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2322_loopback_sample_req_2578_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessL2TagsDaemon_CP_2362_elements(101), ack => phi_stmt_2322_req_1); -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(101) is bound as output of CP function.
    -- CP-element group 102:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	8 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (1) 
      -- CP-element group 102: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2322_entry_trigger
      -- 
    accessL2TagsDaemon_CP_2362_elements(102) <= accessL2TagsDaemon_CP_2362_elements(8);
    -- CP-element group 103:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2322_entry_sample_req
      -- CP-element group 103: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2322_entry_sample_req_ps
      -- 
    phi_stmt_2322_entry_sample_req_2581_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_2322_entry_sample_req_2581_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessL2TagsDaemon_CP_2362_elements(103), ack => phi_stmt_2322_req_0); -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(103) is bound as output of CP function.
    -- CP-element group 104:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: successors 
    -- CP-element group 104:  members (2) 
      -- CP-element group 104: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2322_phi_mux_ack
      -- CP-element group 104: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/phi_stmt_2322_phi_mux_ack_ps
      -- 
    phi_stmt_2322_phi_mux_ack_2584_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 104_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_2322_ack_0, ack => accessL2TagsDaemon_CP_2362_elements(104)); -- 
    -- CP-element group 105:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (4) 
      -- CP-element group 105: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/type_cast_2325_sample_start__ps
      -- CP-element group 105: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/type_cast_2325_sample_completed__ps
      -- CP-element group 105: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/type_cast_2325_sample_start_
      -- CP-element group 105: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/type_cast_2325_sample_completed_
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(105) is bound as output of CP function.
    -- CP-element group 106:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	108 
    -- CP-element group 106:  members (2) 
      -- CP-element group 106: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/type_cast_2325_update_start__ps
      -- CP-element group 106: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/type_cast_2325_update_start_
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(106) is bound as output of CP function.
    -- CP-element group 107:  join  transition  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	108 
    -- CP-element group 107: successors 
    -- CP-element group 107:  members (1) 
      -- CP-element group 107: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/type_cast_2325_update_completed__ps
      -- 
    accessL2TagsDaemon_CP_2362_elements(107) <= accessL2TagsDaemon_CP_2362_elements(108);
    -- CP-element group 108:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: 	106 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	107 
    -- CP-element group 108:  members (1) 
      -- CP-element group 108: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/type_cast_2325_update_completed_
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(108) is a control-delay.
    cp_element_108_delay: control_delay_element  generic map(name => " 108_delay", delay_value => 1)  port map(req => accessL2TagsDaemon_CP_2362_elements(106), ack => accessL2TagsDaemon_CP_2362_elements(108), clk => clk, reset =>reset);
    -- CP-element group 109:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: successors 
    -- CP-element group 109:  members (4) 
      -- CP-element group 109: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/type_cast_2327_sample_start__ps
      -- CP-element group 109: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/type_cast_2327_sample_completed__ps
      -- CP-element group 109: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/type_cast_2327_sample_start_
      -- CP-element group 109: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/type_cast_2327_sample_completed_
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(109) is bound as output of CP function.
    -- CP-element group 110:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	112 
    -- CP-element group 110:  members (2) 
      -- CP-element group 110: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/type_cast_2327_update_start__ps
      -- CP-element group 110: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/type_cast_2327_update_start_
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(110) is bound as output of CP function.
    -- CP-element group 111:  join  transition  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	112 
    -- CP-element group 111: successors 
    -- CP-element group 111:  members (1) 
      -- CP-element group 111: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/type_cast_2327_update_completed__ps
      -- 
    accessL2TagsDaemon_CP_2362_elements(111) <= accessL2TagsDaemon_CP_2362_elements(112);
    -- CP-element group 112:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: 	110 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	111 
    -- CP-element group 112:  members (1) 
      -- CP-element group 112: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/type_cast_2327_update_completed_
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(112) is a control-delay.
    cp_element_112_delay: control_delay_element  generic map(name => " 112_delay", delay_value => 1)  port map(req => accessL2TagsDaemon_CP_2362_elements(110), ack => accessL2TagsDaemon_CP_2362_elements(112), clk => clk, reset =>reset);
    -- CP-element group 113:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	19 
    -- CP-element group 113: 	59 
    -- CP-element group 113: 	40 
    -- CP-element group 113: marked-predecessors 
    -- CP-element group 113: 	115 
    -- CP-element group 113: successors 
    -- CP-element group 113: 	114 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/WPIPE_L2_TAGS_RESPONSE_2482_sample_start_
      -- CP-element group 113: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/WPIPE_L2_TAGS_RESPONSE_2482_Sample/$entry
      -- CP-element group 113: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/WPIPE_L2_TAGS_RESPONSE_2482_Sample/req
      -- 
    req_2610_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2610_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessL2TagsDaemon_CP_2362_elements(113), ack => WPIPE_L2_TAGS_RESPONSE_2482_inst_req_0); -- 
    accessL2TagsDaemon_cp_element_group_113: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 39) := "accessL2TagsDaemon_cp_element_group_113"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= accessL2TagsDaemon_CP_2362_elements(19) & accessL2TagsDaemon_CP_2362_elements(59) & accessL2TagsDaemon_CP_2362_elements(40) & accessL2TagsDaemon_CP_2362_elements(115);
      gj_accessL2TagsDaemon_cp_element_group_113 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessL2TagsDaemon_CP_2362_elements(113), clk => clk, reset => reset); --
    end block;
    -- CP-element group 114:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	113 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	115 
    -- CP-element group 114: marked-successors 
    -- CP-element group 114: 	17 
    -- CP-element group 114: 	55 
    -- CP-element group 114: 	36 
    -- CP-element group 114:  members (6) 
      -- CP-element group 114: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/WPIPE_L2_TAGS_RESPONSE_2482_sample_completed_
      -- CP-element group 114: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/WPIPE_L2_TAGS_RESPONSE_2482_update_start_
      -- CP-element group 114: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/WPIPE_L2_TAGS_RESPONSE_2482_Sample/$exit
      -- CP-element group 114: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/WPIPE_L2_TAGS_RESPONSE_2482_Sample/ack
      -- CP-element group 114: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/WPIPE_L2_TAGS_RESPONSE_2482_Update/$entry
      -- CP-element group 114: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/WPIPE_L2_TAGS_RESPONSE_2482_Update/req
      -- 
    ack_2611_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_L2_TAGS_RESPONSE_2482_inst_ack_0, ack => accessL2TagsDaemon_CP_2362_elements(114)); -- 
    req_2615_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2615_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessL2TagsDaemon_CP_2362_elements(114), ack => WPIPE_L2_TAGS_RESPONSE_2482_inst_req_1); -- 
    -- CP-element group 115:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	114 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115: marked-successors 
    -- CP-element group 115: 	113 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/WPIPE_L2_TAGS_RESPONSE_2482_update_completed_
      -- CP-element group 115: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/WPIPE_L2_TAGS_RESPONSE_2482_Update/$exit
      -- CP-element group 115: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/WPIPE_L2_TAGS_RESPONSE_2482_Update/ack
      -- 
    ack_2616_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 115_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_L2_TAGS_RESPONSE_2482_inst_ack_1, ack => accessL2TagsDaemon_CP_2362_elements(115)); -- 
    -- CP-element group 116:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: 	9 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	10 
    -- CP-element group 116:  members (1) 
      -- CP-element group 116: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group accessL2TagsDaemon_CP_2362_elements(116) is a control-delay.
    cp_element_116_delay: control_delay_element  generic map(name => " 116_delay", delay_value => 1)  port map(req => accessL2TagsDaemon_CP_2362_elements(9), ack => accessL2TagsDaemon_CP_2362_elements(116), clk => clk, reset =>reset);
    -- CP-element group 117:  join  transition  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	12 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117: 	6 
    -- CP-element group 117:  members (1) 
      -- CP-element group 117: 	 branch_block_stmt_2290/do_while_stmt_2291/do_while_stmt_2291_loop_body/$exit
      -- 
    accessL2TagsDaemon_cp_element_group_117: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 39) := "accessL2TagsDaemon_cp_element_group_117"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessL2TagsDaemon_CP_2362_elements(12) & accessL2TagsDaemon_CP_2362_elements(115);
      gj_accessL2TagsDaemon_cp_element_group_117 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessL2TagsDaemon_CP_2362_elements(117), clk => clk, reset => reset); --
    end block;
    -- CP-element group 118:  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	5 
    -- CP-element group 118: successors 
    -- CP-element group 118:  members (2) 
      -- CP-element group 118: 	 branch_block_stmt_2290/do_while_stmt_2291/loop_exit/$exit
      -- CP-element group 118: 	 branch_block_stmt_2290/do_while_stmt_2291/loop_exit/ack
      -- 
    ack_2621_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2291_branch_ack_0, ack => accessL2TagsDaemon_CP_2362_elements(118)); -- 
    -- CP-element group 119:  transition  input  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	5 
    -- CP-element group 119: successors 
    -- CP-element group 119:  members (2) 
      -- CP-element group 119: 	 branch_block_stmt_2290/do_while_stmt_2291/loop_taken/$exit
      -- CP-element group 119: 	 branch_block_stmt_2290/do_while_stmt_2291/loop_taken/ack
      -- 
    ack_2625_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 119_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_2291_branch_ack_1, ack => accessL2TagsDaemon_CP_2362_elements(119)); -- 
    -- CP-element group 120:  transition  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: 	3 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	1 
    -- CP-element group 120:  members (1) 
      -- CP-element group 120: 	 branch_block_stmt_2290/do_while_stmt_2291/$exit
      -- 
    accessL2TagsDaemon_CP_2362_elements(120) <= accessL2TagsDaemon_CP_2362_elements(3);
    accessL2TagsDaemon_do_while_stmt_2291_terminator_2626: loop_terminator -- 
      generic map (name => " accessL2TagsDaemon_do_while_stmt_2291_terminator_2626", max_iterations_in_flight =>15) 
      port map(loop_body_exit => accessL2TagsDaemon_CP_2362_elements(6),loop_continue => accessL2TagsDaemon_CP_2362_elements(119),loop_terminate => accessL2TagsDaemon_CP_2362_elements(118),loop_back => accessL2TagsDaemon_CP_2362_elements(4),loop_exit => accessL2TagsDaemon_CP_2362_elements(3),clk => clk, reset => reset); -- 
    phi_stmt_2293_phi_seq_2436_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= accessL2TagsDaemon_CP_2362_elements(22);
      accessL2TagsDaemon_CP_2362_elements(25)<= src_sample_reqs(0);
      src_sample_acks(0)  <= accessL2TagsDaemon_CP_2362_elements(25);
      accessL2TagsDaemon_CP_2362_elements(26)<= src_update_reqs(0);
      src_update_acks(0)  <= accessL2TagsDaemon_CP_2362_elements(27);
      accessL2TagsDaemon_CP_2362_elements(23) <= phi_mux_reqs(0);
      triggers(1)  <= accessL2TagsDaemon_CP_2362_elements(20);
      accessL2TagsDaemon_CP_2362_elements(29)<= src_sample_reqs(1);
      src_sample_acks(1)  <= accessL2TagsDaemon_CP_2362_elements(33);
      accessL2TagsDaemon_CP_2362_elements(30)<= src_update_reqs(1);
      src_update_acks(1)  <= accessL2TagsDaemon_CP_2362_elements(34);
      accessL2TagsDaemon_CP_2362_elements(21) <= phi_mux_reqs(1);
      phi_stmt_2293_phi_seq_2436 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2293_phi_seq_2436") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => accessL2TagsDaemon_CP_2362_elements(11), 
          phi_sample_ack => accessL2TagsDaemon_CP_2362_elements(18), 
          phi_update_req => accessL2TagsDaemon_CP_2362_elements(14), 
          phi_update_ack => accessL2TagsDaemon_CP_2362_elements(19), 
          phi_mux_ack => accessL2TagsDaemon_CP_2362_elements(24), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2310_phi_seq_2480_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= accessL2TagsDaemon_CP_2362_elements(41);
      accessL2TagsDaemon_CP_2362_elements(46)<= src_sample_reqs(0);
      src_sample_acks(0)  <= accessL2TagsDaemon_CP_2362_elements(48);
      accessL2TagsDaemon_CP_2362_elements(47)<= src_update_reqs(0);
      src_update_acks(0)  <= accessL2TagsDaemon_CP_2362_elements(49);
      accessL2TagsDaemon_CP_2362_elements(42) <= phi_mux_reqs(0);
      triggers(1)  <= accessL2TagsDaemon_CP_2362_elements(43);
      accessL2TagsDaemon_CP_2362_elements(50)<= src_sample_reqs(1);
      src_sample_acks(1)  <= accessL2TagsDaemon_CP_2362_elements(50);
      accessL2TagsDaemon_CP_2362_elements(51)<= src_update_reqs(1);
      src_update_acks(1)  <= accessL2TagsDaemon_CP_2362_elements(52);
      accessL2TagsDaemon_CP_2362_elements(44) <= phi_mux_reqs(1);
      phi_stmt_2310_phi_seq_2480 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2310_phi_seq_2480") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => accessL2TagsDaemon_CP_2362_elements(37), 
          phi_sample_ack => accessL2TagsDaemon_CP_2362_elements(38), 
          phi_update_req => accessL2TagsDaemon_CP_2362_elements(39), 
          phi_update_ack => accessL2TagsDaemon_CP_2362_elements(40), 
          phi_mux_ack => accessL2TagsDaemon_CP_2362_elements(45), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2314_phi_seq_2524_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= accessL2TagsDaemon_CP_2362_elements(60);
      accessL2TagsDaemon_CP_2362_elements(65)<= src_sample_reqs(0);
      src_sample_acks(0)  <= accessL2TagsDaemon_CP_2362_elements(67);
      accessL2TagsDaemon_CP_2362_elements(66)<= src_update_reqs(0);
      src_update_acks(0)  <= accessL2TagsDaemon_CP_2362_elements(68);
      accessL2TagsDaemon_CP_2362_elements(61) <= phi_mux_reqs(0);
      triggers(1)  <= accessL2TagsDaemon_CP_2362_elements(62);
      accessL2TagsDaemon_CP_2362_elements(69)<= src_sample_reqs(1);
      src_sample_acks(1)  <= accessL2TagsDaemon_CP_2362_elements(69);
      accessL2TagsDaemon_CP_2362_elements(70)<= src_update_reqs(1);
      src_update_acks(1)  <= accessL2TagsDaemon_CP_2362_elements(71);
      accessL2TagsDaemon_CP_2362_elements(63) <= phi_mux_reqs(1);
      phi_stmt_2314_phi_seq_2524 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2314_phi_seq_2524") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => accessL2TagsDaemon_CP_2362_elements(56), 
          phi_sample_ack => accessL2TagsDaemon_CP_2362_elements(57), 
          phi_update_req => accessL2TagsDaemon_CP_2362_elements(58), 
          phi_update_ack => accessL2TagsDaemon_CP_2362_elements(59), 
          phi_mux_ack => accessL2TagsDaemon_CP_2362_elements(64), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2318_phi_seq_2568_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= accessL2TagsDaemon_CP_2362_elements(81);
      accessL2TagsDaemon_CP_2362_elements(84)<= src_sample_reqs(0);
      src_sample_acks(0)  <= accessL2TagsDaemon_CP_2362_elements(84);
      accessL2TagsDaemon_CP_2362_elements(85)<= src_update_reqs(0);
      src_update_acks(0)  <= accessL2TagsDaemon_CP_2362_elements(86);
      accessL2TagsDaemon_CP_2362_elements(82) <= phi_mux_reqs(0);
      triggers(1)  <= accessL2TagsDaemon_CP_2362_elements(79);
      accessL2TagsDaemon_CP_2362_elements(88)<= src_sample_reqs(1);
      src_sample_acks(1)  <= accessL2TagsDaemon_CP_2362_elements(92);
      accessL2TagsDaemon_CP_2362_elements(89)<= src_update_reqs(1);
      src_update_acks(1)  <= accessL2TagsDaemon_CP_2362_elements(93);
      accessL2TagsDaemon_CP_2362_elements(80) <= phi_mux_reqs(1);
      phi_stmt_2318_phi_seq_2568 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2318_phi_seq_2568") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => accessL2TagsDaemon_CP_2362_elements(75), 
          phi_sample_ack => accessL2TagsDaemon_CP_2362_elements(76), 
          phi_update_req => accessL2TagsDaemon_CP_2362_elements(77), 
          phi_update_ack => accessL2TagsDaemon_CP_2362_elements(78), 
          phi_mux_ack => accessL2TagsDaemon_CP_2362_elements(83), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_2322_phi_seq_2602_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= accessL2TagsDaemon_CP_2362_elements(102);
      accessL2TagsDaemon_CP_2362_elements(105)<= src_sample_reqs(0);
      src_sample_acks(0)  <= accessL2TagsDaemon_CP_2362_elements(105);
      accessL2TagsDaemon_CP_2362_elements(106)<= src_update_reqs(0);
      src_update_acks(0)  <= accessL2TagsDaemon_CP_2362_elements(107);
      accessL2TagsDaemon_CP_2362_elements(103) <= phi_mux_reqs(0);
      triggers(1)  <= accessL2TagsDaemon_CP_2362_elements(100);
      accessL2TagsDaemon_CP_2362_elements(109)<= src_sample_reqs(1);
      src_sample_acks(1)  <= accessL2TagsDaemon_CP_2362_elements(109);
      accessL2TagsDaemon_CP_2362_elements(110)<= src_update_reqs(1);
      src_update_acks(1)  <= accessL2TagsDaemon_CP_2362_elements(111);
      accessL2TagsDaemon_CP_2362_elements(101) <= phi_mux_reqs(1);
      phi_stmt_2322_phi_seq_2602 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_2322_phi_seq_2602") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => accessL2TagsDaemon_CP_2362_elements(96), 
          phi_sample_ack => accessL2TagsDaemon_CP_2362_elements(97), 
          phi_update_req => accessL2TagsDaemon_CP_2362_elements(98), 
          phi_update_ack => accessL2TagsDaemon_CP_2362_elements(99), 
          phi_mux_ack => accessL2TagsDaemon_CP_2362_elements(104), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_2387_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= accessL2TagsDaemon_CP_2362_elements(7);
        preds(1)  <= accessL2TagsDaemon_CP_2362_elements(8);
        entry_tmerge_2387 : transition_merge -- 
          generic map(name => " entry_tmerge_2387")
          port map (preds => preds, symbol_out => accessL2TagsDaemon_CP_2362_elements(9));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u3_u3_2496_wire : std_logic_vector(2 downto 0);
    signal AND_u1_u1_2555_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_2560_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u1_u22_2478_wire : std_logic_vector(21 downto 0);
    signal CONCAT_u1_u9_2473_wire : std_logic_vector(8 downto 0);
    signal CONCAT_u9_u12_2475_wire : std_logic_vector(11 downto 0);
    signal MUX_2498_wire : std_logic_vector(2 downto 0);
    signal NOT_u1_u1_2493_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_2520_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_2543_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_2545_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_2557_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_2559_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_2572_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_2575_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_2576_wire : std_logic_vector(0 downto 0);
    signal RPIPE_NOBLOCK_L2_TAGS_REQUEST_2321_wire : std_logic_vector(44 downto 0);
    signal access_index_in_set_d_2458 : std_logic_vector(2 downto 0);
    signal call_accessL2TagMemX4096X8_expr_2309_wire : std_logic_vector(242 downto 0);
    signal call_insertIntoSetDirtyDwordMasks_expr_2539_wire : std_logic_vector(63 downto 0);
    signal current_dirty_dword_mask_d_2458 : std_logic_vector(7 downto 0);
    signal dirty_bits_have_been_modified_d_2567 : std_logic_vector(0 downto 0);
    signal init_2322 : std_logic_vector(0 downto 0);
    signal is_hit_d_2458 : std_logic_vector(0 downto 0);
    signal konst_2295_wire_constant : std_logic_vector(242 downto 0);
    signal konst_2313_wire_constant : std_logic_vector(0 downto 0);
    signal konst_2317_wire_constant : std_logic_vector(44 downto 0);
    signal konst_2320_wire_constant : std_logic_vector(44 downto 0);
    signal konst_2335_wire_constant : std_logic_vector(242 downto 0);
    signal konst_2495_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2592_wire_constant : std_logic_vector(0 downto 0);
    signal lwi_has_been_modified_d_2551 : std_logic_vector(0 downto 0);
    signal n_request_d_2331 : std_logic_vector(44 downto 0);
    signal n_request_d_2331_2316_buffered : std_logic_vector(44 downto 0);
    signal next_free_index_on_hit_d_2488 : std_logic_vector(2 downto 0);
    signal read_lwi_d_2439 : std_logic_vector(2 downto 0);
    signal read_set_dirty_dword_masks_d_2447 : std_logic_vector(63 downto 0);
    signal read_set_id_2425 : std_logic_vector(8 downto 0);
    signal read_set_tags_d_2435 : std_logic_vector(167 downto 0);
    signal read_set_valids_d_2443 : std_logic_vector(7 downto 0);
    signal read_write_access_d_2522 : std_logic_vector(0 downto 0);
    signal replace_line_is_valid_d_2458 : std_logic_vector(0 downto 0);
    signal replace_pa_tag_d_2458 : std_logic_vector(20 downto 0);
    signal request_2318 : std_logic_vector(44 downto 0);
    signal request_allocate_on_miss_2369 : std_logic_vector(0 downto 0);
    signal request_allocate_on_miss_d_2410 : std_logic_vector(0 downto 0);
    signal request_counter_2345 : std_logic_vector(7 downto 0);
    signal request_counter_d_2386 : std_logic_vector(7 downto 0);
    signal request_d_2314 : std_logic_vector(44 downto 0);
    signal request_invalidate_2349 : std_logic_vector(0 downto 0);
    signal request_invalidate_d_2390 : std_logic_vector(0 downto 0);
    signal request_pa_dword_id_2361 : std_logic_vector(2 downto 0);
    signal request_pa_dword_id_d_2402 : std_logic_vector(2 downto 0);
    signal request_pa_tag_2357 : std_logic_vector(20 downto 0);
    signal request_pa_tag_d_2398 : std_logic_vector(20 downto 0);
    signal request_rwbar_2353 : std_logic_vector(0 downto 0);
    signal request_rwbar_d_2394 : std_logic_vector(0 downto 0);
    signal request_set_id_2365 : std_logic_vector(8 downto 0);
    signal request_set_id_d_2406 : std_logic_vector(8 downto 0);
    signal request_valid_2341 : std_logic_vector(0 downto 0);
    signal request_valid_d_2382 : std_logic_vector(0 downto 0);
    signal response_d_2480 : std_logic_vector(33 downto 0);
    signal tag_mem_read_2422 : std_logic_vector(0 downto 0);
    signal tag_mem_read_2422_2312_buffered : std_logic_vector(0 downto 0);
    signal tag_mem_read_d_2310 : std_logic_vector(0 downto 0);
    signal tag_mem_response_d_2337 : std_logic_vector(242 downto 0);
    signal tag_mem_response_raw_2293 : std_logic_vector(242 downto 0);
    signal tag_mem_write_d_2578 : std_logic_vector(0 downto 0);
    signal tags_have_been_modified_d_2547 : std_logic_vector(0 downto 0);
    signal type_cast_2325_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_2327_wire_constant : std_logic_vector(0 downto 0);
    signal updated_dirty_dword_mask_d_2516 : std_logic_vector(7 downto 0);
    signal updated_set_dirty_dword_masks_d_2540 : std_logic_vector(63 downto 0);
    signal updated_set_lwi_d_2500 : std_logic_vector(2 downto 0);
    signal updated_set_tags_d_2534 : std_logic_vector(167 downto 0);
    signal updated_set_valids_d_2528 : std_logic_vector(7 downto 0);
    signal valids_have_been_modified_d_2562 : std_logic_vector(0 downto 0);
    signal write_set_id_d_2581 : std_logic_vector(8 downto 0);
    -- 
  begin -- 
    konst_2295_wire_constant <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    konst_2313_wire_constant <= "0";
    konst_2317_wire_constant <= "000000000000000000000000000000000000000000000";
    konst_2320_wire_constant <= "000000000000000000000000000000000000000000000";
    konst_2335_wire_constant <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    konst_2495_wire_constant <= "001";
    konst_2592_wire_constant <= "1";
    type_cast_2325_wire_constant <= "1";
    type_cast_2327_wire_constant <= "0";
    phi_stmt_2293: Block -- phi operator 
      signal idata: std_logic_vector(485 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= konst_2295_wire_constant & call_accessL2TagMemX4096X8_expr_2309_wire;
      req <= phi_stmt_2293_req_0 & phi_stmt_2293_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2293",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 243) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2293_ack_0,
          idata => idata,
          odata => tag_mem_response_raw_2293,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2293
    phi_stmt_2310: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= tag_mem_read_2422_2312_buffered & konst_2313_wire_constant;
      req <= phi_stmt_2310_req_0 & phi_stmt_2310_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2310",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2310_ack_0,
          idata => idata,
          odata => tag_mem_read_d_2310,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2310
    phi_stmt_2314: Block -- phi operator 
      signal idata: std_logic_vector(89 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_request_d_2331_2316_buffered & konst_2317_wire_constant;
      req <= phi_stmt_2314_req_0 & phi_stmt_2314_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2314",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 45) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2314_ack_0,
          idata => idata,
          odata => request_d_2314,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2314
    phi_stmt_2318: Block -- phi operator 
      signal idata: std_logic_vector(89 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= konst_2320_wire_constant & RPIPE_NOBLOCK_L2_TAGS_REQUEST_2321_wire;
      req <= phi_stmt_2318_req_0 & phi_stmt_2318_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2318",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 45) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2318_ack_0,
          idata => idata,
          odata => request_2318,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2318
    phi_stmt_2322: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_2325_wire_constant & type_cast_2327_wire_constant;
      req <= phi_stmt_2322_req_0 & phi_stmt_2322_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_2322",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_2322_ack_0,
          idata => idata,
          odata => init_2322,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_2322
    -- flow-through select operator MUX_2336_inst
    tag_mem_response_d_2337 <= tag_mem_response_raw_2293 when (tag_mem_read_d_2310(0) /=  '0') else konst_2335_wire_constant;
    -- flow-through select operator MUX_2498_inst
    MUX_2498_wire <= ADD_u3_u3_2496_wire when (NOT_u1_u1_2493_wire(0) /=  '0') else read_lwi_d_2439;
    -- flow-through select operator MUX_2499_inst
    updated_set_lwi_d_2500 <= next_free_index_on_hit_d_2488 when (is_hit_d_2458(0) /=  '0') else MUX_2498_wire;
    -- flow-through slice operator slice_2340_inst
    request_valid_2341 <= request_2318(44 downto 44);
    -- flow-through slice operator slice_2344_inst
    request_counter_2345 <= request_2318(43 downto 36);
    -- flow-through slice operator slice_2348_inst
    request_invalidate_2349 <= request_2318(35 downto 35);
    -- flow-through slice operator slice_2352_inst
    request_rwbar_2353 <= request_2318(34 downto 34);
    -- flow-through slice operator slice_2356_inst
    request_pa_tag_2357 <= request_2318(33 downto 13);
    -- flow-through slice operator slice_2360_inst
    request_pa_dword_id_2361 <= request_2318(12 downto 10);
    -- flow-through slice operator slice_2364_inst
    request_set_id_2365 <= request_2318(9 downto 1);
    -- flow-through slice operator slice_2368_inst
    request_allocate_on_miss_2369 <= request_2318(0 downto 0);
    -- flow-through slice operator slice_2381_inst
    request_valid_d_2382 <= request_d_2314(44 downto 44);
    -- flow-through slice operator slice_2385_inst
    request_counter_d_2386 <= request_d_2314(43 downto 36);
    -- flow-through slice operator slice_2389_inst
    request_invalidate_d_2390 <= request_d_2314(35 downto 35);
    -- flow-through slice operator slice_2393_inst
    request_rwbar_d_2394 <= request_d_2314(34 downto 34);
    -- flow-through slice operator slice_2397_inst
    request_pa_tag_d_2398 <= request_d_2314(33 downto 13);
    -- flow-through slice operator slice_2401_inst
    request_pa_dword_id_d_2402 <= request_d_2314(12 downto 10);
    -- flow-through slice operator slice_2405_inst
    request_set_id_d_2406 <= request_d_2314(9 downto 1);
    -- flow-through slice operator slice_2409_inst
    request_allocate_on_miss_d_2410 <= request_d_2314(0 downto 0);
    -- flow-through slice operator slice_2434_inst
    read_set_tags_d_2435 <= tag_mem_response_d_2337(242 downto 75);
    -- flow-through slice operator slice_2438_inst
    read_lwi_d_2439 <= tag_mem_response_d_2337(74 downto 72);
    -- flow-through slice operator slice_2442_inst
    read_set_valids_d_2443 <= tag_mem_response_d_2337(71 downto 64);
    -- flow-through slice operator slice_2446_inst
    read_set_dirty_dword_masks_d_2447 <= tag_mem_response_d_2337(63 downto 0);
    -- interlock W_n_request_d_2329_inst
    process(request_2318) -- 
      variable tmp_var : std_logic_vector(44 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 44 downto 0) := request_2318(44 downto 0);
      n_request_d_2331 <= tmp_var; -- 
    end process;
    -- interlock W_read_set_id_2423_inst
    process(request_set_id_2365) -- 
      variable tmp_var : std_logic_vector(8 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 8 downto 0) := request_set_id_2365(8 downto 0);
      read_set_id_2425 <= tmp_var; -- 
    end process;
    -- interlock W_tag_mem_read_2420_inst
    process(request_valid_2341) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := request_valid_2341(0 downto 0);
      tag_mem_read_2422 <= tmp_var; -- 
    end process;
    -- interlock W_updated_set_dirty_dword_masks_d_2535_inst
    process(call_insertIntoSetDirtyDwordMasks_expr_2539_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 63 downto 0) := call_insertIntoSetDirtyDwordMasks_expr_2539_wire(63 downto 0);
      updated_set_dirty_dword_masks_d_2540 <= tmp_var; -- 
    end process;
    -- interlock W_write_set_id_d_2579_inst
    process(request_set_id_d_2406) -- 
      variable tmp_var : std_logic_vector(8 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 8 downto 0) := request_set_id_d_2406(8 downto 0);
      write_set_id_d_2581 <= tmp_var; -- 
    end process;
    n_request_d_2331_2316_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_request_d_2331_2316_buf_req_0;
      n_request_d_2331_2316_buf_ack_0<= wack(0);
      rreq(0) <= n_request_d_2331_2316_buf_req_1;
      n_request_d_2331_2316_buf_ack_1<= rack(0);
      n_request_d_2331_2316_buf : InterlockBuffer generic map ( -- 
        name => "n_request_d_2331_2316_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 45,
        out_data_width => 45,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_request_d_2331,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_request_d_2331_2316_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    tag_mem_read_2422_2312_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= tag_mem_read_2422_2312_buf_req_0;
      tag_mem_read_2422_2312_buf_ack_0<= wack(0);
      rreq(0) <= tag_mem_read_2422_2312_buf_req_1;
      tag_mem_read_2422_2312_buf_ack_1<= rack(0);
      tag_mem_read_2422_2312_buf : InterlockBuffer generic map ( -- 
        name => "tag_mem_read_2422_2312_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => tag_mem_read_2422,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => tag_mem_read_2422_2312_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_2291_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_2592_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_2291_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_2291_branch_req_0,
          ack0 => do_while_stmt_2291_branch_ack_0,
          ack1 => do_while_stmt_2291_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u3_u3_2496_inst
    process(read_lwi_d_2439) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApIntAdd_proc(read_lwi_d_2439, konst_2495_wire_constant, tmp_var);
      ADD_u3_u3_2496_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2521_inst
    process(request_valid_d_2382, NOT_u1_u1_2520_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(request_valid_d_2382, NOT_u1_u1_2520_wire, tmp_var);
      read_write_access_d_2522 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2546_inst
    process(NOT_u1_u1_2543_wire, NOT_u1_u1_2545_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_2543_wire, NOT_u1_u1_2545_wire, tmp_var);
      tags_have_been_modified_d_2547 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2555_inst
    process(request_invalidate_d_2390, is_hit_d_2458) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(request_invalidate_d_2390, is_hit_d_2458, tmp_var);
      AND_u1_u1_2555_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2560_inst
    process(NOT_u1_u1_2557_wire, NOT_u1_u1_2559_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_2557_wire, NOT_u1_u1_2559_wire, tmp_var);
      AND_u1_u1_2560_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2577_inst
    process(tag_mem_read_d_2310, OR_u1_u1_2576_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(tag_mem_read_d_2310, OR_u1_u1_2576_wire, tmp_var);
      tag_mem_write_d_2578 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u12_u34_2479_inst
    process(CONCAT_u9_u12_2475_wire, CONCAT_u1_u22_2478_wire) -- 
      variable tmp_var : std_logic_vector(33 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u9_u12_2475_wire, CONCAT_u1_u22_2478_wire, tmp_var);
      response_d_2480 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u22_2478_inst
    process(replace_line_is_valid_d_2458, replace_pa_tag_d_2458) -- 
      variable tmp_var : std_logic_vector(21 downto 0); -- 
    begin -- 
      ApConcat_proc(replace_line_is_valid_d_2458, replace_pa_tag_d_2458, tmp_var);
      CONCAT_u1_u22_2478_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u9_2473_inst
    process(is_hit_d_2458, current_dirty_dword_mask_d_2458) -- 
      variable tmp_var : std_logic_vector(8 downto 0); -- 
    begin -- 
      ApConcat_proc(is_hit_d_2458, current_dirty_dword_mask_d_2458, tmp_var);
      CONCAT_u1_u9_2473_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u9_u12_2475_inst
    process(CONCAT_u1_u9_2473_wire, access_index_in_set_d_2458) -- 
      variable tmp_var : std_logic_vector(11 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u9_2473_wire, access_index_in_set_d_2458, tmp_var);
      CONCAT_u9_u12_2475_wire <= tmp_var; --
    end process;
    -- binary operator NEQ_u8_u1_2566_inst
    process(current_dirty_dword_mask_d_2458, updated_dirty_dword_mask_d_2516) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(current_dirty_dword_mask_d_2458, updated_dirty_dword_mask_d_2516, tmp_var);
      dirty_bits_have_been_modified_d_2567 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_2493_inst
    process(request_invalidate_d_2390) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", request_invalidate_d_2390, tmp_var);
      NOT_u1_u1_2493_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_2520_inst
    process(request_invalidate_d_2390) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", request_invalidate_d_2390, tmp_var);
      NOT_u1_u1_2520_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_2543_inst
    process(request_invalidate_d_2390) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", request_invalidate_d_2390, tmp_var);
      NOT_u1_u1_2543_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_2545_inst
    process(is_hit_d_2458) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", is_hit_d_2458, tmp_var);
      NOT_u1_u1_2545_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_2550_inst
    process(request_invalidate_d_2390) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", request_invalidate_d_2390, tmp_var);
      lwi_has_been_modified_d_2551 <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_2557_inst
    process(request_invalidate_d_2390) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", request_invalidate_d_2390, tmp_var);
      NOT_u1_u1_2557_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_2559_inst
    process(is_hit_d_2458) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", is_hit_d_2458, tmp_var);
      NOT_u1_u1_2559_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_2561_inst
    process(AND_u1_u1_2555_wire, AND_u1_u1_2560_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_2555_wire, AND_u1_u1_2560_wire, tmp_var);
      valids_have_been_modified_d_2562 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_2572_inst
    process(tags_have_been_modified_d_2547, lwi_has_been_modified_d_2551) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(tags_have_been_modified_d_2547, lwi_has_been_modified_d_2551, tmp_var);
      OR_u1_u1_2572_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_2575_inst
    process(valids_have_been_modified_d_2562, dirty_bits_have_been_modified_d_2567) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(valids_have_been_modified_d_2562, dirty_bits_have_been_modified_d_2567, tmp_var);
      OR_u1_u1_2575_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_2576_inst
    process(OR_u1_u1_2572_wire, OR_u1_u1_2575_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_2572_wire, OR_u1_u1_2575_wire, tmp_var);
      OR_u1_u1_2576_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_NOBLOCK_L2_TAGS_REQUEST_2321_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(44 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_NOBLOCK_L2_TAGS_REQUEST_2321_inst_req_0;
      RPIPE_NOBLOCK_L2_TAGS_REQUEST_2321_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_NOBLOCK_L2_TAGS_REQUEST_2321_inst_req_1;
      RPIPE_NOBLOCK_L2_TAGS_REQUEST_2321_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_NOBLOCK_L2_TAGS_REQUEST_2321_wire <= data_out(44 downto 0);
      NOBLOCK_L2_TAGS_REQUEST_read_0_gI: SplitGuardInterface generic map(name => "NOBLOCK_L2_TAGS_REQUEST_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      NOBLOCK_L2_TAGS_REQUEST_read_0: InputPort_P2P -- 
        generic map ( name => "NOBLOCK_L2_TAGS_REQUEST_read_0", data_width => 45,    bypass_flag => true,   	nonblocking_read_flag => true,  barrier_flag => false,   queue_depth =>  2)
        port map (-- 
          sample_req => reqL(0) , 
          sample_ack => ackL(0), 
          update_req => reqR(0), 
          update_ack => ackR(0), 
          data => data_out, 
          oreq => NOBLOCK_L2_TAGS_REQUEST_pipe_read_req(0),
          oack => NOBLOCK_L2_TAGS_REQUEST_pipe_read_ack(0),
          odata => NOBLOCK_L2_TAGS_REQUEST_pipe_read_data(44 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_L2_TAGS_RESPONSE_2482_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(33 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_L2_TAGS_RESPONSE_2482_inst_req_0;
      WPIPE_L2_TAGS_RESPONSE_2482_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_L2_TAGS_RESPONSE_2482_inst_req_1;
      WPIPE_L2_TAGS_RESPONSE_2482_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= tag_mem_read_d_2310(0);
      data_in <= response_d_2480;
      L2_TAGS_RESPONSE_write_0_gI: SplitGuardInterface generic map(name => "L2_TAGS_RESPONSE_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      L2_TAGS_RESPONSE_write_0: OutputPortRevised -- 
        generic map ( name => "L2_TAGS_RESPONSE", data_width => 34, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => L2_TAGS_RESPONSE_pipe_write_req(0),
          oack => L2_TAGS_RESPONSE_pipe_write_ack(0),
          odata => L2_TAGS_RESPONSE_pipe_write_data(33 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    operator_accessL2TagMemX4096X8_4866_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      sample_req(0) <= call_accessL2TagMemX4096X8_expr_2309_inst_req_0;
      call_accessL2TagMemX4096X8_expr_2309_inst_ack_0<= sample_ack(0);
      update_req(0) <= call_accessL2TagMemX4096X8_expr_2309_inst_req_1;
      call_accessL2TagMemX4096X8_expr_2309_inst_ack_1<= update_ack(0);
      call_accessL2TagMemX4096X8_expr_2309_inst: accessL2TagMemX4096X8_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        init_flag => init_2322,
        tag_mem_read => tag_mem_read_2422,
        tag_mem_write => tag_mem_write_d_2578,
        read_set_id => read_set_id_2425,
        write_set_id => write_set_id_d_2581,
        tags_have_been_modified => tags_have_been_modified_d_2547,
        lwi_has_been_modified => lwi_has_been_modified_d_2551,
        valids_have_been_modified => valids_have_been_modified_d_2562,
        dirty_bits_have_been_modified => dirty_bits_have_been_modified_d_2567,
        updated_set_tags => updated_set_tags_d_2534,
        updated_set_lwi => updated_set_lwi_d_2500,
        updated_set_valids => updated_set_valids_d_2528,
        updated_set_dirty_dword_masks => updated_set_dirty_dword_masks_d_2540,
        tag_mem_response => call_accessL2TagMemX4096X8_expr_2309_wire,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    volatile_operator_insertIntoSetDirtyDwordMasks_4916: insertIntoSetDirtyDwordMasks_Volatile port map(old_set_mask => read_set_dirty_dword_masks_d_2447, index => access_index_in_set_d_2458, ins_mask => updated_dirty_dword_mask_d_2516, new_set_mask => call_insertIntoSetDirtyDwordMasks_expr_2539_wire); 
    volatile_operator_calculateHits_4899: calculateHits_Volatile port map(set_valids => read_set_valids_d_2443, set_dirty_dword_masks => read_set_dirty_dword_masks_d_2447, set_tags => read_set_tags_d_2435, pa_tag => request_pa_tag_d_2398, replace_index => read_lwi_d_2439, is_hit => is_hit_d_2458, dirty_dword_mask => current_dirty_dword_mask_d_2458, access_index => access_index_in_set_d_2458, replace_line_is_valid => replace_line_is_valid_d_2458, replace_pa_tag => replace_pa_tag_d_2458); 
    volatile_operator_nextFreeIndex_4905: nextFreeIndex_Volatile port map(from_index => access_index_in_set_d_2458, set_valids => read_set_valids_d_2443, next_free_index => next_free_index_on_hit_d_2488); 
    volatile_operator_updateDirtyWordMask_4910: updateDirtyWordMask_Volatile port map(invalidate => request_invalidate_d_2390, read_write_access => tag_mem_read_d_2310, is_hit => is_hit_d_2458, rwbar => request_rwbar_d_2394, dword_id => request_pa_dword_id_d_2402, current_dirty_mask => current_dirty_dword_mask_d_2458, updated_dirty_mask => updated_dirty_dword_mask_d_2516); 
    volatile_operator_updateSetValids_4913: updateSetValids_Volatile port map(invalidate => request_invalidate_d_2390, read_write_access => read_write_access_d_2522, set_valids => read_set_valids_d_2443, access_index => access_index_in_set_d_2458, updated_set_valids => updated_set_valids_d_2528); 
    volatile_operator_updateSetTags_4914: updateSetTags_Volatile port map(read_write_access => read_write_access_d_2522, access_index => access_index_in_set_d_2458, pa_tag => request_pa_tag_d_2398, set_tags => read_set_tags_d_2435, updated_set_tags => updated_set_tags_d_2534); 
    -- 
  end Block; -- data_path
  -- 
end accessL2TagsDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library l2_cache_lib;
use l2_cache_lib.l2_cache_global_package.all;
entity accessSysMem is -- 
  generic (tag_length : integer); 
  port ( -- 
    rwbar : in  std_logic_vector(0 downto 0);
    byte_mask : in  std_logic_vector(7 downto 0);
    addr : in  std_logic_vector(35 downto 0);
    wdata : in  std_logic_vector(63 downto 0);
    rdata : out  std_logic_vector(63 downto 0);
    MEM_TO_L2CACHE_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
    MEM_TO_L2CACHE_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
    MEM_TO_L2CACHE_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
    L2CACHE_TO_MEM_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
    L2CACHE_TO_MEM_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
    L2CACHE_TO_MEM_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity accessSysMem;
architecture accessSysMem_arch of accessSysMem is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 109)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 64)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal rwbar_buffer :  std_logic_vector(0 downto 0);
  signal rwbar_update_enable: Boolean;
  signal byte_mask_buffer :  std_logic_vector(7 downto 0);
  signal byte_mask_update_enable: Boolean;
  signal addr_buffer :  std_logic_vector(35 downto 0);
  signal addr_update_enable: Boolean;
  signal wdata_buffer :  std_logic_vector(63 downto 0);
  signal wdata_update_enable: Boolean;
  -- output port buffer signals
  signal rdata_buffer :  std_logic_vector(63 downto 0);
  signal rdata_update_enable: Boolean;
  signal accessSysMem_CP_2627_start: Boolean;
  signal accessSysMem_CP_2627_symbol: Boolean;
  -- volatile/operator module components. 
  -- links between control-path and data-path
  signal WPIPE_L2CACHE_TO_MEM_REQUEST_2613_inst_req_1 : boolean;
  signal WPIPE_L2CACHE_TO_MEM_REQUEST_2613_inst_ack_0 : boolean;
  signal WPIPE_L2CACHE_TO_MEM_REQUEST_2613_inst_req_0 : boolean;
  signal WPIPE_L2CACHE_TO_MEM_REQUEST_2613_inst_ack_1 : boolean;
  signal RPIPE_MEM_TO_L2CACHE_RESPONSE_2617_inst_req_1 : boolean;
  signal RPIPE_MEM_TO_L2CACHE_RESPONSE_2617_inst_ack_1 : boolean;
  signal RPIPE_MEM_TO_L2CACHE_RESPONSE_2617_inst_ack_0 : boolean;
  signal RPIPE_MEM_TO_L2CACHE_RESPONSE_2617_inst_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "accessSysMem_input_buffer", -- 
      buffer_size => 2,
      bypass_flag => false,
      data_width => tag_length + 109) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= rwbar;
  rwbar_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(8 downto 1) <= byte_mask;
  byte_mask_buffer <= in_buffer_data_out(8 downto 1);
  in_buffer_data_in(44 downto 9) <= addr;
  addr_buffer <= in_buffer_data_out(44 downto 9);
  in_buffer_data_in(108 downto 45) <= wdata;
  wdata_buffer <= in_buffer_data_out(108 downto 45);
  in_buffer_data_in(tag_length + 108 downto 109) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 108 downto 109);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 5) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 1,5 => 15);
    constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1,5 => 15);
    constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 6); -- 
  begin -- 
    preds <= rwbar_update_enable & byte_mask_update_enable & addr_update_enable & wdata_update_enable & in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  accessSysMem_CP_2627_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "accessSysMem_out_buffer", -- 
      buffer_size => 2,
      full_rate => false,
      data_width => tag_length + 64) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(63 downto 0) <= rdata_buffer;
  rdata <= out_buffer_data_out(63 downto 0);
  out_buffer_data_in(tag_length + 63 downto 64) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 63 downto 64);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 15);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessSysMem_CP_2627_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  rdata_update_enable_join: block -- 
    constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
    constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
    constant place_delays: IntegerArray(0 to 0) := (0 => 0);
    constant joinName: string(1 to 24) := "rdata_update_enable_join"; 
    signal preds: BooleanArray(1 to 1); -- 
  begin -- 
    preds(1) <= out_buffer_write_ack_symbol;
    gj_rdata_update_enable_join : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => rdata_update_enable, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 15,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= accessSysMem_CP_2627_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= accessSysMem_CP_2627_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  accessSysMem_CP_2627: Block -- control-path 
    signal accessSysMem_CP_2627_elements: BooleanArray(20 downto 0);
    -- 
  begin -- 
    accessSysMem_CP_2627_elements(0) <= accessSysMem_CP_2627_start;
    accessSysMem_CP_2627_symbol <= accessSysMem_CP_2627_elements(20);
    -- CP-element group 0:  transition  bypass  pipeline-parent 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (1) 
      -- CP-element group 0: 	 $entry
      -- 
    -- CP-element group 1:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	7 
    -- CP-element group 1: 	10 
    -- CP-element group 1:  members (1) 
      -- CP-element group 1: 	 assign_stmt_2612_to_assign_stmt_2622/$entry
      -- 
    accessSysMem_CP_2627_elements(1) <= accessSysMem_CP_2627_elements(0);
    -- CP-element group 2:  join  transition  bypass  pipeline-parent 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: marked-predecessors 
    -- CP-element group 2: 	8 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	15 
    -- CP-element group 2:  members (2) 
      -- CP-element group 2: 	 assign_stmt_2612_to_assign_stmt_2622/rwbar_update_enable_out
      -- CP-element group 2: 	 assign_stmt_2612_to_assign_stmt_2622/rwbar_update_enable
      -- 
    accessSysMem_cp_element_group_2: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "accessSysMem_cp_element_group_2"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessSysMem_CP_2627_elements(8);
      gj_accessSysMem_cp_element_group_2 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessSysMem_CP_2627_elements(2), clk => clk, reset => reset); --
    end block;
    -- CP-element group 3:  join  transition  bypass  pipeline-parent 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: marked-predecessors 
    -- CP-element group 3: 	8 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	16 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 assign_stmt_2612_to_assign_stmt_2622/byte_mask_update_enable
      -- CP-element group 3: 	 assign_stmt_2612_to_assign_stmt_2622/byte_mask_update_enable_out
      -- 
    accessSysMem_cp_element_group_3: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "accessSysMem_cp_element_group_3"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessSysMem_CP_2627_elements(8);
      gj_accessSysMem_cp_element_group_3 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessSysMem_CP_2627_elements(3), clk => clk, reset => reset); --
    end block;
    -- CP-element group 4:  join  transition  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: marked-predecessors 
    -- CP-element group 4: 	8 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	17 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 assign_stmt_2612_to_assign_stmt_2622/addr_update_enable
      -- CP-element group 4: 	 assign_stmt_2612_to_assign_stmt_2622/addr_update_enable_out
      -- 
    accessSysMem_cp_element_group_4: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "accessSysMem_cp_element_group_4"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessSysMem_CP_2627_elements(8);
      gj_accessSysMem_cp_element_group_4 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessSysMem_CP_2627_elements(4), clk => clk, reset => reset); --
    end block;
    -- CP-element group 5:  join  transition  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: marked-predecessors 
    -- CP-element group 5: 	8 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	18 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 assign_stmt_2612_to_assign_stmt_2622/wdata_update_enable_out
      -- CP-element group 5: 	 assign_stmt_2612_to_assign_stmt_2622/wdata_update_enable
      -- 
    accessSysMem_cp_element_group_5: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 31) := "accessSysMem_cp_element_group_5"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= accessSysMem_CP_2627_elements(8);
      gj_accessSysMem_cp_element_group_5 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessSysMem_CP_2627_elements(5), clk => clk, reset => reset); --
    end block;
    -- CP-element group 6:  transition  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: 	19 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	11 
    -- CP-element group 6:  members (2) 
      -- CP-element group 6: 	 assign_stmt_2612_to_assign_stmt_2622/rdata_update_enable_in
      -- CP-element group 6: 	 assign_stmt_2612_to_assign_stmt_2622/rdata_update_enable
      -- 
    accessSysMem_CP_2627_elements(6) <= accessSysMem_CP_2627_elements(19);
    -- CP-element group 7:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	1 
    -- CP-element group 7: marked-predecessors 
    -- CP-element group 7: 	9 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	8 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 assign_stmt_2612_to_assign_stmt_2622/WPIPE_L2CACHE_TO_MEM_REQUEST_2613_sample_start_
      -- CP-element group 7: 	 assign_stmt_2612_to_assign_stmt_2622/WPIPE_L2CACHE_TO_MEM_REQUEST_2613_Sample/req
      -- CP-element group 7: 	 assign_stmt_2612_to_assign_stmt_2622/WPIPE_L2CACHE_TO_MEM_REQUEST_2613_Sample/$entry
      -- 
    req_2650_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2650_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessSysMem_CP_2627_elements(7), ack => WPIPE_L2CACHE_TO_MEM_REQUEST_2613_inst_req_0); -- 
    accessSysMem_cp_element_group_7: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 31) := "accessSysMem_cp_element_group_7"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessSysMem_CP_2627_elements(1) & accessSysMem_CP_2627_elements(9);
      gj_accessSysMem_cp_element_group_7 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessSysMem_CP_2627_elements(7), clk => clk, reset => reset); --
    end block;
    -- CP-element group 8:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	7 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	9 
    -- CP-element group 8: marked-successors 
    -- CP-element group 8: 	2 
    -- CP-element group 8: 	3 
    -- CP-element group 8: 	4 
    -- CP-element group 8: 	5 
    -- CP-element group 8:  members (6) 
      -- CP-element group 8: 	 assign_stmt_2612_to_assign_stmt_2622/WPIPE_L2CACHE_TO_MEM_REQUEST_2613_Sample/$exit
      -- CP-element group 8: 	 assign_stmt_2612_to_assign_stmt_2622/WPIPE_L2CACHE_TO_MEM_REQUEST_2613_Update/req
      -- CP-element group 8: 	 assign_stmt_2612_to_assign_stmt_2622/WPIPE_L2CACHE_TO_MEM_REQUEST_2613_Sample/ack
      -- CP-element group 8: 	 assign_stmt_2612_to_assign_stmt_2622/WPIPE_L2CACHE_TO_MEM_REQUEST_2613_update_start_
      -- CP-element group 8: 	 assign_stmt_2612_to_assign_stmt_2622/WPIPE_L2CACHE_TO_MEM_REQUEST_2613_sample_completed_
      -- CP-element group 8: 	 assign_stmt_2612_to_assign_stmt_2622/WPIPE_L2CACHE_TO_MEM_REQUEST_2613_Update/$entry
      -- 
    ack_2651_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 8_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_L2CACHE_TO_MEM_REQUEST_2613_inst_ack_0, ack => accessSysMem_CP_2627_elements(8)); -- 
    req_2655_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2655_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessSysMem_CP_2627_elements(8), ack => WPIPE_L2CACHE_TO_MEM_REQUEST_2613_inst_req_1); -- 
    -- CP-element group 9:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	8 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	14 
    -- CP-element group 9: marked-successors 
    -- CP-element group 9: 	7 
    -- CP-element group 9:  members (3) 
      -- CP-element group 9: 	 assign_stmt_2612_to_assign_stmt_2622/WPIPE_L2CACHE_TO_MEM_REQUEST_2613_update_completed_
      -- CP-element group 9: 	 assign_stmt_2612_to_assign_stmt_2622/WPIPE_L2CACHE_TO_MEM_REQUEST_2613_Update/$exit
      -- CP-element group 9: 	 assign_stmt_2612_to_assign_stmt_2622/WPIPE_L2CACHE_TO_MEM_REQUEST_2613_Update/ack
      -- 
    ack_2656_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 9_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_L2CACHE_TO_MEM_REQUEST_2613_inst_ack_1, ack => accessSysMem_CP_2627_elements(9)); -- 
    -- CP-element group 10:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	1 
    -- CP-element group 10: marked-predecessors 
    -- CP-element group 10: 	13 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	12 
    -- CP-element group 10:  members (3) 
      -- CP-element group 10: 	 assign_stmt_2612_to_assign_stmt_2622/RPIPE_MEM_TO_L2CACHE_RESPONSE_2617_Sample/rr
      -- CP-element group 10: 	 assign_stmt_2612_to_assign_stmt_2622/RPIPE_MEM_TO_L2CACHE_RESPONSE_2617_Sample/$entry
      -- CP-element group 10: 	 assign_stmt_2612_to_assign_stmt_2622/RPIPE_MEM_TO_L2CACHE_RESPONSE_2617_sample_start_
      -- 
    rr_2664_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2664_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessSysMem_CP_2627_elements(10), ack => RPIPE_MEM_TO_L2CACHE_RESPONSE_2617_inst_req_0); -- 
    accessSysMem_cp_element_group_10: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "accessSysMem_cp_element_group_10"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessSysMem_CP_2627_elements(1) & accessSysMem_CP_2627_elements(13);
      gj_accessSysMem_cp_element_group_10 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessSysMem_CP_2627_elements(10), clk => clk, reset => reset); --
    end block;
    -- CP-element group 11:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	6 
    -- CP-element group 11: 	12 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	13 
    -- CP-element group 11:  members (3) 
      -- CP-element group 11: 	 assign_stmt_2612_to_assign_stmt_2622/RPIPE_MEM_TO_L2CACHE_RESPONSE_2617_Update/$entry
      -- CP-element group 11: 	 assign_stmt_2612_to_assign_stmt_2622/RPIPE_MEM_TO_L2CACHE_RESPONSE_2617_Update/cr
      -- CP-element group 11: 	 assign_stmt_2612_to_assign_stmt_2622/RPIPE_MEM_TO_L2CACHE_RESPONSE_2617_update_start_
      -- 
    cr_2669_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2669_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => accessSysMem_CP_2627_elements(11), ack => RPIPE_MEM_TO_L2CACHE_RESPONSE_2617_inst_req_1); -- 
    accessSysMem_cp_element_group_11: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "accessSysMem_cp_element_group_11"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessSysMem_CP_2627_elements(6) & accessSysMem_CP_2627_elements(12);
      gj_accessSysMem_cp_element_group_11 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessSysMem_CP_2627_elements(11), clk => clk, reset => reset); --
    end block;
    -- CP-element group 12:  transition  input  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	10 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	11 
    -- CP-element group 12:  members (3) 
      -- CP-element group 12: 	 assign_stmt_2612_to_assign_stmt_2622/RPIPE_MEM_TO_L2CACHE_RESPONSE_2617_Sample/ra
      -- CP-element group 12: 	 assign_stmt_2612_to_assign_stmt_2622/RPIPE_MEM_TO_L2CACHE_RESPONSE_2617_Sample/$exit
      -- CP-element group 12: 	 assign_stmt_2612_to_assign_stmt_2622/RPIPE_MEM_TO_L2CACHE_RESPONSE_2617_sample_completed_
      -- 
    ra_2665_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 12_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_MEM_TO_L2CACHE_RESPONSE_2617_inst_ack_0, ack => accessSysMem_CP_2627_elements(12)); -- 
    -- CP-element group 13:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	11 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	14 
    -- CP-element group 13: marked-successors 
    -- CP-element group 13: 	10 
    -- CP-element group 13:  members (3) 
      -- CP-element group 13: 	 assign_stmt_2612_to_assign_stmt_2622/RPIPE_MEM_TO_L2CACHE_RESPONSE_2617_Update/$exit
      -- CP-element group 13: 	 assign_stmt_2612_to_assign_stmt_2622/RPIPE_MEM_TO_L2CACHE_RESPONSE_2617_Update/ca
      -- CP-element group 13: 	 assign_stmt_2612_to_assign_stmt_2622/RPIPE_MEM_TO_L2CACHE_RESPONSE_2617_update_completed_
      -- 
    ca_2670_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 13_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_MEM_TO_L2CACHE_RESPONSE_2617_inst_ack_1, ack => accessSysMem_CP_2627_elements(13)); -- 
    -- CP-element group 14:  join  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	9 
    -- CP-element group 14: 	13 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	20 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 assign_stmt_2612_to_assign_stmt_2622/$exit
      -- 
    accessSysMem_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 32) := "accessSysMem_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= accessSysMem_CP_2627_elements(9) & accessSysMem_CP_2627_elements(13);
      gj_accessSysMem_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => accessSysMem_CP_2627_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  place  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	2 
    -- CP-element group 15: successors 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 rwbar_update_enable
      -- 
    accessSysMem_CP_2627_elements(15) <= accessSysMem_CP_2627_elements(2);
    -- CP-element group 16:  place  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	3 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 byte_mask_update_enable
      -- 
    accessSysMem_CP_2627_elements(16) <= accessSysMem_CP_2627_elements(3);
    -- CP-element group 17:  place  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	4 
    -- CP-element group 17: successors 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 addr_update_enable
      -- 
    accessSysMem_CP_2627_elements(17) <= accessSysMem_CP_2627_elements(4);
    -- CP-element group 18:  place  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	5 
    -- CP-element group 18: successors 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 wdata_update_enable
      -- 
    accessSysMem_CP_2627_elements(18) <= accessSysMem_CP_2627_elements(5);
    -- CP-element group 19:  place  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	6 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 rdata_update_enable
      -- 
    -- CP-element group 20:  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	14 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 $exit
      -- 
    accessSysMem_CP_2627_elements(20) <= accessSysMem_CP_2627_elements(14);
    --  hookup: inputs to control-path 
    accessSysMem_CP_2627_elements(19) <= rdata_update_enable;
    -- hookup: output from control-path 
    addr_update_enable <= accessSysMem_CP_2627_elements(17);
    wdata_update_enable <= accessSysMem_CP_2627_elements(18);
    byte_mask_update_enable <= accessSysMem_CP_2627_elements(16);
    rwbar_update_enable <= accessSysMem_CP_2627_elements(15);
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u1_u2_2605_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u2_u10_2607_wire : std_logic_vector(9 downto 0);
    signal CONCAT_u36_u100_2610_wire : std_logic_vector(99 downto 0);
    signal rdata_plus_err_2618 : std_logic_vector(64 downto 0);
    signal to_sys_bus_2612 : std_logic_vector(109 downto 0);
    signal type_cast_2603_wire_constant : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    type_cast_2603_wire_constant <= "0";
    -- flow-through slice operator slice_2621_inst
    rdata_buffer <= rdata_plus_err_2618(63 downto 0);
    -- binary operator CONCAT_u10_u110_2611_inst
    process(CONCAT_u2_u10_2607_wire, CONCAT_u36_u100_2610_wire) -- 
      variable tmp_var : std_logic_vector(109 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u2_u10_2607_wire, CONCAT_u36_u100_2610_wire, tmp_var);
      to_sys_bus_2612 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_2605_inst
    process(type_cast_2603_wire_constant, rwbar_buffer) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_2603_wire_constant, rwbar_buffer, tmp_var);
      CONCAT_u1_u2_2605_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u2_u10_2607_inst
    process(CONCAT_u1_u2_2605_wire, byte_mask_buffer) -- 
      variable tmp_var : std_logic_vector(9 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_2605_wire, byte_mask_buffer, tmp_var);
      CONCAT_u2_u10_2607_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u36_u100_2610_inst
    process(addr_buffer, wdata_buffer) -- 
      variable tmp_var : std_logic_vector(99 downto 0); -- 
    begin -- 
      ApConcat_proc(addr_buffer, wdata_buffer, tmp_var);
      CONCAT_u36_u100_2610_wire <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_MEM_TO_L2CACHE_RESPONSE_2617_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(64 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_MEM_TO_L2CACHE_RESPONSE_2617_inst_req_0;
      RPIPE_MEM_TO_L2CACHE_RESPONSE_2617_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_MEM_TO_L2CACHE_RESPONSE_2617_inst_req_1;
      RPIPE_MEM_TO_L2CACHE_RESPONSE_2617_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      rdata_plus_err_2618 <= data_out(64 downto 0);
      MEM_TO_L2CACHE_RESPONSE_read_0_gI: SplitGuardInterface generic map(name => "MEM_TO_L2CACHE_RESPONSE_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      MEM_TO_L2CACHE_RESPONSE_read_0: InputPort_P2P -- 
        generic map ( name => "MEM_TO_L2CACHE_RESPONSE_read_0", data_width => 65,    bypass_flag => false,   	nonblocking_read_flag => false,  barrier_flag => false,   queue_depth =>  2)
        port map (-- 
          sample_req => reqL(0) , 
          sample_ack => ackL(0), 
          update_req => reqR(0), 
          update_ack => ackR(0), 
          data => data_out, 
          oreq => MEM_TO_L2CACHE_RESPONSE_pipe_read_req(0),
          oack => MEM_TO_L2CACHE_RESPONSE_pipe_read_ack(0),
          odata => MEM_TO_L2CACHE_RESPONSE_pipe_read_data(64 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared outport operator group (0) : WPIPE_L2CACHE_TO_MEM_REQUEST_2613_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(109 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_L2CACHE_TO_MEM_REQUEST_2613_inst_req_0;
      WPIPE_L2CACHE_TO_MEM_REQUEST_2613_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_L2CACHE_TO_MEM_REQUEST_2613_inst_req_1;
      WPIPE_L2CACHE_TO_MEM_REQUEST_2613_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= to_sys_bus_2612;
      L2CACHE_TO_MEM_REQUEST_write_0_gI: SplitGuardInterface generic map(name => "L2CACHE_TO_MEM_REQUEST_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      L2CACHE_TO_MEM_REQUEST_write_0: OutputPortRevised -- 
        generic map ( name => "L2CACHE_TO_MEM_REQUEST", data_width => 110, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => L2CACHE_TO_MEM_REQUEST_pipe_write_req(0),
          oack => L2CACHE_TO_MEM_REQUEST_pipe_write_ack(0),
          odata => L2CACHE_TO_MEM_REQUEST_pipe_write_data(109 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- 
  end Block; -- data_path
  -- 
end accessSysMem_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library l2_cache_lib;
use l2_cache_lib.l2_cache_global_package.all;
entity calculateHits_Volatile is -- 
  port ( -- 
    set_valids : in  std_logic_vector(7 downto 0);
    set_dirty_dword_masks : in  std_logic_vector(63 downto 0);
    set_tags : in  std_logic_vector(167 downto 0);
    pa_tag : in  std_logic_vector(20 downto 0);
    replace_index : in  std_logic_vector(2 downto 0);
    is_hit : out  std_logic_vector(0 downto 0);
    dirty_dword_mask : out  std_logic_vector(7 downto 0);
    access_index : out  std_logic_vector(2 downto 0);
    replace_line_is_valid : out  std_logic_vector(0 downto 0);
    replace_pa_tag : out  std_logic_vector(20 downto 0)-- 
  );
  -- 
end entity calculateHits_Volatile;
architecture calculateHits_Volatile_arch of calculateHits_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(264-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal set_valids_buffer :  std_logic_vector(7 downto 0);
  signal set_dirty_dword_masks_buffer :  std_logic_vector(63 downto 0);
  signal set_tags_buffer :  std_logic_vector(167 downto 0);
  signal pa_tag_buffer :  std_logic_vector(20 downto 0);
  signal replace_index_buffer :  std_logic_vector(2 downto 0);
  -- output port buffer signals
  signal is_hit_buffer :  std_logic_vector(0 downto 0);
  signal dirty_dword_mask_buffer :  std_logic_vector(7 downto 0);
  signal access_index_buffer :  std_logic_vector(2 downto 0);
  signal replace_line_is_valid_buffer :  std_logic_vector(0 downto 0);
  signal replace_pa_tag_buffer :  std_logic_vector(20 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  set_valids_buffer <= set_valids;
  set_dirty_dword_masks_buffer <= set_dirty_dword_masks;
  set_tags_buffer <= set_tags;
  pa_tag_buffer <= pa_tag;
  replace_index_buffer <= replace_index;
  -- output handling  -------------------------------------------------------
  is_hit <= is_hit_buffer;
  dirty_dword_mask <= dirty_dword_mask_buffer;
  access_index <= access_index_buffer;
  replace_line_is_valid <= replace_line_is_valid_buffer;
  replace_pa_tag <= replace_pa_tag_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal EQ_u21_u1_1490_wire : std_logic_vector(0 downto 0);
    signal EQ_u21_u1_1497_wire : std_logic_vector(0 downto 0);
    signal EQ_u21_u1_1504_wire : std_logic_vector(0 downto 0);
    signal EQ_u21_u1_1511_wire : std_logic_vector(0 downto 0);
    signal EQ_u21_u1_1518_wire : std_logic_vector(0 downto 0);
    signal EQ_u21_u1_1525_wire : std_logic_vector(0 downto 0);
    signal EQ_u21_u1_1532_wire : std_logic_vector(0 downto 0);
    signal EQ_u21_u1_1539_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1343_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1349_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1356_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1362_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1370_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1376_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1383_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1389_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1400_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1406_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1413_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1419_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1427_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1433_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1440_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1446_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1610_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1616_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1623_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1629_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1637_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1643_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1650_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1656_wire : std_logic_vector(0 downto 0);
    signal MUX_1346_wire : std_logic_vector(0 downto 0);
    signal MUX_1352_wire : std_logic_vector(0 downto 0);
    signal MUX_1359_wire : std_logic_vector(0 downto 0);
    signal MUX_1365_wire : std_logic_vector(0 downto 0);
    signal MUX_1373_wire : std_logic_vector(0 downto 0);
    signal MUX_1379_wire : std_logic_vector(0 downto 0);
    signal MUX_1386_wire : std_logic_vector(0 downto 0);
    signal MUX_1392_wire : std_logic_vector(0 downto 0);
    signal MUX_1403_wire : std_logic_vector(20 downto 0);
    signal MUX_1409_wire : std_logic_vector(20 downto 0);
    signal MUX_1416_wire : std_logic_vector(20 downto 0);
    signal MUX_1422_wire : std_logic_vector(20 downto 0);
    signal MUX_1430_wire : std_logic_vector(20 downto 0);
    signal MUX_1436_wire : std_logic_vector(20 downto 0);
    signal MUX_1443_wire : std_logic_vector(20 downto 0);
    signal MUX_1449_wire : std_logic_vector(20 downto 0);
    signal MUX_1564_wire : std_logic_vector(2 downto 0);
    signal MUX_1568_wire : std_logic_vector(2 downto 0);
    signal MUX_1573_wire : std_logic_vector(2 downto 0);
    signal MUX_1577_wire : std_logic_vector(2 downto 0);
    signal MUX_1583_wire : std_logic_vector(2 downto 0);
    signal MUX_1587_wire : std_logic_vector(2 downto 0);
    signal MUX_1592_wire : std_logic_vector(2 downto 0);
    signal MUX_1596_wire : std_logic_vector(2 downto 0);
    signal MUX_1613_wire : std_logic_vector(7 downto 0);
    signal MUX_1619_wire : std_logic_vector(7 downto 0);
    signal MUX_1626_wire : std_logic_vector(7 downto 0);
    signal MUX_1632_wire : std_logic_vector(7 downto 0);
    signal MUX_1640_wire : std_logic_vector(7 downto 0);
    signal MUX_1646_wire : std_logic_vector(7 downto 0);
    signal MUX_1653_wire : std_logic_vector(7 downto 0);
    signal MUX_1659_wire : std_logic_vector(7 downto 0);
    signal OR_u1_u1_1353_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1366_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1367_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1380_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1393_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1394_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1545_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1548_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1549_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1552_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1555_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1556_wire : std_logic_vector(0 downto 0);
    signal OR_u21_u21_1410_wire : std_logic_vector(20 downto 0);
    signal OR_u21_u21_1423_wire : std_logic_vector(20 downto 0);
    signal OR_u21_u21_1424_wire : std_logic_vector(20 downto 0);
    signal OR_u21_u21_1437_wire : std_logic_vector(20 downto 0);
    signal OR_u21_u21_1450_wire : std_logic_vector(20 downto 0);
    signal OR_u21_u21_1451_wire : std_logic_vector(20 downto 0);
    signal OR_u3_u3_1569_wire : std_logic_vector(2 downto 0);
    signal OR_u3_u3_1578_wire : std_logic_vector(2 downto 0);
    signal OR_u3_u3_1579_wire : std_logic_vector(2 downto 0);
    signal OR_u3_u3_1588_wire : std_logic_vector(2 downto 0);
    signal OR_u3_u3_1597_wire : std_logic_vector(2 downto 0);
    signal OR_u3_u3_1598_wire : std_logic_vector(2 downto 0);
    signal OR_u8_u8_1620_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_1633_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_1634_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_1647_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_1660_wire : std_logic_vector(7 downto 0);
    signal OR_u8_u8_1661_wire : std_logic_vector(7 downto 0);
    signal h0_1492 : std_logic_vector(0 downto 0);
    signal h1_1499 : std_logic_vector(0 downto 0);
    signal h2_1506 : std_logic_vector(0 downto 0);
    signal h3_1513 : std_logic_vector(0 downto 0);
    signal h4_1520 : std_logic_vector(0 downto 0);
    signal h5_1527 : std_logic_vector(0 downto 0);
    signal h6_1534 : std_logic_vector(0 downto 0);
    signal h7_1541 : std_logic_vector(0 downto 0);
    signal hit_index_1600 : std_logic_vector(2 downto 0);
    signal konst_1342_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1345_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1348_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1351_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1355_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1358_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1361_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1364_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1369_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1372_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1375_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1378_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1382_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1385_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1388_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1391_wire_constant : std_logic_vector(0 downto 0);
    signal konst_1399_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1402_wire_constant : std_logic_vector(20 downto 0);
    signal konst_1405_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1408_wire_constant : std_logic_vector(20 downto 0);
    signal konst_1412_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1415_wire_constant : std_logic_vector(20 downto 0);
    signal konst_1418_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1421_wire_constant : std_logic_vector(20 downto 0);
    signal konst_1426_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1429_wire_constant : std_logic_vector(20 downto 0);
    signal konst_1432_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1435_wire_constant : std_logic_vector(20 downto 0);
    signal konst_1439_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1442_wire_constant : std_logic_vector(20 downto 0);
    signal konst_1445_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1448_wire_constant : std_logic_vector(20 downto 0);
    signal konst_1563_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1566_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1567_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1571_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1572_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1575_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1576_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1581_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1582_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1585_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1586_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1590_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1591_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1594_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1595_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1609_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1612_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1615_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1618_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1622_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1625_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1628_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1631_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1636_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1639_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1642_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1645_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1649_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1652_wire_constant : std_logic_vector(7 downto 0);
    signal konst_1655_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1658_wire_constant : std_logic_vector(7 downto 0);
    signal m0_1457 : std_logic_vector(7 downto 0);
    signal m1_1461 : std_logic_vector(7 downto 0);
    signal m2_1465 : std_logic_vector(7 downto 0);
    signal m3_1469 : std_logic_vector(7 downto 0);
    signal m4_1473 : std_logic_vector(7 downto 0);
    signal m5_1477 : std_logic_vector(7 downto 0);
    signal m6_1481 : std_logic_vector(7 downto 0);
    signal m7_1485 : std_logic_vector(7 downto 0);
    signal t0_1311 : std_logic_vector(20 downto 0);
    signal t1_1315 : std_logic_vector(20 downto 0);
    signal t2_1319 : std_logic_vector(20 downto 0);
    signal t3_1323 : std_logic_vector(20 downto 0);
    signal t4_1327 : std_logic_vector(20 downto 0);
    signal t5_1331 : std_logic_vector(20 downto 0);
    signal t6_1335 : std_logic_vector(20 downto 0);
    signal t7_1339 : std_logic_vector(20 downto 0);
    signal type_cast_1562_wire_constant : std_logic_vector(2 downto 0);
    signal v0_1279 : std_logic_vector(0 downto 0);
    signal v1_1283 : std_logic_vector(0 downto 0);
    signal v2_1287 : std_logic_vector(0 downto 0);
    signal v3_1291 : std_logic_vector(0 downto 0);
    signal v4_1295 : std_logic_vector(0 downto 0);
    signal v5_1299 : std_logic_vector(0 downto 0);
    signal v6_1303 : std_logic_vector(0 downto 0);
    signal v7_1307 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    konst_1342_wire_constant <= "000";
    konst_1345_wire_constant <= "0";
    konst_1348_wire_constant <= "001";
    konst_1351_wire_constant <= "0";
    konst_1355_wire_constant <= "010";
    konst_1358_wire_constant <= "0";
    konst_1361_wire_constant <= "011";
    konst_1364_wire_constant <= "0";
    konst_1369_wire_constant <= "100";
    konst_1372_wire_constant <= "0";
    konst_1375_wire_constant <= "101";
    konst_1378_wire_constant <= "0";
    konst_1382_wire_constant <= "110";
    konst_1385_wire_constant <= "0";
    konst_1388_wire_constant <= "111";
    konst_1391_wire_constant <= "0";
    konst_1399_wire_constant <= "000";
    konst_1402_wire_constant <= "000000000000000000000";
    konst_1405_wire_constant <= "001";
    konst_1408_wire_constant <= "000000000000000000000";
    konst_1412_wire_constant <= "010";
    konst_1415_wire_constant <= "000000000000000000000";
    konst_1418_wire_constant <= "011";
    konst_1421_wire_constant <= "000000000000000000000";
    konst_1426_wire_constant <= "100";
    konst_1429_wire_constant <= "000000000000000000000";
    konst_1432_wire_constant <= "101";
    konst_1435_wire_constant <= "000000000000000000000";
    konst_1439_wire_constant <= "110";
    konst_1442_wire_constant <= "000000000000000000000";
    konst_1445_wire_constant <= "111";
    konst_1448_wire_constant <= "000000000000000000000";
    konst_1563_wire_constant <= "000";
    konst_1566_wire_constant <= "001";
    konst_1567_wire_constant <= "000";
    konst_1571_wire_constant <= "010";
    konst_1572_wire_constant <= "000";
    konst_1575_wire_constant <= "011";
    konst_1576_wire_constant <= "000";
    konst_1581_wire_constant <= "100";
    konst_1582_wire_constant <= "000";
    konst_1585_wire_constant <= "101";
    konst_1586_wire_constant <= "000";
    konst_1590_wire_constant <= "110";
    konst_1591_wire_constant <= "000";
    konst_1594_wire_constant <= "111";
    konst_1595_wire_constant <= "000";
    konst_1609_wire_constant <= "000";
    konst_1612_wire_constant <= "00000000";
    konst_1615_wire_constant <= "001";
    konst_1618_wire_constant <= "00000000";
    konst_1622_wire_constant <= "010";
    konst_1625_wire_constant <= "00000000";
    konst_1628_wire_constant <= "011";
    konst_1631_wire_constant <= "00000000";
    konst_1636_wire_constant <= "100";
    konst_1639_wire_constant <= "00000000";
    konst_1642_wire_constant <= "101";
    konst_1645_wire_constant <= "00000000";
    konst_1649_wire_constant <= "110";
    konst_1652_wire_constant <= "00000000";
    konst_1655_wire_constant <= "111";
    konst_1658_wire_constant <= "00000000";
    type_cast_1562_wire_constant <= "000";
    -- flow-through select operator MUX_1346_inst
    MUX_1346_wire <= v0_1279 when (EQ_u3_u1_1343_wire(0) /=  '0') else konst_1345_wire_constant;
    -- flow-through select operator MUX_1352_inst
    MUX_1352_wire <= v1_1283 when (EQ_u3_u1_1349_wire(0) /=  '0') else konst_1351_wire_constant;
    -- flow-through select operator MUX_1359_inst
    MUX_1359_wire <= v2_1287 when (EQ_u3_u1_1356_wire(0) /=  '0') else konst_1358_wire_constant;
    -- flow-through select operator MUX_1365_inst
    MUX_1365_wire <= v3_1291 when (EQ_u3_u1_1362_wire(0) /=  '0') else konst_1364_wire_constant;
    -- flow-through select operator MUX_1373_inst
    MUX_1373_wire <= v4_1295 when (EQ_u3_u1_1370_wire(0) /=  '0') else konst_1372_wire_constant;
    -- flow-through select operator MUX_1379_inst
    MUX_1379_wire <= v5_1299 when (EQ_u3_u1_1376_wire(0) /=  '0') else konst_1378_wire_constant;
    -- flow-through select operator MUX_1386_inst
    MUX_1386_wire <= v6_1303 when (EQ_u3_u1_1383_wire(0) /=  '0') else konst_1385_wire_constant;
    -- flow-through select operator MUX_1392_inst
    MUX_1392_wire <= v7_1307 when (EQ_u3_u1_1389_wire(0) /=  '0') else konst_1391_wire_constant;
    -- flow-through select operator MUX_1403_inst
    MUX_1403_wire <= t0_1311 when (EQ_u3_u1_1400_wire(0) /=  '0') else konst_1402_wire_constant;
    -- flow-through select operator MUX_1409_inst
    MUX_1409_wire <= t1_1315 when (EQ_u3_u1_1406_wire(0) /=  '0') else konst_1408_wire_constant;
    -- flow-through select operator MUX_1416_inst
    MUX_1416_wire <= t2_1319 when (EQ_u3_u1_1413_wire(0) /=  '0') else konst_1415_wire_constant;
    -- flow-through select operator MUX_1422_inst
    MUX_1422_wire <= t3_1323 when (EQ_u3_u1_1419_wire(0) /=  '0') else konst_1421_wire_constant;
    -- flow-through select operator MUX_1430_inst
    MUX_1430_wire <= t4_1327 when (EQ_u3_u1_1427_wire(0) /=  '0') else konst_1429_wire_constant;
    -- flow-through select operator MUX_1436_inst
    MUX_1436_wire <= t5_1331 when (EQ_u3_u1_1433_wire(0) /=  '0') else konst_1435_wire_constant;
    -- flow-through select operator MUX_1443_inst
    MUX_1443_wire <= t6_1335 when (EQ_u3_u1_1440_wire(0) /=  '0') else konst_1442_wire_constant;
    -- flow-through select operator MUX_1449_inst
    MUX_1449_wire <= t7_1339 when (EQ_u3_u1_1446_wire(0) /=  '0') else konst_1448_wire_constant;
    -- flow-through select operator MUX_1564_inst
    MUX_1564_wire <= type_cast_1562_wire_constant when (h0_1492(0) /=  '0') else konst_1563_wire_constant;
    -- flow-through select operator MUX_1568_inst
    MUX_1568_wire <= konst_1566_wire_constant when (h1_1499(0) /=  '0') else konst_1567_wire_constant;
    -- flow-through select operator MUX_1573_inst
    MUX_1573_wire <= konst_1571_wire_constant when (h2_1506(0) /=  '0') else konst_1572_wire_constant;
    -- flow-through select operator MUX_1577_inst
    MUX_1577_wire <= konst_1575_wire_constant when (h3_1513(0) /=  '0') else konst_1576_wire_constant;
    -- flow-through select operator MUX_1583_inst
    MUX_1583_wire <= konst_1581_wire_constant when (h4_1520(0) /=  '0') else konst_1582_wire_constant;
    -- flow-through select operator MUX_1587_inst
    MUX_1587_wire <= konst_1585_wire_constant when (h5_1527(0) /=  '0') else konst_1586_wire_constant;
    -- flow-through select operator MUX_1592_inst
    MUX_1592_wire <= konst_1590_wire_constant when (h6_1534(0) /=  '0') else konst_1591_wire_constant;
    -- flow-through select operator MUX_1596_inst
    MUX_1596_wire <= konst_1594_wire_constant when (h7_1541(0) /=  '0') else konst_1595_wire_constant;
    -- flow-through select operator MUX_1605_inst
    access_index_buffer <= hit_index_1600 when (is_hit_buffer(0) /=  '0') else replace_index_buffer;
    -- flow-through select operator MUX_1613_inst
    MUX_1613_wire <= m0_1457 when (EQ_u3_u1_1610_wire(0) /=  '0') else konst_1612_wire_constant;
    -- flow-through select operator MUX_1619_inst
    MUX_1619_wire <= m1_1461 when (EQ_u3_u1_1616_wire(0) /=  '0') else konst_1618_wire_constant;
    -- flow-through select operator MUX_1626_inst
    MUX_1626_wire <= m2_1465 when (EQ_u3_u1_1623_wire(0) /=  '0') else konst_1625_wire_constant;
    -- flow-through select operator MUX_1632_inst
    MUX_1632_wire <= m3_1469 when (EQ_u3_u1_1629_wire(0) /=  '0') else konst_1631_wire_constant;
    -- flow-through select operator MUX_1640_inst
    MUX_1640_wire <= m4_1473 when (EQ_u3_u1_1637_wire(0) /=  '0') else konst_1639_wire_constant;
    -- flow-through select operator MUX_1646_inst
    MUX_1646_wire <= m5_1477 when (EQ_u3_u1_1643_wire(0) /=  '0') else konst_1645_wire_constant;
    -- flow-through select operator MUX_1653_inst
    MUX_1653_wire <= m6_1481 when (EQ_u3_u1_1650_wire(0) /=  '0') else konst_1652_wire_constant;
    -- flow-through select operator MUX_1659_inst
    MUX_1659_wire <= m7_1485 when (EQ_u3_u1_1656_wire(0) /=  '0') else konst_1658_wire_constant;
    -- flow-through slice operator slice_1278_inst
    v0_1279 <= set_valids_buffer(7 downto 7);
    -- flow-through slice operator slice_1282_inst
    v1_1283 <= set_valids_buffer(6 downto 6);
    -- flow-through slice operator slice_1286_inst
    v2_1287 <= set_valids_buffer(5 downto 5);
    -- flow-through slice operator slice_1290_inst
    v3_1291 <= set_valids_buffer(4 downto 4);
    -- flow-through slice operator slice_1294_inst
    v4_1295 <= set_valids_buffer(3 downto 3);
    -- flow-through slice operator slice_1298_inst
    v5_1299 <= set_valids_buffer(2 downto 2);
    -- flow-through slice operator slice_1302_inst
    v6_1303 <= set_valids_buffer(1 downto 1);
    -- flow-through slice operator slice_1306_inst
    v7_1307 <= set_valids_buffer(0 downto 0);
    -- flow-through slice operator slice_1310_inst
    t0_1311 <= set_tags_buffer(167 downto 147);
    -- flow-through slice operator slice_1314_inst
    t1_1315 <= set_tags_buffer(146 downto 126);
    -- flow-through slice operator slice_1318_inst
    t2_1319 <= set_tags_buffer(125 downto 105);
    -- flow-through slice operator slice_1322_inst
    t3_1323 <= set_tags_buffer(104 downto 84);
    -- flow-through slice operator slice_1326_inst
    t4_1327 <= set_tags_buffer(83 downto 63);
    -- flow-through slice operator slice_1330_inst
    t5_1331 <= set_tags_buffer(62 downto 42);
    -- flow-through slice operator slice_1334_inst
    t6_1335 <= set_tags_buffer(41 downto 21);
    -- flow-through slice operator slice_1338_inst
    t7_1339 <= set_tags_buffer(20 downto 0);
    -- flow-through slice operator slice_1456_inst
    m0_1457 <= set_dirty_dword_masks_buffer(63 downto 56);
    -- flow-through slice operator slice_1460_inst
    m1_1461 <= set_dirty_dword_masks_buffer(55 downto 48);
    -- flow-through slice operator slice_1464_inst
    m2_1465 <= set_dirty_dword_masks_buffer(47 downto 40);
    -- flow-through slice operator slice_1468_inst
    m3_1469 <= set_dirty_dword_masks_buffer(39 downto 32);
    -- flow-through slice operator slice_1472_inst
    m4_1473 <= set_dirty_dword_masks_buffer(31 downto 24);
    -- flow-through slice operator slice_1476_inst
    m5_1477 <= set_dirty_dword_masks_buffer(23 downto 16);
    -- flow-through slice operator slice_1480_inst
    m6_1481 <= set_dirty_dword_masks_buffer(15 downto 8);
    -- flow-through slice operator slice_1484_inst
    m7_1485 <= set_dirty_dword_masks_buffer(7 downto 0);
    -- binary operator AND_u1_u1_1491_inst
    process(v0_1279, EQ_u21_u1_1490_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(v0_1279, EQ_u21_u1_1490_wire, tmp_var);
      h0_1492 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1498_inst
    process(v1_1283, EQ_u21_u1_1497_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(v1_1283, EQ_u21_u1_1497_wire, tmp_var);
      h1_1499 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1505_inst
    process(v2_1287, EQ_u21_u1_1504_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(v2_1287, EQ_u21_u1_1504_wire, tmp_var);
      h2_1506 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1512_inst
    process(v3_1291, EQ_u21_u1_1511_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(v3_1291, EQ_u21_u1_1511_wire, tmp_var);
      h3_1513 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1519_inst
    process(v4_1295, EQ_u21_u1_1518_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(v4_1295, EQ_u21_u1_1518_wire, tmp_var);
      h4_1520 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1526_inst
    process(v5_1299, EQ_u21_u1_1525_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(v5_1299, EQ_u21_u1_1525_wire, tmp_var);
      h5_1527 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1533_inst
    process(v6_1303, EQ_u21_u1_1532_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(v6_1303, EQ_u21_u1_1532_wire, tmp_var);
      h6_1534 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1540_inst
    process(v7_1307, EQ_u21_u1_1539_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(v7_1307, EQ_u21_u1_1539_wire, tmp_var);
      h7_1541 <= tmp_var; --
    end process;
    -- binary operator EQ_u21_u1_1490_inst
    process(t0_1311, pa_tag_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(t0_1311, pa_tag_buffer, tmp_var);
      EQ_u21_u1_1490_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u21_u1_1497_inst
    process(t1_1315, pa_tag_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(t1_1315, pa_tag_buffer, tmp_var);
      EQ_u21_u1_1497_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u21_u1_1504_inst
    process(t2_1319, pa_tag_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(t2_1319, pa_tag_buffer, tmp_var);
      EQ_u21_u1_1504_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u21_u1_1511_inst
    process(t3_1323, pa_tag_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(t3_1323, pa_tag_buffer, tmp_var);
      EQ_u21_u1_1511_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u21_u1_1518_inst
    process(t4_1327, pa_tag_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(t4_1327, pa_tag_buffer, tmp_var);
      EQ_u21_u1_1518_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u21_u1_1525_inst
    process(t5_1331, pa_tag_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(t5_1331, pa_tag_buffer, tmp_var);
      EQ_u21_u1_1525_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u21_u1_1532_inst
    process(t6_1335, pa_tag_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(t6_1335, pa_tag_buffer, tmp_var);
      EQ_u21_u1_1532_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u21_u1_1539_inst
    process(t7_1339, pa_tag_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(t7_1339, pa_tag_buffer, tmp_var);
      EQ_u21_u1_1539_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1343_inst
    process(replace_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(replace_index_buffer, konst_1342_wire_constant, tmp_var);
      EQ_u3_u1_1343_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1349_inst
    process(replace_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(replace_index_buffer, konst_1348_wire_constant, tmp_var);
      EQ_u3_u1_1349_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1356_inst
    process(replace_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(replace_index_buffer, konst_1355_wire_constant, tmp_var);
      EQ_u3_u1_1356_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1362_inst
    process(replace_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(replace_index_buffer, konst_1361_wire_constant, tmp_var);
      EQ_u3_u1_1362_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1370_inst
    process(replace_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(replace_index_buffer, konst_1369_wire_constant, tmp_var);
      EQ_u3_u1_1370_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1376_inst
    process(replace_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(replace_index_buffer, konst_1375_wire_constant, tmp_var);
      EQ_u3_u1_1376_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1383_inst
    process(replace_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(replace_index_buffer, konst_1382_wire_constant, tmp_var);
      EQ_u3_u1_1383_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1389_inst
    process(replace_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(replace_index_buffer, konst_1388_wire_constant, tmp_var);
      EQ_u3_u1_1389_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1400_inst
    process(replace_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(replace_index_buffer, konst_1399_wire_constant, tmp_var);
      EQ_u3_u1_1400_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1406_inst
    process(replace_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(replace_index_buffer, konst_1405_wire_constant, tmp_var);
      EQ_u3_u1_1406_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1413_inst
    process(replace_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(replace_index_buffer, konst_1412_wire_constant, tmp_var);
      EQ_u3_u1_1413_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1419_inst
    process(replace_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(replace_index_buffer, konst_1418_wire_constant, tmp_var);
      EQ_u3_u1_1419_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1427_inst
    process(replace_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(replace_index_buffer, konst_1426_wire_constant, tmp_var);
      EQ_u3_u1_1427_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1433_inst
    process(replace_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(replace_index_buffer, konst_1432_wire_constant, tmp_var);
      EQ_u3_u1_1433_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1440_inst
    process(replace_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(replace_index_buffer, konst_1439_wire_constant, tmp_var);
      EQ_u3_u1_1440_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1446_inst
    process(replace_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(replace_index_buffer, konst_1445_wire_constant, tmp_var);
      EQ_u3_u1_1446_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1610_inst
    process(access_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(access_index_buffer, konst_1609_wire_constant, tmp_var);
      EQ_u3_u1_1610_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1616_inst
    process(access_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(access_index_buffer, konst_1615_wire_constant, tmp_var);
      EQ_u3_u1_1616_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1623_inst
    process(access_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(access_index_buffer, konst_1622_wire_constant, tmp_var);
      EQ_u3_u1_1623_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1629_inst
    process(access_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(access_index_buffer, konst_1628_wire_constant, tmp_var);
      EQ_u3_u1_1629_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1637_inst
    process(access_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(access_index_buffer, konst_1636_wire_constant, tmp_var);
      EQ_u3_u1_1637_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1643_inst
    process(access_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(access_index_buffer, konst_1642_wire_constant, tmp_var);
      EQ_u3_u1_1643_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1650_inst
    process(access_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(access_index_buffer, konst_1649_wire_constant, tmp_var);
      EQ_u3_u1_1650_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1656_inst
    process(access_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(access_index_buffer, konst_1655_wire_constant, tmp_var);
      EQ_u3_u1_1656_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1353_inst
    process(MUX_1346_wire, MUX_1352_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1346_wire, MUX_1352_wire, tmp_var);
      OR_u1_u1_1353_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1366_inst
    process(MUX_1359_wire, MUX_1365_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1359_wire, MUX_1365_wire, tmp_var);
      OR_u1_u1_1366_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1367_inst
    process(OR_u1_u1_1353_wire, OR_u1_u1_1366_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_1353_wire, OR_u1_u1_1366_wire, tmp_var);
      OR_u1_u1_1367_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1380_inst
    process(MUX_1373_wire, MUX_1379_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1373_wire, MUX_1379_wire, tmp_var);
      OR_u1_u1_1380_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1393_inst
    process(MUX_1386_wire, MUX_1392_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1386_wire, MUX_1392_wire, tmp_var);
      OR_u1_u1_1393_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1394_inst
    process(OR_u1_u1_1380_wire, OR_u1_u1_1393_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_1380_wire, OR_u1_u1_1393_wire, tmp_var);
      OR_u1_u1_1394_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1395_inst
    process(OR_u1_u1_1367_wire, OR_u1_u1_1394_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_1367_wire, OR_u1_u1_1394_wire, tmp_var);
      replace_line_is_valid_buffer <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1545_inst
    process(h0_1492, h1_1499) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(h0_1492, h1_1499, tmp_var);
      OR_u1_u1_1545_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1548_inst
    process(h2_1506, h3_1513) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(h2_1506, h3_1513, tmp_var);
      OR_u1_u1_1548_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1549_inst
    process(OR_u1_u1_1545_wire, OR_u1_u1_1548_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_1545_wire, OR_u1_u1_1548_wire, tmp_var);
      OR_u1_u1_1549_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1552_inst
    process(h4_1520, h5_1527) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(h4_1520, h5_1527, tmp_var);
      OR_u1_u1_1552_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1555_inst
    process(h6_1534, h7_1541) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(h6_1534, h7_1541, tmp_var);
      OR_u1_u1_1555_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1556_inst
    process(OR_u1_u1_1552_wire, OR_u1_u1_1555_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_1552_wire, OR_u1_u1_1555_wire, tmp_var);
      OR_u1_u1_1556_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_1557_inst
    process(OR_u1_u1_1549_wire, OR_u1_u1_1556_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_1549_wire, OR_u1_u1_1556_wire, tmp_var);
      is_hit_buffer <= tmp_var; --
    end process;
    -- binary operator OR_u21_u21_1410_inst
    process(MUX_1403_wire, MUX_1409_wire) -- 
      variable tmp_var : std_logic_vector(20 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1403_wire, MUX_1409_wire, tmp_var);
      OR_u21_u21_1410_wire <= tmp_var; --
    end process;
    -- binary operator OR_u21_u21_1423_inst
    process(MUX_1416_wire, MUX_1422_wire) -- 
      variable tmp_var : std_logic_vector(20 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1416_wire, MUX_1422_wire, tmp_var);
      OR_u21_u21_1423_wire <= tmp_var; --
    end process;
    -- binary operator OR_u21_u21_1424_inst
    process(OR_u21_u21_1410_wire, OR_u21_u21_1423_wire) -- 
      variable tmp_var : std_logic_vector(20 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u21_u21_1410_wire, OR_u21_u21_1423_wire, tmp_var);
      OR_u21_u21_1424_wire <= tmp_var; --
    end process;
    -- binary operator OR_u21_u21_1437_inst
    process(MUX_1430_wire, MUX_1436_wire) -- 
      variable tmp_var : std_logic_vector(20 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1430_wire, MUX_1436_wire, tmp_var);
      OR_u21_u21_1437_wire <= tmp_var; --
    end process;
    -- binary operator OR_u21_u21_1450_inst
    process(MUX_1443_wire, MUX_1449_wire) -- 
      variable tmp_var : std_logic_vector(20 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1443_wire, MUX_1449_wire, tmp_var);
      OR_u21_u21_1450_wire <= tmp_var; --
    end process;
    -- binary operator OR_u21_u21_1451_inst
    process(OR_u21_u21_1437_wire, OR_u21_u21_1450_wire) -- 
      variable tmp_var : std_logic_vector(20 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u21_u21_1437_wire, OR_u21_u21_1450_wire, tmp_var);
      OR_u21_u21_1451_wire <= tmp_var; --
    end process;
    -- binary operator OR_u21_u21_1452_inst
    process(OR_u21_u21_1424_wire, OR_u21_u21_1451_wire) -- 
      variable tmp_var : std_logic_vector(20 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u21_u21_1424_wire, OR_u21_u21_1451_wire, tmp_var);
      replace_pa_tag_buffer <= tmp_var; --
    end process;
    -- binary operator OR_u3_u3_1569_inst
    process(MUX_1564_wire, MUX_1568_wire) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1564_wire, MUX_1568_wire, tmp_var);
      OR_u3_u3_1569_wire <= tmp_var; --
    end process;
    -- binary operator OR_u3_u3_1578_inst
    process(MUX_1573_wire, MUX_1577_wire) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1573_wire, MUX_1577_wire, tmp_var);
      OR_u3_u3_1578_wire <= tmp_var; --
    end process;
    -- binary operator OR_u3_u3_1579_inst
    process(OR_u3_u3_1569_wire, OR_u3_u3_1578_wire) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u3_u3_1569_wire, OR_u3_u3_1578_wire, tmp_var);
      OR_u3_u3_1579_wire <= tmp_var; --
    end process;
    -- binary operator OR_u3_u3_1588_inst
    process(MUX_1583_wire, MUX_1587_wire) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1583_wire, MUX_1587_wire, tmp_var);
      OR_u3_u3_1588_wire <= tmp_var; --
    end process;
    -- binary operator OR_u3_u3_1597_inst
    process(MUX_1592_wire, MUX_1596_wire) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1592_wire, MUX_1596_wire, tmp_var);
      OR_u3_u3_1597_wire <= tmp_var; --
    end process;
    -- binary operator OR_u3_u3_1598_inst
    process(OR_u3_u3_1588_wire, OR_u3_u3_1597_wire) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u3_u3_1588_wire, OR_u3_u3_1597_wire, tmp_var);
      OR_u3_u3_1598_wire <= tmp_var; --
    end process;
    -- binary operator OR_u3_u3_1599_inst
    process(OR_u3_u3_1579_wire, OR_u3_u3_1598_wire) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u3_u3_1579_wire, OR_u3_u3_1598_wire, tmp_var);
      hit_index_1600 <= tmp_var; --
    end process;
    -- binary operator OR_u8_u8_1620_inst
    process(MUX_1613_wire, MUX_1619_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1613_wire, MUX_1619_wire, tmp_var);
      OR_u8_u8_1620_wire <= tmp_var; --
    end process;
    -- binary operator OR_u8_u8_1633_inst
    process(MUX_1626_wire, MUX_1632_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1626_wire, MUX_1632_wire, tmp_var);
      OR_u8_u8_1633_wire <= tmp_var; --
    end process;
    -- binary operator OR_u8_u8_1634_inst
    process(OR_u8_u8_1620_wire, OR_u8_u8_1633_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u8_u8_1620_wire, OR_u8_u8_1633_wire, tmp_var);
      OR_u8_u8_1634_wire <= tmp_var; --
    end process;
    -- binary operator OR_u8_u8_1647_inst
    process(MUX_1640_wire, MUX_1646_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1640_wire, MUX_1646_wire, tmp_var);
      OR_u8_u8_1647_wire <= tmp_var; --
    end process;
    -- binary operator OR_u8_u8_1660_inst
    process(MUX_1653_wire, MUX_1659_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_1653_wire, MUX_1659_wire, tmp_var);
      OR_u8_u8_1660_wire <= tmp_var; --
    end process;
    -- binary operator OR_u8_u8_1661_inst
    process(OR_u8_u8_1647_wire, OR_u8_u8_1660_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u8_u8_1647_wire, OR_u8_u8_1660_wire, tmp_var);
      OR_u8_u8_1661_wire <= tmp_var; --
    end process;
    -- binary operator OR_u8_u8_1662_inst
    process(OR_u8_u8_1634_wire, OR_u8_u8_1661_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u8_u8_1634_wire, OR_u8_u8_1661_wire, tmp_var);
      dirty_dword_mask_buffer <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end calculateHits_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library l2_cache_lib;
use l2_cache_lib.l2_cache_global_package.all;
entity dwordId_Volatile is -- 
  port ( -- 
    pa : in  std_logic_vector(35 downto 0);
    dword_id : out  std_logic_vector(2 downto 0)-- 
  );
  -- 
end entity dwordId_Volatile;
architecture dwordId_Volatile_arch of dwordId_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(36-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal pa_buffer :  std_logic_vector(35 downto 0);
  -- output port buffer signals
  signal dword_id_buffer :  std_logic_vector(2 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  pa_buffer <= pa;
  -- output handling  -------------------------------------------------------
  dword_id <= dword_id_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    -- 
  begin -- 
    -- flow-through slice operator slice_2629_inst
    dword_id_buffer <= pa_buffer(5 downto 3);
    -- 
  end Block; -- data_path
  -- 
end dwordId_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library l2_cache_lib;
use l2_cache_lib.l2_cache_global_package.all;
entity extractDword_Volatile is -- 
  port ( -- 
    dword_id : in  std_logic_vector(2 downto 0);
    cache_line : in  std_logic_vector(511 downto 0);
    dword : out  std_logic_vector(63 downto 0)-- 
  );
  -- 
end entity extractDword_Volatile;
architecture extractDword_Volatile_arch of extractDword_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(515-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal dword_id_buffer :  std_logic_vector(2 downto 0);
  signal cache_line_buffer :  std_logic_vector(511 downto 0);
  -- output port buffer signals
  signal dword_buffer :  std_logic_vector(63 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  dword_id_buffer <= dword_id;
  cache_line_buffer <= cache_line;
  -- output handling  -------------------------------------------------------
  dword <= dword_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal MUX_2712_wire : std_logic_vector(63 downto 0);
    signal MUX_2716_wire : std_logic_vector(63 downto 0);
    signal MUX_2721_wire : std_logic_vector(63 downto 0);
    signal MUX_2725_wire : std_logic_vector(63 downto 0);
    signal MUX_2731_wire : std_logic_vector(63 downto 0);
    signal MUX_2735_wire : std_logic_vector(63 downto 0);
    signal MUX_2740_wire : std_logic_vector(63 downto 0);
    signal MUX_2744_wire : std_logic_vector(63 downto 0);
    signal OR_u64_u64_2717_wire : std_logic_vector(63 downto 0);
    signal OR_u64_u64_2726_wire : std_logic_vector(63 downto 0);
    signal OR_u64_u64_2727_wire : std_logic_vector(63 downto 0);
    signal OR_u64_u64_2736_wire : std_logic_vector(63 downto 0);
    signal OR_u64_u64_2745_wire : std_logic_vector(63 downto 0);
    signal OR_u64_u64_2746_wire : std_logic_vector(63 downto 0);
    signal d0_2639 : std_logic_vector(63 downto 0);
    signal d1_2643 : std_logic_vector(63 downto 0);
    signal d2_2647 : std_logic_vector(63 downto 0);
    signal d3_2651 : std_logic_vector(63 downto 0);
    signal d4_2655 : std_logic_vector(63 downto 0);
    signal d5_2659 : std_logic_vector(63 downto 0);
    signal d6_2663 : std_logic_vector(63 downto 0);
    signal d7_2667 : std_logic_vector(63 downto 0);
    signal konst_2670_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2675_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2680_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2685_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2690_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2695_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2700_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2705_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2711_wire_constant : std_logic_vector(63 downto 0);
    signal konst_2715_wire_constant : std_logic_vector(63 downto 0);
    signal konst_2720_wire_constant : std_logic_vector(63 downto 0);
    signal konst_2724_wire_constant : std_logic_vector(63 downto 0);
    signal konst_2730_wire_constant : std_logic_vector(63 downto 0);
    signal konst_2734_wire_constant : std_logic_vector(63 downto 0);
    signal konst_2739_wire_constant : std_logic_vector(63 downto 0);
    signal konst_2743_wire_constant : std_logic_vector(63 downto 0);
    signal s0_2672 : std_logic_vector(0 downto 0);
    signal s1_2677 : std_logic_vector(0 downto 0);
    signal s2_2682 : std_logic_vector(0 downto 0);
    signal s3_2687 : std_logic_vector(0 downto 0);
    signal s4_2692 : std_logic_vector(0 downto 0);
    signal s5_2697 : std_logic_vector(0 downto 0);
    signal s6_2702 : std_logic_vector(0 downto 0);
    signal s7_2707 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    konst_2670_wire_constant <= "000";
    konst_2675_wire_constant <= "001";
    konst_2680_wire_constant <= "010";
    konst_2685_wire_constant <= "011";
    konst_2690_wire_constant <= "100";
    konst_2695_wire_constant <= "101";
    konst_2700_wire_constant <= "110";
    konst_2705_wire_constant <= "111";
    konst_2711_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_2715_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_2720_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_2724_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_2730_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_2734_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_2739_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    konst_2743_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    -- flow-through select operator MUX_2712_inst
    MUX_2712_wire <= d0_2639 when (s0_2672(0) /=  '0') else konst_2711_wire_constant;
    -- flow-through select operator MUX_2716_inst
    MUX_2716_wire <= d1_2643 when (s1_2677(0) /=  '0') else konst_2715_wire_constant;
    -- flow-through select operator MUX_2721_inst
    MUX_2721_wire <= d2_2647 when (s2_2682(0) /=  '0') else konst_2720_wire_constant;
    -- flow-through select operator MUX_2725_inst
    MUX_2725_wire <= d3_2651 when (s3_2687(0) /=  '0') else konst_2724_wire_constant;
    -- flow-through select operator MUX_2731_inst
    MUX_2731_wire <= d4_2655 when (s4_2692(0) /=  '0') else konst_2730_wire_constant;
    -- flow-through select operator MUX_2735_inst
    MUX_2735_wire <= d5_2659 when (s5_2697(0) /=  '0') else konst_2734_wire_constant;
    -- flow-through select operator MUX_2740_inst
    MUX_2740_wire <= d6_2663 when (s6_2702(0) /=  '0') else konst_2739_wire_constant;
    -- flow-through select operator MUX_2744_inst
    MUX_2744_wire <= d7_2667 when (s7_2707(0) /=  '0') else konst_2743_wire_constant;
    -- flow-through slice operator slice_2638_inst
    d0_2639 <= cache_line_buffer(511 downto 448);
    -- flow-through slice operator slice_2642_inst
    d1_2643 <= cache_line_buffer(447 downto 384);
    -- flow-through slice operator slice_2646_inst
    d2_2647 <= cache_line_buffer(383 downto 320);
    -- flow-through slice operator slice_2650_inst
    d3_2651 <= cache_line_buffer(319 downto 256);
    -- flow-through slice operator slice_2654_inst
    d4_2655 <= cache_line_buffer(255 downto 192);
    -- flow-through slice operator slice_2658_inst
    d5_2659 <= cache_line_buffer(191 downto 128);
    -- flow-through slice operator slice_2662_inst
    d6_2663 <= cache_line_buffer(127 downto 64);
    -- flow-through slice operator slice_2666_inst
    d7_2667 <= cache_line_buffer(63 downto 0);
    -- binary operator EQ_u3_u1_2671_inst
    process(dword_id_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dword_id_buffer, konst_2670_wire_constant, tmp_var);
      s0_2672 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_2676_inst
    process(dword_id_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dword_id_buffer, konst_2675_wire_constant, tmp_var);
      s1_2677 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_2681_inst
    process(dword_id_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dword_id_buffer, konst_2680_wire_constant, tmp_var);
      s2_2682 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_2686_inst
    process(dword_id_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dword_id_buffer, konst_2685_wire_constant, tmp_var);
      s3_2687 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_2691_inst
    process(dword_id_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dword_id_buffer, konst_2690_wire_constant, tmp_var);
      s4_2692 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_2696_inst
    process(dword_id_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dword_id_buffer, konst_2695_wire_constant, tmp_var);
      s5_2697 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_2701_inst
    process(dword_id_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dword_id_buffer, konst_2700_wire_constant, tmp_var);
      s6_2702 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_2706_inst
    process(dword_id_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dword_id_buffer, konst_2705_wire_constant, tmp_var);
      s7_2707 <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2717_inst
    process(MUX_2712_wire, MUX_2716_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_2712_wire, MUX_2716_wire, tmp_var);
      OR_u64_u64_2717_wire <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2726_inst
    process(MUX_2721_wire, MUX_2725_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_2721_wire, MUX_2725_wire, tmp_var);
      OR_u64_u64_2726_wire <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2727_inst
    process(OR_u64_u64_2717_wire, OR_u64_u64_2726_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u64_u64_2717_wire, OR_u64_u64_2726_wire, tmp_var);
      OR_u64_u64_2727_wire <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2736_inst
    process(MUX_2731_wire, MUX_2735_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_2731_wire, MUX_2735_wire, tmp_var);
      OR_u64_u64_2736_wire <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2745_inst
    process(MUX_2740_wire, MUX_2744_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(MUX_2740_wire, MUX_2744_wire, tmp_var);
      OR_u64_u64_2745_wire <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2746_inst
    process(OR_u64_u64_2736_wire, OR_u64_u64_2745_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u64_u64_2736_wire, OR_u64_u64_2745_wire, tmp_var);
      OR_u64_u64_2746_wire <= tmp_var; --
    end process;
    -- binary operator OR_u64_u64_2747_inst
    process(OR_u64_u64_2727_wire, OR_u64_u64_2746_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u64_u64_2727_wire, OR_u64_u64_2746_wire, tmp_var);
      dword_buffer <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end extractDword_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library l2_cache_lib;
use l2_cache_lib.l2_cache_global_package.all;
entity getNextDirtyOffset_Volatile is -- 
  port ( -- 
    first_time : in  std_logic_vector(0 downto 0);
    last_offset : in  std_logic_vector(2 downto 0);
    dirty_mask : in  std_logic_vector(7 downto 0);
    none_found : out  std_logic_vector(0 downto 0);
    current_offset : out  std_logic_vector(2 downto 0)-- 
  );
  -- 
end entity getNextDirtyOffset_Volatile;
architecture getNextDirtyOffset_Volatile_arch of getNextDirtyOffset_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(12-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal first_time_buffer :  std_logic_vector(0 downto 0);
  signal last_offset_buffer :  std_logic_vector(2 downto 0);
  signal dirty_mask_buffer :  std_logic_vector(7 downto 0);
  -- output port buffer signals
  signal none_found_buffer :  std_logic_vector(0 downto 0);
  signal current_offset_buffer :  std_logic_vector(2 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  first_time_buffer <= first_time;
  last_offset_buffer <= last_offset;
  dirty_mask_buffer <= dirty_mask;
  -- output handling  -------------------------------------------------------
  none_found <= none_found_buffer;
  current_offset <= current_offset_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal ADD_u3_u3_2762_wire : std_logic_vector(2 downto 0);
    signal EQ_u3_u1_2858_wire : std_logic_vector(0 downto 0);
    signal EQ_u8_u1_2855_wire : std_logic_vector(0 downto 0);
    signal MUX_2806_wire : std_logic_vector(2 downto 0);
    signal MUX_2811_wire : std_logic_vector(2 downto 0);
    signal MUX_2816_wire : std_logic_vector(2 downto 0);
    signal MUX_2821_wire : std_logic_vector(2 downto 0);
    signal MUX_2826_wire : std_logic_vector(2 downto 0);
    signal MUX_2831_wire : std_logic_vector(2 downto 0);
    signal MUX_2836_wire : std_logic_vector(2 downto 0);
    signal MUX_2841_wire : std_logic_vector(2 downto 0);
    signal MUX_2843_wire : std_logic_vector(2 downto 0);
    signal MUX_2844_wire : std_logic_vector(2 downto 0);
    signal MUX_2845_wire : std_logic_vector(2 downto 0);
    signal MUX_2846_wire : std_logic_vector(2 downto 0);
    signal MUX_2847_wire : std_logic_vector(2 downto 0);
    signal MUX_2848_wire : std_logic_vector(2 downto 0);
    signal MUX_2849_wire : std_logic_vector(2 downto 0);
    signal SHL_u8_u8_2764_wire : std_logic_vector(7 downto 0);
    signal index_2851 : std_logic_vector(2 downto 0);
    signal konst_2761_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2809_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2810_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2814_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2815_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2819_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2820_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2824_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2825_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2829_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2830_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2834_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2835_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2839_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2840_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2842_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2854_wire_constant : std_logic_vector(7 downto 0);
    signal konst_2857_wire_constant : std_logic_vector(2 downto 0);
    signal s0_2770 : std_logic_vector(0 downto 0);
    signal s1_2774 : std_logic_vector(0 downto 0);
    signal s2_2778 : std_logic_vector(0 downto 0);
    signal s3_2782 : std_logic_vector(0 downto 0);
    signal s4_2786 : std_logic_vector(0 downto 0);
    signal s5_2790 : std_logic_vector(0 downto 0);
    signal s6_2794 : std_logic_vector(0 downto 0);
    signal s7_2798 : std_logic_vector(0 downto 0);
    signal shifted_mask_2766 : std_logic_vector(7 downto 0);
    signal type_cast_2763_wire : std_logic_vector(7 downto 0);
    signal type_cast_2803_wire_constant : std_logic_vector(2 downto 0);
    signal type_cast_2805_wire_constant : std_logic_vector(2 downto 0);
    -- 
  begin -- 
    konst_2761_wire_constant <= "001";
    konst_2809_wire_constant <= "001";
    konst_2810_wire_constant <= "010";
    konst_2814_wire_constant <= "010";
    konst_2815_wire_constant <= "011";
    konst_2819_wire_constant <= "011";
    konst_2820_wire_constant <= "100";
    konst_2824_wire_constant <= "100";
    konst_2825_wire_constant <= "101";
    konst_2829_wire_constant <= "101";
    konst_2830_wire_constant <= "110";
    konst_2834_wire_constant <= "110";
    konst_2835_wire_constant <= "111";
    konst_2839_wire_constant <= "111";
    konst_2840_wire_constant <= "000";
    konst_2842_wire_constant <= "000";
    konst_2854_wire_constant <= "00000000";
    konst_2857_wire_constant <= "111";
    type_cast_2803_wire_constant <= "000";
    type_cast_2805_wire_constant <= "001";
    -- flow-through select operator MUX_2765_inst
    shifted_mask_2766 <= dirty_mask_buffer when (first_time_buffer(0) /=  '0') else SHL_u8_u8_2764_wire;
    -- flow-through select operator MUX_2806_inst
    MUX_2806_wire <= type_cast_2803_wire_constant when (first_time_buffer(0) /=  '0') else type_cast_2805_wire_constant;
    -- flow-through select operator MUX_2811_inst
    MUX_2811_wire <= konst_2809_wire_constant when (first_time_buffer(0) /=  '0') else konst_2810_wire_constant;
    -- flow-through select operator MUX_2816_inst
    MUX_2816_wire <= konst_2814_wire_constant when (first_time_buffer(0) /=  '0') else konst_2815_wire_constant;
    -- flow-through select operator MUX_2821_inst
    MUX_2821_wire <= konst_2819_wire_constant when (first_time_buffer(0) /=  '0') else konst_2820_wire_constant;
    -- flow-through select operator MUX_2826_inst
    MUX_2826_wire <= konst_2824_wire_constant when (first_time_buffer(0) /=  '0') else konst_2825_wire_constant;
    -- flow-through select operator MUX_2831_inst
    MUX_2831_wire <= konst_2829_wire_constant when (first_time_buffer(0) /=  '0') else konst_2830_wire_constant;
    -- flow-through select operator MUX_2836_inst
    MUX_2836_wire <= konst_2834_wire_constant when (first_time_buffer(0) /=  '0') else konst_2835_wire_constant;
    -- flow-through select operator MUX_2841_inst
    MUX_2841_wire <= konst_2839_wire_constant when (first_time_buffer(0) /=  '0') else konst_2840_wire_constant;
    -- flow-through select operator MUX_2843_inst
    MUX_2843_wire <= MUX_2841_wire when (s7_2798(0) /=  '0') else konst_2842_wire_constant;
    -- flow-through select operator MUX_2844_inst
    MUX_2844_wire <= MUX_2836_wire when (s6_2794(0) /=  '0') else MUX_2843_wire;
    -- flow-through select operator MUX_2845_inst
    MUX_2845_wire <= MUX_2831_wire when (s5_2790(0) /=  '0') else MUX_2844_wire;
    -- flow-through select operator MUX_2846_inst
    MUX_2846_wire <= MUX_2826_wire when (s4_2786(0) /=  '0') else MUX_2845_wire;
    -- flow-through select operator MUX_2847_inst
    MUX_2847_wire <= MUX_2821_wire when (s3_2782(0) /=  '0') else MUX_2846_wire;
    -- flow-through select operator MUX_2848_inst
    MUX_2848_wire <= MUX_2816_wire when (s2_2778(0) /=  '0') else MUX_2847_wire;
    -- flow-through select operator MUX_2849_inst
    MUX_2849_wire <= MUX_2811_wire when (s1_2774(0) /=  '0') else MUX_2848_wire;
    -- flow-through select operator MUX_2850_inst
    index_2851 <= MUX_2806_wire when (s0_2770(0) /=  '0') else MUX_2849_wire;
    -- flow-through slice operator slice_2769_inst
    s0_2770 <= shifted_mask_2766(7 downto 7);
    -- flow-through slice operator slice_2773_inst
    s1_2774 <= shifted_mask_2766(6 downto 6);
    -- flow-through slice operator slice_2777_inst
    s2_2778 <= shifted_mask_2766(5 downto 5);
    -- flow-through slice operator slice_2781_inst
    s3_2782 <= shifted_mask_2766(4 downto 4);
    -- flow-through slice operator slice_2785_inst
    s4_2786 <= shifted_mask_2766(3 downto 3);
    -- flow-through slice operator slice_2789_inst
    s5_2790 <= shifted_mask_2766(2 downto 2);
    -- flow-through slice operator slice_2793_inst
    s6_2794 <= shifted_mask_2766(1 downto 1);
    -- flow-through slice operator slice_2797_inst
    s7_2798 <= shifted_mask_2766(0 downto 0);
    -- interlock type_cast_2763_inst
    process(ADD_u3_u3_2762_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 2 downto 0) := ADD_u3_u3_2762_wire(2 downto 0);
      type_cast_2763_wire <= tmp_var; -- 
    end process;
    -- binary operator ADD_u3_u3_2762_inst
    process(last_offset_buffer) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApIntAdd_proc(last_offset_buffer, konst_2761_wire_constant, tmp_var);
      ADD_u3_u3_2762_wire <= tmp_var; --
    end process;
    -- binary operator ADD_u3_u3_2864_inst
    process(last_offset_buffer, index_2851) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApIntAdd_proc(last_offset_buffer, index_2851, tmp_var);
      current_offset_buffer <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_2858_inst
    process(last_offset_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(last_offset_buffer, konst_2857_wire_constant, tmp_var);
      EQ_u3_u1_2858_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u8_u1_2855_inst
    process(shifted_mask_2766) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(shifted_mask_2766, konst_2854_wire_constant, tmp_var);
      EQ_u8_u1_2855_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_2859_inst
    process(EQ_u8_u1_2855_wire, EQ_u3_u1_2858_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(EQ_u8_u1_2855_wire, EQ_u3_u1_2858_wire, tmp_var);
      none_found_buffer <= tmp_var; --
    end process;
    -- binary operator SHL_u8_u8_2764_inst
    process(dirty_mask_buffer, type_cast_2763_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntSHL_proc(dirty_mask_buffer, type_cast_2763_wire, tmp_var);
      SHL_u8_u8_2764_wire <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end getNextDirtyOffset_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library l2_cache_lib;
use l2_cache_lib.l2_cache_global_package.all;
entity insBytes_Volatile is -- 
  port ( -- 
    dword : in  std_logic_vector(63 downto 0);
    bmask : in  std_logic_vector(7 downto 0);
    w_dword : in  std_logic_vector(63 downto 0);
    updated_dword : out  std_logic_vector(63 downto 0)-- 
  );
  -- 
end entity insBytes_Volatile;
architecture insBytes_Volatile_arch of insBytes_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(136-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal dword_buffer :  std_logic_vector(63 downto 0);
  signal bmask_buffer :  std_logic_vector(7 downto 0);
  signal w_dword_buffer :  std_logic_vector(63 downto 0);
  -- output port buffer signals
  signal updated_dword_buffer :  std_logic_vector(63 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  dword_buffer <= dword;
  bmask_buffer <= bmask;
  w_dword_buffer <= w_dword;
  -- output handling  -------------------------------------------------------
  updated_dword <= updated_dword_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u16_u32_316_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_335_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u8_u16_306_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_315_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_325_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_334_wire : std_logic_vector(15 downto 0);
    signal MUX_301_wire : std_logic_vector(7 downto 0);
    signal MUX_305_wire : std_logic_vector(7 downto 0);
    signal MUX_310_wire : std_logic_vector(7 downto 0);
    signal MUX_314_wire : std_logic_vector(7 downto 0);
    signal MUX_320_wire : std_logic_vector(7 downto 0);
    signal MUX_324_wire : std_logic_vector(7 downto 0);
    signal MUX_329_wire : std_logic_vector(7 downto 0);
    signal MUX_333_wire : std_logic_vector(7 downto 0);
    signal b0_204 : std_logic_vector(7 downto 0);
    signal b1_208 : std_logic_vector(7 downto 0);
    signal b2_212 : std_logic_vector(7 downto 0);
    signal b3_216 : std_logic_vector(7 downto 0);
    signal b4_220 : std_logic_vector(7 downto 0);
    signal b5_224 : std_logic_vector(7 downto 0);
    signal b6_228 : std_logic_vector(7 downto 0);
    signal b7_232 : std_logic_vector(7 downto 0);
    signal m0_236 : std_logic_vector(0 downto 0);
    signal m1_240 : std_logic_vector(0 downto 0);
    signal m2_244 : std_logic_vector(0 downto 0);
    signal m3_248 : std_logic_vector(0 downto 0);
    signal m4_252 : std_logic_vector(0 downto 0);
    signal m5_256 : std_logic_vector(0 downto 0);
    signal m6_260 : std_logic_vector(0 downto 0);
    signal m7_264 : std_logic_vector(0 downto 0);
    signal w0_268 : std_logic_vector(7 downto 0);
    signal w1_272 : std_logic_vector(7 downto 0);
    signal w2_276 : std_logic_vector(7 downto 0);
    signal w3_280 : std_logic_vector(7 downto 0);
    signal w4_284 : std_logic_vector(7 downto 0);
    signal w5_288 : std_logic_vector(7 downto 0);
    signal w6_292 : std_logic_vector(7 downto 0);
    signal w7_296 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    -- flow-through select operator MUX_301_inst
    MUX_301_wire <= w0_268 when (m0_236(0) /=  '0') else b0_204;
    -- flow-through select operator MUX_305_inst
    MUX_305_wire <= w1_272 when (m1_240(0) /=  '0') else b1_208;
    -- flow-through select operator MUX_310_inst
    MUX_310_wire <= w2_276 when (m2_244(0) /=  '0') else b2_212;
    -- flow-through select operator MUX_314_inst
    MUX_314_wire <= w3_280 when (m3_248(0) /=  '0') else b3_216;
    -- flow-through select operator MUX_320_inst
    MUX_320_wire <= w4_284 when (m4_252(0) /=  '0') else b4_220;
    -- flow-through select operator MUX_324_inst
    MUX_324_wire <= w5_288 when (m5_256(0) /=  '0') else b5_224;
    -- flow-through select operator MUX_329_inst
    MUX_329_wire <= w6_292 when (m6_260(0) /=  '0') else b6_228;
    -- flow-through select operator MUX_333_inst
    MUX_333_wire <= w7_296 when (m7_264(0) /=  '0') else b7_232;
    -- flow-through slice operator slice_203_inst
    b0_204 <= dword_buffer(63 downto 56);
    -- flow-through slice operator slice_207_inst
    b1_208 <= dword_buffer(55 downto 48);
    -- flow-through slice operator slice_211_inst
    b2_212 <= dword_buffer(47 downto 40);
    -- flow-through slice operator slice_215_inst
    b3_216 <= dword_buffer(39 downto 32);
    -- flow-through slice operator slice_219_inst
    b4_220 <= dword_buffer(31 downto 24);
    -- flow-through slice operator slice_223_inst
    b5_224 <= dword_buffer(23 downto 16);
    -- flow-through slice operator slice_227_inst
    b6_228 <= dword_buffer(15 downto 8);
    -- flow-through slice operator slice_231_inst
    b7_232 <= dword_buffer(7 downto 0);
    -- flow-through slice operator slice_235_inst
    m0_236 <= bmask_buffer(7 downto 7);
    -- flow-through slice operator slice_239_inst
    m1_240 <= bmask_buffer(6 downto 6);
    -- flow-through slice operator slice_243_inst
    m2_244 <= bmask_buffer(5 downto 5);
    -- flow-through slice operator slice_247_inst
    m3_248 <= bmask_buffer(4 downto 4);
    -- flow-through slice operator slice_251_inst
    m4_252 <= bmask_buffer(3 downto 3);
    -- flow-through slice operator slice_255_inst
    m5_256 <= bmask_buffer(2 downto 2);
    -- flow-through slice operator slice_259_inst
    m6_260 <= bmask_buffer(1 downto 1);
    -- flow-through slice operator slice_263_inst
    m7_264 <= bmask_buffer(0 downto 0);
    -- flow-through slice operator slice_267_inst
    w0_268 <= w_dword_buffer(63 downto 56);
    -- flow-through slice operator slice_271_inst
    w1_272 <= w_dword_buffer(55 downto 48);
    -- flow-through slice operator slice_275_inst
    w2_276 <= w_dword_buffer(47 downto 40);
    -- flow-through slice operator slice_279_inst
    w3_280 <= w_dword_buffer(39 downto 32);
    -- flow-through slice operator slice_283_inst
    w4_284 <= w_dword_buffer(31 downto 24);
    -- flow-through slice operator slice_287_inst
    w5_288 <= w_dword_buffer(23 downto 16);
    -- flow-through slice operator slice_291_inst
    w6_292 <= w_dword_buffer(15 downto 8);
    -- flow-through slice operator slice_295_inst
    w7_296 <= w_dword_buffer(7 downto 0);
    -- binary operator CONCAT_u16_u32_316_inst
    process(CONCAT_u8_u16_306_wire, CONCAT_u8_u16_315_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_306_wire, CONCAT_u8_u16_315_wire, tmp_var);
      CONCAT_u16_u32_316_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_335_inst
    process(CONCAT_u8_u16_325_wire, CONCAT_u8_u16_334_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_325_wire, CONCAT_u8_u16_334_wire, tmp_var);
      CONCAT_u16_u32_335_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u32_u64_336_inst
    process(CONCAT_u16_u32_316_wire, CONCAT_u16_u32_335_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u16_u32_316_wire, CONCAT_u16_u32_335_wire, tmp_var);
      updated_dword_buffer <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u16_306_inst
    process(MUX_301_wire, MUX_305_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_301_wire, MUX_305_wire, tmp_var);
      CONCAT_u8_u16_306_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u16_315_inst
    process(MUX_310_wire, MUX_314_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_310_wire, MUX_314_wire, tmp_var);
      CONCAT_u8_u16_315_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u16_325_inst
    process(MUX_320_wire, MUX_324_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_320_wire, MUX_324_wire, tmp_var);
      CONCAT_u8_u16_325_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u16_334_inst
    process(MUX_329_wire, MUX_333_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_329_wire, MUX_333_wire, tmp_var);
      CONCAT_u8_u16_334_wire <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end insBytes_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library l2_cache_lib;
use l2_cache_lib.l2_cache_global_package.all;
entity insertIntoSetDirtyDwordMasks_Volatile is -- 
  port ( -- 
    old_set_mask : in  std_logic_vector(63 downto 0);
    index : in  std_logic_vector(2 downto 0);
    ins_mask : in  std_logic_vector(7 downto 0);
    new_set_mask : out  std_logic_vector(63 downto 0)-- 
  );
  -- 
end entity insertIntoSetDirtyDwordMasks_Volatile;
architecture insertIntoSetDirtyDwordMasks_Volatile_arch of insertIntoSetDirtyDwordMasks_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(75-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal old_set_mask_buffer :  std_logic_vector(63 downto 0);
  signal index_buffer :  std_logic_vector(2 downto 0);
  signal ins_mask_buffer :  std_logic_vector(7 downto 0);
  -- output port buffer signals
  signal new_set_mask_buffer :  std_logic_vector(63 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  old_set_mask_buffer <= old_set_mask;
  index_buffer <= index;
  ins_mask_buffer <= ins_mask;
  -- output handling  -------------------------------------------------------
  new_set_mask <= new_set_mask_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u16_u32_2258_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u16_u32_2285_wire : std_logic_vector(31 downto 0);
    signal CONCAT_u8_u16_2244_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_2257_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_2271_wire : std_logic_vector(15 downto 0);
    signal CONCAT_u8_u16_2284_wire : std_logic_vector(15 downto 0);
    signal EQ_u3_u1_2234_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2240_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2247_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2253_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2261_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2267_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2274_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2280_wire : std_logic_vector(0 downto 0);
    signal MUX_2237_wire : std_logic_vector(7 downto 0);
    signal MUX_2243_wire : std_logic_vector(7 downto 0);
    signal MUX_2250_wire : std_logic_vector(7 downto 0);
    signal MUX_2256_wire : std_logic_vector(7 downto 0);
    signal MUX_2264_wire : std_logic_vector(7 downto 0);
    signal MUX_2270_wire : std_logic_vector(7 downto 0);
    signal MUX_2277_wire : std_logic_vector(7 downto 0);
    signal MUX_2283_wire : std_logic_vector(7 downto 0);
    signal konst_2233_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2239_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2246_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2252_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2260_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2266_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2273_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2279_wire_constant : std_logic_vector(2 downto 0);
    signal o0_2202 : std_logic_vector(7 downto 0);
    signal o1_2206 : std_logic_vector(7 downto 0);
    signal o2_2210 : std_logic_vector(7 downto 0);
    signal o3_2214 : std_logic_vector(7 downto 0);
    signal o4_2218 : std_logic_vector(7 downto 0);
    signal o5_2222 : std_logic_vector(7 downto 0);
    signal o6_2226 : std_logic_vector(7 downto 0);
    signal o7_2230 : std_logic_vector(7 downto 0);
    -- 
  begin -- 
    konst_2233_wire_constant <= "000";
    konst_2239_wire_constant <= "001";
    konst_2246_wire_constant <= "010";
    konst_2252_wire_constant <= "011";
    konst_2260_wire_constant <= "100";
    konst_2266_wire_constant <= "101";
    konst_2273_wire_constant <= "110";
    konst_2279_wire_constant <= "111";
    -- flow-through select operator MUX_2237_inst
    MUX_2237_wire <= ins_mask_buffer when (EQ_u3_u1_2234_wire(0) /=  '0') else o0_2202;
    -- flow-through select operator MUX_2243_inst
    MUX_2243_wire <= ins_mask_buffer when (EQ_u3_u1_2240_wire(0) /=  '0') else o1_2206;
    -- flow-through select operator MUX_2250_inst
    MUX_2250_wire <= ins_mask_buffer when (EQ_u3_u1_2247_wire(0) /=  '0') else o2_2210;
    -- flow-through select operator MUX_2256_inst
    MUX_2256_wire <= ins_mask_buffer when (EQ_u3_u1_2253_wire(0) /=  '0') else o3_2214;
    -- flow-through select operator MUX_2264_inst
    MUX_2264_wire <= ins_mask_buffer when (EQ_u3_u1_2261_wire(0) /=  '0') else o4_2218;
    -- flow-through select operator MUX_2270_inst
    MUX_2270_wire <= ins_mask_buffer when (EQ_u3_u1_2267_wire(0) /=  '0') else o5_2222;
    -- flow-through select operator MUX_2277_inst
    MUX_2277_wire <= ins_mask_buffer when (EQ_u3_u1_2274_wire(0) /=  '0') else o6_2226;
    -- flow-through select operator MUX_2283_inst
    MUX_2283_wire <= ins_mask_buffer when (EQ_u3_u1_2280_wire(0) /=  '0') else o7_2230;
    -- flow-through slice operator slice_2201_inst
    o0_2202 <= old_set_mask_buffer(63 downto 56);
    -- flow-through slice operator slice_2205_inst
    o1_2206 <= old_set_mask_buffer(55 downto 48);
    -- flow-through slice operator slice_2209_inst
    o2_2210 <= old_set_mask_buffer(47 downto 40);
    -- flow-through slice operator slice_2213_inst
    o3_2214 <= old_set_mask_buffer(39 downto 32);
    -- flow-through slice operator slice_2217_inst
    o4_2218 <= old_set_mask_buffer(31 downto 24);
    -- flow-through slice operator slice_2221_inst
    o5_2222 <= old_set_mask_buffer(23 downto 16);
    -- flow-through slice operator slice_2225_inst
    o6_2226 <= old_set_mask_buffer(15 downto 8);
    -- flow-through slice operator slice_2229_inst
    o7_2230 <= old_set_mask_buffer(7 downto 0);
    -- binary operator CONCAT_u16_u32_2258_inst
    process(CONCAT_u8_u16_2244_wire, CONCAT_u8_u16_2257_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_2244_wire, CONCAT_u8_u16_2257_wire, tmp_var);
      CONCAT_u16_u32_2258_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u16_u32_2285_inst
    process(CONCAT_u8_u16_2271_wire, CONCAT_u8_u16_2284_wire) -- 
      variable tmp_var : std_logic_vector(31 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u8_u16_2271_wire, CONCAT_u8_u16_2284_wire, tmp_var);
      CONCAT_u16_u32_2285_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u32_u64_2286_inst
    process(CONCAT_u16_u32_2258_wire, CONCAT_u16_u32_2285_wire) -- 
      variable tmp_var : std_logic_vector(63 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u16_u32_2258_wire, CONCAT_u16_u32_2285_wire, tmp_var);
      new_set_mask_buffer <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u16_2244_inst
    process(MUX_2237_wire, MUX_2243_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_2237_wire, MUX_2243_wire, tmp_var);
      CONCAT_u8_u16_2244_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u16_2257_inst
    process(MUX_2250_wire, MUX_2256_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_2250_wire, MUX_2256_wire, tmp_var);
      CONCAT_u8_u16_2257_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u16_2271_inst
    process(MUX_2264_wire, MUX_2270_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_2264_wire, MUX_2270_wire, tmp_var);
      CONCAT_u8_u16_2271_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u8_u16_2284_inst
    process(MUX_2277_wire, MUX_2283_wire) -- 
      variable tmp_var : std_logic_vector(15 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_2277_wire, MUX_2283_wire, tmp_var);
      CONCAT_u8_u16_2284_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_2234_inst
    process(index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(index_buffer, konst_2233_wire_constant, tmp_var);
      EQ_u3_u1_2234_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_2240_inst
    process(index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(index_buffer, konst_2239_wire_constant, tmp_var);
      EQ_u3_u1_2240_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_2247_inst
    process(index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(index_buffer, konst_2246_wire_constant, tmp_var);
      EQ_u3_u1_2247_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_2253_inst
    process(index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(index_buffer, konst_2252_wire_constant, tmp_var);
      EQ_u3_u1_2253_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_2261_inst
    process(index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(index_buffer, konst_2260_wire_constant, tmp_var);
      EQ_u3_u1_2261_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_2267_inst
    process(index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(index_buffer, konst_2266_wire_constant, tmp_var);
      EQ_u3_u1_2267_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_2274_inst
    process(index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(index_buffer, konst_2273_wire_constant, tmp_var);
      EQ_u3_u1_2274_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_2280_inst
    process(index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(index_buffer, konst_2279_wire_constant, tmp_var);
      EQ_u3_u1_2280_wire <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end insertIntoSetDirtyDwordMasks_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library l2_cache_lib;
use l2_cache_lib.l2_cache_global_package.all;
entity l2CacheDaemon is -- 
  generic (tag_length : integer); 
  port ( -- 
    NOBLOCK_L2_REQUEST_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_L2_REQUEST_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_L2_REQUEST_pipe_read_data : in   std_logic_vector(110 downto 0);
    L2_TAGS_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
    L2_TAGS_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
    L2_TAGS_RESPONSE_pipe_read_data : in   std_logic_vector(33 downto 0);
    NOBLOCK_L2_INVALIDATE_pipe_read_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_L2_INVALIDATE_pipe_read_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_L2_INVALIDATE_pipe_read_data : in   std_logic_vector(30 downto 0);
    NOBLOCK_L2_TAGS_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
    NOBLOCK_L2_TAGS_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
    NOBLOCK_L2_TAGS_REQUEST_pipe_write_data : out  std_logic_vector(44 downto 0);
    L2_RESPONSE_pipe_write_req : out  std_logic_vector(0 downto 0);
    L2_RESPONSE_pipe_write_ack : in   std_logic_vector(0 downto 0);
    L2_RESPONSE_pipe_write_data : out  std_logic_vector(64 downto 0);
    L2_TO_L1_INVALIDATE_pipe_write_req : out  std_logic_vector(0 downto 0);
    L2_TO_L1_INVALIDATE_pipe_write_ack : in   std_logic_vector(0 downto 0);
    L2_TO_L1_INVALIDATE_pipe_write_data : out  std_logic_vector(29 downto 0);
    sys_mem_lock_pipe_write_req : out  std_logic_vector(0 downto 0);
    sys_mem_lock_pipe_write_ack : in   std_logic_vector(0 downto 0);
    sys_mem_lock_pipe_write_data : out  std_logic_vector(0 downto 0);
    readMemoryFromL2_call_reqs : out  std_logic_vector(0 downto 0);
    readMemoryFromL2_call_acks : in   std_logic_vector(0 downto 0);
    readMemoryFromL2_call_data : out  std_logic_vector(29 downto 0);
    readMemoryFromL2_call_tag  :  out  std_logic_vector(0 downto 0);
    readMemoryFromL2_return_reqs : out  std_logic_vector(0 downto 0);
    readMemoryFromL2_return_acks : in   std_logic_vector(0 downto 0);
    readMemoryFromL2_return_data : in   std_logic_vector(511 downto 0);
    readMemoryFromL2_return_tag :  in   std_logic_vector(0 downto 0);
    writeMemoryFromL2_call_reqs : out  std_logic_vector(0 downto 0);
    writeMemoryFromL2_call_acks : in   std_logic_vector(0 downto 0);
    writeMemoryFromL2_call_data : out  std_logic_vector(551 downto 0);
    writeMemoryFromL2_call_tag  :  out  std_logic_vector(0 downto 0);
    writeMemoryFromL2_return_reqs : out  std_logic_vector(0 downto 0);
    writeMemoryFromL2_return_acks : in   std_logic_vector(0 downto 0);
    writeMemoryFromL2_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity l2CacheDaemon;
architecture l2CacheDaemon_arch of l2CacheDaemon is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  -- output port buffer signals
  signal l2CacheDaemon_CP_3229_start: Boolean;
  signal l2CacheDaemon_CP_3229_symbol: Boolean;
  -- volatile/operator module components. 
  -- function library module [accessL2DataMemX4096X512] component not printed.
  component paTag_Volatile is -- 
    port ( -- 
      pa : in  std_logic_vector(35 downto 0);
      pa_tag : out  std_logic_vector(20 downto 0)-- 
    );
    -- 
  end component; 
  component readMemoryFromL2 is -- 
    generic (tag_length : integer); 
    port ( -- 
      line_address : in  std_logic_vector(29 downto 0);
      rline : out  std_logic_vector(511 downto 0);
      sys_mem_lock_pipe_read_req : out  std_logic_vector(0 downto 0);
      sys_mem_lock_pipe_read_ack : in   std_logic_vector(0 downto 0);
      sys_mem_lock_pipe_read_data : in   std_logic_vector(0 downto 0);
      accessSysMem_call_reqs : out  std_logic_vector(0 downto 0);
      accessSysMem_call_acks : in   std_logic_vector(0 downto 0);
      accessSysMem_call_data : out  std_logic_vector(108 downto 0);
      accessSysMem_call_tag  :  out  std_logic_vector(0 downto 0);
      accessSysMem_return_reqs : out  std_logic_vector(0 downto 0);
      accessSysMem_return_acks : in   std_logic_vector(0 downto 0);
      accessSysMem_return_data : in   std_logic_vector(63 downto 0);
      accessSysMem_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component dwordId_Volatile is -- 
    port ( -- 
      pa : in  std_logic_vector(35 downto 0);
      dword_id : out  std_logic_vector(2 downto 0)-- 
    );
    -- 
  end component; 
  component setId_Volatile is -- 
    port ( -- 
      pa : in  std_logic_vector(35 downto 0);
      set_id : out  std_logic_vector(8 downto 0)-- 
    );
    -- 
  end component; 
  component lineAddress_Volatile is -- 
    port ( -- 
      pa : in  std_logic_vector(35 downto 0);
      pa_line_address : out  std_logic_vector(29 downto 0)-- 
    );
    -- 
  end component; 
  component writeMemoryFromL2 is -- 
    generic (tag_length : integer); 
    port ( -- 
      release_lock : in  std_logic_vector(0 downto 0);
      do_write : in  std_logic_vector(0 downto 0);
      dirty_word_mask : in  std_logic_vector(7 downto 0);
      line_address : in  std_logic_vector(29 downto 0);
      wline : in  std_logic_vector(511 downto 0);
      sys_mem_lock_pipe_write_req : out  std_logic_vector(0 downto 0);
      sys_mem_lock_pipe_write_ack : in   std_logic_vector(0 downto 0);
      sys_mem_lock_pipe_write_data : out  std_logic_vector(0 downto 0);
      accessSysMem_call_reqs : out  std_logic_vector(0 downto 0);
      accessSysMem_call_acks : in   std_logic_vector(0 downto 0);
      accessSysMem_call_data : out  std_logic_vector(108 downto 0);
      accessSysMem_call_tag  :  out  std_logic_vector(0 downto 0);
      accessSysMem_return_reqs : out  std_logic_vector(0 downto 0);
      accessSysMem_return_acks : in   std_logic_vector(0 downto 0);
      accessSysMem_return_data : in   std_logic_vector(63 downto 0);
      accessSysMem_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal W_wdata_3403_delayed_9_0_3677_inst_ack_0 : boolean;
  signal W_rwbar_3417_delayed_10_0_3700_inst_req_0 : boolean;
  signal W_byte_mask_3400_delayed_9_0_3668_inst_ack_1 : boolean;
  signal W_pa_dword_id_3402_delayed_9_0_3674_inst_ack_0 : boolean;
  signal W_send_response_3424_delayed_10_0_3713_inst_req_1 : boolean;
  signal W_rwbar_3417_delayed_10_0_3700_inst_ack_1 : boolean;
  signal W_send_response_3424_delayed_10_0_3713_inst_ack_1 : boolean;
  signal W_byte_mask_3400_delayed_9_0_3668_inst_req_1 : boolean;
  signal W_call_write_mem_3437_delayed_5_0_3729_inst_req_0 : boolean;
  signal W_call_write_mem_3437_delayed_5_0_3729_inst_ack_0 : boolean;
  signal WPIPE_L2_RESPONSE_3717_inst_req_0 : boolean;
  signal W_pa_dword_id_3402_delayed_9_0_3674_inst_ack_1 : boolean;
  signal call_stmt_3693_call_req_0 : boolean;
  signal WPIPE_L2_RESPONSE_3717_inst_ack_0 : boolean;
  signal W_line_id_3401_delayed_4_0_3671_inst_req_1 : boolean;
  signal call_stmt_3693_call_req_1 : boolean;
  signal W_send_response_3424_delayed_10_0_3713_inst_req_0 : boolean;
  signal W_wdata_3403_delayed_9_0_3677_inst_req_0 : boolean;
  signal W_rwbar_3417_delayed_10_0_3700_inst_ack_0 : boolean;
  signal call_stmt_3693_call_ack_1 : boolean;
  signal WPIPE_sys_mem_lock_3331_inst_req_1 : boolean;
  signal W_wdata_3403_delayed_9_0_3677_inst_ack_1 : boolean;
  signal WPIPE_L2_RESPONSE_3717_inst_ack_1 : boolean;
  signal WPIPE_sys_mem_lock_3331_inst_ack_1 : boolean;
  signal W_line_id_3401_delayed_4_0_3671_inst_ack_1 : boolean;
  signal W_send_response_3424_delayed_10_0_3713_inst_ack_0 : boolean;
  signal W_pa_dword_id_3402_delayed_9_0_3674_inst_req_0 : boolean;
  signal W_pa_dword_id_3402_delayed_9_0_3674_inst_req_1 : boolean;
  signal WPIPE_L2_RESPONSE_3717_inst_req_1 : boolean;
  signal W_call_write_mem_3437_delayed_5_0_3729_inst_req_1 : boolean;
  signal W_call_write_mem_3437_delayed_5_0_3729_inst_ack_1 : boolean;
  signal WPIPE_sys_mem_lock_3331_inst_ack_0 : boolean;
  signal WPIPE_sys_mem_lock_3331_inst_req_0 : boolean;
  signal do_while_stmt_3336_branch_req_0 : boolean;
  signal W_wdata_3403_delayed_9_0_3677_inst_req_1 : boolean;
  signal W_rwbar_3417_delayed_10_0_3700_inst_req_1 : boolean;
  signal call_stmt_3693_call_ack_0 : boolean;
  signal W_line_id_3401_delayed_4_0_3671_inst_req_0 : boolean;
  signal W_line_id_3401_delayed_4_0_3671_inst_ack_0 : boolean;
  signal W_do_read_line_from_mem_3438_delayed_5_0_3732_inst_req_0 : boolean;
  signal phi_stmt_3338_req_1 : boolean;
  signal phi_stmt_3338_req_0 : boolean;
  signal phi_stmt_3338_ack_0 : boolean;
  signal RPIPE_NOBLOCK_L2_REQUEST_3342_inst_req_0 : boolean;
  signal RPIPE_NOBLOCK_L2_REQUEST_3342_inst_ack_0 : boolean;
  signal RPIPE_NOBLOCK_L2_REQUEST_3342_inst_req_1 : boolean;
  signal RPIPE_NOBLOCK_L2_REQUEST_3342_inst_ack_1 : boolean;
  signal phi_stmt_3343_req_1 : boolean;
  signal phi_stmt_3343_req_0 : boolean;
  signal phi_stmt_3343_ack_0 : boolean;
  signal RPIPE_NOBLOCK_L2_INVALIDATE_3346_inst_req_0 : boolean;
  signal RPIPE_NOBLOCK_L2_INVALIDATE_3346_inst_ack_0 : boolean;
  signal RPIPE_NOBLOCK_L2_INVALIDATE_3346_inst_req_1 : boolean;
  signal RPIPE_NOBLOCK_L2_INVALIDATE_3346_inst_ack_1 : boolean;
  signal phi_stmt_3347_req_1 : boolean;
  signal phi_stmt_3347_req_0 : boolean;
  signal phi_stmt_3347_ack_0 : boolean;
  signal nCOUNTER_3447_3351_buf_req_0 : boolean;
  signal nCOUNTER_3447_3351_buf_ack_0 : boolean;
  signal nCOUNTER_3447_3351_buf_req_1 : boolean;
  signal nCOUNTER_3447_3351_buf_ack_1 : boolean;
  signal WPIPE_L2_TO_L1_INVALIDATE_3397_inst_req_0 : boolean;
  signal WPIPE_L2_TO_L1_INVALIDATE_3397_inst_ack_0 : boolean;
  signal WPIPE_L2_TO_L1_INVALIDATE_3397_inst_req_1 : boolean;
  signal WPIPE_L2_TO_L1_INVALIDATE_3397_inst_ack_1 : boolean;
  signal WPIPE_NOBLOCK_L2_TAGS_REQUEST_3490_inst_req_0 : boolean;
  signal WPIPE_NOBLOCK_L2_TAGS_REQUEST_3490_inst_ack_0 : boolean;
  signal WPIPE_NOBLOCK_L2_TAGS_REQUEST_3490_inst_req_1 : boolean;
  signal WPIPE_NOBLOCK_L2_TAGS_REQUEST_3490_inst_ack_1 : boolean;
  signal W_do_read_line_from_mem_3438_delayed_5_0_3732_inst_ack_0 : boolean;
  signal W_do_tag_access_3276_delayed_4_0_3493_inst_req_0 : boolean;
  signal W_do_tag_access_3276_delayed_4_0_3493_inst_ack_0 : boolean;
  signal W_do_tag_access_3276_delayed_4_0_3493_inst_req_1 : boolean;
  signal W_do_tag_access_3276_delayed_4_0_3493_inst_ack_1 : boolean;
  signal RPIPE_L2_TAGS_RESPONSE_3498_inst_req_0 : boolean;
  signal RPIPE_L2_TAGS_RESPONSE_3498_inst_ack_0 : boolean;
  signal RPIPE_L2_TAGS_RESPONSE_3498_inst_req_1 : boolean;
  signal RPIPE_L2_TAGS_RESPONSE_3498_inst_ack_1 : boolean;
  signal W_access_set_id_3302_delayed_5_0_3520_inst_req_0 : boolean;
  signal W_access_set_id_3302_delayed_5_0_3520_inst_ack_0 : boolean;
  signal W_access_set_id_3302_delayed_5_0_3520_inst_req_1 : boolean;
  signal W_access_set_id_3302_delayed_5_0_3520_inst_ack_1 : boolean;
  signal AND_u1_u1_3539_inst_req_0 : boolean;
  signal AND_u1_u1_3539_inst_ack_0 : boolean;
  signal AND_u1_u1_3539_inst_req_1 : boolean;
  signal AND_u1_u1_3539_inst_ack_1 : boolean;
  signal AND_u1_u1_3551_inst_req_0 : boolean;
  signal AND_u1_u1_3551_inst_ack_0 : boolean;
  signal AND_u1_u1_3551_inst_req_1 : boolean;
  signal AND_u1_u1_3551_inst_ack_1 : boolean;
  signal W_do_tag_access_3331_delayed_5_0_3559_inst_req_0 : boolean;
  signal W_do_tag_access_3331_delayed_5_0_3559_inst_ack_0 : boolean;
  signal W_do_tag_access_3331_delayed_5_0_3559_inst_req_1 : boolean;
  signal W_do_tag_access_3331_delayed_5_0_3559_inst_ack_1 : boolean;
  signal W_inv_valid_3337_delayed_5_0_3562_inst_req_0 : boolean;
  signal W_inv_valid_3337_delayed_5_0_3562_inst_ack_0 : boolean;
  signal W_inv_valid_3337_delayed_5_0_3562_inst_req_1 : boolean;
  signal W_inv_valid_3337_delayed_5_0_3562_inst_ack_1 : boolean;
  signal W_valid_3340_delayed_5_0_3565_inst_req_0 : boolean;
  signal W_valid_3340_delayed_5_0_3565_inst_ack_0 : boolean;
  signal W_valid_3340_delayed_5_0_3565_inst_req_1 : boolean;
  signal W_valid_3340_delayed_5_0_3565_inst_ack_1 : boolean;
  signal W_inv_valid_3366_delayed_5_0_3603_inst_req_0 : boolean;
  signal W_inv_valid_3366_delayed_5_0_3603_inst_ack_0 : boolean;
  signal W_inv_valid_3366_delayed_5_0_3603_inst_req_1 : boolean;
  signal W_inv_valid_3366_delayed_5_0_3603_inst_ack_1 : boolean;
  signal W_inv_pa_line_address_3367_delayed_5_0_3606_inst_req_0 : boolean;
  signal W_inv_pa_line_address_3367_delayed_5_0_3606_inst_ack_0 : boolean;
  signal W_inv_pa_line_address_3367_delayed_5_0_3606_inst_req_1 : boolean;
  signal W_inv_pa_line_address_3367_delayed_5_0_3606_inst_ack_1 : boolean;
  signal OR_u1_u1_3618_inst_req_0 : boolean;
  signal OR_u1_u1_3618_inst_ack_0 : boolean;
  signal OR_u1_u1_3618_inst_req_1 : boolean;
  signal OR_u1_u1_3618_inst_ack_1 : boolean;
  signal W_pa_line_address_3381_delayed_5_0_3627_inst_req_0 : boolean;
  signal W_pa_line_address_3381_delayed_5_0_3627_inst_ack_0 : boolean;
  signal W_pa_line_address_3381_delayed_5_0_3627_inst_req_1 : boolean;
  signal W_pa_line_address_3381_delayed_5_0_3627_inst_ack_1 : boolean;
  signal call_stmt_3633_call_req_0 : boolean;
  signal call_stmt_3633_call_ack_0 : boolean;
  signal call_stmt_3633_call_req_1 : boolean;
  signal call_stmt_3633_call_ack_1 : boolean;
  signal W_access_set_id_3386_delayed_5_0_3634_inst_req_0 : boolean;
  signal W_access_set_id_3386_delayed_5_0_3634_inst_ack_0 : boolean;
  signal W_access_set_id_3386_delayed_5_0_3634_inst_req_1 : boolean;
  signal W_access_set_id_3386_delayed_5_0_3634_inst_ack_1 : boolean;
  signal W_data_read_dword_3391_delayed_5_0_3642_inst_req_0 : boolean;
  signal W_data_read_dword_3391_delayed_5_0_3642_inst_ack_0 : boolean;
  signal W_data_read_dword_3391_delayed_5_0_3642_inst_req_1 : boolean;
  signal W_data_read_dword_3391_delayed_5_0_3642_inst_ack_1 : boolean;
  signal W_access_data_mem_3394_delayed_4_0_3650_inst_req_0 : boolean;
  signal W_access_data_mem_3394_delayed_4_0_3650_inst_ack_0 : boolean;
  signal W_access_data_mem_3394_delayed_4_0_3650_inst_req_1 : boolean;
  signal W_access_data_mem_3394_delayed_4_0_3650_inst_ack_1 : boolean;
  signal W_read_data_line_3395_delayed_4_0_3653_inst_req_0 : boolean;
  signal W_read_data_line_3395_delayed_4_0_3653_inst_ack_0 : boolean;
  signal W_read_data_line_3395_delayed_4_0_3653_inst_req_1 : boolean;
  signal W_read_data_line_3395_delayed_4_0_3653_inst_ack_1 : boolean;
  signal W_data_write_dword_3396_delayed_9_0_3656_inst_req_0 : boolean;
  signal W_data_write_dword_3396_delayed_9_0_3656_inst_ack_0 : boolean;
  signal W_data_write_dword_3396_delayed_9_0_3656_inst_req_1 : boolean;
  signal W_data_write_dword_3396_delayed_9_0_3656_inst_ack_1 : boolean;
  signal W_data_read_dword_3397_delayed_9_0_3659_inst_req_0 : boolean;
  signal W_data_read_dword_3397_delayed_9_0_3659_inst_ack_0 : boolean;
  signal W_data_read_dword_3397_delayed_9_0_3659_inst_req_1 : boolean;
  signal W_data_read_dword_3397_delayed_9_0_3659_inst_ack_1 : boolean;
  signal W_data_write_new_line_3398_delayed_4_0_3662_inst_req_0 : boolean;
  signal W_data_write_new_line_3398_delayed_4_0_3662_inst_ack_0 : boolean;
  signal W_data_write_new_line_3398_delayed_4_0_3662_inst_req_1 : boolean;
  signal W_data_write_new_line_3398_delayed_4_0_3662_inst_ack_1 : boolean;
  signal W_do_write_replaced_line_to_mem_3399_delayed_4_0_3665_inst_req_0 : boolean;
  signal W_do_write_replaced_line_to_mem_3399_delayed_4_0_3665_inst_ack_0 : boolean;
  signal W_do_write_replaced_line_to_mem_3399_delayed_4_0_3665_inst_req_1 : boolean;
  signal W_do_write_replaced_line_to_mem_3399_delayed_4_0_3665_inst_ack_1 : boolean;
  signal W_byte_mask_3400_delayed_9_0_3668_inst_req_0 : boolean;
  signal W_byte_mask_3400_delayed_9_0_3668_inst_ack_0 : boolean;
  signal W_do_read_line_from_mem_3438_delayed_5_0_3732_inst_req_1 : boolean;
  signal W_do_read_line_from_mem_3438_delayed_5_0_3732_inst_ack_1 : boolean;
  signal W_do_write_replaced_line_to_mem_3439_delayed_5_0_3735_inst_req_0 : boolean;
  signal W_do_write_replaced_line_to_mem_3439_delayed_5_0_3735_inst_ack_0 : boolean;
  signal W_do_write_replaced_line_to_mem_3439_delayed_5_0_3735_inst_req_1 : boolean;
  signal W_do_write_replaced_line_to_mem_3439_delayed_5_0_3735_inst_ack_1 : boolean;
  signal W_dirty_word_mask_3440_delayed_5_0_3738_inst_req_0 : boolean;
  signal W_dirty_word_mask_3440_delayed_5_0_3738_inst_ack_0 : boolean;
  signal W_dirty_word_mask_3440_delayed_5_0_3738_inst_req_1 : boolean;
  signal W_dirty_word_mask_3440_delayed_5_0_3738_inst_ack_1 : boolean;
  signal W_write_back_line_address_3441_delayed_5_0_3741_inst_req_0 : boolean;
  signal W_write_back_line_address_3441_delayed_5_0_3741_inst_ack_0 : boolean;
  signal W_write_back_line_address_3441_delayed_5_0_3741_inst_req_1 : boolean;
  signal W_write_back_line_address_3441_delayed_5_0_3741_inst_ack_1 : boolean;
  signal call_stmt_3750_call_req_0 : boolean;
  signal call_stmt_3750_call_ack_0 : boolean;
  signal call_stmt_3750_call_req_1 : boolean;
  signal call_stmt_3750_call_ack_1 : boolean;
  signal do_while_stmt_3336_branch_ack_0 : boolean;
  signal do_while_stmt_3336_branch_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "l2CacheDaemon_input_buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      data_width => tag_length + 0) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(tag_length-1 downto 0) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length-1 downto 0);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  l2CacheDaemon_CP_3229_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "l2CacheDaemon_out_buffer", -- 
      buffer_size => 1,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= l2CacheDaemon_CP_3229_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= l2CacheDaemon_CP_3229_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= l2CacheDaemon_CP_3229_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  l2CacheDaemon_CP_3229: Block -- control-path 
    signal l2CacheDaemon_CP_3229_elements: BooleanArray(226 downto 0);
    -- 
  begin -- 
    l2CacheDaemon_CP_3229_elements(0) <= l2CacheDaemon_CP_3229_start;
    l2CacheDaemon_CP_3229_symbol <= l2CacheDaemon_CP_3229_elements(3);
    -- CP-element group 0:  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 assign_stmt_3334/WPIPE_sys_mem_lock_3331_sample_start_
      -- CP-element group 0: 	 assign_stmt_3334/$entry
      -- CP-element group 0: 	 assign_stmt_3334/WPIPE_sys_mem_lock_3331_Sample/req
      -- CP-element group 0: 	 assign_stmt_3334/WPIPE_sys_mem_lock_3331_Sample/$entry
      -- CP-element group 0: 	 $entry
      -- 
    req_3242_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3242_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(0), ack => WPIPE_sys_mem_lock_3331_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_3334/WPIPE_sys_mem_lock_3331_sample_completed_
      -- CP-element group 1: 	 assign_stmt_3334/WPIPE_sys_mem_lock_3331_Update/req
      -- CP-element group 1: 	 assign_stmt_3334/WPIPE_sys_mem_lock_3331_Update/$entry
      -- CP-element group 1: 	 assign_stmt_3334/WPIPE_sys_mem_lock_3331_Sample/ack
      -- CP-element group 1: 	 assign_stmt_3334/WPIPE_sys_mem_lock_3331_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_3334/WPIPE_sys_mem_lock_3331_update_start_
      -- 
    ack_3243_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_sys_mem_lock_3331_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(1)); -- 
    req_3247_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3247_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(1), ack => WPIPE_sys_mem_lock_3331_inst_req_1); -- 
    -- CP-element group 2:  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	4 
    -- CP-element group 2:  members (7) 
      -- CP-element group 2: 	 branch_block_stmt_3335/branch_block_stmt_3335__entry__
      -- CP-element group 2: 	 branch_block_stmt_3335/$entry
      -- CP-element group 2: 	 assign_stmt_3334/WPIPE_sys_mem_lock_3331_Update/ack
      -- CP-element group 2: 	 assign_stmt_3334/$exit
      -- CP-element group 2: 	 branch_block_stmt_3335/do_while_stmt_3336__entry__
      -- CP-element group 2: 	 assign_stmt_3334/WPIPE_sys_mem_lock_3331_Update/$exit
      -- CP-element group 2: 	 assign_stmt_3334/WPIPE_sys_mem_lock_3331_update_completed_
      -- 
    ack_3248_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_sys_mem_lock_3331_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(2)); -- 
    -- CP-element group 3:  transition  place  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	226 
    -- CP-element group 3: successors 
    -- CP-element group 3:  members (4) 
      -- CP-element group 3: 	 branch_block_stmt_3335/do_while_stmt_3336__exit__
      -- CP-element group 3: 	 branch_block_stmt_3335/branch_block_stmt_3335__exit__
      -- CP-element group 3: 	 $exit
      -- CP-element group 3: 	 branch_block_stmt_3335/$exit
      -- 
    l2CacheDaemon_CP_3229_elements(3) <= l2CacheDaemon_CP_3229_elements(226);
    -- CP-element group 4:  transition  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	10 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336__entry__
      -- CP-element group 4: 	 branch_block_stmt_3335/do_while_stmt_3336/$entry
      -- 
    l2CacheDaemon_CP_3229_elements(4) <= l2CacheDaemon_CP_3229_elements(2);
    -- CP-element group 5:  merge  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	226 
    -- CP-element group 5:  members (1) 
      -- CP-element group 5: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336__exit__
      -- 
    -- Element group l2CacheDaemon_CP_3229_elements(5) is bound as output of CP function.
    -- CP-element group 6:  merge  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_3335/do_while_stmt_3336/loop_back
      -- 
    -- Element group l2CacheDaemon_CP_3229_elements(6) is bound as output of CP function.
    -- CP-element group 7:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	12 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	224 
    -- CP-element group 7: 	225 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_3335/do_while_stmt_3336/condition_done
      -- CP-element group 7: 	 branch_block_stmt_3335/do_while_stmt_3336/loop_exit/$entry
      -- CP-element group 7: 	 branch_block_stmt_3335/do_while_stmt_3336/loop_taken/$entry
      -- 
    l2CacheDaemon_CP_3229_elements(7) <= l2CacheDaemon_CP_3229_elements(12);
    -- CP-element group 8:  branch  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	223 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_3335/do_while_stmt_3336/loop_body_done
      -- 
    l2CacheDaemon_CP_3229_elements(8) <= l2CacheDaemon_CP_3229_elements(223);
    -- CP-element group 9:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	22 
    -- CP-element group 9: 	43 
    -- CP-element group 9: 	64 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/back_edge_to_loop_body
      -- 
    l2CacheDaemon_CP_3229_elements(9) <= l2CacheDaemon_CP_3229_elements(6);
    -- CP-element group 10:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	4 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	24 
    -- CP-element group 10: 	45 
    -- CP-element group 10: 	66 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/first_time_through_loop_body
      -- 
    l2CacheDaemon_CP_3229_elements(10) <= l2CacheDaemon_CP_3229_elements(4);
    -- CP-element group 11:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	18 
    -- CP-element group 11: 	19 
    -- CP-element group 11: 	37 
    -- CP-element group 11: 	38 
    -- CP-element group 11: 	58 
    -- CP-element group 11: 	222 
    -- CP-element group 11: 	59 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/$entry
      -- CP-element group 11: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/loop_body_start
      -- 
    -- Element group l2CacheDaemon_CP_3229_elements(11) is bound as output of CP function.
    -- CP-element group 12:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	15 
    -- CP-element group 12: 	17 
    -- CP-element group 12: 	222 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	7 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/condition_evaluated
      -- 
    condition_evaluated_3270_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_3270_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(12), ack => do_while_stmt_3336_branch_req_0); -- 
    l2CacheDaemon_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "l2CacheDaemon_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(15) & l2CacheDaemon_CP_3229_elements(17) & l2CacheDaemon_CP_3229_elements(222);
      gj_l2CacheDaemon_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	18 
    -- CP-element group 13: 	37 
    -- CP-element group 13: 	58 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	17 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	39 
    -- CP-element group 13: 	60 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3338_sample_start__ps
      -- CP-element group 13: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/aggregated_phi_sample_req
      -- 
    l2CacheDaemon_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "l2CacheDaemon_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(18) & l2CacheDaemon_CP_3229_elements(37) & l2CacheDaemon_CP_3229_elements(58) & l2CacheDaemon_CP_3229_elements(17);
      gj_l2CacheDaemon_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	20 
    -- CP-element group 14: 	40 
    -- CP-element group 14: 	61 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	15 
    -- CP-element group 14: 	223 
    -- CP-element group 14: marked-successors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: 	37 
    -- CP-element group 14: 	58 
    -- CP-element group 14:  members (4) 
      -- CP-element group 14: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3338_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/aggregated_phi_sample_ack
      -- CP-element group 14: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3343_sample_completed_
      -- CP-element group 14: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3347_sample_completed_
      -- 
    l2CacheDaemon_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "l2CacheDaemon_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(20) & l2CacheDaemon_CP_3229_elements(40) & l2CacheDaemon_CP_3229_elements(61);
      gj_l2CacheDaemon_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	14 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	12 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/aggregated_phi_sample_ack_d
      -- 
    -- Element group l2CacheDaemon_CP_3229_elements(15) is a control-delay.
    cp_element_15_delay: control_delay_element  generic map(name => " 15_delay", delay_value => 1)  port map(req => l2CacheDaemon_CP_3229_elements(14), ack => l2CacheDaemon_CP_3229_elements(15), clk => clk, reset =>reset);
    -- CP-element group 16:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	19 
    -- CP-element group 16: 	38 
    -- CP-element group 16: 	59 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	41 
    -- CP-element group 16: 	62 
    -- CP-element group 16:  members (2) 
      -- CP-element group 16: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/aggregated_phi_update_req
      -- CP-element group 16: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3338_update_start__ps
      -- 
    l2CacheDaemon_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "l2CacheDaemon_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(19) & l2CacheDaemon_CP_3229_elements(38) & l2CacheDaemon_CP_3229_elements(59);
      gj_l2CacheDaemon_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	21 
    -- CP-element group 17: 	42 
    -- CP-element group 17: 	63 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	12 
    -- CP-element group 17: marked-successors 
    -- CP-element group 17: 	13 
    -- CP-element group 17:  members (1) 
      -- CP-element group 17: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/aggregated_phi_update_ack
      -- 
    l2CacheDaemon_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "l2CacheDaemon_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(21) & l2CacheDaemon_CP_3229_elements(42) & l2CacheDaemon_CP_3229_elements(63);
      gj_l2CacheDaemon_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	11 
    -- CP-element group 18: marked-predecessors 
    -- CP-element group 18: 	14 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	13 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3338_sample_start_
      -- 
    l2CacheDaemon_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 33) := "l2CacheDaemon_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(11) & l2CacheDaemon_CP_3229_elements(14);
      gj_l2CacheDaemon_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	11 
    -- CP-element group 19: marked-predecessors 
    -- CP-element group 19: 	93 
    -- CP-element group 19: 	81 
    -- CP-element group 19: 	85 
    -- CP-element group 19: 	157 
    -- CP-element group 19: 	101 
    -- CP-element group 19: 	105 
    -- CP-element group 19: 	193 
    -- CP-element group 19: 	189 
    -- CP-element group 19: 	129 
    -- CP-element group 19: 	181 
    -- CP-element group 19: 	125 
    -- CP-element group 19: 	177 
    -- CP-element group 19: 	137 
    -- CP-element group 19: 	141 
    -- CP-element group 19: 	153 
    -- CP-element group 19: 	97 
    -- CP-element group 19: 	169 
    -- CP-element group 19: 	113 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	16 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3338_update_start_
      -- 
    l2CacheDaemon_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 18) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1);
      constant place_markings: IntegerArray(0 to 18)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1,17 => 1,18 => 1);
      constant place_delays: IntegerArray(0 to 18) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0,17 => 0,18 => 0);
      constant joinName: string(1 to 33) := "l2CacheDaemon_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 19); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(11) & l2CacheDaemon_CP_3229_elements(93) & l2CacheDaemon_CP_3229_elements(81) & l2CacheDaemon_CP_3229_elements(85) & l2CacheDaemon_CP_3229_elements(157) & l2CacheDaemon_CP_3229_elements(101) & l2CacheDaemon_CP_3229_elements(105) & l2CacheDaemon_CP_3229_elements(193) & l2CacheDaemon_CP_3229_elements(189) & l2CacheDaemon_CP_3229_elements(129) & l2CacheDaemon_CP_3229_elements(181) & l2CacheDaemon_CP_3229_elements(125) & l2CacheDaemon_CP_3229_elements(177) & l2CacheDaemon_CP_3229_elements(137) & l2CacheDaemon_CP_3229_elements(141) & l2CacheDaemon_CP_3229_elements(153) & l2CacheDaemon_CP_3229_elements(97) & l2CacheDaemon_CP_3229_elements(169) & l2CacheDaemon_CP_3229_elements(113);
      gj_l2CacheDaemon_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 19, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	14 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3338_sample_completed__ps
      -- 
    -- Element group l2CacheDaemon_CP_3229_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	17 
    -- CP-element group 21: 	91 
    -- CP-element group 21: 	80 
    -- CP-element group 21: 	83 
    -- CP-element group 21: 	155 
    -- CP-element group 21: 	103 
    -- CP-element group 21: 	191 
    -- CP-element group 21: 	187 
    -- CP-element group 21: 	127 
    -- CP-element group 21: 	123 
    -- CP-element group 21: 	175 
    -- CP-element group 21: 	179 
    -- CP-element group 21: 	135 
    -- CP-element group 21: 	139 
    -- CP-element group 21: 	151 
    -- CP-element group 21: 	95 
    -- CP-element group 21: 	99 
    -- CP-element group 21: 	167 
    -- CP-element group 21: 	111 
    -- CP-element group 21:  members (2) 
      -- CP-element group 21: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3338_update_completed__ps
      -- CP-element group 21: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3338_update_completed_
      -- 
    -- Element group l2CacheDaemon_CP_3229_elements(21) is bound as output of CP function.
    -- CP-element group 22:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: 	9 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (1) 
      -- CP-element group 22: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3338_loopback_trigger
      -- 
    l2CacheDaemon_CP_3229_elements(22) <= l2CacheDaemon_CP_3229_elements(9);
    -- CP-element group 23:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3338_loopback_sample_req
      -- CP-element group 23: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3338_loopback_sample_req_ps
      -- 
    phi_stmt_3338_loopback_sample_req_3286_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3338_loopback_sample_req_3286_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(23), ack => phi_stmt_3338_req_1); -- 
    -- Element group l2CacheDaemon_CP_3229_elements(23) is bound as output of CP function.
    -- CP-element group 24:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: 	10 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (1) 
      -- CP-element group 24: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3338_entry_trigger
      -- 
    l2CacheDaemon_CP_3229_elements(24) <= l2CacheDaemon_CP_3229_elements(10);
    -- CP-element group 25:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (2) 
      -- CP-element group 25: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3338_entry_sample_req
      -- CP-element group 25: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3338_entry_sample_req_ps
      -- 
    phi_stmt_3338_entry_sample_req_3289_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3338_entry_sample_req_3289_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(25), ack => phi_stmt_3338_req_0); -- 
    -- Element group l2CacheDaemon_CP_3229_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3338_phi_mux_ack
      -- CP-element group 26: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3338_phi_mux_ack_ps
      -- 
    phi_stmt_3338_phi_mux_ack_3292_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3338_ack_0, ack => l2CacheDaemon_CP_3229_elements(26)); -- 
    -- CP-element group 27:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/konst_3340_sample_start__ps
      -- CP-element group 27: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/konst_3340_sample_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/konst_3340_sample_start_
      -- CP-element group 27: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/konst_3340_sample_completed_
      -- 
    -- Element group l2CacheDaemon_CP_3229_elements(27) is bound as output of CP function.
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28: 	30 
    -- CP-element group 28:  members (2) 
      -- CP-element group 28: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/konst_3340_update_start__ps
      -- CP-element group 28: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/konst_3340_update_start_
      -- 
    -- Element group l2CacheDaemon_CP_3229_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: 	30 
    -- CP-element group 29: successors 
    -- CP-element group 29:  members (1) 
      -- CP-element group 29: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/konst_3340_update_completed__ps
      -- 
    l2CacheDaemon_CP_3229_elements(29) <= l2CacheDaemon_CP_3229_elements(30);
    -- CP-element group 30:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	28 
    -- CP-element group 30: successors 
    -- CP-element group 30: 	29 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/konst_3340_update_completed_
      -- 
    -- Element group l2CacheDaemon_CP_3229_elements(30) is a control-delay.
    cp_element_30_delay: control_delay_element  generic map(name => " 30_delay", delay_value => 1)  port map(req => l2CacheDaemon_CP_3229_elements(28), ack => l2CacheDaemon_CP_3229_elements(30), clk => clk, reset =>reset);
    -- CP-element group 31:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	33 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_NOBLOCK_L2_REQUEST_3342_sample_start__ps
      -- 
    -- Element group l2CacheDaemon_CP_3229_elements(31) is bound as output of CP function.
    -- CP-element group 32:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (1) 
      -- CP-element group 32: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_NOBLOCK_L2_REQUEST_3342_update_start__ps
      -- 
    -- Element group l2CacheDaemon_CP_3229_elements(32) is bound as output of CP function.
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: 	31 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	36 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_NOBLOCK_L2_REQUEST_3342_sample_start_
      -- CP-element group 33: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_NOBLOCK_L2_REQUEST_3342_Sample/$entry
      -- CP-element group 33: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_NOBLOCK_L2_REQUEST_3342_Sample/rr
      -- 
    rr_3313_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3313_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(33), ack => RPIPE_NOBLOCK_L2_REQUEST_3342_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "l2CacheDaemon_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(31) & l2CacheDaemon_CP_3229_elements(36);
      gj_l2CacheDaemon_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: 	35 
    -- CP-element group 34: successors 
    -- CP-element group 34: 	36 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_NOBLOCK_L2_REQUEST_3342_update_start_
      -- CP-element group 34: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_NOBLOCK_L2_REQUEST_3342_Update/$entry
      -- CP-element group 34: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_NOBLOCK_L2_REQUEST_3342_Update/cr
      -- 
    cr_3318_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3318_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(34), ack => RPIPE_NOBLOCK_L2_REQUEST_3342_inst_req_1); -- 
    l2CacheDaemon_cp_element_group_34: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "l2CacheDaemon_cp_element_group_34"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(32) & l2CacheDaemon_CP_3229_elements(35);
      gj_l2CacheDaemon_cp_element_group_34 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(34), clk => clk, reset => reset); --
    end block;
    -- CP-element group 35:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	34 
    -- CP-element group 35:  members (4) 
      -- CP-element group 35: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_NOBLOCK_L2_REQUEST_3342_sample_completed__ps
      -- CP-element group 35: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_NOBLOCK_L2_REQUEST_3342_sample_completed_
      -- CP-element group 35: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_NOBLOCK_L2_REQUEST_3342_Sample/$exit
      -- CP-element group 35: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_NOBLOCK_L2_REQUEST_3342_Sample/ra
      -- 
    ra_3314_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_NOBLOCK_L2_REQUEST_3342_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(35)); -- 
    -- CP-element group 36:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	34 
    -- CP-element group 36: successors 
    -- CP-element group 36: marked-successors 
    -- CP-element group 36: 	33 
    -- CP-element group 36:  members (4) 
      -- CP-element group 36: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_NOBLOCK_L2_REQUEST_3342_update_completed__ps
      -- CP-element group 36: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_NOBLOCK_L2_REQUEST_3342_update_completed_
      -- CP-element group 36: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_NOBLOCK_L2_REQUEST_3342_Update/$exit
      -- CP-element group 36: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_NOBLOCK_L2_REQUEST_3342_Update/ca
      -- 
    ca_3319_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 36_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_NOBLOCK_L2_REQUEST_3342_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(36)); -- 
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	11 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	14 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	13 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3343_sample_start_
      -- 
    l2CacheDaemon_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 33) := "l2CacheDaemon_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(11) & l2CacheDaemon_CP_3229_elements(14);
      gj_l2CacheDaemon_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  join  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	11 
    -- CP-element group 38: marked-predecessors 
    -- CP-element group 38: 	93 
    -- CP-element group 38: 	81 
    -- CP-element group 38: 	85 
    -- CP-element group 38: 	157 
    -- CP-element group 38: 	101 
    -- CP-element group 38: 	105 
    -- CP-element group 38: 	109 
    -- CP-element group 38: 	193 
    -- CP-element group 38: 	125 
    -- CP-element group 38: 	117 
    -- CP-element group 38: 	121 
    -- CP-element group 38: 	137 
    -- CP-element group 38: 	141 
    -- CP-element group 38: 	153 
    -- CP-element group 38: 	97 
    -- CP-element group 38: 	78 
    -- CP-element group 38: successors 
    -- CP-element group 38: 	16 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3343_update_start_
      -- 
    l2CacheDaemon_cp_element_group_38: block -- 
      constant place_capacities: IntegerArray(0 to 16) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_markings: IntegerArray(0 to 16)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1,12 => 1,13 => 1,14 => 1,15 => 1,16 => 1);
      constant place_delays: IntegerArray(0 to 16) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0,12 => 0,13 => 0,14 => 0,15 => 0,16 => 0);
      constant joinName: string(1 to 33) := "l2CacheDaemon_cp_element_group_38"; 
      signal preds: BooleanArray(1 to 17); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(11) & l2CacheDaemon_CP_3229_elements(93) & l2CacheDaemon_CP_3229_elements(81) & l2CacheDaemon_CP_3229_elements(85) & l2CacheDaemon_CP_3229_elements(157) & l2CacheDaemon_CP_3229_elements(101) & l2CacheDaemon_CP_3229_elements(105) & l2CacheDaemon_CP_3229_elements(109) & l2CacheDaemon_CP_3229_elements(193) & l2CacheDaemon_CP_3229_elements(125) & l2CacheDaemon_CP_3229_elements(117) & l2CacheDaemon_CP_3229_elements(121) & l2CacheDaemon_CP_3229_elements(137) & l2CacheDaemon_CP_3229_elements(141) & l2CacheDaemon_CP_3229_elements(153) & l2CacheDaemon_CP_3229_elements(97) & l2CacheDaemon_CP_3229_elements(78);
      gj_l2CacheDaemon_cp_element_group_38 : generic_join generic map(name => joinName, number_of_predecessors => 17, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(38), clk => clk, reset => reset); --
    end block;
    -- CP-element group 39:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	13 
    -- CP-element group 39: successors 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3343_sample_start__ps
      -- 
    l2CacheDaemon_CP_3229_elements(39) <= l2CacheDaemon_CP_3229_elements(13);
    -- CP-element group 40:  join  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	14 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3343_sample_completed__ps
      -- 
    -- Element group l2CacheDaemon_CP_3229_elements(40) is bound as output of CP function.
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: 	16 
    -- CP-element group 41: successors 
    -- CP-element group 41:  members (1) 
      -- CP-element group 41: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3343_update_start__ps
      -- 
    l2CacheDaemon_CP_3229_elements(41) <= l2CacheDaemon_CP_3229_elements(16);
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: successors 
    -- CP-element group 42: 	17 
    -- CP-element group 42: 	91 
    -- CP-element group 42: 	80 
    -- CP-element group 42: 	83 
    -- CP-element group 42: 	155 
    -- CP-element group 42: 	103 
    -- CP-element group 42: 	107 
    -- CP-element group 42: 	191 
    -- CP-element group 42: 	123 
    -- CP-element group 42: 	119 
    -- CP-element group 42: 	135 
    -- CP-element group 42: 	139 
    -- CP-element group 42: 	151 
    -- CP-element group 42: 	95 
    -- CP-element group 42: 	99 
    -- CP-element group 42: 	115 
    -- CP-element group 42: 	77 
    -- CP-element group 42:  members (2) 
      -- CP-element group 42: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3343_update_completed_
      -- CP-element group 42: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3343_update_completed__ps
      -- 
    -- Element group l2CacheDaemon_CP_3229_elements(42) is bound as output of CP function.
    -- CP-element group 43:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	9 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (1) 
      -- CP-element group 43: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3343_loopback_trigger
      -- 
    l2CacheDaemon_CP_3229_elements(43) <= l2CacheDaemon_CP_3229_elements(9);
    -- CP-element group 44:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (2) 
      -- CP-element group 44: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3343_loopback_sample_req
      -- CP-element group 44: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3343_loopback_sample_req_ps
      -- 
    phi_stmt_3343_loopback_sample_req_3330_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3343_loopback_sample_req_3330_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(44), ack => phi_stmt_3343_req_1); -- 
    -- Element group l2CacheDaemon_CP_3229_elements(44) is bound as output of CP function.
    -- CP-element group 45:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: 	10 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (1) 
      -- CP-element group 45: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3343_entry_trigger
      -- 
    l2CacheDaemon_CP_3229_elements(45) <= l2CacheDaemon_CP_3229_elements(10);
    -- CP-element group 46:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3343_entry_sample_req
      -- CP-element group 46: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3343_entry_sample_req_ps
      -- 
    phi_stmt_3343_entry_sample_req_3333_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3343_entry_sample_req_3333_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(46), ack => phi_stmt_3343_req_0); -- 
    -- Element group l2CacheDaemon_CP_3229_elements(46) is bound as output of CP function.
    -- CP-element group 47:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (2) 
      -- CP-element group 47: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3343_phi_mux_ack
      -- CP-element group 47: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3343_phi_mux_ack_ps
      -- 
    phi_stmt_3343_phi_mux_ack_3336_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3343_ack_0, ack => l2CacheDaemon_CP_3229_elements(47)); -- 
    -- CP-element group 48:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48:  members (4) 
      -- CP-element group 48: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/konst_3345_sample_start__ps
      -- CP-element group 48: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/konst_3345_sample_completed__ps
      -- CP-element group 48: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/konst_3345_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/konst_3345_sample_completed_
      -- 
    -- Element group l2CacheDaemon_CP_3229_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (2) 
      -- CP-element group 49: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/konst_3345_update_start__ps
      -- CP-element group 49: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/konst_3345_update_start_
      -- 
    -- Element group l2CacheDaemon_CP_3229_elements(49) is bound as output of CP function.
    -- CP-element group 50:  join  transition  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	51 
    -- CP-element group 50: successors 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/konst_3345_update_completed__ps
      -- 
    l2CacheDaemon_CP_3229_elements(50) <= l2CacheDaemon_CP_3229_elements(51);
    -- CP-element group 51:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	50 
    -- CP-element group 51:  members (1) 
      -- CP-element group 51: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/konst_3345_update_completed_
      -- 
    -- Element group l2CacheDaemon_CP_3229_elements(51) is a control-delay.
    cp_element_51_delay: control_delay_element  generic map(name => " 51_delay", delay_value => 1)  port map(req => l2CacheDaemon_CP_3229_elements(49), ack => l2CacheDaemon_CP_3229_elements(51), clk => clk, reset =>reset);
    -- CP-element group 52:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (1) 
      -- CP-element group 52: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_NOBLOCK_L2_INVALIDATE_3346_sample_start__ps
      -- 
    -- Element group l2CacheDaemon_CP_3229_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (1) 
      -- CP-element group 53: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_NOBLOCK_L2_INVALIDATE_3346_update_start__ps
      -- 
    -- Element group l2CacheDaemon_CP_3229_elements(53) is bound as output of CP function.
    -- CP-element group 54:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: marked-predecessors 
    -- CP-element group 54: 	57 
    -- CP-element group 54: successors 
    -- CP-element group 54: 	56 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_NOBLOCK_L2_INVALIDATE_3346_sample_start_
      -- CP-element group 54: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_NOBLOCK_L2_INVALIDATE_3346_Sample/$entry
      -- CP-element group 54: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_NOBLOCK_L2_INVALIDATE_3346_Sample/rr
      -- 
    rr_3357_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3357_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(54), ack => RPIPE_NOBLOCK_L2_INVALIDATE_3346_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_54: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "l2CacheDaemon_cp_element_group_54"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(52) & l2CacheDaemon_CP_3229_elements(57);
      gj_l2CacheDaemon_cp_element_group_54 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(54), clk => clk, reset => reset); --
    end block;
    -- CP-element group 55:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: 	56 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_NOBLOCK_L2_INVALIDATE_3346_update_start_
      -- CP-element group 55: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_NOBLOCK_L2_INVALIDATE_3346_Update/$entry
      -- CP-element group 55: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_NOBLOCK_L2_INVALIDATE_3346_Update/cr
      -- 
    cr_3362_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3362_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(55), ack => RPIPE_NOBLOCK_L2_INVALIDATE_3346_inst_req_1); -- 
    l2CacheDaemon_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "l2CacheDaemon_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(53) & l2CacheDaemon_CP_3229_elements(56);
      gj_l2CacheDaemon_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	54 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	55 
    -- CP-element group 56:  members (4) 
      -- CP-element group 56: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_NOBLOCK_L2_INVALIDATE_3346_sample_completed__ps
      -- CP-element group 56: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_NOBLOCK_L2_INVALIDATE_3346_sample_completed_
      -- CP-element group 56: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_NOBLOCK_L2_INVALIDATE_3346_Sample/$exit
      -- CP-element group 56: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_NOBLOCK_L2_INVALIDATE_3346_Sample/ra
      -- 
    ra_3358_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 56_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_NOBLOCK_L2_INVALIDATE_3346_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(56)); -- 
    -- CP-element group 57:  join  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: marked-successors 
    -- CP-element group 57: 	54 
    -- CP-element group 57:  members (4) 
      -- CP-element group 57: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_NOBLOCK_L2_INVALIDATE_3346_update_completed__ps
      -- CP-element group 57: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_NOBLOCK_L2_INVALIDATE_3346_update_completed_
      -- CP-element group 57: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_NOBLOCK_L2_INVALIDATE_3346_Update/$exit
      -- CP-element group 57: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_NOBLOCK_L2_INVALIDATE_3346_Update/ca
      -- 
    ca_3363_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_NOBLOCK_L2_INVALIDATE_3346_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(57)); -- 
    -- CP-element group 58:  join  transition  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	11 
    -- CP-element group 58: marked-predecessors 
    -- CP-element group 58: 	14 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	13 
    -- CP-element group 58:  members (1) 
      -- CP-element group 58: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3347_sample_start_
      -- 
    l2CacheDaemon_cp_element_group_58: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 33) := "l2CacheDaemon_cp_element_group_58"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(11) & l2CacheDaemon_CP_3229_elements(14);
      gj_l2CacheDaemon_cp_element_group_58 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(58), clk => clk, reset => reset); --
    end block;
    -- CP-element group 59:  join  transition  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	11 
    -- CP-element group 59: marked-predecessors 
    -- CP-element group 59: 	81 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	16 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3347_update_start_
      -- 
    l2CacheDaemon_cp_element_group_59: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "l2CacheDaemon_cp_element_group_59"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(11) & l2CacheDaemon_CP_3229_elements(81);
      gj_l2CacheDaemon_cp_element_group_59 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(59), clk => clk, reset => reset); --
    end block;
    -- CP-element group 60:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	13 
    -- CP-element group 60: successors 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3347_sample_start__ps
      -- 
    l2CacheDaemon_CP_3229_elements(60) <= l2CacheDaemon_CP_3229_elements(13);
    -- CP-element group 61:  join  transition  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	14 
    -- CP-element group 61:  members (1) 
      -- CP-element group 61: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3347_sample_completed__ps
      -- 
    -- Element group l2CacheDaemon_CP_3229_elements(61) is bound as output of CP function.
    -- CP-element group 62:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	16 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (1) 
      -- CP-element group 62: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3347_update_start__ps
      -- 
    l2CacheDaemon_CP_3229_elements(62) <= l2CacheDaemon_CP_3229_elements(16);
    -- CP-element group 63:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	17 
    -- CP-element group 63: 	80 
    -- CP-element group 63:  members (2) 
      -- CP-element group 63: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3347_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3347_update_completed__ps
      -- 
    -- Element group l2CacheDaemon_CP_3229_elements(63) is bound as output of CP function.
    -- CP-element group 64:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	9 
    -- CP-element group 64: successors 
    -- CP-element group 64:  members (1) 
      -- CP-element group 64: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3347_loopback_trigger
      -- 
    l2CacheDaemon_CP_3229_elements(64) <= l2CacheDaemon_CP_3229_elements(9);
    -- CP-element group 65:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (2) 
      -- CP-element group 65: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3347_loopback_sample_req
      -- CP-element group 65: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3347_loopback_sample_req_ps
      -- 
    phi_stmt_3347_loopback_sample_req_3374_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3347_loopback_sample_req_3374_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(65), ack => phi_stmt_3347_req_1); -- 
    -- Element group l2CacheDaemon_CP_3229_elements(65) is bound as output of CP function.
    -- CP-element group 66:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	10 
    -- CP-element group 66: successors 
    -- CP-element group 66:  members (1) 
      -- CP-element group 66: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3347_entry_trigger
      -- 
    l2CacheDaemon_CP_3229_elements(66) <= l2CacheDaemon_CP_3229_elements(10);
    -- CP-element group 67:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: successors 
    -- CP-element group 67:  members (2) 
      -- CP-element group 67: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3347_entry_sample_req
      -- CP-element group 67: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3347_entry_sample_req_ps
      -- 
    phi_stmt_3347_entry_sample_req_3377_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3347_entry_sample_req_3377_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(67), ack => phi_stmt_3347_req_0); -- 
    -- Element group l2CacheDaemon_CP_3229_elements(67) is bound as output of CP function.
    -- CP-element group 68:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: successors 
    -- CP-element group 68:  members (2) 
      -- CP-element group 68: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3347_phi_mux_ack
      -- CP-element group 68: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/phi_stmt_3347_phi_mux_ack_ps
      -- 
    phi_stmt_3347_phi_mux_ack_3380_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 68_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3347_ack_0, ack => l2CacheDaemon_CP_3229_elements(68)); -- 
    -- CP-element group 69:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: successors 
    -- CP-element group 69:  members (4) 
      -- CP-element group 69: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/type_cast_3350_sample_start__ps
      -- CP-element group 69: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/type_cast_3350_sample_completed__ps
      -- CP-element group 69: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/type_cast_3350_sample_start_
      -- CP-element group 69: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/type_cast_3350_sample_completed_
      -- 
    -- Element group l2CacheDaemon_CP_3229_elements(69) is bound as output of CP function.
    -- CP-element group 70:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: successors 
    -- CP-element group 70: 	72 
    -- CP-element group 70:  members (2) 
      -- CP-element group 70: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/type_cast_3350_update_start__ps
      -- CP-element group 70: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/type_cast_3350_update_start_
      -- 
    -- Element group l2CacheDaemon_CP_3229_elements(70) is bound as output of CP function.
    -- CP-element group 71:  join  transition  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	72 
    -- CP-element group 71: successors 
    -- CP-element group 71:  members (1) 
      -- CP-element group 71: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/type_cast_3350_update_completed__ps
      -- 
    l2CacheDaemon_CP_3229_elements(71) <= l2CacheDaemon_CP_3229_elements(72);
    -- CP-element group 72:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	70 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	71 
    -- CP-element group 72:  members (1) 
      -- CP-element group 72: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/type_cast_3350_update_completed_
      -- 
    -- Element group l2CacheDaemon_CP_3229_elements(72) is a control-delay.
    cp_element_72_delay: control_delay_element  generic map(name => " 72_delay", delay_value => 1)  port map(req => l2CacheDaemon_CP_3229_elements(70), ack => l2CacheDaemon_CP_3229_elements(72), clk => clk, reset =>reset);
    -- CP-element group 73:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (4) 
      -- CP-element group 73: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/R_nCOUNTER_3351_sample_start__ps
      -- CP-element group 73: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/R_nCOUNTER_3351_sample_start_
      -- CP-element group 73: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/R_nCOUNTER_3351_Sample/$entry
      -- CP-element group 73: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/R_nCOUNTER_3351_Sample/req
      -- 
    req_3401_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3401_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(73), ack => nCOUNTER_3447_3351_buf_req_0); -- 
    -- Element group l2CacheDaemon_CP_3229_elements(73) is bound as output of CP function.
    -- CP-element group 74:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: successors 
    -- CP-element group 74: 	76 
    -- CP-element group 74:  members (4) 
      -- CP-element group 74: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/R_nCOUNTER_3351_update_start__ps
      -- CP-element group 74: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/R_nCOUNTER_3351_update_start_
      -- CP-element group 74: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/R_nCOUNTER_3351_Update/$entry
      -- CP-element group 74: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/R_nCOUNTER_3351_Update/req
      -- 
    req_3406_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3406_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(74), ack => nCOUNTER_3447_3351_buf_req_1); -- 
    -- Element group l2CacheDaemon_CP_3229_elements(74) is bound as output of CP function.
    -- CP-element group 75:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75:  members (4) 
      -- CP-element group 75: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/R_nCOUNTER_3351_sample_completed__ps
      -- CP-element group 75: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/R_nCOUNTER_3351_sample_completed_
      -- CP-element group 75: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/R_nCOUNTER_3351_Sample/$exit
      -- CP-element group 75: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/R_nCOUNTER_3351_Sample/ack
      -- 
    ack_3402_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_3447_3351_buf_ack_0, ack => l2CacheDaemon_CP_3229_elements(75)); -- 
    -- CP-element group 76:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	74 
    -- CP-element group 76: successors 
    -- CP-element group 76:  members (4) 
      -- CP-element group 76: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/R_nCOUNTER_3351_update_completed__ps
      -- CP-element group 76: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/R_nCOUNTER_3351_update_completed_
      -- CP-element group 76: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/R_nCOUNTER_3351_Update/$exit
      -- CP-element group 76: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/R_nCOUNTER_3351_Update/ack
      -- 
    ack_3407_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 76_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => nCOUNTER_3447_3351_buf_ack_1, ack => l2CacheDaemon_CP_3229_elements(76)); -- 
    -- CP-element group 77:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: 	42 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	79 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	78 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_L2_TO_L1_INVALIDATE_3397_sample_start_
      -- CP-element group 77: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_L2_TO_L1_INVALIDATE_3397_Sample/$entry
      -- CP-element group 77: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_L2_TO_L1_INVALIDATE_3397_Sample/req
      -- 
    req_3416_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3416_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(77), ack => WPIPE_L2_TO_L1_INVALIDATE_3397_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "l2CacheDaemon_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(42) & l2CacheDaemon_CP_3229_elements(79);
      gj_l2CacheDaemon_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	77 
    -- CP-element group 78: successors 
    -- CP-element group 78: 	79 
    -- CP-element group 78: marked-successors 
    -- CP-element group 78: 	38 
    -- CP-element group 78:  members (6) 
      -- CP-element group 78: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_L2_TO_L1_INVALIDATE_3397_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_L2_TO_L1_INVALIDATE_3397_update_start_
      -- CP-element group 78: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_L2_TO_L1_INVALIDATE_3397_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_L2_TO_L1_INVALIDATE_3397_Sample/ack
      -- CP-element group 78: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_L2_TO_L1_INVALIDATE_3397_Update/$entry
      -- CP-element group 78: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_L2_TO_L1_INVALIDATE_3397_Update/req
      -- 
    ack_3417_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_L2_TO_L1_INVALIDATE_3397_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(78)); -- 
    req_3421_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3421_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(78), ack => WPIPE_L2_TO_L1_INVALIDATE_3397_inst_req_1); -- 
    -- CP-element group 79:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	78 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	223 
    -- CP-element group 79: marked-successors 
    -- CP-element group 79: 	77 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_L2_TO_L1_INVALIDATE_3397_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_L2_TO_L1_INVALIDATE_3397_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_L2_TO_L1_INVALIDATE_3397_Update/ack
      -- 
    ack_3422_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_L2_TO_L1_INVALIDATE_3397_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	21 
    -- CP-element group 80: 	42 
    -- CP-element group 80: 	63 
    -- CP-element group 80: marked-predecessors 
    -- CP-element group 80: 	82 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	81 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_NOBLOCK_L2_TAGS_REQUEST_3490_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_NOBLOCK_L2_TAGS_REQUEST_3490_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_NOBLOCK_L2_TAGS_REQUEST_3490_Sample/req
      -- 
    req_3430_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3430_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(80), ack => WPIPE_NOBLOCK_L2_TAGS_REQUEST_3490_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 15,1 => 15,2 => 15,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 33) := "l2CacheDaemon_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(21) & l2CacheDaemon_CP_3229_elements(42) & l2CacheDaemon_CP_3229_elements(63) & l2CacheDaemon_CP_3229_elements(82);
      gj_l2CacheDaemon_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: 	80 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	82 
    -- CP-element group 81: marked-successors 
    -- CP-element group 81: 	19 
    -- CP-element group 81: 	38 
    -- CP-element group 81: 	59 
    -- CP-element group 81:  members (6) 
      -- CP-element group 81: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_NOBLOCK_L2_TAGS_REQUEST_3490_sample_completed_
      -- CP-element group 81: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_NOBLOCK_L2_TAGS_REQUEST_3490_update_start_
      -- CP-element group 81: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_NOBLOCK_L2_TAGS_REQUEST_3490_Sample/$exit
      -- CP-element group 81: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_NOBLOCK_L2_TAGS_REQUEST_3490_Sample/ack
      -- CP-element group 81: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_NOBLOCK_L2_TAGS_REQUEST_3490_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_NOBLOCK_L2_TAGS_REQUEST_3490_Update/req
      -- 
    ack_3431_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 81_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NOBLOCK_L2_TAGS_REQUEST_3490_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(81)); -- 
    req_3435_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3435_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(81), ack => WPIPE_NOBLOCK_L2_TAGS_REQUEST_3490_inst_req_1); -- 
    -- CP-element group 82:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	81 
    -- CP-element group 82: successors 
    -- CP-element group 82: 	223 
    -- CP-element group 82: marked-successors 
    -- CP-element group 82: 	80 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_NOBLOCK_L2_TAGS_REQUEST_3490_update_completed_
      -- CP-element group 82: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_NOBLOCK_L2_TAGS_REQUEST_3490_Update/$exit
      -- CP-element group 82: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_NOBLOCK_L2_TAGS_REQUEST_3490_Update/ack
      -- 
    ack_3436_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_NOBLOCK_L2_TAGS_REQUEST_3490_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(82)); -- 
    -- CP-element group 83:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	21 
    -- CP-element group 83: 	42 
    -- CP-element group 83: marked-predecessors 
    -- CP-element group 83: 	85 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	85 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3495_sample_start_
      -- CP-element group 83: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3495_Sample/$entry
      -- CP-element group 83: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3495_Sample/req
      -- 
    req_3444_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3444_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(83), ack => W_do_tag_access_3276_delayed_4_0_3493_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_83: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 33) := "l2CacheDaemon_cp_element_group_83"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(21) & l2CacheDaemon_CP_3229_elements(42) & l2CacheDaemon_CP_3229_elements(85);
      gj_l2CacheDaemon_cp_element_group_83 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(83), clk => clk, reset => reset); --
    end block;
    -- CP-element group 84:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	89 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3495_update_start_
      -- CP-element group 84: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3495_Update/$entry
      -- CP-element group 84: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3495_Update/req
      -- 
    req_3449_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3449_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(84), ack => W_do_tag_access_3276_delayed_4_0_3493_inst_req_1); -- 
    l2CacheDaemon_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 33) := "l2CacheDaemon_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= l2CacheDaemon_CP_3229_elements(89);
      gj_l2CacheDaemon_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: 	83 
    -- CP-element group 85: successors 
    -- CP-element group 85: marked-successors 
    -- CP-element group 85: 	19 
    -- CP-element group 85: 	38 
    -- CP-element group 85: 	83 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3495_sample_completed_
      -- CP-element group 85: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3495_Sample/$exit
      -- CP-element group 85: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3495_Sample/ack
      -- 
    ack_3445_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 85_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_do_tag_access_3276_delayed_4_0_3493_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(85)); -- 
    -- CP-element group 86:  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: 	87 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3495_update_completed_
      -- CP-element group 86: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3495_Update/$exit
      -- CP-element group 86: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3495_Update/ack
      -- 
    ack_3450_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_do_tag_access_3276_delayed_4_0_3493_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(86)); -- 
    -- CP-element group 87:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	86 
    -- CP-element group 87: marked-predecessors 
    -- CP-element group 87: 	90 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	89 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_L2_TAGS_RESPONSE_3498_sample_start_
      -- CP-element group 87: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_L2_TAGS_RESPONSE_3498_Sample/$entry
      -- CP-element group 87: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_L2_TAGS_RESPONSE_3498_Sample/rr
      -- 
    rr_3458_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3458_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(87), ack => RPIPE_L2_TAGS_RESPONSE_3498_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_87: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 33) := "l2CacheDaemon_cp_element_group_87"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(86) & l2CacheDaemon_CP_3229_elements(90);
      gj_l2CacheDaemon_cp_element_group_87 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(87), clk => clk, reset => reset); --
    end block;
    -- CP-element group 88:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	89 
    -- CP-element group 88: marked-predecessors 
    -- CP-element group 88: 	212 
    -- CP-element group 88: 	216 
    -- CP-element group 88: 	173 
    -- CP-element group 88: 	145 
    -- CP-element group 88: 	204 
    -- CP-element group 88: 	208 
    -- CP-element group 88: 	161 
    -- CP-element group 88: 	200 
    -- CP-element group 88: 	133 
    -- CP-element group 88: 	149 
    -- CP-element group 88: 	165 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_L2_TAGS_RESPONSE_3498_update_start_
      -- CP-element group 88: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_L2_TAGS_RESPONSE_3498_Update/$entry
      -- CP-element group 88: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_L2_TAGS_RESPONSE_3498_Update/cr
      -- 
    cr_3463_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3463_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(88), ack => RPIPE_L2_TAGS_RESPONSE_3498_inst_req_1); -- 
    l2CacheDaemon_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 0);
      constant joinName: string(1 to 33) := "l2CacheDaemon_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(89) & l2CacheDaemon_CP_3229_elements(212) & l2CacheDaemon_CP_3229_elements(216) & l2CacheDaemon_CP_3229_elements(173) & l2CacheDaemon_CP_3229_elements(145) & l2CacheDaemon_CP_3229_elements(204) & l2CacheDaemon_CP_3229_elements(208) & l2CacheDaemon_CP_3229_elements(161) & l2CacheDaemon_CP_3229_elements(200) & l2CacheDaemon_CP_3229_elements(133) & l2CacheDaemon_CP_3229_elements(149) & l2CacheDaemon_CP_3229_elements(165);
      gj_l2CacheDaemon_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: 	87 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	88 
    -- CP-element group 89: marked-successors 
    -- CP-element group 89: 	84 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_L2_TAGS_RESPONSE_3498_sample_completed_
      -- CP-element group 89: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_L2_TAGS_RESPONSE_3498_Sample/$exit
      -- CP-element group 89: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_L2_TAGS_RESPONSE_3498_Sample/ra
      -- 
    ra_3459_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 89_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_L2_TAGS_RESPONSE_3498_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(89)); -- 
    -- CP-element group 90:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90: 	214 
    -- CP-element group 90: 	171 
    -- CP-element group 90: 	143 
    -- CP-element group 90: 	147 
    -- CP-element group 90: 	202 
    -- CP-element group 90: 	206 
    -- CP-element group 90: 	210 
    -- CP-element group 90: 	159 
    -- CP-element group 90: 	163 
    -- CP-element group 90: 	131 
    -- CP-element group 90: 	198 
    -- CP-element group 90: marked-successors 
    -- CP-element group 90: 	87 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_L2_TAGS_RESPONSE_3498_update_completed_
      -- CP-element group 90: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_L2_TAGS_RESPONSE_3498_Update/$exit
      -- CP-element group 90: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/RPIPE_L2_TAGS_RESPONSE_3498_Update/ca
      -- 
    ca_3464_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_L2_TAGS_RESPONSE_3498_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(90)); -- 
    -- CP-element group 91:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	21 
    -- CP-element group 91: 	42 
    -- CP-element group 91: marked-predecessors 
    -- CP-element group 91: 	93 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	93 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3522_sample_start_
      -- CP-element group 91: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3522_Sample/$entry
      -- CP-element group 91: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3522_Sample/req
      -- 
    req_3472_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3472_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(91), ack => W_access_set_id_3302_delayed_5_0_3520_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_91: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 33) := "l2CacheDaemon_cp_element_group_91"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(21) & l2CacheDaemon_CP_3229_elements(42) & l2CacheDaemon_CP_3229_elements(93);
      gj_l2CacheDaemon_cp_element_group_91 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(91), clk => clk, reset => reset); --
    end block;
    -- CP-element group 92:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: marked-predecessors 
    -- CP-element group 92: 	216 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3522_update_start_
      -- CP-element group 92: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3522_Update/$entry
      -- CP-element group 92: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3522_Update/req
      -- 
    req_3477_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3477_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(92), ack => W_access_set_id_3302_delayed_5_0_3520_inst_req_1); -- 
    l2CacheDaemon_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 33) := "l2CacheDaemon_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= l2CacheDaemon_CP_3229_elements(216);
      gj_l2CacheDaemon_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: 	91 
    -- CP-element group 93: successors 
    -- CP-element group 93: marked-successors 
    -- CP-element group 93: 	19 
    -- CP-element group 93: 	38 
    -- CP-element group 93: 	91 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3522_sample_completed_
      -- CP-element group 93: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3522_Sample/$exit
      -- CP-element group 93: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3522_Sample/ack
      -- 
    ack_3473_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 93_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_access_set_id_3302_delayed_5_0_3520_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(93)); -- 
    -- CP-element group 94:  transition  input  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: successors 
    -- CP-element group 94: 	214 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3522_update_completed_
      -- CP-element group 94: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3522_Update/$exit
      -- CP-element group 94: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3522_Update/ack
      -- 
    ack_3478_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_access_set_id_3302_delayed_5_0_3520_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(94)); -- 
    -- CP-element group 95:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	21 
    -- CP-element group 95: 	42 
    -- CP-element group 95: marked-predecessors 
    -- CP-element group 95: 	97 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	97 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/AND_u1_u1_3539_sample_start_
      -- CP-element group 95: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/AND_u1_u1_3539_Sample/$entry
      -- CP-element group 95: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/AND_u1_u1_3539_Sample/rr
      -- 
    rr_3486_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3486_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(95), ack => AND_u1_u1_3539_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_95: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 33) := "l2CacheDaemon_cp_element_group_95"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(21) & l2CacheDaemon_CP_3229_elements(42) & l2CacheDaemon_CP_3229_elements(97);
      gj_l2CacheDaemon_cp_element_group_95 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(95), clk => clk, reset => reset); --
    end block;
    -- CP-element group 96:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: marked-predecessors 
    -- CP-element group 96: 	204 
    -- CP-element group 96: 	200 
    -- CP-element group 96: 	133 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	98 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/AND_u1_u1_3539_update_start_
      -- CP-element group 96: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/AND_u1_u1_3539_Update/$entry
      -- CP-element group 96: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/AND_u1_u1_3539_Update/cr
      -- 
    cr_3491_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3491_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(96), ack => AND_u1_u1_3539_inst_req_1); -- 
    l2CacheDaemon_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 1,1 => 1,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 33) := "l2CacheDaemon_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(204) & l2CacheDaemon_CP_3229_elements(200) & l2CacheDaemon_CP_3229_elements(133);
      gj_l2CacheDaemon_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: 	95 
    -- CP-element group 97: successors 
    -- CP-element group 97: marked-successors 
    -- CP-element group 97: 	19 
    -- CP-element group 97: 	38 
    -- CP-element group 97: 	95 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/AND_u1_u1_3539_sample_completed_
      -- CP-element group 97: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/AND_u1_u1_3539_Sample/$exit
      -- CP-element group 97: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/AND_u1_u1_3539_Sample/ra
      -- 
    ra_3487_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 97_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_3539_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(97)); -- 
    -- CP-element group 98:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	96 
    -- CP-element group 98: successors 
    -- CP-element group 98: 	202 
    -- CP-element group 98: 	131 
    -- CP-element group 98: 	198 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/AND_u1_u1_3539_update_completed_
      -- CP-element group 98: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/AND_u1_u1_3539_Update/$exit
      -- CP-element group 98: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/AND_u1_u1_3539_Update/ca
      -- 
    ca_3492_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_3539_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(98)); -- 
    -- CP-element group 99:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	21 
    -- CP-element group 99: 	42 
    -- CP-element group 99: marked-predecessors 
    -- CP-element group 99: 	101 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	101 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/AND_u1_u1_3551_sample_start_
      -- CP-element group 99: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/AND_u1_u1_3551_Sample/$entry
      -- CP-element group 99: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/AND_u1_u1_3551_Sample/rr
      -- 
    rr_3500_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3500_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(99), ack => AND_u1_u1_3551_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_99: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 33) := "l2CacheDaemon_cp_element_group_99"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(21) & l2CacheDaemon_CP_3229_elements(42) & l2CacheDaemon_CP_3229_elements(101);
      gj_l2CacheDaemon_cp_element_group_99 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(99), clk => clk, reset => reset); --
    end block;
    -- CP-element group 100:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: marked-predecessors 
    -- CP-element group 100: 	145 
    -- CP-element group 100: 	161 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	102 
    -- CP-element group 100:  members (3) 
      -- CP-element group 100: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/AND_u1_u1_3551_update_start_
      -- CP-element group 100: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/AND_u1_u1_3551_Update/$entry
      -- CP-element group 100: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/AND_u1_u1_3551_Update/cr
      -- 
    cr_3505_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3505_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(100), ack => AND_u1_u1_3551_inst_req_1); -- 
    l2CacheDaemon_cp_element_group_100: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_100"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(145) & l2CacheDaemon_CP_3229_elements(161);
      gj_l2CacheDaemon_cp_element_group_100 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(100), clk => clk, reset => reset); --
    end block;
    -- CP-element group 101:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	99 
    -- CP-element group 101: successors 
    -- CP-element group 101: marked-successors 
    -- CP-element group 101: 	19 
    -- CP-element group 101: 	38 
    -- CP-element group 101: 	99 
    -- CP-element group 101:  members (3) 
      -- CP-element group 101: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/AND_u1_u1_3551_sample_completed_
      -- CP-element group 101: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/AND_u1_u1_3551_Sample/$exit
      -- CP-element group 101: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/AND_u1_u1_3551_Sample/ra
      -- 
    ra_3501_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 101_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_3551_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(101)); -- 
    -- CP-element group 102:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	100 
    -- CP-element group 102: successors 
    -- CP-element group 102: 	143 
    -- CP-element group 102: 	159 
    -- CP-element group 102:  members (3) 
      -- CP-element group 102: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/AND_u1_u1_3551_update_completed_
      -- CP-element group 102: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/AND_u1_u1_3551_Update/$exit
      -- CP-element group 102: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/AND_u1_u1_3551_Update/ca
      -- 
    ca_3506_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => AND_u1_u1_3551_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(102)); -- 
    -- CP-element group 103:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	21 
    -- CP-element group 103: 	42 
    -- CP-element group 103: marked-predecessors 
    -- CP-element group 103: 	105 
    -- CP-element group 103: successors 
    -- CP-element group 103: 	105 
    -- CP-element group 103:  members (3) 
      -- CP-element group 103: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3561_sample_start_
      -- CP-element group 103: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3561_Sample/$entry
      -- CP-element group 103: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3561_Sample/req
      -- 
    req_3514_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3514_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(103), ack => W_do_tag_access_3331_delayed_5_0_3559_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_103: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_103"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(21) & l2CacheDaemon_CP_3229_elements(42) & l2CacheDaemon_CP_3229_elements(105);
      gj_l2CacheDaemon_cp_element_group_103 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(103), clk => clk, reset => reset); --
    end block;
    -- CP-element group 104:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: marked-predecessors 
    -- CP-element group 104: 	145 
    -- CP-element group 104: 	208 
    -- CP-element group 104: 	200 
    -- CP-element group 104: 	149 
    -- CP-element group 104: 	165 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	106 
    -- CP-element group 104:  members (3) 
      -- CP-element group 104: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3561_update_start_
      -- CP-element group 104: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3561_Update/$entry
      -- CP-element group 104: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3561_Update/req
      -- 
    req_3519_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3519_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(104), ack => W_do_tag_access_3331_delayed_5_0_3559_inst_req_1); -- 
    l2CacheDaemon_cp_element_group_104: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_104"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(145) & l2CacheDaemon_CP_3229_elements(208) & l2CacheDaemon_CP_3229_elements(200) & l2CacheDaemon_CP_3229_elements(149) & l2CacheDaemon_CP_3229_elements(165);
      gj_l2CacheDaemon_cp_element_group_104 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(104), clk => clk, reset => reset); --
    end block;
    -- CP-element group 105:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	103 
    -- CP-element group 105: successors 
    -- CP-element group 105: marked-successors 
    -- CP-element group 105: 	19 
    -- CP-element group 105: 	38 
    -- CP-element group 105: 	103 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3561_sample_completed_
      -- CP-element group 105: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3561_Sample/$exit
      -- CP-element group 105: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3561_Sample/ack
      -- 
    ack_3515_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_do_tag_access_3331_delayed_5_0_3559_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(105)); -- 
    -- CP-element group 106:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	104 
    -- CP-element group 106: successors 
    -- CP-element group 106: 	143 
    -- CP-element group 106: 	147 
    -- CP-element group 106: 	206 
    -- CP-element group 106: 	163 
    -- CP-element group 106: 	198 
    -- CP-element group 106:  members (3) 
      -- CP-element group 106: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3561_update_completed_
      -- CP-element group 106: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3561_Update/$exit
      -- CP-element group 106: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3561_Update/ack
      -- 
    ack_3520_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_do_tag_access_3331_delayed_5_0_3559_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(106)); -- 
    -- CP-element group 107:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 107: predecessors 
    -- CP-element group 107: 	42 
    -- CP-element group 107: marked-predecessors 
    -- CP-element group 107: 	109 
    -- CP-element group 107: successors 
    -- CP-element group 107: 	109 
    -- CP-element group 107:  members (3) 
      -- CP-element group 107: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3564_sample_start_
      -- CP-element group 107: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3564_Sample/$entry
      -- CP-element group 107: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3564_Sample/req
      -- 
    req_3528_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3528_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(107), ack => W_inv_valid_3337_delayed_5_0_3562_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_107: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_107"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(42) & l2CacheDaemon_CP_3229_elements(109);
      gj_l2CacheDaemon_cp_element_group_107 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(107), clk => clk, reset => reset); --
    end block;
    -- CP-element group 108:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 108: predecessors 
    -- CP-element group 108: marked-predecessors 
    -- CP-element group 108: 	145 
    -- CP-element group 108: 	208 
    -- CP-element group 108: 	200 
    -- CP-element group 108: 	149 
    -- CP-element group 108: 	165 
    -- CP-element group 108: successors 
    -- CP-element group 108: 	110 
    -- CP-element group 108:  members (3) 
      -- CP-element group 108: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3564_update_start_
      -- CP-element group 108: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3564_Update/$entry
      -- CP-element group 108: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3564_Update/req
      -- 
    req_3533_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3533_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(108), ack => W_inv_valid_3337_delayed_5_0_3562_inst_req_1); -- 
    l2CacheDaemon_cp_element_group_108: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_108"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(145) & l2CacheDaemon_CP_3229_elements(208) & l2CacheDaemon_CP_3229_elements(200) & l2CacheDaemon_CP_3229_elements(149) & l2CacheDaemon_CP_3229_elements(165);
      gj_l2CacheDaemon_cp_element_group_108 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(108), clk => clk, reset => reset); --
    end block;
    -- CP-element group 109:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 109: predecessors 
    -- CP-element group 109: 	107 
    -- CP-element group 109: successors 
    -- CP-element group 109: marked-successors 
    -- CP-element group 109: 	38 
    -- CP-element group 109: 	107 
    -- CP-element group 109:  members (3) 
      -- CP-element group 109: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3564_sample_completed_
      -- CP-element group 109: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3564_Sample/$exit
      -- CP-element group 109: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3564_Sample/ack
      -- 
    ack_3529_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 109_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_inv_valid_3337_delayed_5_0_3562_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(109)); -- 
    -- CP-element group 110:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 110: predecessors 
    -- CP-element group 110: 	108 
    -- CP-element group 110: successors 
    -- CP-element group 110: 	143 
    -- CP-element group 110: 	147 
    -- CP-element group 110: 	206 
    -- CP-element group 110: 	163 
    -- CP-element group 110: 	198 
    -- CP-element group 110:  members (3) 
      -- CP-element group 110: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3564_update_completed_
      -- CP-element group 110: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3564_Update/$exit
      -- CP-element group 110: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3564_Update/ack
      -- 
    ack_3534_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 110_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_inv_valid_3337_delayed_5_0_3562_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(110)); -- 
    -- CP-element group 111:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 111: predecessors 
    -- CP-element group 111: 	21 
    -- CP-element group 111: marked-predecessors 
    -- CP-element group 111: 	113 
    -- CP-element group 111: successors 
    -- CP-element group 111: 	113 
    -- CP-element group 111:  members (3) 
      -- CP-element group 111: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3567_sample_start_
      -- CP-element group 111: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3567_Sample/$entry
      -- CP-element group 111: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3567_Sample/req
      -- 
    req_3542_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3542_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(111), ack => W_valid_3340_delayed_5_0_3565_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_111: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_111"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(21) & l2CacheDaemon_CP_3229_elements(113);
      gj_l2CacheDaemon_cp_element_group_111 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(111), clk => clk, reset => reset); --
    end block;
    -- CP-element group 112:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 112: predecessors 
    -- CP-element group 112: marked-predecessors 
    -- CP-element group 112: 	145 
    -- CP-element group 112: 	208 
    -- CP-element group 112: 	200 
    -- CP-element group 112: 	149 
    -- CP-element group 112: 	165 
    -- CP-element group 112: successors 
    -- CP-element group 112: 	114 
    -- CP-element group 112:  members (3) 
      -- CP-element group 112: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3567_update_start_
      -- CP-element group 112: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3567_Update/$entry
      -- CP-element group 112: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3567_Update/req
      -- 
    req_3547_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3547_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(112), ack => W_valid_3340_delayed_5_0_3565_inst_req_1); -- 
    l2CacheDaemon_cp_element_group_112: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_112"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(145) & l2CacheDaemon_CP_3229_elements(208) & l2CacheDaemon_CP_3229_elements(200) & l2CacheDaemon_CP_3229_elements(149) & l2CacheDaemon_CP_3229_elements(165);
      gj_l2CacheDaemon_cp_element_group_112 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(112), clk => clk, reset => reset); --
    end block;
    -- CP-element group 113:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 113: predecessors 
    -- CP-element group 113: 	111 
    -- CP-element group 113: successors 
    -- CP-element group 113: marked-successors 
    -- CP-element group 113: 	19 
    -- CP-element group 113: 	111 
    -- CP-element group 113:  members (3) 
      -- CP-element group 113: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3567_sample_completed_
      -- CP-element group 113: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3567_Sample/$exit
      -- CP-element group 113: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3567_Sample/ack
      -- 
    ack_3543_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 113_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_valid_3340_delayed_5_0_3565_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(113)); -- 
    -- CP-element group 114:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 114: predecessors 
    -- CP-element group 114: 	112 
    -- CP-element group 114: successors 
    -- CP-element group 114: 	143 
    -- CP-element group 114: 	147 
    -- CP-element group 114: 	206 
    -- CP-element group 114: 	163 
    -- CP-element group 114: 	198 
    -- CP-element group 114:  members (3) 
      -- CP-element group 114: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3567_update_completed_
      -- CP-element group 114: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3567_Update/$exit
      -- CP-element group 114: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3567_Update/ack
      -- 
    ack_3548_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 114_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_valid_3340_delayed_5_0_3565_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(114)); -- 
    -- CP-element group 115:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 115: predecessors 
    -- CP-element group 115: 	42 
    -- CP-element group 115: marked-predecessors 
    -- CP-element group 115: 	117 
    -- CP-element group 115: successors 
    -- CP-element group 115: 	117 
    -- CP-element group 115:  members (3) 
      -- CP-element group 115: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3605_sample_start_
      -- CP-element group 115: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3605_Sample/$entry
      -- CP-element group 115: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3605_Sample/req
      -- 
    req_3556_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3556_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(115), ack => W_inv_valid_3366_delayed_5_0_3603_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_115: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_115"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(42) & l2CacheDaemon_CP_3229_elements(117);
      gj_l2CacheDaemon_cp_element_group_115 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(115), clk => clk, reset => reset); --
    end block;
    -- CP-element group 116:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 116: predecessors 
    -- CP-element group 116: marked-predecessors 
    -- CP-element group 116: 	216 
    -- CP-element group 116: successors 
    -- CP-element group 116: 	118 
    -- CP-element group 116:  members (3) 
      -- CP-element group 116: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3605_update_start_
      -- CP-element group 116: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3605_Update/$entry
      -- CP-element group 116: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3605_Update/req
      -- 
    req_3561_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3561_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(116), ack => W_inv_valid_3366_delayed_5_0_3603_inst_req_1); -- 
    l2CacheDaemon_cp_element_group_116: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_116"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= l2CacheDaemon_CP_3229_elements(216);
      gj_l2CacheDaemon_cp_element_group_116 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(116), clk => clk, reset => reset); --
    end block;
    -- CP-element group 117:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 117: predecessors 
    -- CP-element group 117: 	115 
    -- CP-element group 117: successors 
    -- CP-element group 117: marked-successors 
    -- CP-element group 117: 	38 
    -- CP-element group 117: 	115 
    -- CP-element group 117:  members (3) 
      -- CP-element group 117: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3605_sample_completed_
      -- CP-element group 117: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3605_Sample/$exit
      -- CP-element group 117: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3605_Sample/ack
      -- 
    ack_3557_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 117_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_inv_valid_3366_delayed_5_0_3603_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(117)); -- 
    -- CP-element group 118:  transition  input  bypass  pipeline-parent 
    -- CP-element group 118: predecessors 
    -- CP-element group 118: 	116 
    -- CP-element group 118: successors 
    -- CP-element group 118: 	214 
    -- CP-element group 118:  members (3) 
      -- CP-element group 118: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3605_update_completed_
      -- CP-element group 118: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3605_Update/$exit
      -- CP-element group 118: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3605_Update/ack
      -- 
    ack_3562_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 118_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_inv_valid_3366_delayed_5_0_3603_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(118)); -- 
    -- CP-element group 119:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 119: predecessors 
    -- CP-element group 119: 	42 
    -- CP-element group 119: marked-predecessors 
    -- CP-element group 119: 	121 
    -- CP-element group 119: successors 
    -- CP-element group 119: 	121 
    -- CP-element group 119:  members (3) 
      -- CP-element group 119: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3608_sample_start_
      -- CP-element group 119: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3608_Sample/$entry
      -- CP-element group 119: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3608_Sample/req
      -- 
    req_3570_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3570_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(119), ack => W_inv_pa_line_address_3367_delayed_5_0_3606_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_119: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_119"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(42) & l2CacheDaemon_CP_3229_elements(121);
      gj_l2CacheDaemon_cp_element_group_119 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(119), clk => clk, reset => reset); --
    end block;
    -- CP-element group 120:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 120: predecessors 
    -- CP-element group 120: marked-predecessors 
    -- CP-element group 120: 	216 
    -- CP-element group 120: successors 
    -- CP-element group 120: 	122 
    -- CP-element group 120:  members (3) 
      -- CP-element group 120: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3608_update_start_
      -- CP-element group 120: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3608_Update/$entry
      -- CP-element group 120: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3608_Update/req
      -- 
    req_3575_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3575_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(120), ack => W_inv_pa_line_address_3367_delayed_5_0_3606_inst_req_1); -- 
    l2CacheDaemon_cp_element_group_120: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_120"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= l2CacheDaemon_CP_3229_elements(216);
      gj_l2CacheDaemon_cp_element_group_120 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(120), clk => clk, reset => reset); --
    end block;
    -- CP-element group 121:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 121: predecessors 
    -- CP-element group 121: 	119 
    -- CP-element group 121: successors 
    -- CP-element group 121: marked-successors 
    -- CP-element group 121: 	38 
    -- CP-element group 121: 	119 
    -- CP-element group 121:  members (3) 
      -- CP-element group 121: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3608_sample_completed_
      -- CP-element group 121: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3608_Sample/$exit
      -- CP-element group 121: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3608_Sample/ack
      -- 
    ack_3571_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 121_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_inv_pa_line_address_3367_delayed_5_0_3606_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(121)); -- 
    -- CP-element group 122:  transition  input  bypass  pipeline-parent 
    -- CP-element group 122: predecessors 
    -- CP-element group 122: 	120 
    -- CP-element group 122: successors 
    -- CP-element group 122: 	214 
    -- CP-element group 122:  members (3) 
      -- CP-element group 122: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3608_update_completed_
      -- CP-element group 122: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3608_Update/$exit
      -- CP-element group 122: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3608_Update/ack
      -- 
    ack_3576_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 122_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_inv_pa_line_address_3367_delayed_5_0_3606_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(122)); -- 
    -- CP-element group 123:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 123: predecessors 
    -- CP-element group 123: 	21 
    -- CP-element group 123: 	42 
    -- CP-element group 123: marked-predecessors 
    -- CP-element group 123: 	125 
    -- CP-element group 123: successors 
    -- CP-element group 123: 	125 
    -- CP-element group 123:  members (3) 
      -- CP-element group 123: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/OR_u1_u1_3618_sample_start_
      -- CP-element group 123: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/OR_u1_u1_3618_Sample/$entry
      -- CP-element group 123: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/OR_u1_u1_3618_Sample/rr
      -- 
    rr_3584_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3584_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(123), ack => OR_u1_u1_3618_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_123: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_123"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(21) & l2CacheDaemon_CP_3229_elements(42) & l2CacheDaemon_CP_3229_elements(125);
      gj_l2CacheDaemon_cp_element_group_123 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(123), clk => clk, reset => reset); --
    end block;
    -- CP-element group 124:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 124: predecessors 
    -- CP-element group 124: marked-predecessors 
    -- CP-element group 124: 	145 
    -- CP-element group 124: successors 
    -- CP-element group 124: 	126 
    -- CP-element group 124:  members (3) 
      -- CP-element group 124: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/OR_u1_u1_3618_update_start_
      -- CP-element group 124: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/OR_u1_u1_3618_Update/$entry
      -- CP-element group 124: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/OR_u1_u1_3618_Update/cr
      -- 
    cr_3589_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3589_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(124), ack => OR_u1_u1_3618_inst_req_1); -- 
    l2CacheDaemon_cp_element_group_124: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_124"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= l2CacheDaemon_CP_3229_elements(145);
      gj_l2CacheDaemon_cp_element_group_124 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(124), clk => clk, reset => reset); --
    end block;
    -- CP-element group 125:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 125: predecessors 
    -- CP-element group 125: 	123 
    -- CP-element group 125: successors 
    -- CP-element group 125: marked-successors 
    -- CP-element group 125: 	19 
    -- CP-element group 125: 	38 
    -- CP-element group 125: 	123 
    -- CP-element group 125:  members (3) 
      -- CP-element group 125: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/OR_u1_u1_3618_sample_completed_
      -- CP-element group 125: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/OR_u1_u1_3618_Sample/$exit
      -- CP-element group 125: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/OR_u1_u1_3618_Sample/ra
      -- 
    ra_3585_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 125_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u1_u1_3618_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(125)); -- 
    -- CP-element group 126:  transition  input  bypass  pipeline-parent 
    -- CP-element group 126: predecessors 
    -- CP-element group 126: 	124 
    -- CP-element group 126: successors 
    -- CP-element group 126: 	143 
    -- CP-element group 126:  members (3) 
      -- CP-element group 126: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/OR_u1_u1_3618_update_completed_
      -- CP-element group 126: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/OR_u1_u1_3618_Update/$exit
      -- CP-element group 126: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/OR_u1_u1_3618_Update/ca
      -- 
    ca_3590_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 126_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => OR_u1_u1_3618_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(126)); -- 
    -- CP-element group 127:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 127: predecessors 
    -- CP-element group 127: 	21 
    -- CP-element group 127: marked-predecessors 
    -- CP-element group 127: 	129 
    -- CP-element group 127: successors 
    -- CP-element group 127: 	129 
    -- CP-element group 127:  members (3) 
      -- CP-element group 127: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3629_sample_start_
      -- CP-element group 127: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3629_Sample/$entry
      -- CP-element group 127: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3629_Sample/req
      -- 
    req_3598_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3598_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(127), ack => W_pa_line_address_3381_delayed_5_0_3627_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_127: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_127"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(21) & l2CacheDaemon_CP_3229_elements(129);
      gj_l2CacheDaemon_cp_element_group_127 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(127), clk => clk, reset => reset); --
    end block;
    -- CP-element group 128:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 128: predecessors 
    -- CP-element group 128: marked-predecessors 
    -- CP-element group 128: 	133 
    -- CP-element group 128: successors 
    -- CP-element group 128: 	130 
    -- CP-element group 128:  members (3) 
      -- CP-element group 128: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3629_update_start_
      -- CP-element group 128: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3629_Update/$entry
      -- CP-element group 128: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3629_Update/req
      -- 
    req_3603_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3603_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(128), ack => W_pa_line_address_3381_delayed_5_0_3627_inst_req_1); -- 
    l2CacheDaemon_cp_element_group_128: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_128"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= l2CacheDaemon_CP_3229_elements(133);
      gj_l2CacheDaemon_cp_element_group_128 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(128), clk => clk, reset => reset); --
    end block;
    -- CP-element group 129:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 129: predecessors 
    -- CP-element group 129: 	127 
    -- CP-element group 129: successors 
    -- CP-element group 129: marked-successors 
    -- CP-element group 129: 	19 
    -- CP-element group 129: 	127 
    -- CP-element group 129:  members (3) 
      -- CP-element group 129: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3629_sample_completed_
      -- CP-element group 129: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3629_Sample/$exit
      -- CP-element group 129: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3629_Sample/ack
      -- 
    ack_3599_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 129_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_pa_line_address_3381_delayed_5_0_3627_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(129)); -- 
    -- CP-element group 130:  transition  input  bypass  pipeline-parent 
    -- CP-element group 130: predecessors 
    -- CP-element group 130: 	128 
    -- CP-element group 130: successors 
    -- CP-element group 130: 	131 
    -- CP-element group 130:  members (3) 
      -- CP-element group 130: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3629_update_completed_
      -- CP-element group 130: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3629_Update/$exit
      -- CP-element group 130: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3629_Update/ack
      -- 
    ack_3604_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 130_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_pa_line_address_3381_delayed_5_0_3627_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(130)); -- 
    -- CP-element group 131:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 131: predecessors 
    -- CP-element group 131: 	90 
    -- CP-element group 131: 	130 
    -- CP-element group 131: 	98 
    -- CP-element group 131: marked-predecessors 
    -- CP-element group 131: 	133 
    -- CP-element group 131: successors 
    -- CP-element group 131: 	133 
    -- CP-element group 131:  members (3) 
      -- CP-element group 131: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3633_sample_start_
      -- CP-element group 131: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3633_Sample/$entry
      -- CP-element group 131: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3633_Sample/crr
      -- 
    crr_3612_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3612_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(131), ack => call_stmt_3633_call_req_0); -- 
    l2CacheDaemon_cp_element_group_131: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_131"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(90) & l2CacheDaemon_CP_3229_elements(130) & l2CacheDaemon_CP_3229_elements(98) & l2CacheDaemon_CP_3229_elements(133);
      gj_l2CacheDaemon_cp_element_group_131 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(131), clk => clk, reset => reset); --
    end block;
    -- CP-element group 132:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 132: predecessors 
    -- CP-element group 132: marked-predecessors 
    -- CP-element group 132: 	185 
    -- CP-element group 132: successors 
    -- CP-element group 132: 	134 
    -- CP-element group 132:  members (3) 
      -- CP-element group 132: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3633_update_start_
      -- CP-element group 132: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3633_Update/$entry
      -- CP-element group 132: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3633_Update/ccr
      -- 
    ccr_3617_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3617_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(132), ack => call_stmt_3633_call_req_1); -- 
    l2CacheDaemon_cp_element_group_132: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_132"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= l2CacheDaemon_CP_3229_elements(185);
      gj_l2CacheDaemon_cp_element_group_132 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(132), clk => clk, reset => reset); --
    end block;
    -- CP-element group 133:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 133: predecessors 
    -- CP-element group 133: 	131 
    -- CP-element group 133: successors 
    -- CP-element group 133: marked-successors 
    -- CP-element group 133: 	88 
    -- CP-element group 133: 	128 
    -- CP-element group 133: 	131 
    -- CP-element group 133: 	96 
    -- CP-element group 133:  members (3) 
      -- CP-element group 133: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3633_sample_completed_
      -- CP-element group 133: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3633_Sample/$exit
      -- CP-element group 133: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3633_Sample/cra
      -- 
    cra_3613_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 133_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_3633_call_ack_0, ack => l2CacheDaemon_CP_3229_elements(133)); -- 
    -- CP-element group 134:  transition  input  bypass  pipeline-parent 
    -- CP-element group 134: predecessors 
    -- CP-element group 134: 	132 
    -- CP-element group 134: successors 
    -- CP-element group 134: 	183 
    -- CP-element group 134:  members (3) 
      -- CP-element group 134: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3633_update_completed_
      -- CP-element group 134: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3633_Update/$exit
      -- CP-element group 134: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3633_Update/cca
      -- 
    cca_3618_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 134_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_3633_call_ack_1, ack => l2CacheDaemon_CP_3229_elements(134)); -- 
    -- CP-element group 135:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 135: predecessors 
    -- CP-element group 135: 	21 
    -- CP-element group 135: 	42 
    -- CP-element group 135: marked-predecessors 
    -- CP-element group 135: 	137 
    -- CP-element group 135: successors 
    -- CP-element group 135: 	137 
    -- CP-element group 135:  members (3) 
      -- CP-element group 135: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3636_sample_start_
      -- CP-element group 135: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3636_Sample/$entry
      -- CP-element group 135: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3636_Sample/req
      -- 
    req_3626_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3626_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(135), ack => W_access_set_id_3386_delayed_5_0_3634_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_135: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_135"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(21) & l2CacheDaemon_CP_3229_elements(42) & l2CacheDaemon_CP_3229_elements(137);
      gj_l2CacheDaemon_cp_element_group_135 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(135), clk => clk, reset => reset); --
    end block;
    -- CP-element group 136:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 136: predecessors 
    -- CP-element group 136: marked-predecessors 
    -- CP-element group 136: 	173 
    -- CP-element group 136: successors 
    -- CP-element group 136: 	138 
    -- CP-element group 136:  members (3) 
      -- CP-element group 136: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3636_update_start_
      -- CP-element group 136: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3636_Update/$entry
      -- CP-element group 136: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3636_Update/req
      -- 
    req_3631_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3631_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(136), ack => W_access_set_id_3386_delayed_5_0_3634_inst_req_1); -- 
    l2CacheDaemon_cp_element_group_136: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_136"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= l2CacheDaemon_CP_3229_elements(173);
      gj_l2CacheDaemon_cp_element_group_136 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(136), clk => clk, reset => reset); --
    end block;
    -- CP-element group 137:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 137: predecessors 
    -- CP-element group 137: 	135 
    -- CP-element group 137: successors 
    -- CP-element group 137: marked-successors 
    -- CP-element group 137: 	19 
    -- CP-element group 137: 	38 
    -- CP-element group 137: 	135 
    -- CP-element group 137:  members (3) 
      -- CP-element group 137: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3636_sample_completed_
      -- CP-element group 137: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3636_Sample/$exit
      -- CP-element group 137: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3636_Sample/ack
      -- 
    ack_3627_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 137_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_access_set_id_3386_delayed_5_0_3634_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(137)); -- 
    -- CP-element group 138:  transition  input  bypass  pipeline-parent 
    -- CP-element group 138: predecessors 
    -- CP-element group 138: 	136 
    -- CP-element group 138: successors 
    -- CP-element group 138: 	171 
    -- CP-element group 138:  members (3) 
      -- CP-element group 138: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3636_update_completed_
      -- CP-element group 138: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3636_Update/$exit
      -- CP-element group 138: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3636_Update/ack
      -- 
    ack_3632_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 138_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_access_set_id_3386_delayed_5_0_3634_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(138)); -- 
    -- CP-element group 139:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 139: predecessors 
    -- CP-element group 139: 	21 
    -- CP-element group 139: 	42 
    -- CP-element group 139: marked-predecessors 
    -- CP-element group 139: 	141 
    -- CP-element group 139: successors 
    -- CP-element group 139: 	141 
    -- CP-element group 139:  members (3) 
      -- CP-element group 139: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3644_sample_start_
      -- CP-element group 139: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3644_Sample/$entry
      -- CP-element group 139: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3644_Sample/req
      -- 
    req_3640_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3640_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(139), ack => W_data_read_dword_3391_delayed_5_0_3642_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_139: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_139"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(21) & l2CacheDaemon_CP_3229_elements(42) & l2CacheDaemon_CP_3229_elements(141);
      gj_l2CacheDaemon_cp_element_group_139 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(139), clk => clk, reset => reset); --
    end block;
    -- CP-element group 140:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 140: predecessors 
    -- CP-element group 140: marked-predecessors 
    -- CP-element group 140: 	149 
    -- CP-element group 140: successors 
    -- CP-element group 140: 	142 
    -- CP-element group 140:  members (3) 
      -- CP-element group 140: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3644_update_start_
      -- CP-element group 140: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3644_Update/$entry
      -- CP-element group 140: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3644_Update/req
      -- 
    req_3645_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3645_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(140), ack => W_data_read_dword_3391_delayed_5_0_3642_inst_req_1); -- 
    l2CacheDaemon_cp_element_group_140: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_140"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= l2CacheDaemon_CP_3229_elements(149);
      gj_l2CacheDaemon_cp_element_group_140 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(140), clk => clk, reset => reset); --
    end block;
    -- CP-element group 141:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 141: predecessors 
    -- CP-element group 141: 	139 
    -- CP-element group 141: successors 
    -- CP-element group 141: marked-successors 
    -- CP-element group 141: 	19 
    -- CP-element group 141: 	38 
    -- CP-element group 141: 	139 
    -- CP-element group 141:  members (3) 
      -- CP-element group 141: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3644_sample_completed_
      -- CP-element group 141: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3644_Sample/$exit
      -- CP-element group 141: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3644_Sample/ack
      -- 
    ack_3641_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 141_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_read_dword_3391_delayed_5_0_3642_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(141)); -- 
    -- CP-element group 142:  transition  input  bypass  pipeline-parent 
    -- CP-element group 142: predecessors 
    -- CP-element group 142: 	140 
    -- CP-element group 142: successors 
    -- CP-element group 142: 	147 
    -- CP-element group 142:  members (3) 
      -- CP-element group 142: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3644_update_completed_
      -- CP-element group 142: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3644_Update/$exit
      -- CP-element group 142: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3644_Update/ack
      -- 
    ack_3646_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 142_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_read_dword_3391_delayed_5_0_3642_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(142)); -- 
    -- CP-element group 143:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 143: predecessors 
    -- CP-element group 143: 	90 
    -- CP-element group 143: 	102 
    -- CP-element group 143: 	106 
    -- CP-element group 143: 	110 
    -- CP-element group 143: 	126 
    -- CP-element group 143: 	114 
    -- CP-element group 143: marked-predecessors 
    -- CP-element group 143: 	145 
    -- CP-element group 143: successors 
    -- CP-element group 143: 	145 
    -- CP-element group 143:  members (3) 
      -- CP-element group 143: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3652_sample_start_
      -- CP-element group 143: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3652_Sample/$entry
      -- CP-element group 143: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3652_Sample/req
      -- 
    req_3654_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3654_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(143), ack => W_access_data_mem_3394_delayed_4_0_3650_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_143: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_143"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(90) & l2CacheDaemon_CP_3229_elements(102) & l2CacheDaemon_CP_3229_elements(106) & l2CacheDaemon_CP_3229_elements(110) & l2CacheDaemon_CP_3229_elements(126) & l2CacheDaemon_CP_3229_elements(114) & l2CacheDaemon_CP_3229_elements(145);
      gj_l2CacheDaemon_cp_element_group_143 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(143), clk => clk, reset => reset); --
    end block;
    -- CP-element group 144:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 144: predecessors 
    -- CP-element group 144: marked-predecessors 
    -- CP-element group 144: 	185 
    -- CP-element group 144: successors 
    -- CP-element group 144: 	146 
    -- CP-element group 144:  members (3) 
      -- CP-element group 144: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3652_update_start_
      -- CP-element group 144: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3652_Update/$entry
      -- CP-element group 144: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3652_Update/req
      -- 
    req_3659_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3659_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(144), ack => W_access_data_mem_3394_delayed_4_0_3650_inst_req_1); -- 
    l2CacheDaemon_cp_element_group_144: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_144"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= l2CacheDaemon_CP_3229_elements(185);
      gj_l2CacheDaemon_cp_element_group_144 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(144), clk => clk, reset => reset); --
    end block;
    -- CP-element group 145:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 145: predecessors 
    -- CP-element group 145: 	143 
    -- CP-element group 145: successors 
    -- CP-element group 145: marked-successors 
    -- CP-element group 145: 	88 
    -- CP-element group 145: 	143 
    -- CP-element group 145: 	104 
    -- CP-element group 145: 	108 
    -- CP-element group 145: 	124 
    -- CP-element group 145: 	100 
    -- CP-element group 145: 	112 
    -- CP-element group 145:  members (3) 
      -- CP-element group 145: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3652_sample_completed_
      -- CP-element group 145: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3652_Sample/$exit
      -- CP-element group 145: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3652_Sample/ack
      -- 
    ack_3655_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 145_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_access_data_mem_3394_delayed_4_0_3650_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(145)); -- 
    -- CP-element group 146:  transition  input  bypass  pipeline-parent 
    -- CP-element group 146: predecessors 
    -- CP-element group 146: 	144 
    -- CP-element group 146: successors 
    -- CP-element group 146: 	183 
    -- CP-element group 146:  members (3) 
      -- CP-element group 146: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3652_update_completed_
      -- CP-element group 146: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3652_Update/$exit
      -- CP-element group 146: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3652_Update/ack
      -- 
    ack_3660_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 146_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_access_data_mem_3394_delayed_4_0_3650_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(146)); -- 
    -- CP-element group 147:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 147: predecessors 
    -- CP-element group 147: 	90 
    -- CP-element group 147: 	106 
    -- CP-element group 147: 	110 
    -- CP-element group 147: 	142 
    -- CP-element group 147: 	114 
    -- CP-element group 147: marked-predecessors 
    -- CP-element group 147: 	149 
    -- CP-element group 147: successors 
    -- CP-element group 147: 	149 
    -- CP-element group 147:  members (3) 
      -- CP-element group 147: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3655_sample_start_
      -- CP-element group 147: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3655_Sample/$entry
      -- CP-element group 147: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3655_Sample/req
      -- 
    req_3668_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3668_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(147), ack => W_read_data_line_3395_delayed_4_0_3653_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_147: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_147"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(90) & l2CacheDaemon_CP_3229_elements(106) & l2CacheDaemon_CP_3229_elements(110) & l2CacheDaemon_CP_3229_elements(142) & l2CacheDaemon_CP_3229_elements(114) & l2CacheDaemon_CP_3229_elements(149);
      gj_l2CacheDaemon_cp_element_group_147 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(147), clk => clk, reset => reset); --
    end block;
    -- CP-element group 148:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 148: predecessors 
    -- CP-element group 148: marked-predecessors 
    -- CP-element group 148: 	185 
    -- CP-element group 148: successors 
    -- CP-element group 148: 	150 
    -- CP-element group 148:  members (3) 
      -- CP-element group 148: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3655_update_start_
      -- CP-element group 148: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3655_Update/$entry
      -- CP-element group 148: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3655_Update/req
      -- 
    req_3673_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3673_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(148), ack => W_read_data_line_3395_delayed_4_0_3653_inst_req_1); -- 
    l2CacheDaemon_cp_element_group_148: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_148"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= l2CacheDaemon_CP_3229_elements(185);
      gj_l2CacheDaemon_cp_element_group_148 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(148), clk => clk, reset => reset); --
    end block;
    -- CP-element group 149:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 149: predecessors 
    -- CP-element group 149: 	147 
    -- CP-element group 149: successors 
    -- CP-element group 149: marked-successors 
    -- CP-element group 149: 	88 
    -- CP-element group 149: 	147 
    -- CP-element group 149: 	104 
    -- CP-element group 149: 	108 
    -- CP-element group 149: 	140 
    -- CP-element group 149: 	112 
    -- CP-element group 149:  members (3) 
      -- CP-element group 149: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3655_sample_completed_
      -- CP-element group 149: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3655_Sample/$exit
      -- CP-element group 149: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3655_Sample/ack
      -- 
    ack_3669_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 149_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_data_line_3395_delayed_4_0_3653_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(149)); -- 
    -- CP-element group 150:  transition  input  bypass  pipeline-parent 
    -- CP-element group 150: predecessors 
    -- CP-element group 150: 	148 
    -- CP-element group 150: successors 
    -- CP-element group 150: 	183 
    -- CP-element group 150:  members (3) 
      -- CP-element group 150: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3655_update_completed_
      -- CP-element group 150: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3655_Update/$exit
      -- CP-element group 150: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3655_Update/ack
      -- 
    ack_3674_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 150_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_read_data_line_3395_delayed_4_0_3653_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(150)); -- 
    -- CP-element group 151:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 151: predecessors 
    -- CP-element group 151: 	21 
    -- CP-element group 151: 	42 
    -- CP-element group 151: marked-predecessors 
    -- CP-element group 151: 	153 
    -- CP-element group 151: successors 
    -- CP-element group 151: 	153 
    -- CP-element group 151:  members (3) 
      -- CP-element group 151: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3658_sample_start_
      -- CP-element group 151: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3658_Sample/$entry
      -- CP-element group 151: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3658_Sample/req
      -- 
    req_3682_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3682_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(151), ack => W_data_write_dword_3396_delayed_9_0_3656_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_151: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_151"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(21) & l2CacheDaemon_CP_3229_elements(42) & l2CacheDaemon_CP_3229_elements(153);
      gj_l2CacheDaemon_cp_element_group_151 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(151), clk => clk, reset => reset); --
    end block;
    -- CP-element group 152:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 152: predecessors 
    -- CP-element group 152: marked-predecessors 
    -- CP-element group 152: 	185 
    -- CP-element group 152: successors 
    -- CP-element group 152: 	154 
    -- CP-element group 152:  members (3) 
      -- CP-element group 152: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3658_update_start_
      -- CP-element group 152: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3658_Update/$entry
      -- CP-element group 152: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3658_Update/req
      -- 
    req_3687_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3687_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(152), ack => W_data_write_dword_3396_delayed_9_0_3656_inst_req_1); -- 
    l2CacheDaemon_cp_element_group_152: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_152"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= l2CacheDaemon_CP_3229_elements(185);
      gj_l2CacheDaemon_cp_element_group_152 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(152), clk => clk, reset => reset); --
    end block;
    -- CP-element group 153:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 153: predecessors 
    -- CP-element group 153: 	151 
    -- CP-element group 153: successors 
    -- CP-element group 153: marked-successors 
    -- CP-element group 153: 	19 
    -- CP-element group 153: 	38 
    -- CP-element group 153: 	151 
    -- CP-element group 153:  members (3) 
      -- CP-element group 153: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3658_sample_completed_
      -- CP-element group 153: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3658_Sample/$exit
      -- CP-element group 153: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3658_Sample/ack
      -- 
    ack_3683_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 153_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_write_dword_3396_delayed_9_0_3656_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(153)); -- 
    -- CP-element group 154:  transition  input  bypass  pipeline-parent 
    -- CP-element group 154: predecessors 
    -- CP-element group 154: 	152 
    -- CP-element group 154: successors 
    -- CP-element group 154: 	183 
    -- CP-element group 154:  members (3) 
      -- CP-element group 154: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3658_update_completed_
      -- CP-element group 154: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3658_Update/$exit
      -- CP-element group 154: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3658_Update/ack
      -- 
    ack_3688_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 154_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_write_dword_3396_delayed_9_0_3656_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(154)); -- 
    -- CP-element group 155:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 155: predecessors 
    -- CP-element group 155: 	21 
    -- CP-element group 155: 	42 
    -- CP-element group 155: marked-predecessors 
    -- CP-element group 155: 	157 
    -- CP-element group 155: successors 
    -- CP-element group 155: 	157 
    -- CP-element group 155:  members (3) 
      -- CP-element group 155: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3661_sample_start_
      -- CP-element group 155: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3661_Sample/$entry
      -- CP-element group 155: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3661_Sample/req
      -- 
    req_3696_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3696_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(155), ack => W_data_read_dword_3397_delayed_9_0_3659_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_155: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_155"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(21) & l2CacheDaemon_CP_3229_elements(42) & l2CacheDaemon_CP_3229_elements(157);
      gj_l2CacheDaemon_cp_element_group_155 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(155), clk => clk, reset => reset); --
    end block;
    -- CP-element group 156:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 156: predecessors 
    -- CP-element group 156: marked-predecessors 
    -- CP-element group 156: 	185 
    -- CP-element group 156: successors 
    -- CP-element group 156: 	158 
    -- CP-element group 156:  members (3) 
      -- CP-element group 156: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3661_update_start_
      -- CP-element group 156: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3661_Update/$entry
      -- CP-element group 156: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3661_Update/req
      -- 
    req_3701_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3701_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(156), ack => W_data_read_dword_3397_delayed_9_0_3659_inst_req_1); -- 
    l2CacheDaemon_cp_element_group_156: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_156"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= l2CacheDaemon_CP_3229_elements(185);
      gj_l2CacheDaemon_cp_element_group_156 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(156), clk => clk, reset => reset); --
    end block;
    -- CP-element group 157:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 157: predecessors 
    -- CP-element group 157: 	155 
    -- CP-element group 157: successors 
    -- CP-element group 157: marked-successors 
    -- CP-element group 157: 	19 
    -- CP-element group 157: 	38 
    -- CP-element group 157: 	155 
    -- CP-element group 157:  members (3) 
      -- CP-element group 157: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3661_sample_completed_
      -- CP-element group 157: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3661_Sample/$exit
      -- CP-element group 157: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3661_Sample/ack
      -- 
    ack_3697_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 157_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_read_dword_3397_delayed_9_0_3659_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(157)); -- 
    -- CP-element group 158:  transition  input  bypass  pipeline-parent 
    -- CP-element group 158: predecessors 
    -- CP-element group 158: 	156 
    -- CP-element group 158: successors 
    -- CP-element group 158: 	183 
    -- CP-element group 158:  members (3) 
      -- CP-element group 158: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3661_update_completed_
      -- CP-element group 158: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3661_Update/$exit
      -- CP-element group 158: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3661_Update/ack
      -- 
    ack_3702_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 158_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_read_dword_3397_delayed_9_0_3659_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(158)); -- 
    -- CP-element group 159:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 159: predecessors 
    -- CP-element group 159: 	90 
    -- CP-element group 159: 	102 
    -- CP-element group 159: marked-predecessors 
    -- CP-element group 159: 	161 
    -- CP-element group 159: successors 
    -- CP-element group 159: 	161 
    -- CP-element group 159:  members (3) 
      -- CP-element group 159: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3664_sample_start_
      -- CP-element group 159: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3664_Sample/$entry
      -- CP-element group 159: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3664_Sample/req
      -- 
    req_3710_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3710_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(159), ack => W_data_write_new_line_3398_delayed_4_0_3662_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_159: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_159"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(90) & l2CacheDaemon_CP_3229_elements(102) & l2CacheDaemon_CP_3229_elements(161);
      gj_l2CacheDaemon_cp_element_group_159 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(159), clk => clk, reset => reset); --
    end block;
    -- CP-element group 160:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 160: predecessors 
    -- CP-element group 160: marked-predecessors 
    -- CP-element group 160: 	185 
    -- CP-element group 160: successors 
    -- CP-element group 160: 	162 
    -- CP-element group 160:  members (3) 
      -- CP-element group 160: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3664_update_start_
      -- CP-element group 160: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3664_Update/$entry
      -- CP-element group 160: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3664_Update/req
      -- 
    req_3715_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3715_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(160), ack => W_data_write_new_line_3398_delayed_4_0_3662_inst_req_1); -- 
    l2CacheDaemon_cp_element_group_160: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_160"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= l2CacheDaemon_CP_3229_elements(185);
      gj_l2CacheDaemon_cp_element_group_160 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(160), clk => clk, reset => reset); --
    end block;
    -- CP-element group 161:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 161: predecessors 
    -- CP-element group 161: 	159 
    -- CP-element group 161: successors 
    -- CP-element group 161: marked-successors 
    -- CP-element group 161: 	88 
    -- CP-element group 161: 	159 
    -- CP-element group 161: 	100 
    -- CP-element group 161:  members (3) 
      -- CP-element group 161: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3664_sample_completed_
      -- CP-element group 161: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3664_Sample/$exit
      -- CP-element group 161: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3664_Sample/ack
      -- 
    ack_3711_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 161_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_write_new_line_3398_delayed_4_0_3662_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(161)); -- 
    -- CP-element group 162:  transition  input  bypass  pipeline-parent 
    -- CP-element group 162: predecessors 
    -- CP-element group 162: 	160 
    -- CP-element group 162: successors 
    -- CP-element group 162: 	183 
    -- CP-element group 162:  members (3) 
      -- CP-element group 162: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3664_update_completed_
      -- CP-element group 162: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3664_Update/$exit
      -- CP-element group 162: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3664_Update/ack
      -- 
    ack_3716_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 162_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_data_write_new_line_3398_delayed_4_0_3662_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(162)); -- 
    -- CP-element group 163:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 163: predecessors 
    -- CP-element group 163: 	90 
    -- CP-element group 163: 	106 
    -- CP-element group 163: 	110 
    -- CP-element group 163: 	114 
    -- CP-element group 163: marked-predecessors 
    -- CP-element group 163: 	165 
    -- CP-element group 163: successors 
    -- CP-element group 163: 	165 
    -- CP-element group 163:  members (3) 
      -- CP-element group 163: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3667_sample_start_
      -- CP-element group 163: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3667_Sample/$entry
      -- CP-element group 163: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3667_Sample/req
      -- 
    req_3724_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3724_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(163), ack => W_do_write_replaced_line_to_mem_3399_delayed_4_0_3665_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_163: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_163"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(90) & l2CacheDaemon_CP_3229_elements(106) & l2CacheDaemon_CP_3229_elements(110) & l2CacheDaemon_CP_3229_elements(114) & l2CacheDaemon_CP_3229_elements(165);
      gj_l2CacheDaemon_cp_element_group_163 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(163), clk => clk, reset => reset); --
    end block;
    -- CP-element group 164:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 164: predecessors 
    -- CP-element group 164: marked-predecessors 
    -- CP-element group 164: 	185 
    -- CP-element group 164: successors 
    -- CP-element group 164: 	166 
    -- CP-element group 164:  members (3) 
      -- CP-element group 164: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3667_update_start_
      -- CP-element group 164: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3667_Update/$entry
      -- CP-element group 164: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3667_Update/req
      -- 
    req_3729_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3729_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(164), ack => W_do_write_replaced_line_to_mem_3399_delayed_4_0_3665_inst_req_1); -- 
    l2CacheDaemon_cp_element_group_164: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_164"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= l2CacheDaemon_CP_3229_elements(185);
      gj_l2CacheDaemon_cp_element_group_164 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(164), clk => clk, reset => reset); --
    end block;
    -- CP-element group 165:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 165: predecessors 
    -- CP-element group 165: 	163 
    -- CP-element group 165: successors 
    -- CP-element group 165: marked-successors 
    -- CP-element group 165: 	88 
    -- CP-element group 165: 	104 
    -- CP-element group 165: 	163 
    -- CP-element group 165: 	108 
    -- CP-element group 165: 	112 
    -- CP-element group 165:  members (3) 
      -- CP-element group 165: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3667_sample_completed_
      -- CP-element group 165: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3667_Sample/$exit
      -- CP-element group 165: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3667_Sample/ack
      -- 
    ack_3725_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 165_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_do_write_replaced_line_to_mem_3399_delayed_4_0_3665_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(165)); -- 
    -- CP-element group 166:  transition  input  bypass  pipeline-parent 
    -- CP-element group 166: predecessors 
    -- CP-element group 166: 	164 
    -- CP-element group 166: successors 
    -- CP-element group 166: 	183 
    -- CP-element group 166:  members (3) 
      -- CP-element group 166: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3667_update_completed_
      -- CP-element group 166: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3667_Update/$exit
      -- CP-element group 166: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3667_Update/ack
      -- 
    ack_3730_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 166_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_do_write_replaced_line_to_mem_3399_delayed_4_0_3665_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(166)); -- 
    -- CP-element group 167:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 167: predecessors 
    -- CP-element group 167: 	21 
    -- CP-element group 167: marked-predecessors 
    -- CP-element group 167: 	169 
    -- CP-element group 167: successors 
    -- CP-element group 167: 	169 
    -- CP-element group 167:  members (3) 
      -- CP-element group 167: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3670_sample_start_
      -- CP-element group 167: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3670_Sample/$entry
      -- CP-element group 167: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3670_Sample/req
      -- 
    req_3738_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3738_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(167), ack => W_byte_mask_3400_delayed_9_0_3668_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_167: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_167"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(21) & l2CacheDaemon_CP_3229_elements(169);
      gj_l2CacheDaemon_cp_element_group_167 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(167), clk => clk, reset => reset); --
    end block;
    -- CP-element group 168:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 168: predecessors 
    -- CP-element group 168: marked-predecessors 
    -- CP-element group 168: 	185 
    -- CP-element group 168: successors 
    -- CP-element group 168: 	170 
    -- CP-element group 168:  members (3) 
      -- CP-element group 168: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3670_Update/req
      -- CP-element group 168: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3670_Update/$entry
      -- CP-element group 168: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3670_update_start_
      -- 
    req_3743_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3743_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(168), ack => W_byte_mask_3400_delayed_9_0_3668_inst_req_1); -- 
    l2CacheDaemon_cp_element_group_168: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_168"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= l2CacheDaemon_CP_3229_elements(185);
      gj_l2CacheDaemon_cp_element_group_168 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(168), clk => clk, reset => reset); --
    end block;
    -- CP-element group 169:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 169: predecessors 
    -- CP-element group 169: 	167 
    -- CP-element group 169: successors 
    -- CP-element group 169: marked-successors 
    -- CP-element group 169: 	19 
    -- CP-element group 169: 	167 
    -- CP-element group 169:  members (3) 
      -- CP-element group 169: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3670_sample_completed_
      -- CP-element group 169: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3670_Sample/$exit
      -- CP-element group 169: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3670_Sample/ack
      -- 
    ack_3739_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 169_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_byte_mask_3400_delayed_9_0_3668_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(169)); -- 
    -- CP-element group 170:  transition  input  bypass  pipeline-parent 
    -- CP-element group 170: predecessors 
    -- CP-element group 170: 	168 
    -- CP-element group 170: successors 
    -- CP-element group 170: 	183 
    -- CP-element group 170:  members (3) 
      -- CP-element group 170: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3670_Update/ack
      -- CP-element group 170: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3670_Update/$exit
      -- CP-element group 170: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3670_update_completed_
      -- 
    ack_3744_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 170_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_byte_mask_3400_delayed_9_0_3668_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(170)); -- 
    -- CP-element group 171:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 171: predecessors 
    -- CP-element group 171: 	90 
    -- CP-element group 171: 	138 
    -- CP-element group 171: marked-predecessors 
    -- CP-element group 171: 	173 
    -- CP-element group 171: successors 
    -- CP-element group 171: 	173 
    -- CP-element group 171:  members (3) 
      -- CP-element group 171: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3673_Sample/$entry
      -- CP-element group 171: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3673_sample_start_
      -- CP-element group 171: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3673_Sample/req
      -- 
    req_3752_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3752_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(171), ack => W_line_id_3401_delayed_4_0_3671_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_171: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_171"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(90) & l2CacheDaemon_CP_3229_elements(138) & l2CacheDaemon_CP_3229_elements(173);
      gj_l2CacheDaemon_cp_element_group_171 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(171), clk => clk, reset => reset); --
    end block;
    -- CP-element group 172:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 172: predecessors 
    -- CP-element group 172: marked-predecessors 
    -- CP-element group 172: 	185 
    -- CP-element group 172: successors 
    -- CP-element group 172: 	174 
    -- CP-element group 172:  members (3) 
      -- CP-element group 172: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3673_Update/req
      -- CP-element group 172: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3673_Update/$entry
      -- CP-element group 172: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3673_update_start_
      -- 
    req_3757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(172), ack => W_line_id_3401_delayed_4_0_3671_inst_req_1); -- 
    l2CacheDaemon_cp_element_group_172: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_172"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= l2CacheDaemon_CP_3229_elements(185);
      gj_l2CacheDaemon_cp_element_group_172 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(172), clk => clk, reset => reset); --
    end block;
    -- CP-element group 173:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 173: predecessors 
    -- CP-element group 173: 	171 
    -- CP-element group 173: successors 
    -- CP-element group 173: marked-successors 
    -- CP-element group 173: 	88 
    -- CP-element group 173: 	171 
    -- CP-element group 173: 	136 
    -- CP-element group 173:  members (3) 
      -- CP-element group 173: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3673_Sample/$exit
      -- CP-element group 173: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3673_sample_completed_
      -- CP-element group 173: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3673_Sample/ack
      -- 
    ack_3753_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 173_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_line_id_3401_delayed_4_0_3671_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(173)); -- 
    -- CP-element group 174:  transition  input  bypass  pipeline-parent 
    -- CP-element group 174: predecessors 
    -- CP-element group 174: 	172 
    -- CP-element group 174: successors 
    -- CP-element group 174: 	183 
    -- CP-element group 174:  members (3) 
      -- CP-element group 174: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3673_update_completed_
      -- CP-element group 174: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3673_Update/ack
      -- CP-element group 174: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3673_Update/$exit
      -- 
    ack_3758_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 174_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_line_id_3401_delayed_4_0_3671_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(174)); -- 
    -- CP-element group 175:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 175: predecessors 
    -- CP-element group 175: 	21 
    -- CP-element group 175: marked-predecessors 
    -- CP-element group 175: 	177 
    -- CP-element group 175: successors 
    -- CP-element group 175: 	177 
    -- CP-element group 175:  members (3) 
      -- CP-element group 175: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3676_Sample/$entry
      -- CP-element group 175: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3676_Sample/req
      -- CP-element group 175: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3676_sample_start_
      -- 
    req_3766_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3766_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(175), ack => W_pa_dword_id_3402_delayed_9_0_3674_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_175: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_175"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(21) & l2CacheDaemon_CP_3229_elements(177);
      gj_l2CacheDaemon_cp_element_group_175 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(175), clk => clk, reset => reset); --
    end block;
    -- CP-element group 176:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 176: predecessors 
    -- CP-element group 176: marked-predecessors 
    -- CP-element group 176: 	185 
    -- CP-element group 176: successors 
    -- CP-element group 176: 	178 
    -- CP-element group 176:  members (3) 
      -- CP-element group 176: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3676_Update/$entry
      -- CP-element group 176: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3676_update_start_
      -- CP-element group 176: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3676_Update/req
      -- 
    req_3771_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3771_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(176), ack => W_pa_dword_id_3402_delayed_9_0_3674_inst_req_1); -- 
    l2CacheDaemon_cp_element_group_176: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_176"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= l2CacheDaemon_CP_3229_elements(185);
      gj_l2CacheDaemon_cp_element_group_176 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(176), clk => clk, reset => reset); --
    end block;
    -- CP-element group 177:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 177: predecessors 
    -- CP-element group 177: 	175 
    -- CP-element group 177: successors 
    -- CP-element group 177: marked-successors 
    -- CP-element group 177: 	19 
    -- CP-element group 177: 	175 
    -- CP-element group 177:  members (3) 
      -- CP-element group 177: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3676_Sample/ack
      -- CP-element group 177: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3676_Sample/$exit
      -- CP-element group 177: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3676_sample_completed_
      -- 
    ack_3767_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 177_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_pa_dword_id_3402_delayed_9_0_3674_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(177)); -- 
    -- CP-element group 178:  transition  input  bypass  pipeline-parent 
    -- CP-element group 178: predecessors 
    -- CP-element group 178: 	176 
    -- CP-element group 178: successors 
    -- CP-element group 178: 	183 
    -- CP-element group 178:  members (3) 
      -- CP-element group 178: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3676_Update/$exit
      -- CP-element group 178: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3676_Update/ack
      -- CP-element group 178: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3676_update_completed_
      -- 
    ack_3772_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 178_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_pa_dword_id_3402_delayed_9_0_3674_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(178)); -- 
    -- CP-element group 179:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 179: predecessors 
    -- CP-element group 179: 	21 
    -- CP-element group 179: marked-predecessors 
    -- CP-element group 179: 	181 
    -- CP-element group 179: successors 
    -- CP-element group 179: 	181 
    -- CP-element group 179:  members (3) 
      -- CP-element group 179: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3679_Sample/req
      -- CP-element group 179: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3679_Sample/$entry
      -- CP-element group 179: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3679_sample_start_
      -- 
    req_3780_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3780_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(179), ack => W_wdata_3403_delayed_9_0_3677_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_179: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_179"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(21) & l2CacheDaemon_CP_3229_elements(181);
      gj_l2CacheDaemon_cp_element_group_179 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(179), clk => clk, reset => reset); --
    end block;
    -- CP-element group 180:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 180: predecessors 
    -- CP-element group 180: marked-predecessors 
    -- CP-element group 180: 	185 
    -- CP-element group 180: successors 
    -- CP-element group 180: 	182 
    -- CP-element group 180:  members (3) 
      -- CP-element group 180: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3679_Update/$entry
      -- CP-element group 180: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3679_update_start_
      -- CP-element group 180: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3679_Update/req
      -- 
    req_3785_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3785_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(180), ack => W_wdata_3403_delayed_9_0_3677_inst_req_1); -- 
    l2CacheDaemon_cp_element_group_180: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_180"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= l2CacheDaemon_CP_3229_elements(185);
      gj_l2CacheDaemon_cp_element_group_180 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(180), clk => clk, reset => reset); --
    end block;
    -- CP-element group 181:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 181: predecessors 
    -- CP-element group 181: 	179 
    -- CP-element group 181: successors 
    -- CP-element group 181: marked-successors 
    -- CP-element group 181: 	19 
    -- CP-element group 181: 	179 
    -- CP-element group 181:  members (3) 
      -- CP-element group 181: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3679_Sample/ack
      -- CP-element group 181: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3679_Sample/$exit
      -- CP-element group 181: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3679_sample_completed_
      -- 
    ack_3781_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 181_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_wdata_3403_delayed_9_0_3677_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(181)); -- 
    -- CP-element group 182:  transition  input  bypass  pipeline-parent 
    -- CP-element group 182: predecessors 
    -- CP-element group 182: 	180 
    -- CP-element group 182: successors 
    -- CP-element group 182: 	183 
    -- CP-element group 182:  members (3) 
      -- CP-element group 182: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3679_Update/ack
      -- CP-element group 182: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3679_update_completed_
      -- CP-element group 182: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3679_Update/$exit
      -- 
    ack_3786_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 182_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_wdata_3403_delayed_9_0_3677_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(182)); -- 
    -- CP-element group 183:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 183: predecessors 
    -- CP-element group 183: 	170 
    -- CP-element group 183: 	174 
    -- CP-element group 183: 	146 
    -- CP-element group 183: 	154 
    -- CP-element group 183: 	158 
    -- CP-element group 183: 	162 
    -- CP-element group 183: 	182 
    -- CP-element group 183: 	178 
    -- CP-element group 183: 	134 
    -- CP-element group 183: 	150 
    -- CP-element group 183: 	166 
    -- CP-element group 183: marked-predecessors 
    -- CP-element group 183: 	185 
    -- CP-element group 183: successors 
    -- CP-element group 183: 	185 
    -- CP-element group 183:  members (3) 
      -- CP-element group 183: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3693_sample_start_
      -- CP-element group 183: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3693_Sample/crr
      -- CP-element group 183: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3693_Sample/$entry
      -- 
    crr_3794_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3794_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(183), ack => call_stmt_3693_call_req_0); -- 
    l2CacheDaemon_cp_element_group_183: block -- 
      constant place_capacities: IntegerArray(0 to 11) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1,10 => 1,11 => 1);
      constant place_markings: IntegerArray(0 to 11)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 1);
      constant place_delays: IntegerArray(0 to 11) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0,10 => 0,11 => 1);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_183"; 
      signal preds: BooleanArray(1 to 12); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(170) & l2CacheDaemon_CP_3229_elements(174) & l2CacheDaemon_CP_3229_elements(146) & l2CacheDaemon_CP_3229_elements(154) & l2CacheDaemon_CP_3229_elements(158) & l2CacheDaemon_CP_3229_elements(162) & l2CacheDaemon_CP_3229_elements(182) & l2CacheDaemon_CP_3229_elements(178) & l2CacheDaemon_CP_3229_elements(134) & l2CacheDaemon_CP_3229_elements(150) & l2CacheDaemon_CP_3229_elements(166) & l2CacheDaemon_CP_3229_elements(185);
      gj_l2CacheDaemon_cp_element_group_183 : generic_join generic map(name => joinName, number_of_predecessors => 12, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(183), clk => clk, reset => reset); --
    end block;
    -- CP-element group 184:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 184: predecessors 
    -- CP-element group 184: marked-predecessors 
    -- CP-element group 184: 	220 
    -- CP-element group 184: 	196 
    -- CP-element group 184: successors 
    -- CP-element group 184: 	186 
    -- CP-element group 184:  members (3) 
      -- CP-element group 184: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3693_update_start_
      -- CP-element group 184: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3693_Update/ccr
      -- CP-element group 184: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3693_Update/$entry
      -- 
    ccr_3799_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3799_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(184), ack => call_stmt_3693_call_req_1); -- 
    l2CacheDaemon_cp_element_group_184: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_184"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(220) & l2CacheDaemon_CP_3229_elements(196);
      gj_l2CacheDaemon_cp_element_group_184 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(184), clk => clk, reset => reset); --
    end block;
    -- CP-element group 185:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 185: predecessors 
    -- CP-element group 185: 	183 
    -- CP-element group 185: successors 
    -- CP-element group 185: marked-successors 
    -- CP-element group 185: 	172 
    -- CP-element group 185: 	144 
    -- CP-element group 185: 	148 
    -- CP-element group 185: 	156 
    -- CP-element group 185: 	160 
    -- CP-element group 185: 	164 
    -- CP-element group 185: 	132 
    -- CP-element group 185: 	183 
    -- CP-element group 185: 	176 
    -- CP-element group 185: 	180 
    -- CP-element group 185: 	152 
    -- CP-element group 185: 	168 
    -- CP-element group 185:  members (3) 
      -- CP-element group 185: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3693_sample_completed_
      -- CP-element group 185: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3693_Sample/$exit
      -- CP-element group 185: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3693_Sample/cra
      -- 
    cra_3795_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 185_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_3693_call_ack_0, ack => l2CacheDaemon_CP_3229_elements(185)); -- 
    -- CP-element group 186:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 186: predecessors 
    -- CP-element group 186: 	184 
    -- CP-element group 186: successors 
    -- CP-element group 186: 	218 
    -- CP-element group 186: 	195 
    -- CP-element group 186:  members (3) 
      -- CP-element group 186: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3693_update_completed_
      -- CP-element group 186: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3693_Update/$exit
      -- CP-element group 186: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3693_Update/cca
      -- 
    cca_3800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 186_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_3693_call_ack_1, ack => l2CacheDaemon_CP_3229_elements(186)); -- 
    -- CP-element group 187:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 187: predecessors 
    -- CP-element group 187: 	21 
    -- CP-element group 187: marked-predecessors 
    -- CP-element group 187: 	189 
    -- CP-element group 187: successors 
    -- CP-element group 187: 	189 
    -- CP-element group 187:  members (3) 
      -- CP-element group 187: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3702_Sample/req
      -- CP-element group 187: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3702_Sample/$entry
      -- CP-element group 187: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3702_sample_start_
      -- 
    req_3808_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3808_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(187), ack => W_rwbar_3417_delayed_10_0_3700_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_187: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_187"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(21) & l2CacheDaemon_CP_3229_elements(189);
      gj_l2CacheDaemon_cp_element_group_187 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(187), clk => clk, reset => reset); --
    end block;
    -- CP-element group 188:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 188: predecessors 
    -- CP-element group 188: marked-predecessors 
    -- CP-element group 188: 	196 
    -- CP-element group 188: successors 
    -- CP-element group 188: 	190 
    -- CP-element group 188:  members (3) 
      -- CP-element group 188: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3702_update_start_
      -- CP-element group 188: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3702_Update/$entry
      -- CP-element group 188: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3702_Update/req
      -- 
    req_3813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(188), ack => W_rwbar_3417_delayed_10_0_3700_inst_req_1); -- 
    l2CacheDaemon_cp_element_group_188: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_188"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= l2CacheDaemon_CP_3229_elements(196);
      gj_l2CacheDaemon_cp_element_group_188 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(188), clk => clk, reset => reset); --
    end block;
    -- CP-element group 189:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 189: predecessors 
    -- CP-element group 189: 	187 
    -- CP-element group 189: successors 
    -- CP-element group 189: marked-successors 
    -- CP-element group 189: 	19 
    -- CP-element group 189: 	187 
    -- CP-element group 189:  members (3) 
      -- CP-element group 189: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3702_sample_completed_
      -- CP-element group 189: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3702_Sample/$exit
      -- CP-element group 189: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3702_Sample/ack
      -- 
    ack_3809_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 189_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_3417_delayed_10_0_3700_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(189)); -- 
    -- CP-element group 190:  transition  input  bypass  pipeline-parent 
    -- CP-element group 190: predecessors 
    -- CP-element group 190: 	188 
    -- CP-element group 190: successors 
    -- CP-element group 190: 	195 
    -- CP-element group 190:  members (3) 
      -- CP-element group 190: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3702_Update/ack
      -- CP-element group 190: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3702_update_completed_
      -- CP-element group 190: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3702_Update/$exit
      -- 
    ack_3814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 190_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_rwbar_3417_delayed_10_0_3700_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(190)); -- 
    -- CP-element group 191:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 191: predecessors 
    -- CP-element group 191: 	21 
    -- CP-element group 191: 	42 
    -- CP-element group 191: marked-predecessors 
    -- CP-element group 191: 	193 
    -- CP-element group 191: successors 
    -- CP-element group 191: 	193 
    -- CP-element group 191:  members (3) 
      -- CP-element group 191: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3715_Sample/$entry
      -- CP-element group 191: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3715_Sample/req
      -- CP-element group 191: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3715_sample_start_
      -- 
    req_3822_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3822_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(191), ack => W_send_response_3424_delayed_10_0_3713_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_191: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_191"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(21) & l2CacheDaemon_CP_3229_elements(42) & l2CacheDaemon_CP_3229_elements(193);
      gj_l2CacheDaemon_cp_element_group_191 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(191), clk => clk, reset => reset); --
    end block;
    -- CP-element group 192:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 192: predecessors 
    -- CP-element group 192: marked-predecessors 
    -- CP-element group 192: 	196 
    -- CP-element group 192: successors 
    -- CP-element group 192: 	194 
    -- CP-element group 192:  members (3) 
      -- CP-element group 192: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3715_Update/$entry
      -- CP-element group 192: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3715_update_start_
      -- CP-element group 192: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3715_Update/req
      -- 
    req_3827_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3827_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(192), ack => W_send_response_3424_delayed_10_0_3713_inst_req_1); -- 
    l2CacheDaemon_cp_element_group_192: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_192"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= l2CacheDaemon_CP_3229_elements(196);
      gj_l2CacheDaemon_cp_element_group_192 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(192), clk => clk, reset => reset); --
    end block;
    -- CP-element group 193:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 193: predecessors 
    -- CP-element group 193: 	191 
    -- CP-element group 193: successors 
    -- CP-element group 193: marked-successors 
    -- CP-element group 193: 	19 
    -- CP-element group 193: 	38 
    -- CP-element group 193: 	191 
    -- CP-element group 193:  members (3) 
      -- CP-element group 193: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3715_Sample/$exit
      -- CP-element group 193: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3715_Sample/ack
      -- CP-element group 193: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3715_sample_completed_
      -- 
    ack_3823_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 193_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send_response_3424_delayed_10_0_3713_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(193)); -- 
    -- CP-element group 194:  transition  input  bypass  pipeline-parent 
    -- CP-element group 194: predecessors 
    -- CP-element group 194: 	192 
    -- CP-element group 194: successors 
    -- CP-element group 194: 	195 
    -- CP-element group 194:  members (3) 
      -- CP-element group 194: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3715_Update/$exit
      -- CP-element group 194: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3715_Update/ack
      -- CP-element group 194: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3715_update_completed_
      -- 
    ack_3828_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 194_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_send_response_3424_delayed_10_0_3713_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(194)); -- 
    -- CP-element group 195:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 195: predecessors 
    -- CP-element group 195: 	194 
    -- CP-element group 195: 	186 
    -- CP-element group 195: 	190 
    -- CP-element group 195: marked-predecessors 
    -- CP-element group 195: 	197 
    -- CP-element group 195: successors 
    -- CP-element group 195: 	196 
    -- CP-element group 195:  members (3) 
      -- CP-element group 195: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_L2_RESPONSE_3717_Sample/$entry
      -- CP-element group 195: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_L2_RESPONSE_3717_Sample/req
      -- CP-element group 195: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_L2_RESPONSE_3717_sample_start_
      -- 
    req_3836_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3836_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(195), ack => WPIPE_L2_RESPONSE_3717_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_195: block -- 
      constant place_capacities: IntegerArray(0 to 3) := (0 => 1,1 => 1,2 => 1,3 => 1);
      constant place_markings: IntegerArray(0 to 3)  := (0 => 0,1 => 0,2 => 0,3 => 1);
      constant place_delays: IntegerArray(0 to 3) := (0 => 0,1 => 0,2 => 0,3 => 0);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_195"; 
      signal preds: BooleanArray(1 to 4); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(194) & l2CacheDaemon_CP_3229_elements(186) & l2CacheDaemon_CP_3229_elements(190) & l2CacheDaemon_CP_3229_elements(197);
      gj_l2CacheDaemon_cp_element_group_195 : generic_join generic map(name => joinName, number_of_predecessors => 4, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(195), clk => clk, reset => reset); --
    end block;
    -- CP-element group 196:  fork  transition  input  output  bypass  pipeline-parent 
    -- CP-element group 196: predecessors 
    -- CP-element group 196: 	195 
    -- CP-element group 196: successors 
    -- CP-element group 196: 	197 
    -- CP-element group 196: marked-successors 
    -- CP-element group 196: 	192 
    -- CP-element group 196: 	188 
    -- CP-element group 196: 	184 
    -- CP-element group 196:  members (6) 
      -- CP-element group 196: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_L2_RESPONSE_3717_Update/$entry
      -- CP-element group 196: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_L2_RESPONSE_3717_update_start_
      -- CP-element group 196: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_L2_RESPONSE_3717_Sample/ack
      -- CP-element group 196: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_L2_RESPONSE_3717_Sample/$exit
      -- CP-element group 196: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_L2_RESPONSE_3717_Update/req
      -- CP-element group 196: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_L2_RESPONSE_3717_sample_completed_
      -- 
    ack_3837_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 196_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_L2_RESPONSE_3717_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(196)); -- 
    req_3841_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3841_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(196), ack => WPIPE_L2_RESPONSE_3717_inst_req_1); -- 
    -- CP-element group 197:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 197: predecessors 
    -- CP-element group 197: 	196 
    -- CP-element group 197: successors 
    -- CP-element group 197: 	223 
    -- CP-element group 197: marked-successors 
    -- CP-element group 197: 	195 
    -- CP-element group 197:  members (3) 
      -- CP-element group 197: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_L2_RESPONSE_3717_Update/$exit
      -- CP-element group 197: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_L2_RESPONSE_3717_Update/ack
      -- CP-element group 197: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/WPIPE_L2_RESPONSE_3717_update_completed_
      -- 
    ack_3842_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 197_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_L2_RESPONSE_3717_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(197)); -- 
    -- CP-element group 198:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 198: predecessors 
    -- CP-element group 198: 	90 
    -- CP-element group 198: 	106 
    -- CP-element group 198: 	110 
    -- CP-element group 198: 	98 
    -- CP-element group 198: 	114 
    -- CP-element group 198: marked-predecessors 
    -- CP-element group 198: 	200 
    -- CP-element group 198: successors 
    -- CP-element group 198: 	200 
    -- CP-element group 198:  members (3) 
      -- CP-element group 198: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3731_sample_start_
      -- CP-element group 198: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3731_Sample/req
      -- CP-element group 198: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3731_Sample/$entry
      -- 
    req_3850_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3850_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(198), ack => W_call_write_mem_3437_delayed_5_0_3729_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_198: block -- 
      constant place_capacities: IntegerArray(0 to 5) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1);
      constant place_markings: IntegerArray(0 to 5)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant place_delays: IntegerArray(0 to 5) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 1);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_198"; 
      signal preds: BooleanArray(1 to 6); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(90) & l2CacheDaemon_CP_3229_elements(106) & l2CacheDaemon_CP_3229_elements(110) & l2CacheDaemon_CP_3229_elements(98) & l2CacheDaemon_CP_3229_elements(114) & l2CacheDaemon_CP_3229_elements(200);
      gj_l2CacheDaemon_cp_element_group_198 : generic_join generic map(name => joinName, number_of_predecessors => 6, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(198), clk => clk, reset => reset); --
    end block;
    -- CP-element group 199:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 199: predecessors 
    -- CP-element group 199: marked-predecessors 
    -- CP-element group 199: 	220 
    -- CP-element group 199: successors 
    -- CP-element group 199: 	201 
    -- CP-element group 199:  members (3) 
      -- CP-element group 199: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3731_Update/req
      -- CP-element group 199: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3731_update_start_
      -- CP-element group 199: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3731_Update/$entry
      -- 
    req_3855_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3855_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(199), ack => W_call_write_mem_3437_delayed_5_0_3729_inst_req_1); -- 
    l2CacheDaemon_cp_element_group_199: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_199"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= l2CacheDaemon_CP_3229_elements(220);
      gj_l2CacheDaemon_cp_element_group_199 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(199), clk => clk, reset => reset); --
    end block;
    -- CP-element group 200:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 200: predecessors 
    -- CP-element group 200: 	198 
    -- CP-element group 200: successors 
    -- CP-element group 200: marked-successors 
    -- CP-element group 200: 	88 
    -- CP-element group 200: 	104 
    -- CP-element group 200: 	108 
    -- CP-element group 200: 	198 
    -- CP-element group 200: 	96 
    -- CP-element group 200: 	112 
    -- CP-element group 200:  members (3) 
      -- CP-element group 200: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3731_Sample/ack
      -- CP-element group 200: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3731_sample_completed_
      -- CP-element group 200: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3731_Sample/$exit
      -- 
    ack_3851_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 200_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_call_write_mem_3437_delayed_5_0_3729_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(200)); -- 
    -- CP-element group 201:  transition  input  bypass  pipeline-parent 
    -- CP-element group 201: predecessors 
    -- CP-element group 201: 	199 
    -- CP-element group 201: successors 
    -- CP-element group 201: 	218 
    -- CP-element group 201:  members (3) 
      -- CP-element group 201: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3731_Update/ack
      -- CP-element group 201: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3731_Update/$exit
      -- CP-element group 201: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3731_update_completed_
      -- 
    ack_3856_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 201_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_call_write_mem_3437_delayed_5_0_3729_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(201)); -- 
    -- CP-element group 202:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 202: predecessors 
    -- CP-element group 202: 	90 
    -- CP-element group 202: 	98 
    -- CP-element group 202: marked-predecessors 
    -- CP-element group 202: 	204 
    -- CP-element group 202: successors 
    -- CP-element group 202: 	204 
    -- CP-element group 202:  members (3) 
      -- CP-element group 202: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3734_sample_start_
      -- CP-element group 202: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3734_Sample/$entry
      -- CP-element group 202: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3734_Sample/req
      -- 
    req_3864_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3864_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(202), ack => W_do_read_line_from_mem_3438_delayed_5_0_3732_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_202: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_202"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(90) & l2CacheDaemon_CP_3229_elements(98) & l2CacheDaemon_CP_3229_elements(204);
      gj_l2CacheDaemon_cp_element_group_202 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(202), clk => clk, reset => reset); --
    end block;
    -- CP-element group 203:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 203: predecessors 
    -- CP-element group 203: marked-predecessors 
    -- CP-element group 203: 	220 
    -- CP-element group 203: successors 
    -- CP-element group 203: 	205 
    -- CP-element group 203:  members (3) 
      -- CP-element group 203: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3734_update_start_
      -- CP-element group 203: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3734_Update/$entry
      -- CP-element group 203: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3734_Update/req
      -- 
    req_3869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(203), ack => W_do_read_line_from_mem_3438_delayed_5_0_3732_inst_req_1); -- 
    l2CacheDaemon_cp_element_group_203: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_203"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= l2CacheDaemon_CP_3229_elements(220);
      gj_l2CacheDaemon_cp_element_group_203 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(203), clk => clk, reset => reset); --
    end block;
    -- CP-element group 204:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 204: predecessors 
    -- CP-element group 204: 	202 
    -- CP-element group 204: successors 
    -- CP-element group 204: marked-successors 
    -- CP-element group 204: 	88 
    -- CP-element group 204: 	202 
    -- CP-element group 204: 	96 
    -- CP-element group 204:  members (3) 
      -- CP-element group 204: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3734_sample_completed_
      -- CP-element group 204: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3734_Sample/$exit
      -- CP-element group 204: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3734_Sample/ack
      -- 
    ack_3865_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 204_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_do_read_line_from_mem_3438_delayed_5_0_3732_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(204)); -- 
    -- CP-element group 205:  transition  input  bypass  pipeline-parent 
    -- CP-element group 205: predecessors 
    -- CP-element group 205: 	203 
    -- CP-element group 205: successors 
    -- CP-element group 205: 	218 
    -- CP-element group 205:  members (3) 
      -- CP-element group 205: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3734_update_completed_
      -- CP-element group 205: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3734_Update/$exit
      -- CP-element group 205: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3734_Update/ack
      -- 
    ack_3870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 205_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_do_read_line_from_mem_3438_delayed_5_0_3732_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(205)); -- 
    -- CP-element group 206:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 206: predecessors 
    -- CP-element group 206: 	90 
    -- CP-element group 206: 	106 
    -- CP-element group 206: 	110 
    -- CP-element group 206: 	114 
    -- CP-element group 206: marked-predecessors 
    -- CP-element group 206: 	208 
    -- CP-element group 206: successors 
    -- CP-element group 206: 	208 
    -- CP-element group 206:  members (3) 
      -- CP-element group 206: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3737_sample_start_
      -- CP-element group 206: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3737_Sample/$entry
      -- CP-element group 206: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3737_Sample/req
      -- 
    req_3878_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3878_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(206), ack => W_do_write_replaced_line_to_mem_3439_delayed_5_0_3735_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_206: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_206"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(90) & l2CacheDaemon_CP_3229_elements(106) & l2CacheDaemon_CP_3229_elements(110) & l2CacheDaemon_CP_3229_elements(114) & l2CacheDaemon_CP_3229_elements(208);
      gj_l2CacheDaemon_cp_element_group_206 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(206), clk => clk, reset => reset); --
    end block;
    -- CP-element group 207:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 207: predecessors 
    -- CP-element group 207: marked-predecessors 
    -- CP-element group 207: 	220 
    -- CP-element group 207: successors 
    -- CP-element group 207: 	209 
    -- CP-element group 207:  members (3) 
      -- CP-element group 207: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3737_update_start_
      -- CP-element group 207: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3737_Update/$entry
      -- CP-element group 207: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3737_Update/req
      -- 
    req_3883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(207), ack => W_do_write_replaced_line_to_mem_3439_delayed_5_0_3735_inst_req_1); -- 
    l2CacheDaemon_cp_element_group_207: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_207"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= l2CacheDaemon_CP_3229_elements(220);
      gj_l2CacheDaemon_cp_element_group_207 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(207), clk => clk, reset => reset); --
    end block;
    -- CP-element group 208:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 208: predecessors 
    -- CP-element group 208: 	206 
    -- CP-element group 208: successors 
    -- CP-element group 208: marked-successors 
    -- CP-element group 208: 	88 
    -- CP-element group 208: 	206 
    -- CP-element group 208: 	104 
    -- CP-element group 208: 	108 
    -- CP-element group 208: 	112 
    -- CP-element group 208:  members (3) 
      -- CP-element group 208: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3737_sample_completed_
      -- CP-element group 208: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3737_Sample/$exit
      -- CP-element group 208: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3737_Sample/ack
      -- 
    ack_3879_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 208_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_do_write_replaced_line_to_mem_3439_delayed_5_0_3735_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(208)); -- 
    -- CP-element group 209:  transition  input  bypass  pipeline-parent 
    -- CP-element group 209: predecessors 
    -- CP-element group 209: 	207 
    -- CP-element group 209: successors 
    -- CP-element group 209: 	218 
    -- CP-element group 209:  members (3) 
      -- CP-element group 209: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3737_update_completed_
      -- CP-element group 209: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3737_Update/$exit
      -- CP-element group 209: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3737_Update/ack
      -- 
    ack_3884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 209_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_do_write_replaced_line_to_mem_3439_delayed_5_0_3735_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(209)); -- 
    -- CP-element group 210:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 210: predecessors 
    -- CP-element group 210: 	90 
    -- CP-element group 210: marked-predecessors 
    -- CP-element group 210: 	212 
    -- CP-element group 210: successors 
    -- CP-element group 210: 	212 
    -- CP-element group 210:  members (3) 
      -- CP-element group 210: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3740_sample_start_
      -- CP-element group 210: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3740_Sample/$entry
      -- CP-element group 210: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3740_Sample/req
      -- 
    req_3892_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3892_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(210), ack => W_dirty_word_mask_3440_delayed_5_0_3738_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_210: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_210"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(90) & l2CacheDaemon_CP_3229_elements(212);
      gj_l2CacheDaemon_cp_element_group_210 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(210), clk => clk, reset => reset); --
    end block;
    -- CP-element group 211:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 211: predecessors 
    -- CP-element group 211: marked-predecessors 
    -- CP-element group 211: 	220 
    -- CP-element group 211: successors 
    -- CP-element group 211: 	213 
    -- CP-element group 211:  members (3) 
      -- CP-element group 211: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3740_update_start_
      -- CP-element group 211: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3740_Update/$entry
      -- CP-element group 211: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3740_Update/req
      -- 
    req_3897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(211), ack => W_dirty_word_mask_3440_delayed_5_0_3738_inst_req_1); -- 
    l2CacheDaemon_cp_element_group_211: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_211"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= l2CacheDaemon_CP_3229_elements(220);
      gj_l2CacheDaemon_cp_element_group_211 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(211), clk => clk, reset => reset); --
    end block;
    -- CP-element group 212:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 212: predecessors 
    -- CP-element group 212: 	210 
    -- CP-element group 212: successors 
    -- CP-element group 212: marked-successors 
    -- CP-element group 212: 	88 
    -- CP-element group 212: 	210 
    -- CP-element group 212:  members (3) 
      -- CP-element group 212: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3740_sample_completed_
      -- CP-element group 212: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3740_Sample/$exit
      -- CP-element group 212: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3740_Sample/ack
      -- 
    ack_3893_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 212_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_dirty_word_mask_3440_delayed_5_0_3738_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(212)); -- 
    -- CP-element group 213:  transition  input  bypass  pipeline-parent 
    -- CP-element group 213: predecessors 
    -- CP-element group 213: 	211 
    -- CP-element group 213: successors 
    -- CP-element group 213: 	218 
    -- CP-element group 213:  members (3) 
      -- CP-element group 213: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3740_update_completed_
      -- CP-element group 213: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3740_Update/$exit
      -- CP-element group 213: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3740_Update/ack
      -- 
    ack_3898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 213_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_dirty_word_mask_3440_delayed_5_0_3738_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(213)); -- 
    -- CP-element group 214:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 214: predecessors 
    -- CP-element group 214: 	90 
    -- CP-element group 214: 	94 
    -- CP-element group 214: 	122 
    -- CP-element group 214: 	118 
    -- CP-element group 214: marked-predecessors 
    -- CP-element group 214: 	216 
    -- CP-element group 214: successors 
    -- CP-element group 214: 	216 
    -- CP-element group 214:  members (3) 
      -- CP-element group 214: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3743_sample_start_
      -- CP-element group 214: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3743_Sample/$entry
      -- CP-element group 214: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3743_Sample/req
      -- 
    req_3906_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3906_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(214), ack => W_write_back_line_address_3441_delayed_5_0_3741_inst_req_0); -- 
    l2CacheDaemon_cp_element_group_214: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 1);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_214"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(90) & l2CacheDaemon_CP_3229_elements(94) & l2CacheDaemon_CP_3229_elements(122) & l2CacheDaemon_CP_3229_elements(118) & l2CacheDaemon_CP_3229_elements(216);
      gj_l2CacheDaemon_cp_element_group_214 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(214), clk => clk, reset => reset); --
    end block;
    -- CP-element group 215:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 215: predecessors 
    -- CP-element group 215: marked-predecessors 
    -- CP-element group 215: 	220 
    -- CP-element group 215: successors 
    -- CP-element group 215: 	217 
    -- CP-element group 215:  members (3) 
      -- CP-element group 215: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3743_update_start_
      -- CP-element group 215: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3743_Update/$entry
      -- CP-element group 215: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3743_Update/req
      -- 
    req_3911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(215), ack => W_write_back_line_address_3441_delayed_5_0_3741_inst_req_1); -- 
    l2CacheDaemon_cp_element_group_215: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_215"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= l2CacheDaemon_CP_3229_elements(220);
      gj_l2CacheDaemon_cp_element_group_215 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(215), clk => clk, reset => reset); --
    end block;
    -- CP-element group 216:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 216: predecessors 
    -- CP-element group 216: 	214 
    -- CP-element group 216: successors 
    -- CP-element group 216: marked-successors 
    -- CP-element group 216: 	92 
    -- CP-element group 216: 	214 
    -- CP-element group 216: 	88 
    -- CP-element group 216: 	120 
    -- CP-element group 216: 	116 
    -- CP-element group 216:  members (3) 
      -- CP-element group 216: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3743_sample_completed_
      -- CP-element group 216: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3743_Sample/$exit
      -- CP-element group 216: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3743_Sample/ack
      -- 
    ack_3907_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 216_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_back_line_address_3441_delayed_5_0_3741_inst_ack_0, ack => l2CacheDaemon_CP_3229_elements(216)); -- 
    -- CP-element group 217:  transition  input  bypass  pipeline-parent 
    -- CP-element group 217: predecessors 
    -- CP-element group 217: 	215 
    -- CP-element group 217: successors 
    -- CP-element group 217: 	218 
    -- CP-element group 217:  members (3) 
      -- CP-element group 217: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3743_update_completed_
      -- CP-element group 217: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3743_Update/$exit
      -- CP-element group 217: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/assign_stmt_3743_Update/ack
      -- 
    ack_3912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 217_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_write_back_line_address_3441_delayed_5_0_3741_inst_ack_1, ack => l2CacheDaemon_CP_3229_elements(217)); -- 
    -- CP-element group 218:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 218: predecessors 
    -- CP-element group 218: 	213 
    -- CP-element group 218: 	217 
    -- CP-element group 218: 	201 
    -- CP-element group 218: 	205 
    -- CP-element group 218: 	209 
    -- CP-element group 218: 	186 
    -- CP-element group 218: marked-predecessors 
    -- CP-element group 218: 	220 
    -- CP-element group 218: successors 
    -- CP-element group 218: 	220 
    -- CP-element group 218:  members (3) 
      -- CP-element group 218: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3750_sample_start_
      -- CP-element group 218: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3750_Sample/$entry
      -- CP-element group 218: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3750_Sample/crr
      -- 
    crr_3920_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3920_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(218), ack => call_stmt_3750_call_req_0); -- 
    l2CacheDaemon_cp_element_group_218: block -- 
      constant place_capacities: IntegerArray(0 to 6) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1);
      constant place_markings: IntegerArray(0 to 6)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
      constant place_delays: IntegerArray(0 to 6) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 1);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_218"; 
      signal preds: BooleanArray(1 to 7); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(213) & l2CacheDaemon_CP_3229_elements(217) & l2CacheDaemon_CP_3229_elements(201) & l2CacheDaemon_CP_3229_elements(205) & l2CacheDaemon_CP_3229_elements(209) & l2CacheDaemon_CP_3229_elements(186) & l2CacheDaemon_CP_3229_elements(220);
      gj_l2CacheDaemon_cp_element_group_218 : generic_join generic map(name => joinName, number_of_predecessors => 7, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(218), clk => clk, reset => reset); --
    end block;
    -- CP-element group 219:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 219: predecessors 
    -- CP-element group 219: marked-predecessors 
    -- CP-element group 219: 	221 
    -- CP-element group 219: successors 
    -- CP-element group 219: 	221 
    -- CP-element group 219:  members (3) 
      -- CP-element group 219: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3750_update_start_
      -- CP-element group 219: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3750_Update/$entry
      -- CP-element group 219: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3750_Update/ccr
      -- 
    ccr_3925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => l2CacheDaemon_CP_3229_elements(219), ack => call_stmt_3750_call_req_1); -- 
    l2CacheDaemon_cp_element_group_219: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_219"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= l2CacheDaemon_CP_3229_elements(221);
      gj_l2CacheDaemon_cp_element_group_219 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(219), clk => clk, reset => reset); --
    end block;
    -- CP-element group 220:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 220: predecessors 
    -- CP-element group 220: 	218 
    -- CP-element group 220: successors 
    -- CP-element group 220: marked-successors 
    -- CP-element group 220: 	215 
    -- CP-element group 220: 	218 
    -- CP-element group 220: 	203 
    -- CP-element group 220: 	207 
    -- CP-element group 220: 	211 
    -- CP-element group 220: 	184 
    -- CP-element group 220: 	199 
    -- CP-element group 220:  members (3) 
      -- CP-element group 220: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3750_sample_completed_
      -- CP-element group 220: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3750_Sample/$exit
      -- CP-element group 220: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3750_Sample/cra
      -- 
    cra_3921_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 220_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_3750_call_ack_0, ack => l2CacheDaemon_CP_3229_elements(220)); -- 
    -- CP-element group 221:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 221: predecessors 
    -- CP-element group 221: 	219 
    -- CP-element group 221: successors 
    -- CP-element group 221: 	223 
    -- CP-element group 221: marked-successors 
    -- CP-element group 221: 	219 
    -- CP-element group 221:  members (3) 
      -- CP-element group 221: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3750_update_completed_
      -- CP-element group 221: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3750_Update/$exit
      -- CP-element group 221: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/call_stmt_3750_Update/cca
      -- 
    cca_3926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 221_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_3750_call_ack_1, ack => l2CacheDaemon_CP_3229_elements(221)); -- 
    -- CP-element group 222:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 222: predecessors 
    -- CP-element group 222: 	11 
    -- CP-element group 222: successors 
    -- CP-element group 222: 	12 
    -- CP-element group 222:  members (1) 
      -- CP-element group 222: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group l2CacheDaemon_CP_3229_elements(222) is a control-delay.
    cp_element_222_delay: control_delay_element  generic map(name => " 222_delay", delay_value => 1)  port map(req => l2CacheDaemon_CP_3229_elements(11), ack => l2CacheDaemon_CP_3229_elements(222), clk => clk, reset =>reset);
    -- CP-element group 223:  join  transition  bypass  pipeline-parent 
    -- CP-element group 223: predecessors 
    -- CP-element group 223: 	14 
    -- CP-element group 223: 	79 
    -- CP-element group 223: 	82 
    -- CP-element group 223: 	221 
    -- CP-element group 223: 	197 
    -- CP-element group 223: successors 
    -- CP-element group 223: 	8 
    -- CP-element group 223:  members (1) 
      -- CP-element group 223: 	 branch_block_stmt_3335/do_while_stmt_3336/do_while_stmt_3336_loop_body/$exit
      -- 
    l2CacheDaemon_cp_element_group_223: block -- 
      constant place_capacities: IntegerArray(0 to 4) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15);
      constant place_markings: IntegerArray(0 to 4)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant place_delays: IntegerArray(0 to 4) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0);
      constant joinName: string(1 to 34) := "l2CacheDaemon_cp_element_group_223"; 
      signal preds: BooleanArray(1 to 5); -- 
    begin -- 
      preds <= l2CacheDaemon_CP_3229_elements(14) & l2CacheDaemon_CP_3229_elements(79) & l2CacheDaemon_CP_3229_elements(82) & l2CacheDaemon_CP_3229_elements(221) & l2CacheDaemon_CP_3229_elements(197);
      gj_l2CacheDaemon_cp_element_group_223 : generic_join generic map(name => joinName, number_of_predecessors => 5, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(223), clk => clk, reset => reset); --
    end block;
    -- CP-element group 224:  transition  input  bypass  pipeline-parent 
    -- CP-element group 224: predecessors 
    -- CP-element group 224: 	7 
    -- CP-element group 224: successors 
    -- CP-element group 224:  members (2) 
      -- CP-element group 224: 	 branch_block_stmt_3335/do_while_stmt_3336/loop_exit/$exit
      -- CP-element group 224: 	 branch_block_stmt_3335/do_while_stmt_3336/loop_exit/ack
      -- 
    ack_3931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 224_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_3336_branch_ack_0, ack => l2CacheDaemon_CP_3229_elements(224)); -- 
    -- CP-element group 225:  transition  input  bypass  pipeline-parent 
    -- CP-element group 225: predecessors 
    -- CP-element group 225: 	7 
    -- CP-element group 225: successors 
    -- CP-element group 225:  members (2) 
      -- CP-element group 225: 	 branch_block_stmt_3335/do_while_stmt_3336/loop_taken/$exit
      -- CP-element group 225: 	 branch_block_stmt_3335/do_while_stmt_3336/loop_taken/ack
      -- 
    ack_3935_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 225_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_3336_branch_ack_1, ack => l2CacheDaemon_CP_3229_elements(225)); -- 
    -- CP-element group 226:  transition  bypass  pipeline-parent 
    -- CP-element group 226: predecessors 
    -- CP-element group 226: 	5 
    -- CP-element group 226: successors 
    -- CP-element group 226: 	3 
    -- CP-element group 226:  members (1) 
      -- CP-element group 226: 	 branch_block_stmt_3335/do_while_stmt_3336/$exit
      -- 
    l2CacheDaemon_CP_3229_elements(226) <= l2CacheDaemon_CP_3229_elements(5);
    l2CacheDaemon_do_while_stmt_3336_terminator_3936: loop_terminator -- 
      generic map (name => " l2CacheDaemon_do_while_stmt_3336_terminator_3936", max_iterations_in_flight =>15) 
      port map(loop_body_exit => l2CacheDaemon_CP_3229_elements(8),loop_continue => l2CacheDaemon_CP_3229_elements(225),loop_terminate => l2CacheDaemon_CP_3229_elements(224),loop_back => l2CacheDaemon_CP_3229_elements(6),loop_exit => l2CacheDaemon_CP_3229_elements(5),clk => clk, reset => reset); -- 
    phi_stmt_3338_phi_seq_3320_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= l2CacheDaemon_CP_3229_elements(24);
      l2CacheDaemon_CP_3229_elements(27)<= src_sample_reqs(0);
      src_sample_acks(0)  <= l2CacheDaemon_CP_3229_elements(27);
      l2CacheDaemon_CP_3229_elements(28)<= src_update_reqs(0);
      src_update_acks(0)  <= l2CacheDaemon_CP_3229_elements(29);
      l2CacheDaemon_CP_3229_elements(25) <= phi_mux_reqs(0);
      triggers(1)  <= l2CacheDaemon_CP_3229_elements(22);
      l2CacheDaemon_CP_3229_elements(31)<= src_sample_reqs(1);
      src_sample_acks(1)  <= l2CacheDaemon_CP_3229_elements(35);
      l2CacheDaemon_CP_3229_elements(32)<= src_update_reqs(1);
      src_update_acks(1)  <= l2CacheDaemon_CP_3229_elements(36);
      l2CacheDaemon_CP_3229_elements(23) <= phi_mux_reqs(1);
      phi_stmt_3338_phi_seq_3320 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_3338_phi_seq_3320") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => l2CacheDaemon_CP_3229_elements(13), 
          phi_sample_ack => l2CacheDaemon_CP_3229_elements(20), 
          phi_update_req => l2CacheDaemon_CP_3229_elements(16), 
          phi_update_ack => l2CacheDaemon_CP_3229_elements(21), 
          phi_mux_ack => l2CacheDaemon_CP_3229_elements(26), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_3343_phi_seq_3364_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= l2CacheDaemon_CP_3229_elements(45);
      l2CacheDaemon_CP_3229_elements(48)<= src_sample_reqs(0);
      src_sample_acks(0)  <= l2CacheDaemon_CP_3229_elements(48);
      l2CacheDaemon_CP_3229_elements(49)<= src_update_reqs(0);
      src_update_acks(0)  <= l2CacheDaemon_CP_3229_elements(50);
      l2CacheDaemon_CP_3229_elements(46) <= phi_mux_reqs(0);
      triggers(1)  <= l2CacheDaemon_CP_3229_elements(43);
      l2CacheDaemon_CP_3229_elements(52)<= src_sample_reqs(1);
      src_sample_acks(1)  <= l2CacheDaemon_CP_3229_elements(56);
      l2CacheDaemon_CP_3229_elements(53)<= src_update_reqs(1);
      src_update_acks(1)  <= l2CacheDaemon_CP_3229_elements(57);
      l2CacheDaemon_CP_3229_elements(44) <= phi_mux_reqs(1);
      phi_stmt_3343_phi_seq_3364 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_3343_phi_seq_3364") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => l2CacheDaemon_CP_3229_elements(39), 
          phi_sample_ack => l2CacheDaemon_CP_3229_elements(40), 
          phi_update_req => l2CacheDaemon_CP_3229_elements(41), 
          phi_update_ack => l2CacheDaemon_CP_3229_elements(42), 
          phi_mux_ack => l2CacheDaemon_CP_3229_elements(47), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_3347_phi_seq_3408_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= l2CacheDaemon_CP_3229_elements(66);
      l2CacheDaemon_CP_3229_elements(69)<= src_sample_reqs(0);
      src_sample_acks(0)  <= l2CacheDaemon_CP_3229_elements(69);
      l2CacheDaemon_CP_3229_elements(70)<= src_update_reqs(0);
      src_update_acks(0)  <= l2CacheDaemon_CP_3229_elements(71);
      l2CacheDaemon_CP_3229_elements(67) <= phi_mux_reqs(0);
      triggers(1)  <= l2CacheDaemon_CP_3229_elements(64);
      l2CacheDaemon_CP_3229_elements(73)<= src_sample_reqs(1);
      src_sample_acks(1)  <= l2CacheDaemon_CP_3229_elements(75);
      l2CacheDaemon_CP_3229_elements(74)<= src_update_reqs(1);
      src_update_acks(1)  <= l2CacheDaemon_CP_3229_elements(76);
      l2CacheDaemon_CP_3229_elements(65) <= phi_mux_reqs(1);
      phi_stmt_3347_phi_seq_3408 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_3347_phi_seq_3408") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => l2CacheDaemon_CP_3229_elements(60), 
          phi_sample_ack => l2CacheDaemon_CP_3229_elements(61), 
          phi_update_req => l2CacheDaemon_CP_3229_elements(62), 
          phi_update_ack => l2CacheDaemon_CP_3229_elements(63), 
          phi_mux_ack => l2CacheDaemon_CP_3229_elements(68), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_3271_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= l2CacheDaemon_CP_3229_elements(9);
        preds(1)  <= l2CacheDaemon_CP_3229_elements(10);
        entry_tmerge_3271 : transition_merge -- 
          generic map(name => " entry_tmerge_3271")
          port map (preds => preds, symbol_out => l2CacheDaemon_CP_3229_elements(11));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal ADD_u8_u8_3444_wire : std_logic_vector(7 downto 0);
    signal AND_u1_u1_3316_3316_delayed_5_0_3540 : std_logic_vector(0 downto 0);
    signal AND_u1_u1_3325_3325_delayed_5_0_3552 : std_logic_vector(0 downto 0);
    signal AND_u1_u1_3441_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_3571_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_3577_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_3581_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_3583_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_3590_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_3598_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u1_u2_3478_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u9_3475_wire : std_logic_vector(8 downto 0);
    signal CONCAT_u21_u24_3482_wire : std_logic_vector(23 downto 0);
    signal CONCAT_u24_u34_3486_wire : std_logic_vector(33 downto 0);
    signal CONCAT_u9_u10_3485_wire : std_logic_vector(9 downto 0);
    signal CONCAT_u9_u11_3479_wire : std_logic_vector(10 downto 0);
    signal COUNTER_3347 : std_logic_vector(7 downto 0);
    signal MUX_3710_wire : std_logic_vector(63 downto 0);
    signal NEQ_u8_u1_3574_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_3402_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_3408_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_3410_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_3439_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_3467_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_3537_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_3544_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_3549_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_3556_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_3580_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_3588_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_3596_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_3600_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_3377_3377_delayed_5_0_3619 : std_logic_vector(0 downto 0);
    signal OR_u1_u1_3582_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_3623_wire : std_logic_vector(0 downto 0);
    signal RPIPE_NOBLOCK_L2_INVALIDATE_3346_wire : std_logic_vector(30 downto 0);
    signal RPIPE_NOBLOCK_L2_REQUEST_3342_wire : std_logic_vector(110 downto 0);
    signal access_data_mem_3394_delayed_4_0_3652 : std_logic_vector(0 downto 0);
    signal access_data_mem_3626 : std_logic_vector(0 downto 0);
    signal access_index_in_set_3511 : std_logic_vector(2 downto 0);
    signal access_set_id_3302_delayed_5_0_3522 : std_logic_vector(8 downto 0);
    signal access_set_id_3386_delayed_5_0_3636 : std_logic_vector(8 downto 0);
    signal access_set_id_3453 : std_logic_vector(8 downto 0);
    signal access_tag_3459 : std_logic_vector(20 downto 0);
    signal access_tags_command_3488 : std_logic_vector(44 downto 0);
    signal access_tags_resp_3499 : std_logic_vector(33 downto 0);
    signal allocate_on_miss_3470 : std_logic_vector(0 downto 0);
    signal byte_mask_3368 : std_logic_vector(7 downto 0);
    signal byte_mask_3400_delayed_9_0_3670 : std_logic_vector(7 downto 0);
    signal call_dwordId_expr_3431_wire : std_logic_vector(2 downto 0);
    signal call_lineAddress_expr_3423_wire : std_logic_vector(29 downto 0);
    signal call_paTag_expr_3435_wire : std_logic_vector(20 downto 0);
    signal call_setId_expr_3427_wire : std_logic_vector(8 downto 0);
    signal call_write_mem_3437_delayed_5_0_3731 : std_logic_vector(0 downto 0);
    signal call_write_mem_3728 : std_logic_vector(0 downto 0);
    signal data_read_dword_3391_delayed_5_0_3644 : std_logic_vector(0 downto 0);
    signal data_read_dword_3397_delayed_9_0_3661 : std_logic_vector(0 downto 0);
    signal data_read_dword_3593 : std_logic_vector(0 downto 0);
    signal data_write_dword_3396_delayed_9_0_3658 : std_logic_vector(0 downto 0);
    signal data_write_dword_3602 : std_logic_vector(0 downto 0);
    signal data_write_new_line_3398_delayed_4_0_3664 : std_logic_vector(0 downto 0);
    signal data_write_new_line_3558 : std_logic_vector(0 downto 0);
    signal dirty_word_mask_3440_delayed_5_0_3740 : std_logic_vector(7 downto 0);
    signal dirty_word_mask_3507 : std_logic_vector(7 downto 0);
    signal do_read_line_from_mem_3438_delayed_5_0_3734 : std_logic_vector(0 downto 0);
    signal do_read_line_from_mem_3546 : std_logic_vector(0 downto 0);
    signal do_tag_access_3276_delayed_4_0_3495 : std_logic_vector(0 downto 0);
    signal do_tag_access_3331_delayed_5_0_3561 : std_logic_vector(0 downto 0);
    signal do_tag_access_3464 : std_logic_vector(0 downto 0);
    signal do_write_replaced_line_to_mem_3399_delayed_4_0_3667 : std_logic_vector(0 downto 0);
    signal do_write_replaced_line_to_mem_3439_delayed_5_0_3737 : std_logic_vector(0 downto 0);
    signal do_write_replaced_line_to_mem_3585 : std_logic_vector(0 downto 0);
    signal get_req_3412 : std_logic_vector(0 downto 0);
    signal inv_pa_line_address_3367_delayed_5_0_3608 : std_logic_vector(29 downto 0);
    signal inv_pa_line_address_3392 : std_logic_vector(29 downto 0);
    signal inv_set_id_3420 : std_logic_vector(8 downto 0);
    signal inv_tag_3416 : std_logic_vector(20 downto 0);
    signal inv_valid_3337_delayed_5_0_3564 : std_logic_vector(0 downto 0);
    signal inv_valid_3366_delayed_5_0_3605 : std_logic_vector(0 downto 0);
    signal inv_valid_3388 : std_logic_vector(0 downto 0);
    signal invalidate_request_3343 : std_logic_vector(30 downto 0);
    signal is_hit_3503 : std_logic_vector(0 downto 0);
    signal konst_3340_wire_constant : std_logic_vector(110 downto 0);
    signal konst_3345_wire_constant : std_logic_vector(30 downto 0);
    signal konst_3443_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3573_wire_constant : std_logic_vector(7 downto 0);
    signal konst_3756_wire_constant : std_logic_vector(0 downto 0);
    signal l2_cache_request_3338 : std_logic_vector(110 downto 0);
    signal l2_resp_3712 : std_logic_vector(64 downto 0);
    signal line_id_3401_delayed_4_0_3673 : std_logic_vector(11 downto 0);
    signal line_id_3641 : std_logic_vector(11 downto 0);
    signal lock_3360 : std_logic_vector(0 downto 0);
    signal nCOUNTER_3447 : std_logic_vector(7 downto 0);
    signal nCOUNTER_3447_3351_buffered : std_logic_vector(7 downto 0);
    signal pa_3372 : std_logic_vector(35 downto 0);
    signal pa_dword_id_3402_delayed_9_0_3676 : std_logic_vector(2 downto 0);
    signal pa_dword_id_3432 : std_logic_vector(2 downto 0);
    signal pa_line_address_3381_delayed_5_0_3629 : std_logic_vector(29 downto 0);
    signal pa_line_address_3424 : std_logic_vector(29 downto 0);
    signal pa_mem_cache_line_3633 : std_logic_vector(511 downto 0);
    signal pa_set_id_3428 : std_logic_vector(8 downto 0);
    signal pa_tag_3436 : std_logic_vector(20 downto 0);
    signal read_data_line_3395_delayed_4_0_3655 : std_logic_vector(0 downto 0);
    signal read_data_line_3649 : std_logic_vector(0 downto 0);
    signal read_dword_from_data_3693 : std_logic_vector(63 downto 0);
    signal replace_line_is_valid_3515 : std_logic_vector(0 downto 0);
    signal replace_pa_line_address_3527 : std_logic_vector(29 downto 0);
    signal replace_pa_tag_3519 : std_logic_vector(20 downto 0);
    signal rwbar_3364 : std_logic_vector(0 downto 0);
    signal rwbar_3417_delayed_10_0_3702 : std_logic_vector(0 downto 0);
    signal send_response_3405 : std_logic_vector(0 downto 0);
    signal send_response_3424_delayed_10_0_3715 : std_logic_vector(0 downto 0);
    signal type_cast_3333_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_3350_wire_constant : std_logic_vector(7 downto 0);
    signal type_cast_3473_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_3705_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_3709_wire_constant : std_logic_vector(63 downto 0);
    signal valid_3340_delayed_5_0_3567 : std_logic_vector(0 downto 0);
    signal valid_3356 : std_logic_vector(0 downto 0);
    signal wdata_3376 : std_logic_vector(63 downto 0);
    signal wdata_3403_delayed_9_0_3679 : std_logic_vector(63 downto 0);
    signal write_back_line_address_3441_delayed_5_0_3743 : std_logic_vector(29 downto 0);
    signal write_back_line_address_3614 : std_logic_vector(29 downto 0);
    signal writeback_line_from_data_3693 : std_logic_vector(511 downto 0);
    -- 
  begin -- 
    konst_3340_wire_constant <= "000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000000";
    konst_3345_wire_constant <= "0000000000000000000000000000000";
    konst_3443_wire_constant <= "00000001";
    konst_3573_wire_constant <= "00000000";
    konst_3756_wire_constant <= "1";
    type_cast_3333_wire_constant <= "1";
    type_cast_3350_wire_constant <= "00000000";
    type_cast_3473_wire_constant <= "1";
    type_cast_3705_wire_constant <= "0";
    type_cast_3709_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_3338: Block -- phi operator 
      signal idata: std_logic_vector(221 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= konst_3340_wire_constant & RPIPE_NOBLOCK_L2_REQUEST_3342_wire;
      req <= phi_stmt_3338_req_0 & phi_stmt_3338_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3338",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 111) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3338_ack_0,
          idata => idata,
          odata => l2_cache_request_3338,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3338
    phi_stmt_3343: Block -- phi operator 
      signal idata: std_logic_vector(61 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= konst_3345_wire_constant & RPIPE_NOBLOCK_L2_INVALIDATE_3346_wire;
      req <= phi_stmt_3343_req_0 & phi_stmt_3343_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3343",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 31) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3343_ack_0,
          idata => idata,
          odata => invalidate_request_3343,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3343
    phi_stmt_3347: Block -- phi operator 
      signal idata: std_logic_vector(15 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3350_wire_constant & nCOUNTER_3447_3351_buffered;
      req <= phi_stmt_3347_req_0 & phi_stmt_3347_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3347",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 8) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3347_ack_0,
          idata => idata,
          odata => COUNTER_3347,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3347
    -- flow-through select operator MUX_3446_inst
    nCOUNTER_3447 <= ADD_u8_u8_3444_wire when (AND_u1_u1_3441_wire(0) /=  '0') else COUNTER_3347;
    -- flow-through select operator MUX_3452_inst
    access_set_id_3453 <= inv_set_id_3420 when (inv_valid_3388(0) /=  '0') else pa_set_id_3428;
    -- flow-through select operator MUX_3458_inst
    access_tag_3459 <= inv_tag_3416 when (inv_valid_3388(0) /=  '0') else pa_tag_3436;
    -- flow-through select operator MUX_3613_inst
    write_back_line_address_3614 <= inv_pa_line_address_3367_delayed_5_0_3608 when (inv_valid_3366_delayed_5_0_3605(0) /=  '0') else replace_pa_line_address_3527;
    -- flow-through select operator MUX_3710_inst
    MUX_3710_wire <= read_dword_from_data_3693 when (rwbar_3417_delayed_10_0_3702(0) /=  '0') else type_cast_3709_wire_constant;
    -- flow-through slice operator slice_3355_inst
    valid_3356 <= l2_cache_request_3338(110 downto 110);
    -- flow-through slice operator slice_3359_inst
    lock_3360 <= l2_cache_request_3338(109 downto 109);
    -- flow-through slice operator slice_3363_inst
    rwbar_3364 <= l2_cache_request_3338(108 downto 108);
    -- flow-through slice operator slice_3367_inst
    byte_mask_3368 <= l2_cache_request_3338(107 downto 100);
    -- flow-through slice operator slice_3371_inst
    pa_3372 <= l2_cache_request_3338(99 downto 64);
    -- flow-through slice operator slice_3375_inst
    wdata_3376 <= l2_cache_request_3338(63 downto 0);
    -- flow-through slice operator slice_3387_inst
    inv_valid_3388 <= invalidate_request_3343(30 downto 30);
    -- flow-through slice operator slice_3391_inst
    inv_pa_line_address_3392 <= invalidate_request_3343(29 downto 0);
    -- flow-through slice operator slice_3415_inst
    inv_tag_3416 <= inv_pa_line_address_3392(29 downto 9);
    -- flow-through slice operator slice_3419_inst
    inv_set_id_3420 <= inv_pa_line_address_3392(8 downto 0);
    -- flow-through slice operator slice_3502_inst
    is_hit_3503 <= access_tags_resp_3499(33 downto 33);
    -- flow-through slice operator slice_3506_inst
    dirty_word_mask_3507 <= access_tags_resp_3499(32 downto 25);
    -- flow-through slice operator slice_3510_inst
    access_index_in_set_3511 <= access_tags_resp_3499(24 downto 22);
    -- flow-through slice operator slice_3514_inst
    replace_line_is_valid_3515 <= access_tags_resp_3499(21 downto 21);
    -- flow-through slice operator slice_3518_inst
    replace_pa_tag_3519 <= access_tags_resp_3499(20 downto 0);
    W_access_data_mem_3394_delayed_4_0_3650_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_access_data_mem_3394_delayed_4_0_3650_inst_req_0;
      W_access_data_mem_3394_delayed_4_0_3650_inst_ack_0<= wack(0);
      rreq(0) <= W_access_data_mem_3394_delayed_4_0_3650_inst_req_1;
      W_access_data_mem_3394_delayed_4_0_3650_inst_ack_1<= rack(0);
      W_access_data_mem_3394_delayed_4_0_3650_inst : InterlockBuffer generic map ( -- 
        name => "W_access_data_mem_3394_delayed_4_0_3650_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => access_data_mem_3626,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => access_data_mem_3394_delayed_4_0_3652,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_access_set_id_3302_delayed_5_0_3520_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_access_set_id_3302_delayed_5_0_3520_inst_req_0;
      W_access_set_id_3302_delayed_5_0_3520_inst_ack_0<= wack(0);
      rreq(0) <= W_access_set_id_3302_delayed_5_0_3520_inst_req_1;
      W_access_set_id_3302_delayed_5_0_3520_inst_ack_1<= rack(0);
      W_access_set_id_3302_delayed_5_0_3520_inst : InterlockBuffer generic map ( -- 
        name => "W_access_set_id_3302_delayed_5_0_3520_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 9,
        out_data_width => 9,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => access_set_id_3453,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => access_set_id_3302_delayed_5_0_3522,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_access_set_id_3386_delayed_5_0_3634_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_access_set_id_3386_delayed_5_0_3634_inst_req_0;
      W_access_set_id_3386_delayed_5_0_3634_inst_ack_0<= wack(0);
      rreq(0) <= W_access_set_id_3386_delayed_5_0_3634_inst_req_1;
      W_access_set_id_3386_delayed_5_0_3634_inst_ack_1<= rack(0);
      W_access_set_id_3386_delayed_5_0_3634_inst : InterlockBuffer generic map ( -- 
        name => "W_access_set_id_3386_delayed_5_0_3634_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 9,
        out_data_width => 9,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => access_set_id_3453,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => access_set_id_3386_delayed_5_0_3636,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_byte_mask_3400_delayed_9_0_3668_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_byte_mask_3400_delayed_9_0_3668_inst_req_0;
      W_byte_mask_3400_delayed_9_0_3668_inst_ack_0<= wack(0);
      rreq(0) <= W_byte_mask_3400_delayed_9_0_3668_inst_req_1;
      W_byte_mask_3400_delayed_9_0_3668_inst_ack_1<= rack(0);
      W_byte_mask_3400_delayed_9_0_3668_inst : InterlockBuffer generic map ( -- 
        name => "W_byte_mask_3400_delayed_9_0_3668_inst",
        buffer_size => 9,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => byte_mask_3368,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => byte_mask_3400_delayed_9_0_3670,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_call_write_mem_3437_delayed_5_0_3729_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_call_write_mem_3437_delayed_5_0_3729_inst_req_0;
      W_call_write_mem_3437_delayed_5_0_3729_inst_ack_0<= wack(0);
      rreq(0) <= W_call_write_mem_3437_delayed_5_0_3729_inst_req_1;
      W_call_write_mem_3437_delayed_5_0_3729_inst_ack_1<= rack(0);
      W_call_write_mem_3437_delayed_5_0_3729_inst : InterlockBuffer generic map ( -- 
        name => "W_call_write_mem_3437_delayed_5_0_3729_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => call_write_mem_3728,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => call_write_mem_3437_delayed_5_0_3731,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_data_read_dword_3391_delayed_5_0_3642_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_data_read_dword_3391_delayed_5_0_3642_inst_req_0;
      W_data_read_dword_3391_delayed_5_0_3642_inst_ack_0<= wack(0);
      rreq(0) <= W_data_read_dword_3391_delayed_5_0_3642_inst_req_1;
      W_data_read_dword_3391_delayed_5_0_3642_inst_ack_1<= rack(0);
      W_data_read_dword_3391_delayed_5_0_3642_inst : InterlockBuffer generic map ( -- 
        name => "W_data_read_dword_3391_delayed_5_0_3642_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => data_read_dword_3593,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => data_read_dword_3391_delayed_5_0_3644,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_data_read_dword_3397_delayed_9_0_3659_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_data_read_dword_3397_delayed_9_0_3659_inst_req_0;
      W_data_read_dword_3397_delayed_9_0_3659_inst_ack_0<= wack(0);
      rreq(0) <= W_data_read_dword_3397_delayed_9_0_3659_inst_req_1;
      W_data_read_dword_3397_delayed_9_0_3659_inst_ack_1<= rack(0);
      W_data_read_dword_3397_delayed_9_0_3659_inst : InterlockBuffer generic map ( -- 
        name => "W_data_read_dword_3397_delayed_9_0_3659_inst",
        buffer_size => 9,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => data_read_dword_3593,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => data_read_dword_3397_delayed_9_0_3661,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_data_write_dword_3396_delayed_9_0_3656_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_data_write_dword_3396_delayed_9_0_3656_inst_req_0;
      W_data_write_dword_3396_delayed_9_0_3656_inst_ack_0<= wack(0);
      rreq(0) <= W_data_write_dword_3396_delayed_9_0_3656_inst_req_1;
      W_data_write_dword_3396_delayed_9_0_3656_inst_ack_1<= rack(0);
      W_data_write_dword_3396_delayed_9_0_3656_inst : InterlockBuffer generic map ( -- 
        name => "W_data_write_dword_3396_delayed_9_0_3656_inst",
        buffer_size => 9,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => data_write_dword_3602,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => data_write_dword_3396_delayed_9_0_3658,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_data_write_new_line_3398_delayed_4_0_3662_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_data_write_new_line_3398_delayed_4_0_3662_inst_req_0;
      W_data_write_new_line_3398_delayed_4_0_3662_inst_ack_0<= wack(0);
      rreq(0) <= W_data_write_new_line_3398_delayed_4_0_3662_inst_req_1;
      W_data_write_new_line_3398_delayed_4_0_3662_inst_ack_1<= rack(0);
      W_data_write_new_line_3398_delayed_4_0_3662_inst : InterlockBuffer generic map ( -- 
        name => "W_data_write_new_line_3398_delayed_4_0_3662_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => data_write_new_line_3558,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => data_write_new_line_3398_delayed_4_0_3664,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_dirty_word_mask_3440_delayed_5_0_3738_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_dirty_word_mask_3440_delayed_5_0_3738_inst_req_0;
      W_dirty_word_mask_3440_delayed_5_0_3738_inst_ack_0<= wack(0);
      rreq(0) <= W_dirty_word_mask_3440_delayed_5_0_3738_inst_req_1;
      W_dirty_word_mask_3440_delayed_5_0_3738_inst_ack_1<= rack(0);
      W_dirty_word_mask_3440_delayed_5_0_3738_inst : InterlockBuffer generic map ( -- 
        name => "W_dirty_word_mask_3440_delayed_5_0_3738_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => dirty_word_mask_3507,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => dirty_word_mask_3440_delayed_5_0_3740,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_do_read_line_from_mem_3438_delayed_5_0_3732_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_do_read_line_from_mem_3438_delayed_5_0_3732_inst_req_0;
      W_do_read_line_from_mem_3438_delayed_5_0_3732_inst_ack_0<= wack(0);
      rreq(0) <= W_do_read_line_from_mem_3438_delayed_5_0_3732_inst_req_1;
      W_do_read_line_from_mem_3438_delayed_5_0_3732_inst_ack_1<= rack(0);
      W_do_read_line_from_mem_3438_delayed_5_0_3732_inst : InterlockBuffer generic map ( -- 
        name => "W_do_read_line_from_mem_3438_delayed_5_0_3732_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => do_read_line_from_mem_3546,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => do_read_line_from_mem_3438_delayed_5_0_3734,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_do_tag_access_3276_delayed_4_0_3493_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_do_tag_access_3276_delayed_4_0_3493_inst_req_0;
      W_do_tag_access_3276_delayed_4_0_3493_inst_ack_0<= wack(0);
      rreq(0) <= W_do_tag_access_3276_delayed_4_0_3493_inst_req_1;
      W_do_tag_access_3276_delayed_4_0_3493_inst_ack_1<= rack(0);
      W_do_tag_access_3276_delayed_4_0_3493_inst : InterlockBuffer generic map ( -- 
        name => "W_do_tag_access_3276_delayed_4_0_3493_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => do_tag_access_3464,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => do_tag_access_3276_delayed_4_0_3495,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_do_tag_access_3331_delayed_5_0_3559_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_do_tag_access_3331_delayed_5_0_3559_inst_req_0;
      W_do_tag_access_3331_delayed_5_0_3559_inst_ack_0<= wack(0);
      rreq(0) <= W_do_tag_access_3331_delayed_5_0_3559_inst_req_1;
      W_do_tag_access_3331_delayed_5_0_3559_inst_ack_1<= rack(0);
      W_do_tag_access_3331_delayed_5_0_3559_inst : InterlockBuffer generic map ( -- 
        name => "W_do_tag_access_3331_delayed_5_0_3559_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => do_tag_access_3464,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => do_tag_access_3331_delayed_5_0_3561,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_do_write_replaced_line_to_mem_3399_delayed_4_0_3665_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_do_write_replaced_line_to_mem_3399_delayed_4_0_3665_inst_req_0;
      W_do_write_replaced_line_to_mem_3399_delayed_4_0_3665_inst_ack_0<= wack(0);
      rreq(0) <= W_do_write_replaced_line_to_mem_3399_delayed_4_0_3665_inst_req_1;
      W_do_write_replaced_line_to_mem_3399_delayed_4_0_3665_inst_ack_1<= rack(0);
      W_do_write_replaced_line_to_mem_3399_delayed_4_0_3665_inst : InterlockBuffer generic map ( -- 
        name => "W_do_write_replaced_line_to_mem_3399_delayed_4_0_3665_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => do_write_replaced_line_to_mem_3585,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => do_write_replaced_line_to_mem_3399_delayed_4_0_3667,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_do_write_replaced_line_to_mem_3439_delayed_5_0_3735_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_do_write_replaced_line_to_mem_3439_delayed_5_0_3735_inst_req_0;
      W_do_write_replaced_line_to_mem_3439_delayed_5_0_3735_inst_ack_0<= wack(0);
      rreq(0) <= W_do_write_replaced_line_to_mem_3439_delayed_5_0_3735_inst_req_1;
      W_do_write_replaced_line_to_mem_3439_delayed_5_0_3735_inst_ack_1<= rack(0);
      W_do_write_replaced_line_to_mem_3439_delayed_5_0_3735_inst : InterlockBuffer generic map ( -- 
        name => "W_do_write_replaced_line_to_mem_3439_delayed_5_0_3735_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => do_write_replaced_line_to_mem_3585,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => do_write_replaced_line_to_mem_3439_delayed_5_0_3737,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_inv_pa_line_address_3367_delayed_5_0_3606_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_inv_pa_line_address_3367_delayed_5_0_3606_inst_req_0;
      W_inv_pa_line_address_3367_delayed_5_0_3606_inst_ack_0<= wack(0);
      rreq(0) <= W_inv_pa_line_address_3367_delayed_5_0_3606_inst_req_1;
      W_inv_pa_line_address_3367_delayed_5_0_3606_inst_ack_1<= rack(0);
      W_inv_pa_line_address_3367_delayed_5_0_3606_inst : InterlockBuffer generic map ( -- 
        name => "W_inv_pa_line_address_3367_delayed_5_0_3606_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 30,
        out_data_width => 30,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inv_pa_line_address_3392,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inv_pa_line_address_3367_delayed_5_0_3608,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_inv_valid_3337_delayed_5_0_3562_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_inv_valid_3337_delayed_5_0_3562_inst_req_0;
      W_inv_valid_3337_delayed_5_0_3562_inst_ack_0<= wack(0);
      rreq(0) <= W_inv_valid_3337_delayed_5_0_3562_inst_req_1;
      W_inv_valid_3337_delayed_5_0_3562_inst_ack_1<= rack(0);
      W_inv_valid_3337_delayed_5_0_3562_inst : InterlockBuffer generic map ( -- 
        name => "W_inv_valid_3337_delayed_5_0_3562_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inv_valid_3388,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inv_valid_3337_delayed_5_0_3564,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_inv_valid_3366_delayed_5_0_3603_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_inv_valid_3366_delayed_5_0_3603_inst_req_0;
      W_inv_valid_3366_delayed_5_0_3603_inst_ack_0<= wack(0);
      rreq(0) <= W_inv_valid_3366_delayed_5_0_3603_inst_req_1;
      W_inv_valid_3366_delayed_5_0_3603_inst_ack_1<= rack(0);
      W_inv_valid_3366_delayed_5_0_3603_inst : InterlockBuffer generic map ( -- 
        name => "W_inv_valid_3366_delayed_5_0_3603_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => inv_valid_3388,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => inv_valid_3366_delayed_5_0_3605,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_line_id_3401_delayed_4_0_3671_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_line_id_3401_delayed_4_0_3671_inst_req_0;
      W_line_id_3401_delayed_4_0_3671_inst_ack_0<= wack(0);
      rreq(0) <= W_line_id_3401_delayed_4_0_3671_inst_req_1;
      W_line_id_3401_delayed_4_0_3671_inst_ack_1<= rack(0);
      W_line_id_3401_delayed_4_0_3671_inst : InterlockBuffer generic map ( -- 
        name => "W_line_id_3401_delayed_4_0_3671_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 12,
        out_data_width => 12,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => line_id_3641,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => line_id_3401_delayed_4_0_3673,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_pa_dword_id_3402_delayed_9_0_3674_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_pa_dword_id_3402_delayed_9_0_3674_inst_req_0;
      W_pa_dword_id_3402_delayed_9_0_3674_inst_ack_0<= wack(0);
      rreq(0) <= W_pa_dword_id_3402_delayed_9_0_3674_inst_req_1;
      W_pa_dword_id_3402_delayed_9_0_3674_inst_ack_1<= rack(0);
      W_pa_dword_id_3402_delayed_9_0_3674_inst : InterlockBuffer generic map ( -- 
        name => "W_pa_dword_id_3402_delayed_9_0_3674_inst",
        buffer_size => 9,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 3,
        out_data_width => 3,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => pa_dword_id_3432,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pa_dword_id_3402_delayed_9_0_3676,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_pa_dword_id_3429_inst
    process(call_dwordId_expr_3431_wire) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 2 downto 0) := call_dwordId_expr_3431_wire(2 downto 0);
      pa_dword_id_3432 <= tmp_var; -- 
    end process;
    W_pa_line_address_3381_delayed_5_0_3627_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_pa_line_address_3381_delayed_5_0_3627_inst_req_0;
      W_pa_line_address_3381_delayed_5_0_3627_inst_ack_0<= wack(0);
      rreq(0) <= W_pa_line_address_3381_delayed_5_0_3627_inst_req_1;
      W_pa_line_address_3381_delayed_5_0_3627_inst_ack_1<= rack(0);
      W_pa_line_address_3381_delayed_5_0_3627_inst : InterlockBuffer generic map ( -- 
        name => "W_pa_line_address_3381_delayed_5_0_3627_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 30,
        out_data_width => 30,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => pa_line_address_3424,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => pa_line_address_3381_delayed_5_0_3629,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    -- interlock W_pa_line_address_3421_inst
    process(call_lineAddress_expr_3423_wire) -- 
      variable tmp_var : std_logic_vector(29 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 29 downto 0) := call_lineAddress_expr_3423_wire(29 downto 0);
      pa_line_address_3424 <= tmp_var; -- 
    end process;
    -- interlock W_pa_set_id_3425_inst
    process(call_setId_expr_3427_wire) -- 
      variable tmp_var : std_logic_vector(8 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 8 downto 0) := call_setId_expr_3427_wire(8 downto 0);
      pa_set_id_3428 <= tmp_var; -- 
    end process;
    -- interlock W_pa_tag_3433_inst
    process(call_paTag_expr_3435_wire) -- 
      variable tmp_var : std_logic_vector(20 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 20 downto 0) := call_paTag_expr_3435_wire(20 downto 0);
      pa_tag_3436 <= tmp_var; -- 
    end process;
    W_read_data_line_3395_delayed_4_0_3653_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_read_data_line_3395_delayed_4_0_3653_inst_req_0;
      W_read_data_line_3395_delayed_4_0_3653_inst_ack_0<= wack(0);
      rreq(0) <= W_read_data_line_3395_delayed_4_0_3653_inst_req_1;
      W_read_data_line_3395_delayed_4_0_3653_inst_ack_1<= rack(0);
      W_read_data_line_3395_delayed_4_0_3653_inst : InterlockBuffer generic map ( -- 
        name => "W_read_data_line_3395_delayed_4_0_3653_inst",
        buffer_size => 4,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => read_data_line_3649,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => read_data_line_3395_delayed_4_0_3655,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_rwbar_3417_delayed_10_0_3700_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_rwbar_3417_delayed_10_0_3700_inst_req_0;
      W_rwbar_3417_delayed_10_0_3700_inst_ack_0<= wack(0);
      rreq(0) <= W_rwbar_3417_delayed_10_0_3700_inst_req_1;
      W_rwbar_3417_delayed_10_0_3700_inst_ack_1<= rack(0);
      W_rwbar_3417_delayed_10_0_3700_inst : InterlockBuffer generic map ( -- 
        name => "W_rwbar_3417_delayed_10_0_3700_inst",
        buffer_size => 10,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rwbar_3364,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => rwbar_3417_delayed_10_0_3702,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_send_response_3424_delayed_10_0_3713_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_send_response_3424_delayed_10_0_3713_inst_req_0;
      W_send_response_3424_delayed_10_0_3713_inst_ack_0<= wack(0);
      rreq(0) <= W_send_response_3424_delayed_10_0_3713_inst_req_1;
      W_send_response_3424_delayed_10_0_3713_inst_ack_1<= rack(0);
      W_send_response_3424_delayed_10_0_3713_inst : InterlockBuffer generic map ( -- 
        name => "W_send_response_3424_delayed_10_0_3713_inst",
        buffer_size => 10,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => send_response_3405,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => send_response_3424_delayed_10_0_3715,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_valid_3340_delayed_5_0_3565_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_valid_3340_delayed_5_0_3565_inst_req_0;
      W_valid_3340_delayed_5_0_3565_inst_ack_0<= wack(0);
      rreq(0) <= W_valid_3340_delayed_5_0_3565_inst_req_1;
      W_valid_3340_delayed_5_0_3565_inst_ack_1<= rack(0);
      W_valid_3340_delayed_5_0_3565_inst : InterlockBuffer generic map ( -- 
        name => "W_valid_3340_delayed_5_0_3565_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => valid_3356,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => valid_3340_delayed_5_0_3567,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_wdata_3403_delayed_9_0_3677_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_wdata_3403_delayed_9_0_3677_inst_req_0;
      W_wdata_3403_delayed_9_0_3677_inst_ack_0<= wack(0);
      rreq(0) <= W_wdata_3403_delayed_9_0_3677_inst_req_1;
      W_wdata_3403_delayed_9_0_3677_inst_ack_1<= rack(0);
      W_wdata_3403_delayed_9_0_3677_inst : InterlockBuffer generic map ( -- 
        name => "W_wdata_3403_delayed_9_0_3677_inst",
        buffer_size => 9,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => wdata_3376,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => wdata_3403_delayed_9_0_3679,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_write_back_line_address_3441_delayed_5_0_3741_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_write_back_line_address_3441_delayed_5_0_3741_inst_req_0;
      W_write_back_line_address_3441_delayed_5_0_3741_inst_ack_0<= wack(0);
      rreq(0) <= W_write_back_line_address_3441_delayed_5_0_3741_inst_req_1;
      W_write_back_line_address_3441_delayed_5_0_3741_inst_ack_1<= rack(0);
      W_write_back_line_address_3441_delayed_5_0_3741_inst : InterlockBuffer generic map ( -- 
        name => "W_write_back_line_address_3441_delayed_5_0_3741_inst",
        buffer_size => 5,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 30,
        out_data_width => 30,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => write_back_line_address_3614,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => write_back_line_address_3441_delayed_5_0_3743,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    nCOUNTER_3447_3351_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= nCOUNTER_3447_3351_buf_req_0;
      nCOUNTER_3447_3351_buf_ack_0<= wack(0);
      rreq(0) <= nCOUNTER_3447_3351_buf_req_1;
      nCOUNTER_3447_3351_buf_ack_1<= rack(0);
      nCOUNTER_3447_3351_buf : InterlockBuffer generic map ( -- 
        name => "nCOUNTER_3447_3351_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 8,
        out_data_width => 8,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => nCOUNTER_3447,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => nCOUNTER_3447_3351_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_3336_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= konst_3756_wire_constant;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_3336_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_3336_branch_req_0,
          ack0 => do_while_stmt_3336_branch_ack_0,
          ack1 => do_while_stmt_3336_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u8_u8_3444_inst
    process(COUNTER_3347) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntAdd_proc(COUNTER_3347, konst_3443_wire_constant, tmp_var);
      ADD_u8_u8_3444_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_3404_inst
    process(NOT_u1_u1_3402_wire, valid_3356) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_3402_wire, valid_3356, tmp_var);
      send_response_3405 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_3441_inst
    process(NOT_u1_u1_3439_wire, valid_3356) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_3439_wire, valid_3356, tmp_var);
      AND_u1_u1_3441_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_3469_inst
    process(NOT_u1_u1_3467_wire, valid_3356) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_3467_wire, valid_3356, tmp_var);
      allocate_on_miss_3470 <= tmp_var; --
    end process;
    -- shared split operator group (4) : AND_u1_u1_3539_inst 
    ApIntAnd_group_4: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 5);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= NOT_u1_u1_3537_wire & valid_3356;
      AND_u1_u1_3316_3316_delayed_5_0_3540 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u1_u1_3539_inst_req_0;
      AND_u1_u1_3539_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u1_u1_3539_inst_req_1;
      AND_u1_u1_3539_inst_ack_1 <= ackR_unguarded(0);
      ApIntAnd_group_4_gI: SplitGuardInterface generic map(name => "ApIntAnd_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_4",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 1, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 5,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 4
    -- binary operator AND_u1_u1_3545_inst
    process(AND_u1_u1_3316_3316_delayed_5_0_3540, NOT_u1_u1_3544_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_3316_3316_delayed_5_0_3540, NOT_u1_u1_3544_wire, tmp_var);
      do_read_line_from_mem_3546 <= tmp_var; --
    end process;
    -- shared split operator group (6) : AND_u1_u1_3551_inst 
    ApIntAnd_group_6: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 5);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= NOT_u1_u1_3549_wire & valid_3356;
      AND_u1_u1_3325_3325_delayed_5_0_3552 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= AND_u1_u1_3551_inst_req_0;
      AND_u1_u1_3551_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= AND_u1_u1_3551_inst_req_1;
      AND_u1_u1_3551_inst_ack_1 <= ackR_unguarded(0);
      ApIntAnd_group_6_gI: SplitGuardInterface generic map(name => "ApIntAnd_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntAnd",
          name => "ApIntAnd_group_6",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 1, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 5,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 6
    -- binary operator AND_u1_u1_3557_inst
    process(AND_u1_u1_3325_3325_delayed_5_0_3552, NOT_u1_u1_3556_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_3325_3325_delayed_5_0_3552, NOT_u1_u1_3556_wire, tmp_var);
      data_write_new_line_3558 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_3571_inst
    process(do_tag_access_3331_delayed_5_0_3561, replace_line_is_valid_3515) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(do_tag_access_3331_delayed_5_0_3561, replace_line_is_valid_3515, tmp_var);
      AND_u1_u1_3571_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_3577_inst
    process(inv_valid_3337_delayed_5_0_3564, is_hit_3503) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(inv_valid_3337_delayed_5_0_3564, is_hit_3503, tmp_var);
      AND_u1_u1_3577_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_3581_inst
    process(valid_3340_delayed_5_0_3567, NOT_u1_u1_3580_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(valid_3340_delayed_5_0_3567, NOT_u1_u1_3580_wire, tmp_var);
      AND_u1_u1_3581_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_3583_inst
    process(NEQ_u8_u1_3574_wire, OR_u1_u1_3582_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NEQ_u8_u1_3574_wire, OR_u1_u1_3582_wire, tmp_var);
      AND_u1_u1_3583_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_3584_inst
    process(AND_u1_u1_3571_wire, AND_u1_u1_3583_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_3571_wire, AND_u1_u1_3583_wire, tmp_var);
      do_write_replaced_line_to_mem_3585 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_3590_inst
    process(NOT_u1_u1_3588_wire, valid_3356) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_3588_wire, valid_3356, tmp_var);
      AND_u1_u1_3590_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_3592_inst
    process(AND_u1_u1_3590_wire, rwbar_3364) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_3590_wire, rwbar_3364, tmp_var);
      data_read_dword_3593 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_3598_inst
    process(NOT_u1_u1_3596_wire, valid_3356) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_3596_wire, valid_3356, tmp_var);
      AND_u1_u1_3598_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_3601_inst
    process(AND_u1_u1_3598_wire, NOT_u1_u1_3600_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(AND_u1_u1_3598_wire, NOT_u1_u1_3600_wire, tmp_var);
      data_write_dword_3602 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u11_u45_3487_inst
    process(CONCAT_u9_u11_3479_wire, CONCAT_u24_u34_3486_wire) -- 
      variable tmp_var : std_logic_vector(44 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u9_u11_3479_wire, CONCAT_u24_u34_3486_wire, tmp_var);
      access_tags_command_3488 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_3478_inst
    process(inv_valid_3388, rwbar_3364) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(inv_valid_3388, rwbar_3364, tmp_var);
      CONCAT_u1_u2_3478_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u65_3711_inst
    process(type_cast_3705_wire_constant, MUX_3710_wire) -- 
      variable tmp_var : std_logic_vector(64 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_3705_wire_constant, MUX_3710_wire, tmp_var);
      l2_resp_3712 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u9_3475_inst
    process(type_cast_3473_wire_constant, COUNTER_3347) -- 
      variable tmp_var : std_logic_vector(8 downto 0); -- 
    begin -- 
      ApConcat_proc(type_cast_3473_wire_constant, COUNTER_3347, tmp_var);
      CONCAT_u1_u9_3475_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u21_u24_3482_inst
    process(access_tag_3459, pa_dword_id_3432) -- 
      variable tmp_var : std_logic_vector(23 downto 0); -- 
    begin -- 
      ApConcat_proc(access_tag_3459, pa_dword_id_3432, tmp_var);
      CONCAT_u21_u24_3482_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u21_u30_3526_inst
    process(replace_pa_tag_3519, access_set_id_3302_delayed_5_0_3522) -- 
      variable tmp_var : std_logic_vector(29 downto 0); -- 
    begin -- 
      ApConcat_proc(replace_pa_tag_3519, access_set_id_3302_delayed_5_0_3522, tmp_var);
      replace_pa_line_address_3527 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u24_u34_3486_inst
    process(CONCAT_u21_u24_3482_wire, CONCAT_u9_u10_3485_wire) -- 
      variable tmp_var : std_logic_vector(33 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u21_u24_3482_wire, CONCAT_u9_u10_3485_wire, tmp_var);
      CONCAT_u24_u34_3486_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u3_u12_3640_inst
    process(access_index_in_set_3511, access_set_id_3386_delayed_5_0_3636) -- 
      variable tmp_var : std_logic_vector(11 downto 0); -- 
    begin -- 
      ApConcat_proc(access_index_in_set_3511, access_set_id_3386_delayed_5_0_3636, tmp_var);
      line_id_3641 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u9_u10_3485_inst
    process(access_set_id_3453, allocate_on_miss_3470) -- 
      variable tmp_var : std_logic_vector(9 downto 0); -- 
    begin -- 
      ApConcat_proc(access_set_id_3453, allocate_on_miss_3470, tmp_var);
      CONCAT_u9_u10_3485_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u9_u11_3479_inst
    process(CONCAT_u1_u9_3475_wire, CONCAT_u1_u2_3478_wire) -- 
      variable tmp_var : std_logic_vector(10 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u9_3475_wire, CONCAT_u1_u2_3478_wire, tmp_var);
      CONCAT_u9_u11_3479_wire <= tmp_var; --
    end process;
    -- binary operator NEQ_u8_u1_3574_inst
    process(dirty_word_mask_3507) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntNe_proc(dirty_word_mask_3507, konst_3573_wire_constant, tmp_var);
      NEQ_u8_u1_3574_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_3402_inst
    process(inv_valid_3388) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", inv_valid_3388, tmp_var);
      NOT_u1_u1_3402_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_3408_inst
    process(inv_valid_3388) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", inv_valid_3388, tmp_var);
      NOT_u1_u1_3408_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_3410_inst
    process(valid_3356) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", valid_3356, tmp_var);
      NOT_u1_u1_3410_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_3439_inst
    process(inv_valid_3388) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", inv_valid_3388, tmp_var);
      NOT_u1_u1_3439_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_3467_inst
    process(inv_valid_3388) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", inv_valid_3388, tmp_var);
      NOT_u1_u1_3467_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_3537_inst
    process(inv_valid_3388) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", inv_valid_3388, tmp_var);
      NOT_u1_u1_3537_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_3544_inst
    process(is_hit_3503) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", is_hit_3503, tmp_var);
      NOT_u1_u1_3544_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_3549_inst
    process(inv_valid_3388) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", inv_valid_3388, tmp_var);
      NOT_u1_u1_3549_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_3556_inst
    process(is_hit_3503) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", is_hit_3503, tmp_var);
      NOT_u1_u1_3556_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_3580_inst
    process(is_hit_3503) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", is_hit_3503, tmp_var);
      NOT_u1_u1_3580_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_3588_inst
    process(inv_valid_3388) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", inv_valid_3388, tmp_var);
      NOT_u1_u1_3588_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_3596_inst
    process(inv_valid_3388) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", inv_valid_3388, tmp_var);
      NOT_u1_u1_3596_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_3600_inst
    process(rwbar_3364) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", rwbar_3364, tmp_var);
      NOT_u1_u1_3600_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_3411_inst
    process(NOT_u1_u1_3408_wire, NOT_u1_u1_3410_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(NOT_u1_u1_3408_wire, NOT_u1_u1_3410_wire, tmp_var);
      get_req_3412 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_3463_inst
    process(inv_valid_3388, valid_3356) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(inv_valid_3388, valid_3356, tmp_var);
      do_tag_access_3464 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_3582_inst
    process(AND_u1_u1_3577_wire, AND_u1_u1_3581_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(AND_u1_u1_3577_wire, AND_u1_u1_3581_wire, tmp_var);
      OR_u1_u1_3582_wire <= tmp_var; --
    end process;
    -- shared split operator group (44) : OR_u1_u1_3618_inst 
    ApIntOr_group_44: Block -- 
      signal data_in: std_logic_vector(1 downto 0);
      signal data_out: std_logic_vector(0 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 5);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= data_read_dword_3593 & data_write_dword_3602;
      OR_u1_u1_3377_3377_delayed_5_0_3619 <= data_out(0 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= OR_u1_u1_3618_inst_req_0;
      OR_u1_u1_3618_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= OR_u1_u1_3618_inst_req_1;
      OR_u1_u1_3618_inst_ack_1 <= ackR_unguarded(0);
      ApIntOr_group_44_gI: SplitGuardInterface generic map(name => "ApIntOr_group_44_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApIntOr",
          name => "ApIntOr_group_44",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 1,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 1, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 1,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 5,
          flow_through => false,
          full_rate  => true,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 44
    -- binary operator OR_u1_u1_3623_inst
    process(do_write_replaced_line_to_mem_3585, data_write_new_line_3558) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(do_write_replaced_line_to_mem_3585, data_write_new_line_3558, tmp_var);
      OR_u1_u1_3623_wire <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_3625_inst
    process(OR_u1_u1_3623_wire, OR_u1_u1_3377_3377_delayed_5_0_3619) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(OR_u1_u1_3623_wire, OR_u1_u1_3377_3377_delayed_5_0_3619, tmp_var);
      access_data_mem_3626 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_3648_inst
    process(do_write_replaced_line_to_mem_3585, data_read_dword_3391_delayed_5_0_3644) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(do_write_replaced_line_to_mem_3585, data_read_dword_3391_delayed_5_0_3644, tmp_var);
      read_data_line_3649 <= tmp_var; --
    end process;
    -- binary operator OR_u1_u1_3727_inst
    process(do_write_replaced_line_to_mem_3585, do_read_line_from_mem_3546) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(do_write_replaced_line_to_mem_3585, do_read_line_from_mem_3546, tmp_var);
      call_write_mem_3728 <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_L2_TAGS_RESPONSE_3498_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(33 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_L2_TAGS_RESPONSE_3498_inst_req_0;
      RPIPE_L2_TAGS_RESPONSE_3498_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_L2_TAGS_RESPONSE_3498_inst_req_1;
      RPIPE_L2_TAGS_RESPONSE_3498_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= do_tag_access_3276_delayed_4_0_3495(0);
      access_tags_resp_3499 <= data_out(33 downto 0);
      L2_TAGS_RESPONSE_read_0_gI: SplitGuardInterface generic map(name => "L2_TAGS_RESPONSE_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      L2_TAGS_RESPONSE_read_0: InputPort_P2P -- 
        generic map ( name => "L2_TAGS_RESPONSE_read_0", data_width => 34,    bypass_flag => true,   	nonblocking_read_flag => false,  barrier_flag => false,   queue_depth =>  2)
        port map (-- 
          sample_req => reqL(0) , 
          sample_ack => ackL(0), 
          update_req => reqR(0), 
          update_ack => ackR(0), 
          data => data_out, 
          oreq => L2_TAGS_RESPONSE_pipe_read_req(0),
          oack => L2_TAGS_RESPONSE_pipe_read_ack(0),
          odata => L2_TAGS_RESPONSE_pipe_read_data(33 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared inport operator group (1) : RPIPE_NOBLOCK_L2_INVALIDATE_3346_inst 
    InportGroup_1: Block -- 
      signal data_out: std_logic_vector(30 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_NOBLOCK_L2_INVALIDATE_3346_inst_req_0;
      RPIPE_NOBLOCK_L2_INVALIDATE_3346_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_NOBLOCK_L2_INVALIDATE_3346_inst_req_1;
      RPIPE_NOBLOCK_L2_INVALIDATE_3346_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      RPIPE_NOBLOCK_L2_INVALIDATE_3346_wire <= data_out(30 downto 0);
      NOBLOCK_L2_INVALIDATE_read_1_gI: SplitGuardInterface generic map(name => "NOBLOCK_L2_INVALIDATE_read_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      NOBLOCK_L2_INVALIDATE_read_1: InputPortRevised -- 
        generic map ( name => "NOBLOCK_L2_INVALIDATE_read_1", data_width => 31,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => true,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => NOBLOCK_L2_INVALIDATE_pipe_read_req(0),
          oack => NOBLOCK_L2_INVALIDATE_pipe_read_ack(0),
          odata => NOBLOCK_L2_INVALIDATE_pipe_read_data(30 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 1
    -- shared inport operator group (2) : RPIPE_NOBLOCK_L2_REQUEST_3342_inst 
    InportGroup_2: Block -- 
      signal data_out: std_logic_vector(110 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_NOBLOCK_L2_REQUEST_3342_inst_req_0;
      RPIPE_NOBLOCK_L2_REQUEST_3342_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_NOBLOCK_L2_REQUEST_3342_inst_req_1;
      RPIPE_NOBLOCK_L2_REQUEST_3342_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= get_req_3412(0);
      RPIPE_NOBLOCK_L2_REQUEST_3342_wire <= data_out(110 downto 0);
      NOBLOCK_L2_REQUEST_read_2_gI: SplitGuardInterface generic map(name => "NOBLOCK_L2_REQUEST_read_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      NOBLOCK_L2_REQUEST_read_2: InputPort_P2P -- 
        generic map ( name => "NOBLOCK_L2_REQUEST_read_2", data_width => 111,    bypass_flag => false,   	nonblocking_read_flag => true,  barrier_flag => false,   queue_depth =>  2)
        port map (-- 
          sample_req => reqL(0) , 
          sample_ack => ackL(0), 
          update_req => reqR(0), 
          update_ack => ackR(0), 
          data => data_out, 
          oreq => NOBLOCK_L2_REQUEST_pipe_read_req(0),
          oack => NOBLOCK_L2_REQUEST_pipe_read_ack(0),
          odata => NOBLOCK_L2_REQUEST_pipe_read_data(110 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 2
    -- shared outport operator group (0) : WPIPE_L2_RESPONSE_3717_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(64 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_L2_RESPONSE_3717_inst_req_0;
      WPIPE_L2_RESPONSE_3717_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_L2_RESPONSE_3717_inst_req_1;
      WPIPE_L2_RESPONSE_3717_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= send_response_3424_delayed_10_0_3715(0);
      data_in <= l2_resp_3712;
      L2_RESPONSE_write_0_gI: SplitGuardInterface generic map(name => "L2_RESPONSE_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      L2_RESPONSE_write_0: OutputPortRevised -- 
        generic map ( name => "L2_RESPONSE", data_width => 65, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => L2_RESPONSE_pipe_write_req(0),
          oack => L2_RESPONSE_pipe_write_ack(0),
          odata => L2_RESPONSE_pipe_write_data(64 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    -- shared outport operator group (1) : WPIPE_L2_TO_L1_INVALIDATE_3397_inst 
    OutportGroup_1: Block -- 
      signal data_in: std_logic_vector(29 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_L2_TO_L1_INVALIDATE_3397_inst_req_0;
      WPIPE_L2_TO_L1_INVALIDATE_3397_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_L2_TO_L1_INVALIDATE_3397_inst_req_1;
      WPIPE_L2_TO_L1_INVALIDATE_3397_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= inv_valid_3388(0);
      data_in <= inv_pa_line_address_3392;
      L2_TO_L1_INVALIDATE_write_1_gI: SplitGuardInterface generic map(name => "L2_TO_L1_INVALIDATE_write_1_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      L2_TO_L1_INVALIDATE_write_1: OutputPortRevised -- 
        generic map ( name => "L2_TO_L1_INVALIDATE", data_width => 30, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => L2_TO_L1_INVALIDATE_pipe_write_req(0),
          oack => L2_TO_L1_INVALIDATE_pipe_write_ack(0),
          odata => L2_TO_L1_INVALIDATE_pipe_write_data(29 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 1
    -- shared outport operator group (2) : WPIPE_NOBLOCK_L2_TAGS_REQUEST_3490_inst 
    OutportGroup_2: Block -- 
      signal data_in: std_logic_vector(44 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_NOBLOCK_L2_TAGS_REQUEST_3490_inst_req_0;
      WPIPE_NOBLOCK_L2_TAGS_REQUEST_3490_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_NOBLOCK_L2_TAGS_REQUEST_3490_inst_req_1;
      WPIPE_NOBLOCK_L2_TAGS_REQUEST_3490_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= do_tag_access_3464(0);
      data_in <= access_tags_command_3488;
      NOBLOCK_L2_TAGS_REQUEST_write_2_gI: SplitGuardInterface generic map(name => "NOBLOCK_L2_TAGS_REQUEST_write_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      NOBLOCK_L2_TAGS_REQUEST_write_2: OutputPortRevised -- 
        generic map ( name => "NOBLOCK_L2_TAGS_REQUEST", data_width => 45, num_reqs => 1, input_buffering => inBUFs, full_rate => true,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => NOBLOCK_L2_TAGS_REQUEST_pipe_write_req(0),
          oack => NOBLOCK_L2_TAGS_REQUEST_pipe_write_ack(0),
          odata => NOBLOCK_L2_TAGS_REQUEST_pipe_write_data(44 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 2
    -- shared outport operator group (3) : WPIPE_sys_mem_lock_3331_inst 
    OutportGroup_3: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_sys_mem_lock_3331_inst_req_0;
      WPIPE_sys_mem_lock_3331_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_sys_mem_lock_3331_inst_req_1;
      WPIPE_sys_mem_lock_3331_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <=  '1';
      data_in <= type_cast_3333_wire_constant;
      sys_mem_lock_write_3_gI: SplitGuardInterface generic map(name => "sys_mem_lock_write_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      sys_mem_lock_write_3: OutputPortRevised -- 
        generic map ( name => "sys_mem_lock", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => sys_mem_lock_pipe_write_req(0),
          oack => sys_mem_lock_pipe_write_ack(0),
          odata => sys_mem_lock_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 3
    volatile_operator_dwordId_6962: dwordId_Volatile port map(pa => pa_3372, dword_id => call_dwordId_expr_3431_wire); 
    volatile_operator_lineAddress_6958: lineAddress_Volatile port map(pa => pa_3372, pa_line_address => call_lineAddress_expr_3423_wire); 
    volatile_operator_paTag_6964: paTag_Volatile port map(pa => pa_3372, pa_tag => call_paTag_expr_3435_wire); 
    volatile_operator_setId_6960: setId_Volatile port map(pa => pa_3372, set_id => call_setId_expr_3427_wire); 
    -- shared call operator group (4) : call_stmt_3633_call 
    readMemoryFromL2_call_group_4: Block -- 
      signal data_in: std_logic_vector(29 downto 0);
      signal data_out: std_logic_vector(511 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_3633_call_req_0;
      call_stmt_3633_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_3633_call_req_1;
      call_stmt_3633_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= do_read_line_from_mem_3546(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      readMemoryFromL2_call_group_4_gI: SplitGuardInterface generic map(name => "readMemoryFromL2_call_group_4_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= pa_line_address_3381_delayed_5_0_3629;
      pa_mem_cache_line_3633 <= data_out(511 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 30,
        owidth => 30,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => readMemoryFromL2_call_reqs(0),
          ackR => readMemoryFromL2_call_acks(0),
          dataR => readMemoryFromL2_call_data(29 downto 0),
          tagR => readMemoryFromL2_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 512,
          owidth => 512,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => readMemoryFromL2_return_acks(0), -- cross-over
          ackL => readMemoryFromL2_return_reqs(0), -- cross-over
          dataL => readMemoryFromL2_return_data(511 downto 0),
          tagL => readMemoryFromL2_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 4
    operator_accessL2DataMemX4096X512_7039_block : block -- 
      signal sample_req, sample_ack, update_req, update_ack: BooleanArray(0 downto 0); 
      signal sample_req_ug, sample_ack_ug, update_req_ug, update_ack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      sample_req_ug(0) <= call_stmt_3693_call_req_0;
      call_stmt_3693_call_ack_0<= sample_ack_ug(0);
      update_req_ug(0) <= call_stmt_3693_call_req_1;
      call_stmt_3693_call_ack_1<= update_ack_ug(0);
      guard_vector(0) <=  access_data_mem_3394_delayed_4_0_3652(0);
      call_stmt_3693_call_gI: SplitGuardInterface generic map(name => "call_stmt_3693_call_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_ug,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_ug,
        cr_in => update_req_ug,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_ug,
        guards => guard_vector); -- 
      call_stmt_3693_call: accessL2DataMemX4096X512_Operator  port map ( -- 
        sample_req => sample_req(0), 
        sample_ack => sample_ack(0), 
        update_req => update_req(0), 
        update_ack => update_ack(0), 
        read_data_line => read_data_line_3395_delayed_4_0_3655,
        data_write_dword => data_write_dword_3396_delayed_9_0_3658,
        data_read_dword => data_read_dword_3397_delayed_9_0_3661,
        data_write_new_line => data_write_new_line_3398_delayed_4_0_3664,
        do_write_replaced_line_to_mem => do_write_replaced_line_to_mem_3399_delayed_4_0_3667,
        byte_mask => byte_mask_3400_delayed_9_0_3670,
        line_id => line_id_3401_delayed_4_0_3673,
        pa_dword_id => pa_dword_id_3402_delayed_9_0_3676,
        w_dword => wdata_3403_delayed_9_0_3679,
        line_to_be_inserted => pa_mem_cache_line_3633,
        read_dword_from_data => read_dword_from_data_3693,
        writeback_line_from_data => writeback_line_from_data_3693,
        clk => clk, reset => reset  
        -- 
      );-- 
    end block;
    -- shared call operator group (6) : call_stmt_3750_call 
    writeMemoryFromL2_call_group_6: Block -- 
      signal data_in: std_logic_vector(551 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs: IntegerArray(0 downto 0) := (others => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 4);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_3750_call_req_0;
      call_stmt_3750_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_3750_call_req_1;
      call_stmt_3750_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <= call_write_mem_3437_delayed_5_0_3731(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      writeMemoryFromL2_call_group_6_gI: SplitGuardInterface generic map(name => "writeMemoryFromL2_call_group_6_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= do_read_line_from_mem_3438_delayed_5_0_3734 & do_write_replaced_line_to_mem_3439_delayed_5_0_3737 & dirty_word_mask_3440_delayed_5_0_3740 & write_back_line_address_3441_delayed_5_0_3743 & writeback_line_from_data_3693;
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 552,
        owidth => 552,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => writeMemoryFromL2_call_reqs(0),
          ackR => writeMemoryFromL2_call_acks(0),
          dataR => writeMemoryFromL2_call_data(551 downto 0),
          tagR => writeMemoryFromL2_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseNoData -- 
        generic map ( -- 
          detailed_buffering_per_output => outBUFs, 
          twidth => 1,
          name => "OutputDemuxBaseNoData",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          reqL => writeMemoryFromL2_return_acks(0), -- cross-over
          ackL => writeMemoryFromL2_return_reqs(0), -- cross-over
          tagL => writeMemoryFromL2_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 6
    -- 
  end Block; -- data_path
  -- 
end l2CacheDaemon_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library l2_cache_lib;
use l2_cache_lib.l2_cache_global_package.all;
entity lineAddress_Volatile is -- 
  port ( -- 
    pa : in  std_logic_vector(35 downto 0);
    pa_line_address : out  std_logic_vector(29 downto 0)-- 
  );
  -- 
end entity lineAddress_Volatile;
architecture lineAddress_Volatile_arch of lineAddress_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(36-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal pa_buffer :  std_logic_vector(35 downto 0);
  -- output port buffer signals
  signal pa_line_address_buffer :  std_logic_vector(29 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  pa_buffer <= pa;
  -- output handling  -------------------------------------------------------
  pa_line_address <= pa_line_address_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    -- 
  begin -- 
    -- flow-through slice operator slice_3049_inst
    pa_line_address_buffer <= pa_buffer(35 downto 6);
    -- 
  end Block; -- data_path
  -- 
end lineAddress_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library l2_cache_lib;
use l2_cache_lib.l2_cache_global_package.all;
entity nextFreeIndex_Volatile is -- 
  port ( -- 
    from_index : in  std_logic_vector(2 downto 0);
    set_valids : in  std_logic_vector(7 downto 0);
    next_free_index : out  std_logic_vector(2 downto 0)-- 
  );
  -- 
end entity nextFreeIndex_Volatile;
architecture nextFreeIndex_Volatile_arch of nextFreeIndex_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(11-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal from_index_buffer :  std_logic_vector(2 downto 0);
  signal set_valids_buffer :  std_logic_vector(7 downto 0);
  -- output port buffer signals
  signal next_free_index_buffer :  std_logic_vector(2 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  from_index_buffer <= from_index;
  set_valids_buffer <= set_valids;
  -- output handling  -------------------------------------------------------
  next_free_index <= next_free_index_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal MUX_1727_wire : std_logic_vector(2 downto 0);
    signal MUX_1728_wire : std_logic_vector(2 downto 0);
    signal MUX_1729_wire : std_logic_vector(2 downto 0);
    signal MUX_1730_wire : std_logic_vector(2 downto 0);
    signal MUX_1731_wire : std_logic_vector(2 downto 0);
    signal MUX_1732_wire : std_logic_vector(2 downto 0);
    signal NOT_u1_u1_1705_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1709_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1712_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1715_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1718_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1721_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1724_wire : std_logic_vector(0 downto 0);
    signal konst_1710_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1713_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1716_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1719_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1722_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1725_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1726_wire_constant : std_logic_vector(2 downto 0);
    signal offset_1734 : std_logic_vector(2 downto 0);
    signal rset_valids_1674 : std_logic_vector(7 downto 0);
    signal type_cast_1672_wire : std_logic_vector(7 downto 0);
    signal type_cast_1707_wire_constant : std_logic_vector(2 downto 0);
    signal v1_1678 : std_logic_vector(0 downto 0);
    signal v2_1682 : std_logic_vector(0 downto 0);
    signal v3_1686 : std_logic_vector(0 downto 0);
    signal v4_1690 : std_logic_vector(0 downto 0);
    signal v5_1694 : std_logic_vector(0 downto 0);
    signal v6_1698 : std_logic_vector(0 downto 0);
    signal v7_1702 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    konst_1710_wire_constant <= "010";
    konst_1713_wire_constant <= "011";
    konst_1716_wire_constant <= "100";
    konst_1719_wire_constant <= "101";
    konst_1722_wire_constant <= "110";
    konst_1725_wire_constant <= "111";
    konst_1726_wire_constant <= "001";
    type_cast_1707_wire_constant <= "001";
    -- flow-through select operator MUX_1727_inst
    MUX_1727_wire <= konst_1725_wire_constant when (NOT_u1_u1_1724_wire(0) /=  '0') else konst_1726_wire_constant;
    -- flow-through select operator MUX_1728_inst
    MUX_1728_wire <= konst_1722_wire_constant when (NOT_u1_u1_1721_wire(0) /=  '0') else MUX_1727_wire;
    -- flow-through select operator MUX_1729_inst
    MUX_1729_wire <= konst_1719_wire_constant when (NOT_u1_u1_1718_wire(0) /=  '0') else MUX_1728_wire;
    -- flow-through select operator MUX_1730_inst
    MUX_1730_wire <= konst_1716_wire_constant when (NOT_u1_u1_1715_wire(0) /=  '0') else MUX_1729_wire;
    -- flow-through select operator MUX_1731_inst
    MUX_1731_wire <= konst_1713_wire_constant when (NOT_u1_u1_1712_wire(0) /=  '0') else MUX_1730_wire;
    -- flow-through select operator MUX_1732_inst
    MUX_1732_wire <= konst_1710_wire_constant when (NOT_u1_u1_1709_wire(0) /=  '0') else MUX_1731_wire;
    -- flow-through select operator MUX_1733_inst
    offset_1734 <= type_cast_1707_wire_constant when (NOT_u1_u1_1705_wire(0) /=  '0') else MUX_1732_wire;
    -- flow-through slice operator slice_1677_inst
    v1_1678 <= rset_valids_1674(6 downto 6);
    -- flow-through slice operator slice_1681_inst
    v2_1682 <= rset_valids_1674(5 downto 5);
    -- flow-through slice operator slice_1685_inst
    v3_1686 <= rset_valids_1674(4 downto 4);
    -- flow-through slice operator slice_1689_inst
    v4_1690 <= rset_valids_1674(3 downto 3);
    -- flow-through slice operator slice_1693_inst
    v5_1694 <= rset_valids_1674(2 downto 2);
    -- flow-through slice operator slice_1697_inst
    v6_1698 <= rset_valids_1674(1 downto 1);
    -- flow-through slice operator slice_1701_inst
    v7_1702 <= rset_valids_1674(0 downto 0);
    -- interlock type_cast_1672_inst
    process(from_index_buffer) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 2 downto 0) := from_index_buffer(2 downto 0);
      type_cast_1672_wire <= tmp_var; -- 
    end process;
    -- binary operator ADD_u3_u3_1738_inst
    process(from_index_buffer, offset_1734) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApIntAdd_proc(from_index_buffer, offset_1734, tmp_var);
      next_free_index_buffer <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1705_inst
    process(v1_1678) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", v1_1678, tmp_var);
      NOT_u1_u1_1705_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1709_inst
    process(v2_1682) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", v2_1682, tmp_var);
      NOT_u1_u1_1709_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1712_inst
    process(v3_1686) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", v3_1686, tmp_var);
      NOT_u1_u1_1712_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1715_inst
    process(v4_1690) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", v4_1690, tmp_var);
      NOT_u1_u1_1715_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1718_inst
    process(v5_1694) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", v5_1694, tmp_var);
      NOT_u1_u1_1718_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1721_inst
    process(v6_1698) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", v6_1698, tmp_var);
      NOT_u1_u1_1721_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1724_inst
    process(v7_1702) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", v7_1702, tmp_var);
      NOT_u1_u1_1724_wire <= tmp_var; -- 
    end process;
    -- binary operator ROL_u8_u8_1673_inst
    process(set_valids_buffer, type_cast_1672_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApIntROL_proc(set_valids_buffer, type_cast_1672_wire, tmp_var);
      rset_valids_1674 <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end nextFreeIndex_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library l2_cache_lib;
use l2_cache_lib.l2_cache_global_package.all;
entity paTag_Volatile is -- 
  port ( -- 
    pa : in  std_logic_vector(35 downto 0);
    pa_tag : out  std_logic_vector(20 downto 0)-- 
  );
  -- 
end entity paTag_Volatile;
architecture paTag_Volatile_arch of paTag_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(36-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal pa_buffer :  std_logic_vector(35 downto 0);
  -- output port buffer signals
  signal pa_tag_buffer :  std_logic_vector(20 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  pa_buffer <= pa;
  -- output handling  -------------------------------------------------------
  pa_tag <= pa_tag_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    -- 
  begin -- 
    -- flow-through slice operator slice_3065_inst
    pa_tag_buffer <= pa_buffer(35 downto 15);
    -- 
  end Block; -- data_path
  -- 
end paTag_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library l2_cache_lib;
use l2_cache_lib.l2_cache_global_package.all;
entity readMemoryFromL2 is -- 
  generic (tag_length : integer); 
  port ( -- 
    line_address : in  std_logic_vector(29 downto 0);
    rline : out  std_logic_vector(511 downto 0);
    sys_mem_lock_pipe_read_req : out  std_logic_vector(0 downto 0);
    sys_mem_lock_pipe_read_ack : in   std_logic_vector(0 downto 0);
    sys_mem_lock_pipe_read_data : in   std_logic_vector(0 downto 0);
    accessSysMem_call_reqs : out  std_logic_vector(0 downto 0);
    accessSysMem_call_acks : in   std_logic_vector(0 downto 0);
    accessSysMem_call_data : out  std_logic_vector(108 downto 0);
    accessSysMem_call_tag  :  out  std_logic_vector(0 downto 0);
    accessSysMem_return_reqs : out  std_logic_vector(0 downto 0);
    accessSysMem_return_acks : in   std_logic_vector(0 downto 0);
    accessSysMem_return_data : in   std_logic_vector(63 downto 0);
    accessSysMem_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity readMemoryFromL2;
architecture readMemoryFromL2_arch of readMemoryFromL2 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 30)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 512)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal line_address_buffer :  std_logic_vector(29 downto 0);
  signal line_address_update_enable: Boolean;
  -- output port buffer signals
  signal rline_buffer :  std_logic_vector(511 downto 0);
  signal rline_update_enable: Boolean;
  signal readMemoryFromL2_CP_2700_start: Boolean;
  signal readMemoryFromL2_CP_2700_symbol: Boolean;
  -- volatile/operator module components. 
  component accessSysMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      byte_mask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEM_TO_L2CACHE_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEM_TO_L2CACHE_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEM_TO_L2CACHE_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      L2CACHE_TO_MEM_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      L2CACHE_TO_MEM_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      L2CACHE_TO_MEM_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- links between control-path and data-path
  signal W_s0_2928_delayed_8_0_3121_inst_ack_1 : boolean;
  signal W_r0_3125_inst_ack_1 : boolean;
  signal do_while_stmt_3077_branch_req_0 : boolean;
  signal W_r0_3125_inst_ack_0 : boolean;
  signal phi_stmt_3079_ack_0 : boolean;
  signal phi_stmt_3079_req_1 : boolean;
  signal call_stmt_3112_call_req_0 : boolean;
  signal call_stmt_3112_call_ack_0 : boolean;
  signal RPIPE_sys_mem_lock_3074_inst_req_0 : boolean;
  signal W_r0_3125_inst_req_0 : boolean;
  signal RPIPE_sys_mem_lock_3074_inst_ack_0 : boolean;
  signal RPIPE_sys_mem_lock_3074_inst_ack_1 : boolean;
  signal call_stmt_3112_call_req_1 : boolean;
  signal call_stmt_3112_call_ack_1 : boolean;
  signal W_s0_2928_delayed_8_0_3121_inst_req_0 : boolean;
  signal RPIPE_sys_mem_lock_3074_inst_req_1 : boolean;
  signal n_DWORD_ID_3094_3081_buf_ack_0 : boolean;
  signal W_r1_3137_inst_ack_0 : boolean;
  signal n_DWORD_ID_3094_3081_buf_req_1 : boolean;
  signal n_DWORD_ID_3094_3081_buf_ack_1 : boolean;
  signal W_s0_2928_delayed_8_0_3121_inst_ack_0 : boolean;
  signal W_s0_2928_delayed_8_0_3121_inst_req_1 : boolean;
  signal W_r1_3137_inst_req_1 : boolean;
  signal n_DWORD_ID_3094_3081_buf_req_0 : boolean;
  signal W_r0_3125_inst_req_1 : boolean;
  signal W_s1_2937_delayed_8_0_3133_inst_ack_1 : boolean;
  signal W_s4_2964_delayed_8_0_3169_inst_req_0 : boolean;
  signal W_s4_2964_delayed_8_0_3169_inst_ack_0 : boolean;
  signal W_s1_2937_delayed_8_0_3133_inst_req_1 : boolean;
  signal phi_stmt_3079_req_0 : boolean;
  signal W_r1_3137_inst_ack_1 : boolean;
  signal W_r1_3137_inst_req_0 : boolean;
  signal W_r3_3161_inst_req_1 : boolean;
  signal W_r3_3161_inst_ack_1 : boolean;
  signal W_r3_3161_inst_req_0 : boolean;
  signal W_r3_3161_inst_ack_0 : boolean;
  signal W_r2_3149_inst_ack_1 : boolean;
  signal W_r2_3149_inst_req_1 : boolean;
  signal W_r2_3149_inst_ack_0 : boolean;
  signal W_r2_3149_inst_req_0 : boolean;
  signal W_s1_2937_delayed_8_0_3133_inst_ack_0 : boolean;
  signal W_s2_2946_delayed_8_0_3145_inst_ack_1 : boolean;
  signal W_s1_2937_delayed_8_0_3133_inst_req_0 : boolean;
  signal W_s2_2946_delayed_8_0_3145_inst_req_1 : boolean;
  signal W_s2_2946_delayed_8_0_3145_inst_req_0 : boolean;
  signal W_s4_2964_delayed_8_0_3169_inst_req_1 : boolean;
  signal W_s4_2964_delayed_8_0_3169_inst_ack_1 : boolean;
  signal W_s2_2946_delayed_8_0_3145_inst_ack_0 : boolean;
  signal W_s3_2955_delayed_8_0_3157_inst_ack_1 : boolean;
  signal W_s3_2955_delayed_8_0_3157_inst_req_1 : boolean;
  signal W_s3_2955_delayed_8_0_3157_inst_ack_0 : boolean;
  signal W_s3_2955_delayed_8_0_3157_inst_req_0 : boolean;
  signal W_r4_3173_inst_req_0 : boolean;
  signal W_r4_3173_inst_ack_0 : boolean;
  signal W_r4_3173_inst_req_1 : boolean;
  signal W_r4_3173_inst_ack_1 : boolean;
  signal W_s5_2973_delayed_8_0_3181_inst_req_0 : boolean;
  signal W_s5_2973_delayed_8_0_3181_inst_ack_0 : boolean;
  signal W_s5_2973_delayed_8_0_3181_inst_req_1 : boolean;
  signal W_s5_2973_delayed_8_0_3181_inst_ack_1 : boolean;
  signal W_r5_3185_inst_req_0 : boolean;
  signal W_r5_3185_inst_ack_0 : boolean;
  signal W_r5_3185_inst_req_1 : boolean;
  signal W_r5_3185_inst_ack_1 : boolean;
  signal W_s6_2982_delayed_8_0_3193_inst_req_0 : boolean;
  signal W_s6_2982_delayed_8_0_3193_inst_ack_0 : boolean;
  signal W_s6_2982_delayed_8_0_3193_inst_req_1 : boolean;
  signal W_s6_2982_delayed_8_0_3193_inst_ack_1 : boolean;
  signal W_r6_3197_inst_req_0 : boolean;
  signal W_r6_3197_inst_ack_0 : boolean;
  signal W_r6_3197_inst_req_1 : boolean;
  signal W_r6_3197_inst_ack_1 : boolean;
  signal W_s7_2991_delayed_8_0_3205_inst_req_0 : boolean;
  signal W_s7_2991_delayed_8_0_3205_inst_ack_0 : boolean;
  signal W_s7_2991_delayed_8_0_3205_inst_req_1 : boolean;
  signal W_s7_2991_delayed_8_0_3205_inst_ack_1 : boolean;
  signal W_r7_3209_inst_req_0 : boolean;
  signal W_r7_3209_inst_ack_0 : boolean;
  signal W_r7_3209_inst_req_1 : boolean;
  signal W_r7_3209_inst_ack_1 : boolean;
  signal do_while_stmt_3077_branch_ack_0 : boolean;
  signal do_while_stmt_3077_branch_ack_1 : boolean;
  signal CONCAT_u256_u512_3230_inst_req_0 : boolean;
  signal CONCAT_u256_u512_3230_inst_ack_0 : boolean;
  signal CONCAT_u256_u512_3230_inst_req_1 : boolean;
  signal CONCAT_u256_u512_3230_inst_ack_1 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "readMemoryFromL2_input_buffer", -- 
      buffer_size => 0,
      bypass_flag => true,
      data_width => tag_length + 30) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(29 downto 0) <= line_address;
  line_address_buffer <= in_buffer_data_out(29 downto 0);
  in_buffer_data_in(tag_length + 29 downto 30) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 29 downto 30);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  readMemoryFromL2_CP_2700_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "readMemoryFromL2_out_buffer", -- 
      buffer_size => 0,
      full_rate => false,
      data_width => tag_length + 512) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(511 downto 0) <= rline_buffer;
  rline <= out_buffer_data_out(511 downto 0);
  out_buffer_data_in(tag_length + 511 downto 512) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length + 511 downto 512);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= readMemoryFromL2_CP_2700_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= readMemoryFromL2_CP_2700_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= readMemoryFromL2_CP_2700_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  readMemoryFromL2_CP_2700: Block -- control-path 
    signal readMemoryFromL2_CP_2700_elements: BooleanArray(106 downto 0);
    -- 
  begin -- 
    readMemoryFromL2_CP_2700_elements(0) <= readMemoryFromL2_CP_2700_start;
    readMemoryFromL2_CP_2700_symbol <= readMemoryFromL2_CP_2700_elements(106);
    -- CP-element group 0:  transition  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	1 
    -- CP-element group 0:  members (5) 
      -- CP-element group 0: 	 assign_stmt_3075/RPIPE_sys_mem_lock_3074_Sample/$entry
      -- CP-element group 0: 	 assign_stmt_3075/$entry
      -- CP-element group 0: 	 assign_stmt_3075/RPIPE_sys_mem_lock_3074_Sample/rr
      -- CP-element group 0: 	 assign_stmt_3075/RPIPE_sys_mem_lock_3074_sample_start_
      -- CP-element group 0: 	 $entry
      -- 
    rr_2713_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_2713_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(0), ack => RPIPE_sys_mem_lock_3074_inst_req_0); -- 
    -- CP-element group 1:  transition  input  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	0 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	2 
    -- CP-element group 1:  members (6) 
      -- CP-element group 1: 	 assign_stmt_3075/RPIPE_sys_mem_lock_3074_sample_completed_
      -- CP-element group 1: 	 assign_stmt_3075/RPIPE_sys_mem_lock_3074_update_start_
      -- CP-element group 1: 	 assign_stmt_3075/RPIPE_sys_mem_lock_3074_Sample/$exit
      -- CP-element group 1: 	 assign_stmt_3075/RPIPE_sys_mem_lock_3074_Sample/ra
      -- CP-element group 1: 	 assign_stmt_3075/RPIPE_sys_mem_lock_3074_Update/$entry
      -- CP-element group 1: 	 assign_stmt_3075/RPIPE_sys_mem_lock_3074_Update/cr
      -- 
    ra_2714_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 1_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_sys_mem_lock_3074_inst_ack_0, ack => readMemoryFromL2_CP_2700_elements(1)); -- 
    cr_2718_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_2718_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(1), ack => RPIPE_sys_mem_lock_3074_inst_req_1); -- 
    -- CP-element group 2:  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	1 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	4 
    -- CP-element group 2:  members (7) 
      -- CP-element group 2: 	 assign_stmt_3075/RPIPE_sys_mem_lock_3074_update_completed_
      -- CP-element group 2: 	 assign_stmt_3075/RPIPE_sys_mem_lock_3074_Update/ca
      -- CP-element group 2: 	 assign_stmt_3075/$exit
      -- CP-element group 2: 	 branch_block_stmt_3076/do_while_stmt_3077__entry__
      -- CP-element group 2: 	 branch_block_stmt_3076/$entry
      -- CP-element group 2: 	 assign_stmt_3075/RPIPE_sys_mem_lock_3074_Update/$exit
      -- CP-element group 2: 	 branch_block_stmt_3076/branch_block_stmt_3076__entry__
      -- 
    ca_2719_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => RPIPE_sys_mem_lock_3074_inst_ack_1, ack => readMemoryFromL2_CP_2700_elements(2)); -- 
    -- CP-element group 3:  fork  transition  place  output  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	104 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	105 
    -- CP-element group 3: 	106 
    -- CP-element group 3:  members (10) 
      -- CP-element group 3: 	 branch_block_stmt_3076/$exit
      -- CP-element group 3: 	 branch_block_stmt_3076/do_while_stmt_3077__exit__
      -- CP-element group 3: 	 branch_block_stmt_3076/branch_block_stmt_3076__exit__
      -- CP-element group 3: 	 assign_stmt_3231/$entry
      -- CP-element group 3: 	 assign_stmt_3231/CONCAT_u256_u512_3230_sample_start_
      -- CP-element group 3: 	 assign_stmt_3231/CONCAT_u256_u512_3230_update_start_
      -- CP-element group 3: 	 assign_stmt_3231/CONCAT_u256_u512_3230_Sample/$entry
      -- CP-element group 3: 	 assign_stmt_3231/CONCAT_u256_u512_3230_Sample/rr
      -- CP-element group 3: 	 assign_stmt_3231/CONCAT_u256_u512_3230_Update/$entry
      -- CP-element group 3: 	 assign_stmt_3231/CONCAT_u256_u512_3230_Update/cr
      -- 
    rr_3050_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " rr_3050_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(3), ack => CONCAT_u256_u512_3230_inst_req_0); -- 
    cr_3055_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " cr_3055_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(3), ack => CONCAT_u256_u512_3230_inst_req_1); -- 
    readMemoryFromL2_CP_2700_elements(3) <= readMemoryFromL2_CP_2700_elements(104);
    -- CP-element group 4:  transition  place  bypass  pipeline-parent 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	2 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	10 
    -- CP-element group 4:  members (2) 
      -- CP-element group 4: 	 branch_block_stmt_3076/do_while_stmt_3077/$entry
      -- CP-element group 4: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077__entry__
      -- 
    readMemoryFromL2_CP_2700_elements(4) <= readMemoryFromL2_CP_2700_elements(2);
    -- CP-element group 5:  merge  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	104 
    -- CP-element group 5:  members (1) 
      -- CP-element group 5: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077__exit__
      -- 
    -- Element group readMemoryFromL2_CP_2700_elements(5) is bound as output of CP function.
    -- CP-element group 6:  merge  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	9 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_3076/do_while_stmt_3077/loop_back
      -- 
    -- Element group readMemoryFromL2_CP_2700_elements(6) is bound as output of CP function.
    -- CP-element group 7:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: 	12 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	102 
    -- CP-element group 7: 	103 
    -- CP-element group 7:  members (3) 
      -- CP-element group 7: 	 branch_block_stmt_3076/do_while_stmt_3077/condition_done
      -- CP-element group 7: 	 branch_block_stmt_3076/do_while_stmt_3077/loop_exit/$entry
      -- CP-element group 7: 	 branch_block_stmt_3076/do_while_stmt_3077/loop_taken/$entry
      -- 
    readMemoryFromL2_CP_2700_elements(7) <= readMemoryFromL2_CP_2700_elements(12);
    -- CP-element group 8:  branch  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	101 
    -- CP-element group 8: successors 
    -- CP-element group 8:  members (1) 
      -- CP-element group 8: 	 branch_block_stmt_3076/do_while_stmt_3077/loop_body_done
      -- 
    readMemoryFromL2_CP_2700_elements(8) <= readMemoryFromL2_CP_2700_elements(101);
    -- CP-element group 9:  transition  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	6 
    -- CP-element group 9: successors 
    -- CP-element group 9: 	19 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/back_edge_to_loop_body
      -- 
    readMemoryFromL2_CP_2700_elements(9) <= readMemoryFromL2_CP_2700_elements(6);
    -- CP-element group 10:  transition  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	4 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	21 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/first_time_through_loop_body
      -- 
    readMemoryFromL2_CP_2700_elements(10) <= readMemoryFromL2_CP_2700_elements(4);
    -- CP-element group 11:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	15 
    -- CP-element group 11: 	16 
    -- CP-element group 11: 	100 
    -- CP-element group 11:  members (2) 
      -- CP-element group 11: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/$entry
      -- CP-element group 11: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/loop_body_start
      -- 
    -- Element group readMemoryFromL2_CP_2700_elements(11) is bound as output of CP function.
    -- CP-element group 12:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: 	14 
    -- CP-element group 12: 	18 
    -- CP-element group 12: 	100 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	7 
    -- CP-element group 12:  members (1) 
      -- CP-element group 12: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/condition_evaluated
      -- 
    condition_evaluated_2741_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_2741_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(12), ack => do_while_stmt_3077_branch_req_0); -- 
    readMemoryFromL2_cp_element_group_12: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_12"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= readMemoryFromL2_CP_2700_elements(14) & readMemoryFromL2_CP_2700_elements(18) & readMemoryFromL2_CP_2700_elements(100);
      gj_readMemoryFromL2_cp_element_group_12 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(12), clk => clk, reset => reset); --
    end block;
    -- CP-element group 13:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	15 
    -- CP-element group 13: marked-predecessors 
    -- CP-element group 13: 	18 
    -- CP-element group 13: successors 
    -- CP-element group 13:  members (2) 
      -- CP-element group 13: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/aggregated_phi_sample_req
      -- CP-element group 13: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/phi_stmt_3079_sample_start__ps
      -- 
    readMemoryFromL2_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readMemoryFromL2_CP_2700_elements(15) & readMemoryFromL2_CP_2700_elements(18);
      gj_readMemoryFromL2_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	17 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	12 
    -- CP-element group 14:  members (1) 
      -- CP-element group 14: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/aggregated_phi_sample_ack_d
      -- 
    -- Element group readMemoryFromL2_CP_2700_elements(14) is a control-delay.
    cp_element_14_delay: control_delay_element  generic map(name => " 14_delay", delay_value => 1)  port map(req => readMemoryFromL2_CP_2700_elements(17), ack => readMemoryFromL2_CP_2700_elements(14), clk => clk, reset =>reset);
    -- CP-element group 15:  join  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	11 
    -- CP-element group 15: marked-predecessors 
    -- CP-element group 15: 	17 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	13 
    -- CP-element group 15:  members (1) 
      -- CP-element group 15: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/phi_stmt_3079_sample_start_
      -- 
    readMemoryFromL2_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readMemoryFromL2_CP_2700_elements(11) & readMemoryFromL2_CP_2700_elements(17);
      gj_readMemoryFromL2_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	11 
    -- CP-element group 16: marked-predecessors 
    -- CP-element group 16: 	34 
    -- CP-element group 16: 	38 
    -- CP-element group 16: 	46 
    -- CP-element group 16: 	54 
    -- CP-element group 16: 	62 
    -- CP-element group 16: 	70 
    -- CP-element group 16: 	78 
    -- CP-element group 16: 	86 
    -- CP-element group 16: 	94 
    -- CP-element group 16: successors 
    -- CP-element group 16:  members (3) 
      -- CP-element group 16: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/phi_stmt_3079_update_start__ps
      -- CP-element group 16: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/phi_stmt_3079_update_start_
      -- CP-element group 16: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/aggregated_phi_update_req
      -- 
    readMemoryFromL2_cp_element_group_16: block -- 
      constant place_capacities: IntegerArray(0 to 9) := (0 => 15,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_markings: IntegerArray(0 to 9)  := (0 => 0,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1,8 => 1,9 => 1);
      constant place_delays: IntegerArray(0 to 9) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0,9 => 0);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_16"; 
      signal preds: BooleanArray(1 to 10); -- 
    begin -- 
      preds <= readMemoryFromL2_CP_2700_elements(11) & readMemoryFromL2_CP_2700_elements(34) & readMemoryFromL2_CP_2700_elements(38) & readMemoryFromL2_CP_2700_elements(46) & readMemoryFromL2_CP_2700_elements(54) & readMemoryFromL2_CP_2700_elements(62) & readMemoryFromL2_CP_2700_elements(70) & readMemoryFromL2_CP_2700_elements(78) & readMemoryFromL2_CP_2700_elements(86) & readMemoryFromL2_CP_2700_elements(94);
      gj_readMemoryFromL2_cp_element_group_16 : generic_join generic map(name => joinName, number_of_predecessors => 10, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(16), clk => clk, reset => reset); --
    end block;
    -- CP-element group 17:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	14 
    -- CP-element group 17: 	101 
    -- CP-element group 17: marked-successors 
    -- CP-element group 17: 	15 
    -- CP-element group 17:  members (3) 
      -- CP-element group 17: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/aggregated_phi_sample_ack
      -- CP-element group 17: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/phi_stmt_3079_sample_completed__ps
      -- CP-element group 17: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/phi_stmt_3079_sample_completed_
      -- 
    -- Element group readMemoryFromL2_CP_2700_elements(17) is bound as output of CP function.
    -- CP-element group 18:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	12 
    -- CP-element group 18: 	32 
    -- CP-element group 18: 	36 
    -- CP-element group 18: 	44 
    -- CP-element group 18: 	52 
    -- CP-element group 18: 	60 
    -- CP-element group 18: 	68 
    -- CP-element group 18: 	76 
    -- CP-element group 18: 	84 
    -- CP-element group 18: 	92 
    -- CP-element group 18: marked-successors 
    -- CP-element group 18: 	13 
    -- CP-element group 18:  members (3) 
      -- CP-element group 18: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/phi_stmt_3079_update_completed__ps
      -- CP-element group 18: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/phi_stmt_3079_update_completed_
      -- CP-element group 18: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/aggregated_phi_update_ack
      -- 
    -- Element group readMemoryFromL2_CP_2700_elements(18) is bound as output of CP function.
    -- CP-element group 19:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	9 
    -- CP-element group 19: successors 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/phi_stmt_3079_loopback_trigger
      -- 
    readMemoryFromL2_CP_2700_elements(19) <= readMemoryFromL2_CP_2700_elements(9);
    -- CP-element group 20:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: successors 
    -- CP-element group 20:  members (2) 
      -- CP-element group 20: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/phi_stmt_3079_loopback_sample_req_ps
      -- CP-element group 20: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/phi_stmt_3079_loopback_sample_req
      -- 
    phi_stmt_3079_loopback_sample_req_2757_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3079_loopback_sample_req_2757_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(20), ack => phi_stmt_3079_req_0); -- 
    -- Element group readMemoryFromL2_CP_2700_elements(20) is bound as output of CP function.
    -- CP-element group 21:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: 	10 
    -- CP-element group 21: successors 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/phi_stmt_3079_entry_trigger
      -- 
    readMemoryFromL2_CP_2700_elements(21) <= readMemoryFromL2_CP_2700_elements(10);
    -- CP-element group 22:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/phi_stmt_3079_entry_sample_req
      -- CP-element group 22: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/phi_stmt_3079_entry_sample_req_ps
      -- 
    phi_stmt_3079_entry_sample_req_2760_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3079_entry_sample_req_2760_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(22), ack => phi_stmt_3079_req_1); -- 
    -- Element group readMemoryFromL2_CP_2700_elements(22) is bound as output of CP function.
    -- CP-element group 23:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (2) 
      -- CP-element group 23: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/phi_stmt_3079_phi_mux_ack_ps
      -- CP-element group 23: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/phi_stmt_3079_phi_mux_ack
      -- 
    phi_stmt_3079_phi_mux_ack_2763_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 23_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3079_ack_0, ack => readMemoryFromL2_CP_2700_elements(23)); -- 
    -- CP-element group 24:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24: 	26 
    -- CP-element group 24:  members (4) 
      -- CP-element group 24: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/R_n_DWORD_ID_3081_sample_start__ps
      -- CP-element group 24: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/R_n_DWORD_ID_3081_Sample/$entry
      -- CP-element group 24: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/R_n_DWORD_ID_3081_sample_start_
      -- CP-element group 24: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/R_n_DWORD_ID_3081_Sample/req
      -- 
    req_2776_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2776_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(24), ack => n_DWORD_ID_3094_3081_buf_req_0); -- 
    -- Element group readMemoryFromL2_CP_2700_elements(24) is bound as output of CP function.
    -- CP-element group 25:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: successors 
    -- CP-element group 25: 	27 
    -- CP-element group 25:  members (4) 
      -- CP-element group 25: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/R_n_DWORD_ID_3081_update_start__ps
      -- CP-element group 25: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/R_n_DWORD_ID_3081_Update/$entry
      -- CP-element group 25: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/R_n_DWORD_ID_3081_Update/req
      -- CP-element group 25: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/R_n_DWORD_ID_3081_update_start_
      -- 
    req_2781_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2781_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(25), ack => n_DWORD_ID_3094_3081_buf_req_1); -- 
    -- Element group readMemoryFromL2_CP_2700_elements(25) is bound as output of CP function.
    -- CP-element group 26:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: 	24 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (4) 
      -- CP-element group 26: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/R_n_DWORD_ID_3081_sample_completed__ps
      -- CP-element group 26: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/R_n_DWORD_ID_3081_Sample/ack
      -- CP-element group 26: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/R_n_DWORD_ID_3081_sample_completed_
      -- CP-element group 26: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/R_n_DWORD_ID_3081_Sample/$exit
      -- 
    ack_2777_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 26_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_DWORD_ID_3094_3081_buf_ack_0, ack => readMemoryFromL2_CP_2700_elements(26)); -- 
    -- CP-element group 27:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: 	25 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (4) 
      -- CP-element group 27: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/R_n_DWORD_ID_3081_Update/$exit
      -- CP-element group 27: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/R_n_DWORD_ID_3081_update_completed__ps
      -- CP-element group 27: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/R_n_DWORD_ID_3081_Update/ack
      -- CP-element group 27: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/R_n_DWORD_ID_3081_update_completed_
      -- 
    ack_2782_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => n_DWORD_ID_3094_3081_buf_ack_1, ack => readMemoryFromL2_CP_2700_elements(27)); -- 
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/type_cast_3083_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/type_cast_3083_sample_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/type_cast_3083_sample_completed_
      -- CP-element group 28: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/type_cast_3083_sample_start_
      -- 
    -- Element group readMemoryFromL2_CP_2700_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/type_cast_3083_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/type_cast_3083_update_start_
      -- 
    -- Element group readMemoryFromL2_CP_2700_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/type_cast_3083_update_completed__ps
      -- 
    readMemoryFromL2_CP_2700_elements(30) <= readMemoryFromL2_CP_2700_elements(31);
    -- CP-element group 31:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	30 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/type_cast_3083_update_completed_
      -- 
    -- Element group readMemoryFromL2_CP_2700_elements(31) is a control-delay.
    cp_element_31_delay: control_delay_element  generic map(name => " 31_delay", delay_value => 1)  port map(req => readMemoryFromL2_CP_2700_elements(29), ack => readMemoryFromL2_CP_2700_elements(31), clk => clk, reset =>reset);
    -- CP-element group 32:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: 	18 
    -- CP-element group 32: marked-predecessors 
    -- CP-element group 32: 	34 
    -- CP-element group 32: successors 
    -- CP-element group 32: 	34 
    -- CP-element group 32:  members (3) 
      -- CP-element group 32: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/call_stmt_3112_Sample/$entry
      -- CP-element group 32: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/call_stmt_3112_Sample/crr
      -- CP-element group 32: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/call_stmt_3112_sample_start_
      -- 
    crr_2799_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_2799_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(32), ack => call_stmt_3112_call_req_0); -- 
    readMemoryFromL2_cp_element_group_32: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_32"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readMemoryFromL2_CP_2700_elements(18) & readMemoryFromL2_CP_2700_elements(34);
      gj_readMemoryFromL2_cp_element_group_32 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(32), clk => clk, reset => reset); --
    end block;
    -- CP-element group 33:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: marked-predecessors 
    -- CP-element group 33: 	42 
    -- CP-element group 33: 	50 
    -- CP-element group 33: 	58 
    -- CP-element group 33: 	66 
    -- CP-element group 33: 	74 
    -- CP-element group 33: 	82 
    -- CP-element group 33: 	90 
    -- CP-element group 33: 	98 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (3) 
      -- CP-element group 33: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/call_stmt_3112_update_start_
      -- CP-element group 33: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/call_stmt_3112_Update/$entry
      -- CP-element group 33: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/call_stmt_3112_Update/ccr
      -- 
    ccr_2804_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_2804_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(33), ack => call_stmt_3112_call_req_1); -- 
    readMemoryFromL2_cp_element_group_33: block -- 
      constant place_capacities: IntegerArray(0 to 7) := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_markings: IntegerArray(0 to 7)  := (0 => 1,1 => 1,2 => 1,3 => 1,4 => 1,5 => 1,6 => 1,7 => 1);
      constant place_delays: IntegerArray(0 to 7) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_33"; 
      signal preds: BooleanArray(1 to 8); -- 
    begin -- 
      preds <= readMemoryFromL2_CP_2700_elements(42) & readMemoryFromL2_CP_2700_elements(50) & readMemoryFromL2_CP_2700_elements(58) & readMemoryFromL2_CP_2700_elements(66) & readMemoryFromL2_CP_2700_elements(74) & readMemoryFromL2_CP_2700_elements(82) & readMemoryFromL2_CP_2700_elements(90) & readMemoryFromL2_CP_2700_elements(98);
      gj_readMemoryFromL2_cp_element_group_33 : generic_join generic map(name => joinName, number_of_predecessors => 8, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(33), clk => clk, reset => reset); --
    end block;
    -- CP-element group 34:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	32 
    -- CP-element group 34: successors 
    -- CP-element group 34: marked-successors 
    -- CP-element group 34: 	16 
    -- CP-element group 34: 	32 
    -- CP-element group 34:  members (3) 
      -- CP-element group 34: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/call_stmt_3112_Sample/$exit
      -- CP-element group 34: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/call_stmt_3112_Sample/cra
      -- CP-element group 34: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/call_stmt_3112_sample_completed_
      -- 
    cra_2800_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 34_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_3112_call_ack_0, ack => readMemoryFromL2_CP_2700_elements(34)); -- 
    -- CP-element group 35:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	40 
    -- CP-element group 35: 	48 
    -- CP-element group 35: 	56 
    -- CP-element group 35: 	64 
    -- CP-element group 35: 	72 
    -- CP-element group 35: 	80 
    -- CP-element group 35: 	88 
    -- CP-element group 35: 	96 
    -- CP-element group 35:  members (3) 
      -- CP-element group 35: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/call_stmt_3112_update_completed_
      -- CP-element group 35: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/call_stmt_3112_Update/$exit
      -- CP-element group 35: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/call_stmt_3112_Update/cca
      -- 
    cca_2805_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 35_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_3112_call_ack_1, ack => readMemoryFromL2_CP_2700_elements(35)); -- 
    -- CP-element group 36:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	18 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	38 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	38 
    -- CP-element group 36:  members (3) 
      -- CP-element group 36: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3123_Sample/$entry
      -- CP-element group 36: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3123_Sample/req
      -- CP-element group 36: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3123_sample_start_
      -- 
    req_2813_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2813_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(36), ack => W_s0_2928_delayed_8_0_3121_inst_req_0); -- 
    readMemoryFromL2_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readMemoryFromL2_CP_2700_elements(18) & readMemoryFromL2_CP_2700_elements(38);
      gj_readMemoryFromL2_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	42 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	39 
    -- CP-element group 37:  members (3) 
      -- CP-element group 37: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3123_update_start_
      -- CP-element group 37: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3123_Update/req
      -- CP-element group 37: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3123_Update/$entry
      -- 
    req_2818_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2818_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(37), ack => W_s0_2928_delayed_8_0_3121_inst_req_1); -- 
    readMemoryFromL2_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= readMemoryFromL2_CP_2700_elements(42);
      gj_readMemoryFromL2_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	36 
    -- CP-element group 38: successors 
    -- CP-element group 38: marked-successors 
    -- CP-element group 38: 	16 
    -- CP-element group 38: 	36 
    -- CP-element group 38:  members (3) 
      -- CP-element group 38: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3123_sample_completed_
      -- CP-element group 38: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3123_Sample/$exit
      -- CP-element group 38: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3123_Sample/ack
      -- 
    ack_2814_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 38_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_s0_2928_delayed_8_0_3121_inst_ack_0, ack => readMemoryFromL2_CP_2700_elements(38)); -- 
    -- CP-element group 39:  transition  input  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: 	37 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	40 
    -- CP-element group 39:  members (3) 
      -- CP-element group 39: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3123_Update/ack
      -- CP-element group 39: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3123_Update/$exit
      -- CP-element group 39: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3123_update_completed_
      -- 
    ack_2819_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 39_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_s0_2928_delayed_8_0_3121_inst_ack_1, ack => readMemoryFromL2_CP_2700_elements(39)); -- 
    -- CP-element group 40:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	35 
    -- CP-element group 40: 	39 
    -- CP-element group 40: marked-predecessors 
    -- CP-element group 40: 	42 
    -- CP-element group 40: successors 
    -- CP-element group 40: 	42 
    -- CP-element group 40:  members (3) 
      -- CP-element group 40: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3127_sample_start_
      -- CP-element group 40: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3127_Sample/$entry
      -- CP-element group 40: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3127_Sample/req
      -- 
    req_2827_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2827_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(40), ack => W_r0_3125_inst_req_0); -- 
    readMemoryFromL2_cp_element_group_40: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_40"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= readMemoryFromL2_CP_2700_elements(35) & readMemoryFromL2_CP_2700_elements(39) & readMemoryFromL2_CP_2700_elements(42);
      gj_readMemoryFromL2_cp_element_group_40 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(40), clk => clk, reset => reset); --
    end block;
    -- CP-element group 41:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: marked-predecessors 
    -- CP-element group 41: 	43 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	43 
    -- CP-element group 41:  members (3) 
      -- CP-element group 41: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3127_update_start_
      -- CP-element group 41: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3127_Update/req
      -- CP-element group 41: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3127_Update/$entry
      -- 
    req_2832_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2832_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(41), ack => W_r0_3125_inst_req_1); -- 
    readMemoryFromL2_cp_element_group_41: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_41"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= readMemoryFromL2_CP_2700_elements(43);
      gj_readMemoryFromL2_cp_element_group_41 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(41), clk => clk, reset => reset); --
    end block;
    -- CP-element group 42:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	40 
    -- CP-element group 42: successors 
    -- CP-element group 42: marked-successors 
    -- CP-element group 42: 	33 
    -- CP-element group 42: 	37 
    -- CP-element group 42: 	40 
    -- CP-element group 42:  members (3) 
      -- CP-element group 42: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3127_Sample/ack
      -- CP-element group 42: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3127_sample_completed_
      -- CP-element group 42: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3127_Sample/$exit
      -- 
    ack_2828_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 42_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_r0_3125_inst_ack_0, ack => readMemoryFromL2_CP_2700_elements(42)); -- 
    -- CP-element group 43:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: 	41 
    -- CP-element group 43: successors 
    -- CP-element group 43: 	101 
    -- CP-element group 43: marked-successors 
    -- CP-element group 43: 	41 
    -- CP-element group 43:  members (3) 
      -- CP-element group 43: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3127_Update/$exit
      -- CP-element group 43: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3127_Update/ack
      -- CP-element group 43: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3127_update_completed_
      -- 
    ack_2833_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 43_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_r0_3125_inst_ack_1, ack => readMemoryFromL2_CP_2700_elements(43)); -- 
    -- CP-element group 44:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	18 
    -- CP-element group 44: marked-predecessors 
    -- CP-element group 44: 	46 
    -- CP-element group 44: successors 
    -- CP-element group 44: 	46 
    -- CP-element group 44:  members (3) 
      -- CP-element group 44: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3135_sample_start_
      -- CP-element group 44: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3135_Sample/req
      -- CP-element group 44: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3135_Sample/$entry
      -- 
    req_2841_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2841_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(44), ack => W_s1_2937_delayed_8_0_3133_inst_req_0); -- 
    readMemoryFromL2_cp_element_group_44: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_44"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readMemoryFromL2_CP_2700_elements(18) & readMemoryFromL2_CP_2700_elements(46);
      gj_readMemoryFromL2_cp_element_group_44 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(44), clk => clk, reset => reset); --
    end block;
    -- CP-element group 45:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: marked-predecessors 
    -- CP-element group 45: 	50 
    -- CP-element group 45: successors 
    -- CP-element group 45: 	47 
    -- CP-element group 45:  members (3) 
      -- CP-element group 45: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3135_Update/req
      -- CP-element group 45: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3135_Update/$entry
      -- CP-element group 45: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3135_update_start_
      -- 
    req_2846_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2846_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(45), ack => W_s1_2937_delayed_8_0_3133_inst_req_1); -- 
    readMemoryFromL2_cp_element_group_45: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_45"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= readMemoryFromL2_CP_2700_elements(50);
      gj_readMemoryFromL2_cp_element_group_45 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(45), clk => clk, reset => reset); --
    end block;
    -- CP-element group 46:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: 	44 
    -- CP-element group 46: successors 
    -- CP-element group 46: marked-successors 
    -- CP-element group 46: 	16 
    -- CP-element group 46: 	44 
    -- CP-element group 46:  members (3) 
      -- CP-element group 46: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3135_sample_completed_
      -- CP-element group 46: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3135_Sample/ack
      -- CP-element group 46: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3135_Sample/$exit
      -- 
    ack_2842_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_s1_2937_delayed_8_0_3133_inst_ack_0, ack => readMemoryFromL2_CP_2700_elements(46)); -- 
    -- CP-element group 47:  transition  input  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: 	45 
    -- CP-element group 47: successors 
    -- CP-element group 47: 	48 
    -- CP-element group 47:  members (3) 
      -- CP-element group 47: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3135_Update/ack
      -- CP-element group 47: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3135_Update/$exit
      -- CP-element group 47: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3135_update_completed_
      -- 
    ack_2847_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 47_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_s1_2937_delayed_8_0_3133_inst_ack_1, ack => readMemoryFromL2_CP_2700_elements(47)); -- 
    -- CP-element group 48:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: 	35 
    -- CP-element group 48: 	47 
    -- CP-element group 48: marked-predecessors 
    -- CP-element group 48: 	50 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (3) 
      -- CP-element group 48: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3139_Sample/$entry
      -- CP-element group 48: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3139_sample_start_
      -- CP-element group 48: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3139_Sample/req
      -- 
    req_2855_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2855_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(48), ack => W_r1_3137_inst_req_0); -- 
    readMemoryFromL2_cp_element_group_48: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_48"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= readMemoryFromL2_CP_2700_elements(35) & readMemoryFromL2_CP_2700_elements(47) & readMemoryFromL2_CP_2700_elements(50);
      gj_readMemoryFromL2_cp_element_group_48 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(48), clk => clk, reset => reset); --
    end block;
    -- CP-element group 49:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: marked-predecessors 
    -- CP-element group 49: 	51 
    -- CP-element group 49: successors 
    -- CP-element group 49: 	51 
    -- CP-element group 49:  members (3) 
      -- CP-element group 49: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3139_update_start_
      -- CP-element group 49: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3139_Update/req
      -- CP-element group 49: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3139_Update/$entry
      -- 
    req_2860_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2860_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(49), ack => W_r1_3137_inst_req_1); -- 
    readMemoryFromL2_cp_element_group_49: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_49"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= readMemoryFromL2_CP_2700_elements(51);
      gj_readMemoryFromL2_cp_element_group_49 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(49), clk => clk, reset => reset); --
    end block;
    -- CP-element group 50:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50: marked-successors 
    -- CP-element group 50: 	33 
    -- CP-element group 50: 	45 
    -- CP-element group 50: 	48 
    -- CP-element group 50:  members (3) 
      -- CP-element group 50: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3139_sample_completed_
      -- CP-element group 50: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3139_Sample/ack
      -- CP-element group 50: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3139_Sample/$exit
      -- 
    ack_2856_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 50_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_r1_3137_inst_ack_0, ack => readMemoryFromL2_CP_2700_elements(50)); -- 
    -- CP-element group 51:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: 	49 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	101 
    -- CP-element group 51: marked-successors 
    -- CP-element group 51: 	49 
    -- CP-element group 51:  members (3) 
      -- CP-element group 51: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3139_Update/$exit
      -- CP-element group 51: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3139_update_completed_
      -- CP-element group 51: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3139_Update/ack
      -- 
    ack_2861_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 51_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_r1_3137_inst_ack_1, ack => readMemoryFromL2_CP_2700_elements(51)); -- 
    -- CP-element group 52:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: 	18 
    -- CP-element group 52: marked-predecessors 
    -- CP-element group 52: 	54 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (3) 
      -- CP-element group 52: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3147_Sample/$entry
      -- CP-element group 52: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3147_sample_start_
      -- CP-element group 52: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3147_Sample/req
      -- 
    req_2869_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2869_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(52), ack => W_s2_2946_delayed_8_0_3145_inst_req_0); -- 
    readMemoryFromL2_cp_element_group_52: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_52"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readMemoryFromL2_CP_2700_elements(18) & readMemoryFromL2_CP_2700_elements(54);
      gj_readMemoryFromL2_cp_element_group_52 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(52), clk => clk, reset => reset); --
    end block;
    -- CP-element group 53:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: marked-predecessors 
    -- CP-element group 53: 	58 
    -- CP-element group 53: successors 
    -- CP-element group 53: 	55 
    -- CP-element group 53:  members (3) 
      -- CP-element group 53: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3147_update_start_
      -- CP-element group 53: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3147_Update/req
      -- CP-element group 53: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3147_Update/$entry
      -- 
    req_2874_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2874_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(53), ack => W_s2_2946_delayed_8_0_3145_inst_req_1); -- 
    readMemoryFromL2_cp_element_group_53: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_53"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= readMemoryFromL2_CP_2700_elements(58);
      gj_readMemoryFromL2_cp_element_group_53 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(53), clk => clk, reset => reset); --
    end block;
    -- CP-element group 54:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54: marked-successors 
    -- CP-element group 54: 	16 
    -- CP-element group 54: 	52 
    -- CP-element group 54:  members (3) 
      -- CP-element group 54: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3147_Sample/$exit
      -- CP-element group 54: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3147_sample_completed_
      -- CP-element group 54: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3147_Sample/ack
      -- 
    ack_2870_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_s2_2946_delayed_8_0_3145_inst_ack_0, ack => readMemoryFromL2_CP_2700_elements(54)); -- 
    -- CP-element group 55:  transition  input  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	53 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	56 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3147_update_completed_
      -- CP-element group 55: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3147_Update/ack
      -- CP-element group 55: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3147_Update/$exit
      -- 
    ack_2875_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 55_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_s2_2946_delayed_8_0_3145_inst_ack_1, ack => readMemoryFromL2_CP_2700_elements(55)); -- 
    -- CP-element group 56:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: 	35 
    -- CP-element group 56: 	55 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	58 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3151_Sample/req
      -- CP-element group 56: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3151_Sample/$entry
      -- CP-element group 56: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3151_sample_start_
      -- 
    req_2883_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2883_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(56), ack => W_r2_3149_inst_req_0); -- 
    readMemoryFromL2_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= readMemoryFromL2_CP_2700_elements(35) & readMemoryFromL2_CP_2700_elements(55) & readMemoryFromL2_CP_2700_elements(58);
      gj_readMemoryFromL2_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: marked-predecessors 
    -- CP-element group 57: 	59 
    -- CP-element group 57: successors 
    -- CP-element group 57: 	59 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3151_Update/req
      -- CP-element group 57: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3151_Update/$entry
      -- CP-element group 57: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3151_update_start_
      -- 
    req_2888_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2888_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(57), ack => W_r2_3149_inst_req_1); -- 
    readMemoryFromL2_cp_element_group_57: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_57"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= readMemoryFromL2_CP_2700_elements(59);
      gj_readMemoryFromL2_cp_element_group_57 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(57), clk => clk, reset => reset); --
    end block;
    -- CP-element group 58:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	33 
    -- CP-element group 58: 	53 
    -- CP-element group 58: 	56 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3151_Sample/ack
      -- CP-element group 58: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3151_Sample/$exit
      -- CP-element group 58: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3151_sample_completed_
      -- 
    ack_2884_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_r2_3149_inst_ack_0, ack => readMemoryFromL2_CP_2700_elements(58)); -- 
    -- CP-element group 59:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	57 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	101 
    -- CP-element group 59: marked-successors 
    -- CP-element group 59: 	57 
    -- CP-element group 59:  members (3) 
      -- CP-element group 59: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3151_Update/ack
      -- CP-element group 59: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3151_Update/$exit
      -- CP-element group 59: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3151_update_completed_
      -- 
    ack_2889_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 59_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_r2_3149_inst_ack_1, ack => readMemoryFromL2_CP_2700_elements(59)); -- 
    -- CP-element group 60:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	18 
    -- CP-element group 60: marked-predecessors 
    -- CP-element group 60: 	62 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	62 
    -- CP-element group 60:  members (3) 
      -- CP-element group 60: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3159_sample_start_
      -- CP-element group 60: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3159_Sample/req
      -- CP-element group 60: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3159_Sample/$entry
      -- 
    req_2897_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2897_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(60), ack => W_s3_2955_delayed_8_0_3157_inst_req_0); -- 
    readMemoryFromL2_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readMemoryFromL2_CP_2700_elements(18) & readMemoryFromL2_CP_2700_elements(62);
      gj_readMemoryFromL2_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: marked-predecessors 
    -- CP-element group 61: 	66 
    -- CP-element group 61: successors 
    -- CP-element group 61: 	63 
    -- CP-element group 61:  members (3) 
      -- CP-element group 61: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3159_update_start_
      -- CP-element group 61: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3159_Update/req
      -- CP-element group 61: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3159_Update/$entry
      -- 
    req_2902_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2902_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(61), ack => W_s3_2955_delayed_8_0_3157_inst_req_1); -- 
    readMemoryFromL2_cp_element_group_61: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_61"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= readMemoryFromL2_CP_2700_elements(66);
      gj_readMemoryFromL2_cp_element_group_61 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(61), clk => clk, reset => reset); --
    end block;
    -- CP-element group 62:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	60 
    -- CP-element group 62: successors 
    -- CP-element group 62: marked-successors 
    -- CP-element group 62: 	16 
    -- CP-element group 62: 	60 
    -- CP-element group 62:  members (3) 
      -- CP-element group 62: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3159_sample_completed_
      -- CP-element group 62: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3159_Sample/ack
      -- CP-element group 62: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3159_Sample/$exit
      -- 
    ack_2898_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_s3_2955_delayed_8_0_3157_inst_ack_0, ack => readMemoryFromL2_CP_2700_elements(62)); -- 
    -- CP-element group 63:  transition  input  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	61 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	64 
    -- CP-element group 63:  members (3) 
      -- CP-element group 63: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3159_update_completed_
      -- CP-element group 63: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3159_Update/ack
      -- CP-element group 63: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3159_Update/$exit
      -- 
    ack_2903_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 63_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_s3_2955_delayed_8_0_3157_inst_ack_1, ack => readMemoryFromL2_CP_2700_elements(63)); -- 
    -- CP-element group 64:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	35 
    -- CP-element group 64: 	63 
    -- CP-element group 64: marked-predecessors 
    -- CP-element group 64: 	66 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	66 
    -- CP-element group 64:  members (3) 
      -- CP-element group 64: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3163_Sample/req
      -- CP-element group 64: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3163_Sample/$entry
      -- CP-element group 64: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3163_sample_start_
      -- 
    req_2911_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2911_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(64), ack => W_r3_3161_inst_req_0); -- 
    readMemoryFromL2_cp_element_group_64: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_64"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= readMemoryFromL2_CP_2700_elements(35) & readMemoryFromL2_CP_2700_elements(63) & readMemoryFromL2_CP_2700_elements(66);
      gj_readMemoryFromL2_cp_element_group_64 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(64), clk => clk, reset => reset); --
    end block;
    -- CP-element group 65:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: marked-predecessors 
    -- CP-element group 65: 	67 
    -- CP-element group 65: successors 
    -- CP-element group 65: 	67 
    -- CP-element group 65:  members (3) 
      -- CP-element group 65: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3163_Update/req
      -- CP-element group 65: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3163_Update/$entry
      -- CP-element group 65: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3163_update_start_
      -- 
    req_2916_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2916_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(65), ack => W_r3_3161_inst_req_1); -- 
    readMemoryFromL2_cp_element_group_65: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_65"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= readMemoryFromL2_CP_2700_elements(67);
      gj_readMemoryFromL2_cp_element_group_65 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(65), clk => clk, reset => reset); --
    end block;
    -- CP-element group 66:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 66: predecessors 
    -- CP-element group 66: 	64 
    -- CP-element group 66: successors 
    -- CP-element group 66: marked-successors 
    -- CP-element group 66: 	33 
    -- CP-element group 66: 	61 
    -- CP-element group 66: 	64 
    -- CP-element group 66:  members (3) 
      -- CP-element group 66: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3163_Sample/ack
      -- CP-element group 66: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3163_Sample/$exit
      -- CP-element group 66: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3163_sample_completed_
      -- 
    ack_2912_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 66_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_r3_3161_inst_ack_0, ack => readMemoryFromL2_CP_2700_elements(66)); -- 
    -- CP-element group 67:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 67: predecessors 
    -- CP-element group 67: 	65 
    -- CP-element group 67: successors 
    -- CP-element group 67: 	101 
    -- CP-element group 67: marked-successors 
    -- CP-element group 67: 	65 
    -- CP-element group 67:  members (3) 
      -- CP-element group 67: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3163_Update/ack
      -- CP-element group 67: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3163_Update/$exit
      -- CP-element group 67: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3163_update_completed_
      -- 
    ack_2917_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 67_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_r3_3161_inst_ack_1, ack => readMemoryFromL2_CP_2700_elements(67)); -- 
    -- CP-element group 68:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 68: predecessors 
    -- CP-element group 68: 	18 
    -- CP-element group 68: marked-predecessors 
    -- CP-element group 68: 	70 
    -- CP-element group 68: successors 
    -- CP-element group 68: 	70 
    -- CP-element group 68:  members (3) 
      -- CP-element group 68: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3171_Sample/req
      -- CP-element group 68: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3171_Sample/$entry
      -- CP-element group 68: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3171_sample_start_
      -- 
    req_2925_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2925_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(68), ack => W_s4_2964_delayed_8_0_3169_inst_req_0); -- 
    readMemoryFromL2_cp_element_group_68: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_68"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readMemoryFromL2_CP_2700_elements(18) & readMemoryFromL2_CP_2700_elements(70);
      gj_readMemoryFromL2_cp_element_group_68 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(68), clk => clk, reset => reset); --
    end block;
    -- CP-element group 69:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 69: predecessors 
    -- CP-element group 69: marked-predecessors 
    -- CP-element group 69: 	74 
    -- CP-element group 69: successors 
    -- CP-element group 69: 	71 
    -- CP-element group 69:  members (3) 
      -- CP-element group 69: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3171_update_start_
      -- CP-element group 69: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3171_Update/$entry
      -- CP-element group 69: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3171_Update/req
      -- 
    req_2930_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2930_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(69), ack => W_s4_2964_delayed_8_0_3169_inst_req_1); -- 
    readMemoryFromL2_cp_element_group_69: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_69"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= readMemoryFromL2_CP_2700_elements(74);
      gj_readMemoryFromL2_cp_element_group_69 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(69), clk => clk, reset => reset); --
    end block;
    -- CP-element group 70:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 70: predecessors 
    -- CP-element group 70: 	68 
    -- CP-element group 70: successors 
    -- CP-element group 70: marked-successors 
    -- CP-element group 70: 	16 
    -- CP-element group 70: 	68 
    -- CP-element group 70:  members (3) 
      -- CP-element group 70: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3171_Sample/ack
      -- CP-element group 70: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3171_Sample/$exit
      -- CP-element group 70: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3171_sample_completed_
      -- 
    ack_2926_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 70_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_s4_2964_delayed_8_0_3169_inst_ack_0, ack => readMemoryFromL2_CP_2700_elements(70)); -- 
    -- CP-element group 71:  transition  input  bypass  pipeline-parent 
    -- CP-element group 71: predecessors 
    -- CP-element group 71: 	69 
    -- CP-element group 71: successors 
    -- CP-element group 71: 	72 
    -- CP-element group 71:  members (3) 
      -- CP-element group 71: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3171_update_completed_
      -- CP-element group 71: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3171_Update/$exit
      -- CP-element group 71: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3171_Update/ack
      -- 
    ack_2931_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 71_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_s4_2964_delayed_8_0_3169_inst_ack_1, ack => readMemoryFromL2_CP_2700_elements(71)); -- 
    -- CP-element group 72:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 72: predecessors 
    -- CP-element group 72: 	35 
    -- CP-element group 72: 	71 
    -- CP-element group 72: marked-predecessors 
    -- CP-element group 72: 	74 
    -- CP-element group 72: successors 
    -- CP-element group 72: 	74 
    -- CP-element group 72:  members (3) 
      -- CP-element group 72: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3175_Sample/$entry
      -- CP-element group 72: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3175_sample_start_
      -- CP-element group 72: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3175_Sample/req
      -- 
    req_2939_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2939_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(72), ack => W_r4_3173_inst_req_0); -- 
    readMemoryFromL2_cp_element_group_72: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_72"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= readMemoryFromL2_CP_2700_elements(35) & readMemoryFromL2_CP_2700_elements(71) & readMemoryFromL2_CP_2700_elements(74);
      gj_readMemoryFromL2_cp_element_group_72 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(72), clk => clk, reset => reset); --
    end block;
    -- CP-element group 73:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 73: predecessors 
    -- CP-element group 73: marked-predecessors 
    -- CP-element group 73: 	75 
    -- CP-element group 73: successors 
    -- CP-element group 73: 	75 
    -- CP-element group 73:  members (3) 
      -- CP-element group 73: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3175_update_start_
      -- CP-element group 73: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3175_Update/$entry
      -- CP-element group 73: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3175_Update/req
      -- 
    req_2944_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2944_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(73), ack => W_r4_3173_inst_req_1); -- 
    readMemoryFromL2_cp_element_group_73: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_73"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= readMemoryFromL2_CP_2700_elements(75);
      gj_readMemoryFromL2_cp_element_group_73 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(73), clk => clk, reset => reset); --
    end block;
    -- CP-element group 74:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 74: predecessors 
    -- CP-element group 74: 	72 
    -- CP-element group 74: successors 
    -- CP-element group 74: marked-successors 
    -- CP-element group 74: 	33 
    -- CP-element group 74: 	69 
    -- CP-element group 74: 	72 
    -- CP-element group 74:  members (3) 
      -- CP-element group 74: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3175_sample_completed_
      -- CP-element group 74: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3175_Sample/$exit
      -- CP-element group 74: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3175_Sample/ack
      -- 
    ack_2940_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 74_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_r4_3173_inst_ack_0, ack => readMemoryFromL2_CP_2700_elements(74)); -- 
    -- CP-element group 75:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 75: predecessors 
    -- CP-element group 75: 	73 
    -- CP-element group 75: successors 
    -- CP-element group 75: 	101 
    -- CP-element group 75: marked-successors 
    -- CP-element group 75: 	73 
    -- CP-element group 75:  members (3) 
      -- CP-element group 75: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3175_update_completed_
      -- CP-element group 75: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3175_Update/$exit
      -- CP-element group 75: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3175_Update/ack
      -- 
    ack_2945_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 75_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_r4_3173_inst_ack_1, ack => readMemoryFromL2_CP_2700_elements(75)); -- 
    -- CP-element group 76:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 76: predecessors 
    -- CP-element group 76: 	18 
    -- CP-element group 76: marked-predecessors 
    -- CP-element group 76: 	78 
    -- CP-element group 76: successors 
    -- CP-element group 76: 	78 
    -- CP-element group 76:  members (3) 
      -- CP-element group 76: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3183_sample_start_
      -- CP-element group 76: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3183_Sample/$entry
      -- CP-element group 76: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3183_Sample/req
      -- 
    req_2953_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2953_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(76), ack => W_s5_2973_delayed_8_0_3181_inst_req_0); -- 
    readMemoryFromL2_cp_element_group_76: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_76"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readMemoryFromL2_CP_2700_elements(18) & readMemoryFromL2_CP_2700_elements(78);
      gj_readMemoryFromL2_cp_element_group_76 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(76), clk => clk, reset => reset); --
    end block;
    -- CP-element group 77:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 77: predecessors 
    -- CP-element group 77: marked-predecessors 
    -- CP-element group 77: 	82 
    -- CP-element group 77: successors 
    -- CP-element group 77: 	79 
    -- CP-element group 77:  members (3) 
      -- CP-element group 77: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3183_update_start_
      -- CP-element group 77: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3183_Update/$entry
      -- CP-element group 77: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3183_Update/req
      -- 
    req_2958_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2958_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(77), ack => W_s5_2973_delayed_8_0_3181_inst_req_1); -- 
    readMemoryFromL2_cp_element_group_77: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_77"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= readMemoryFromL2_CP_2700_elements(82);
      gj_readMemoryFromL2_cp_element_group_77 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(77), clk => clk, reset => reset); --
    end block;
    -- CP-element group 78:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 78: predecessors 
    -- CP-element group 78: 	76 
    -- CP-element group 78: successors 
    -- CP-element group 78: marked-successors 
    -- CP-element group 78: 	16 
    -- CP-element group 78: 	76 
    -- CP-element group 78:  members (3) 
      -- CP-element group 78: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3183_sample_completed_
      -- CP-element group 78: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3183_Sample/$exit
      -- CP-element group 78: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3183_Sample/ack
      -- 
    ack_2954_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 78_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_s5_2973_delayed_8_0_3181_inst_ack_0, ack => readMemoryFromL2_CP_2700_elements(78)); -- 
    -- CP-element group 79:  transition  input  bypass  pipeline-parent 
    -- CP-element group 79: predecessors 
    -- CP-element group 79: 	77 
    -- CP-element group 79: successors 
    -- CP-element group 79: 	80 
    -- CP-element group 79:  members (3) 
      -- CP-element group 79: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3183_update_completed_
      -- CP-element group 79: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3183_Update/$exit
      -- CP-element group 79: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3183_Update/ack
      -- 
    ack_2959_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 79_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_s5_2973_delayed_8_0_3181_inst_ack_1, ack => readMemoryFromL2_CP_2700_elements(79)); -- 
    -- CP-element group 80:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 80: predecessors 
    -- CP-element group 80: 	35 
    -- CP-element group 80: 	79 
    -- CP-element group 80: marked-predecessors 
    -- CP-element group 80: 	82 
    -- CP-element group 80: successors 
    -- CP-element group 80: 	82 
    -- CP-element group 80:  members (3) 
      -- CP-element group 80: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3187_sample_start_
      -- CP-element group 80: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3187_Sample/$entry
      -- CP-element group 80: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3187_Sample/req
      -- 
    req_2967_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2967_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(80), ack => W_r5_3185_inst_req_0); -- 
    readMemoryFromL2_cp_element_group_80: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_80"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= readMemoryFromL2_CP_2700_elements(35) & readMemoryFromL2_CP_2700_elements(79) & readMemoryFromL2_CP_2700_elements(82);
      gj_readMemoryFromL2_cp_element_group_80 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(80), clk => clk, reset => reset); --
    end block;
    -- CP-element group 81:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 81: predecessors 
    -- CP-element group 81: marked-predecessors 
    -- CP-element group 81: 	83 
    -- CP-element group 81: successors 
    -- CP-element group 81: 	83 
    -- CP-element group 81:  members (3) 
      -- CP-element group 81: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3187_update_start_
      -- CP-element group 81: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3187_Update/$entry
      -- CP-element group 81: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3187_Update/req
      -- 
    req_2972_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2972_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(81), ack => W_r5_3185_inst_req_1); -- 
    readMemoryFromL2_cp_element_group_81: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_81"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= readMemoryFromL2_CP_2700_elements(83);
      gj_readMemoryFromL2_cp_element_group_81 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(81), clk => clk, reset => reset); --
    end block;
    -- CP-element group 82:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 82: predecessors 
    -- CP-element group 82: 	80 
    -- CP-element group 82: successors 
    -- CP-element group 82: marked-successors 
    -- CP-element group 82: 	33 
    -- CP-element group 82: 	77 
    -- CP-element group 82: 	80 
    -- CP-element group 82:  members (3) 
      -- CP-element group 82: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3187_sample_completed_
      -- CP-element group 82: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3187_Sample/$exit
      -- CP-element group 82: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3187_Sample/ack
      -- 
    ack_2968_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 82_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_r5_3185_inst_ack_0, ack => readMemoryFromL2_CP_2700_elements(82)); -- 
    -- CP-element group 83:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 83: predecessors 
    -- CP-element group 83: 	81 
    -- CP-element group 83: successors 
    -- CP-element group 83: 	101 
    -- CP-element group 83: marked-successors 
    -- CP-element group 83: 	81 
    -- CP-element group 83:  members (3) 
      -- CP-element group 83: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3187_update_completed_
      -- CP-element group 83: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3187_Update/$exit
      -- CP-element group 83: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3187_Update/ack
      -- 
    ack_2973_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 83_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_r5_3185_inst_ack_1, ack => readMemoryFromL2_CP_2700_elements(83)); -- 
    -- CP-element group 84:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 84: predecessors 
    -- CP-element group 84: 	18 
    -- CP-element group 84: marked-predecessors 
    -- CP-element group 84: 	86 
    -- CP-element group 84: successors 
    -- CP-element group 84: 	86 
    -- CP-element group 84:  members (3) 
      -- CP-element group 84: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3195_sample_start_
      -- CP-element group 84: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3195_Sample/$entry
      -- CP-element group 84: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3195_Sample/req
      -- 
    req_2981_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2981_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(84), ack => W_s6_2982_delayed_8_0_3193_inst_req_0); -- 
    readMemoryFromL2_cp_element_group_84: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_84"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readMemoryFromL2_CP_2700_elements(18) & readMemoryFromL2_CP_2700_elements(86);
      gj_readMemoryFromL2_cp_element_group_84 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(84), clk => clk, reset => reset); --
    end block;
    -- CP-element group 85:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 85: predecessors 
    -- CP-element group 85: marked-predecessors 
    -- CP-element group 85: 	90 
    -- CP-element group 85: successors 
    -- CP-element group 85: 	87 
    -- CP-element group 85:  members (3) 
      -- CP-element group 85: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3195_update_start_
      -- CP-element group 85: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3195_Update/$entry
      -- CP-element group 85: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3195_Update/req
      -- 
    req_2986_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2986_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(85), ack => W_s6_2982_delayed_8_0_3193_inst_req_1); -- 
    readMemoryFromL2_cp_element_group_85: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_85"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= readMemoryFromL2_CP_2700_elements(90);
      gj_readMemoryFromL2_cp_element_group_85 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(85), clk => clk, reset => reset); --
    end block;
    -- CP-element group 86:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 86: predecessors 
    -- CP-element group 86: 	84 
    -- CP-element group 86: successors 
    -- CP-element group 86: marked-successors 
    -- CP-element group 86: 	16 
    -- CP-element group 86: 	84 
    -- CP-element group 86:  members (3) 
      -- CP-element group 86: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3195_sample_completed_
      -- CP-element group 86: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3195_Sample/$exit
      -- CP-element group 86: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3195_Sample/ack
      -- 
    ack_2982_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 86_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_s6_2982_delayed_8_0_3193_inst_ack_0, ack => readMemoryFromL2_CP_2700_elements(86)); -- 
    -- CP-element group 87:  transition  input  bypass  pipeline-parent 
    -- CP-element group 87: predecessors 
    -- CP-element group 87: 	85 
    -- CP-element group 87: successors 
    -- CP-element group 87: 	88 
    -- CP-element group 87:  members (3) 
      -- CP-element group 87: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3195_update_completed_
      -- CP-element group 87: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3195_Update/$exit
      -- CP-element group 87: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3195_Update/ack
      -- 
    ack_2987_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 87_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_s6_2982_delayed_8_0_3193_inst_ack_1, ack => readMemoryFromL2_CP_2700_elements(87)); -- 
    -- CP-element group 88:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 88: predecessors 
    -- CP-element group 88: 	35 
    -- CP-element group 88: 	87 
    -- CP-element group 88: marked-predecessors 
    -- CP-element group 88: 	90 
    -- CP-element group 88: successors 
    -- CP-element group 88: 	90 
    -- CP-element group 88:  members (3) 
      -- CP-element group 88: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3199_sample_start_
      -- CP-element group 88: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3199_Sample/$entry
      -- CP-element group 88: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3199_Sample/req
      -- 
    req_2995_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_2995_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(88), ack => W_r6_3197_inst_req_0); -- 
    readMemoryFromL2_cp_element_group_88: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_88"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= readMemoryFromL2_CP_2700_elements(35) & readMemoryFromL2_CP_2700_elements(87) & readMemoryFromL2_CP_2700_elements(90);
      gj_readMemoryFromL2_cp_element_group_88 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(88), clk => clk, reset => reset); --
    end block;
    -- CP-element group 89:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 89: predecessors 
    -- CP-element group 89: marked-predecessors 
    -- CP-element group 89: 	91 
    -- CP-element group 89: successors 
    -- CP-element group 89: 	91 
    -- CP-element group 89:  members (3) 
      -- CP-element group 89: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3199_update_start_
      -- CP-element group 89: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3199_Update/$entry
      -- CP-element group 89: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3199_Update/req
      -- 
    req_3000_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3000_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(89), ack => W_r6_3197_inst_req_1); -- 
    readMemoryFromL2_cp_element_group_89: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_89"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= readMemoryFromL2_CP_2700_elements(91);
      gj_readMemoryFromL2_cp_element_group_89 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(89), clk => clk, reset => reset); --
    end block;
    -- CP-element group 90:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 90: predecessors 
    -- CP-element group 90: 	88 
    -- CP-element group 90: successors 
    -- CP-element group 90: marked-successors 
    -- CP-element group 90: 	33 
    -- CP-element group 90: 	85 
    -- CP-element group 90: 	88 
    -- CP-element group 90:  members (3) 
      -- CP-element group 90: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3199_sample_completed_
      -- CP-element group 90: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3199_Sample/$exit
      -- CP-element group 90: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3199_Sample/ack
      -- 
    ack_2996_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 90_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_r6_3197_inst_ack_0, ack => readMemoryFromL2_CP_2700_elements(90)); -- 
    -- CP-element group 91:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 91: predecessors 
    -- CP-element group 91: 	89 
    -- CP-element group 91: successors 
    -- CP-element group 91: 	101 
    -- CP-element group 91: marked-successors 
    -- CP-element group 91: 	89 
    -- CP-element group 91:  members (3) 
      -- CP-element group 91: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3199_update_completed_
      -- CP-element group 91: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3199_Update/$exit
      -- CP-element group 91: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3199_Update/ack
      -- 
    ack_3001_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 91_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_r6_3197_inst_ack_1, ack => readMemoryFromL2_CP_2700_elements(91)); -- 
    -- CP-element group 92:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 92: predecessors 
    -- CP-element group 92: 	18 
    -- CP-element group 92: marked-predecessors 
    -- CP-element group 92: 	94 
    -- CP-element group 92: successors 
    -- CP-element group 92: 	94 
    -- CP-element group 92:  members (3) 
      -- CP-element group 92: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3207_sample_start_
      -- CP-element group 92: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3207_Sample/$entry
      -- CP-element group 92: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3207_Sample/req
      -- 
    req_3009_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3009_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(92), ack => W_s7_2991_delayed_8_0_3205_inst_req_0); -- 
    readMemoryFromL2_cp_element_group_92: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_92"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= readMemoryFromL2_CP_2700_elements(18) & readMemoryFromL2_CP_2700_elements(94);
      gj_readMemoryFromL2_cp_element_group_92 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(92), clk => clk, reset => reset); --
    end block;
    -- CP-element group 93:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 93: predecessors 
    -- CP-element group 93: marked-predecessors 
    -- CP-element group 93: 	98 
    -- CP-element group 93: successors 
    -- CP-element group 93: 	95 
    -- CP-element group 93:  members (3) 
      -- CP-element group 93: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3207_update_start_
      -- CP-element group 93: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3207_Update/$entry
      -- CP-element group 93: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3207_Update/req
      -- 
    req_3014_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3014_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(93), ack => W_s7_2991_delayed_8_0_3205_inst_req_1); -- 
    readMemoryFromL2_cp_element_group_93: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_93"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= readMemoryFromL2_CP_2700_elements(98);
      gj_readMemoryFromL2_cp_element_group_93 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(93), clk => clk, reset => reset); --
    end block;
    -- CP-element group 94:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 94: predecessors 
    -- CP-element group 94: 	92 
    -- CP-element group 94: successors 
    -- CP-element group 94: marked-successors 
    -- CP-element group 94: 	16 
    -- CP-element group 94: 	92 
    -- CP-element group 94:  members (3) 
      -- CP-element group 94: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3207_sample_completed_
      -- CP-element group 94: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3207_Sample/$exit
      -- CP-element group 94: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3207_Sample/ack
      -- 
    ack_3010_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 94_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_s7_2991_delayed_8_0_3205_inst_ack_0, ack => readMemoryFromL2_CP_2700_elements(94)); -- 
    -- CP-element group 95:  transition  input  bypass  pipeline-parent 
    -- CP-element group 95: predecessors 
    -- CP-element group 95: 	93 
    -- CP-element group 95: successors 
    -- CP-element group 95: 	96 
    -- CP-element group 95:  members (3) 
      -- CP-element group 95: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3207_update_completed_
      -- CP-element group 95: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3207_Update/$exit
      -- CP-element group 95: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3207_Update/ack
      -- 
    ack_3015_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 95_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_s7_2991_delayed_8_0_3205_inst_ack_1, ack => readMemoryFromL2_CP_2700_elements(95)); -- 
    -- CP-element group 96:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 96: predecessors 
    -- CP-element group 96: 	35 
    -- CP-element group 96: 	95 
    -- CP-element group 96: marked-predecessors 
    -- CP-element group 96: 	98 
    -- CP-element group 96: successors 
    -- CP-element group 96: 	98 
    -- CP-element group 96:  members (3) 
      -- CP-element group 96: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3211_sample_start_
      -- CP-element group 96: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3211_Sample/$entry
      -- CP-element group 96: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3211_Sample/req
      -- 
    req_3023_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3023_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(96), ack => W_r7_3209_inst_req_0); -- 
    readMemoryFromL2_cp_element_group_96: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_96"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= readMemoryFromL2_CP_2700_elements(35) & readMemoryFromL2_CP_2700_elements(95) & readMemoryFromL2_CP_2700_elements(98);
      gj_readMemoryFromL2_cp_element_group_96 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(96), clk => clk, reset => reset); --
    end block;
    -- CP-element group 97:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 97: predecessors 
    -- CP-element group 97: marked-predecessors 
    -- CP-element group 97: 	99 
    -- CP-element group 97: successors 
    -- CP-element group 97: 	99 
    -- CP-element group 97:  members (3) 
      -- CP-element group 97: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3211_update_start_
      -- CP-element group 97: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3211_Update/$entry
      -- CP-element group 97: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3211_Update/req
      -- 
    req_3028_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3028_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => readMemoryFromL2_CP_2700_elements(97), ack => W_r7_3209_inst_req_1); -- 
    readMemoryFromL2_cp_element_group_97: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 36) := "readMemoryFromL2_cp_element_group_97"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= readMemoryFromL2_CP_2700_elements(99);
      gj_readMemoryFromL2_cp_element_group_97 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(97), clk => clk, reset => reset); --
    end block;
    -- CP-element group 98:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 98: predecessors 
    -- CP-element group 98: 	96 
    -- CP-element group 98: successors 
    -- CP-element group 98: marked-successors 
    -- CP-element group 98: 	33 
    -- CP-element group 98: 	93 
    -- CP-element group 98: 	96 
    -- CP-element group 98:  members (3) 
      -- CP-element group 98: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3211_sample_completed_
      -- CP-element group 98: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3211_Sample/$exit
      -- CP-element group 98: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3211_Sample/ack
      -- 
    ack_3024_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 98_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_r7_3209_inst_ack_0, ack => readMemoryFromL2_CP_2700_elements(98)); -- 
    -- CP-element group 99:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 99: predecessors 
    -- CP-element group 99: 	97 
    -- CP-element group 99: successors 
    -- CP-element group 99: 	101 
    -- CP-element group 99: marked-successors 
    -- CP-element group 99: 	97 
    -- CP-element group 99:  members (3) 
      -- CP-element group 99: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3211_update_completed_
      -- CP-element group 99: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3211_Update/$exit
      -- CP-element group 99: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/assign_stmt_3211_Update/ack
      -- 
    ack_3029_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 99_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => W_r7_3209_inst_ack_1, ack => readMemoryFromL2_CP_2700_elements(99)); -- 
    -- CP-element group 100:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 100: predecessors 
    -- CP-element group 100: 	11 
    -- CP-element group 100: successors 
    -- CP-element group 100: 	12 
    -- CP-element group 100:  members (1) 
      -- CP-element group 100: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group readMemoryFromL2_CP_2700_elements(100) is a control-delay.
    cp_element_100_delay: control_delay_element  generic map(name => " 100_delay", delay_value => 1)  port map(req => readMemoryFromL2_CP_2700_elements(11), ack => readMemoryFromL2_CP_2700_elements(100), clk => clk, reset =>reset);
    -- CP-element group 101:  join  transition  bypass  pipeline-parent 
    -- CP-element group 101: predecessors 
    -- CP-element group 101: 	17 
    -- CP-element group 101: 	43 
    -- CP-element group 101: 	51 
    -- CP-element group 101: 	59 
    -- CP-element group 101: 	67 
    -- CP-element group 101: 	75 
    -- CP-element group 101: 	83 
    -- CP-element group 101: 	91 
    -- CP-element group 101: 	99 
    -- CP-element group 101: successors 
    -- CP-element group 101: 	8 
    -- CP-element group 101:  members (1) 
      -- CP-element group 101: 	 branch_block_stmt_3076/do_while_stmt_3077/do_while_stmt_3077_loop_body/$exit
      -- 
    readMemoryFromL2_cp_element_group_101: block -- 
      constant place_capacities: IntegerArray(0 to 8) := (0 => 15,1 => 15,2 => 15,3 => 15,4 => 15,5 => 15,6 => 15,7 => 15,8 => 15);
      constant place_markings: IntegerArray(0 to 8)  := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant place_delays: IntegerArray(0 to 8) := (0 => 0,1 => 0,2 => 0,3 => 0,4 => 0,5 => 0,6 => 0,7 => 0,8 => 0);
      constant joinName: string(1 to 37) := "readMemoryFromL2_cp_element_group_101"; 
      signal preds: BooleanArray(1 to 9); -- 
    begin -- 
      preds <= readMemoryFromL2_CP_2700_elements(17) & readMemoryFromL2_CP_2700_elements(43) & readMemoryFromL2_CP_2700_elements(51) & readMemoryFromL2_CP_2700_elements(59) & readMemoryFromL2_CP_2700_elements(67) & readMemoryFromL2_CP_2700_elements(75) & readMemoryFromL2_CP_2700_elements(83) & readMemoryFromL2_CP_2700_elements(91) & readMemoryFromL2_CP_2700_elements(99);
      gj_readMemoryFromL2_cp_element_group_101 : generic_join generic map(name => joinName, number_of_predecessors => 9, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(101), clk => clk, reset => reset); --
    end block;
    -- CP-element group 102:  transition  input  bypass  pipeline-parent 
    -- CP-element group 102: predecessors 
    -- CP-element group 102: 	7 
    -- CP-element group 102: successors 
    -- CP-element group 102:  members (2) 
      -- CP-element group 102: 	 branch_block_stmt_3076/do_while_stmt_3077/loop_exit/$exit
      -- CP-element group 102: 	 branch_block_stmt_3076/do_while_stmt_3077/loop_exit/ack
      -- 
    ack_3034_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 102_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_3077_branch_ack_0, ack => readMemoryFromL2_CP_2700_elements(102)); -- 
    -- CP-element group 103:  transition  input  bypass  pipeline-parent 
    -- CP-element group 103: predecessors 
    -- CP-element group 103: 	7 
    -- CP-element group 103: successors 
    -- CP-element group 103:  members (2) 
      -- CP-element group 103: 	 branch_block_stmt_3076/do_while_stmt_3077/loop_taken/$exit
      -- CP-element group 103: 	 branch_block_stmt_3076/do_while_stmt_3077/loop_taken/ack
      -- 
    ack_3038_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 103_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_3077_branch_ack_1, ack => readMemoryFromL2_CP_2700_elements(103)); -- 
    -- CP-element group 104:  transition  bypass  pipeline-parent 
    -- CP-element group 104: predecessors 
    -- CP-element group 104: 	5 
    -- CP-element group 104: successors 
    -- CP-element group 104: 	3 
    -- CP-element group 104:  members (1) 
      -- CP-element group 104: 	 branch_block_stmt_3076/do_while_stmt_3077/$exit
      -- 
    readMemoryFromL2_CP_2700_elements(104) <= readMemoryFromL2_CP_2700_elements(5);
    -- CP-element group 105:  transition  input  bypass 
    -- CP-element group 105: predecessors 
    -- CP-element group 105: 	3 
    -- CP-element group 105: successors 
    -- CP-element group 105:  members (3) 
      -- CP-element group 105: 	 assign_stmt_3231/CONCAT_u256_u512_3230_sample_completed_
      -- CP-element group 105: 	 assign_stmt_3231/CONCAT_u256_u512_3230_Sample/$exit
      -- CP-element group 105: 	 assign_stmt_3231/CONCAT_u256_u512_3230_Sample/ra
      -- 
    ra_3051_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 105_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u256_u512_3230_inst_ack_0, ack => readMemoryFromL2_CP_2700_elements(105)); -- 
    -- CP-element group 106:  transition  input  bypass 
    -- CP-element group 106: predecessors 
    -- CP-element group 106: 	3 
    -- CP-element group 106: successors 
    -- CP-element group 106:  members (5) 
      -- CP-element group 106: 	 $exit
      -- CP-element group 106: 	 assign_stmt_3231/$exit
      -- CP-element group 106: 	 assign_stmt_3231/CONCAT_u256_u512_3230_update_completed_
      -- CP-element group 106: 	 assign_stmt_3231/CONCAT_u256_u512_3230_Update/$exit
      -- CP-element group 106: 	 assign_stmt_3231/CONCAT_u256_u512_3230_Update/ca
      -- 
    ca_3056_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 106_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => CONCAT_u256_u512_3230_inst_ack_1, ack => readMemoryFromL2_CP_2700_elements(106)); -- 
    readMemoryFromL2_do_while_stmt_3077_terminator_3039: loop_terminator -- 
      generic map (name => " readMemoryFromL2_do_while_stmt_3077_terminator_3039", max_iterations_in_flight =>15) 
      port map(loop_body_exit => readMemoryFromL2_CP_2700_elements(8),loop_continue => readMemoryFromL2_CP_2700_elements(103),loop_terminate => readMemoryFromL2_CP_2700_elements(102),loop_back => readMemoryFromL2_CP_2700_elements(6),loop_exit => readMemoryFromL2_CP_2700_elements(5),clk => clk, reset => reset); -- 
    phi_stmt_3079_phi_seq_2791_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= readMemoryFromL2_CP_2700_elements(19);
      readMemoryFromL2_CP_2700_elements(24)<= src_sample_reqs(0);
      src_sample_acks(0)  <= readMemoryFromL2_CP_2700_elements(26);
      readMemoryFromL2_CP_2700_elements(25)<= src_update_reqs(0);
      src_update_acks(0)  <= readMemoryFromL2_CP_2700_elements(27);
      readMemoryFromL2_CP_2700_elements(20) <= phi_mux_reqs(0);
      triggers(1)  <= readMemoryFromL2_CP_2700_elements(21);
      readMemoryFromL2_CP_2700_elements(28)<= src_sample_reqs(1);
      src_sample_acks(1)  <= readMemoryFromL2_CP_2700_elements(28);
      readMemoryFromL2_CP_2700_elements(29)<= src_update_reqs(1);
      src_update_acks(1)  <= readMemoryFromL2_CP_2700_elements(30);
      readMemoryFromL2_CP_2700_elements(22) <= phi_mux_reqs(1);
      phi_stmt_3079_phi_seq_2791 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_3079_phi_seq_2791") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => readMemoryFromL2_CP_2700_elements(13), 
          phi_sample_ack => readMemoryFromL2_CP_2700_elements(17), 
          phi_update_req => readMemoryFromL2_CP_2700_elements(16), 
          phi_update_ack => readMemoryFromL2_CP_2700_elements(18), 
          phi_mux_ack => readMemoryFromL2_CP_2700_elements(23), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_2742_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= readMemoryFromL2_CP_2700_elements(9);
        preds(1)  <= readMemoryFromL2_CP_2700_elements(10);
        entry_tmerge_2742 : transition_merge -- 
          generic map(name => " entry_tmerge_2742")
          port map (preds => preds, symbol_out => readMemoryFromL2_CP_2700_elements(11));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u128_u256_3222_wire : std_logic_vector(255 downto 0);
    signal CONCAT_u128_u256_3229_wire : std_logic_vector(255 downto 0);
    signal CONCAT_u30_u33_3098_wire : std_logic_vector(32 downto 0);
    signal CONCAT_u64_u128_3218_wire : std_logic_vector(127 downto 0);
    signal CONCAT_u64_u128_3221_wire : std_logic_vector(127 downto 0);
    signal CONCAT_u64_u128_3225_wire : std_logic_vector(127 downto 0);
    signal CONCAT_u64_u128_3228_wire : std_logic_vector(127 downto 0);
    signal DWORD_ID_3079 : std_logic_vector(2 downto 0);
    signal NOT_u8_u8_3107_wire_constant : std_logic_vector(7 downto 0);
    signal acquired_lock_3075 : std_logic_vector(0 downto 0);
    signal continue_flag_3089 : std_logic_vector(0 downto 0);
    signal konst_3087_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3092_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3118_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3130_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3142_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3154_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3166_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3178_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3190_wire_constant : std_logic_vector(2 downto 0);
    signal konst_3202_wire_constant : std_logic_vector(2 downto 0);
    signal n_DWORD_ID_3094 : std_logic_vector(2 downto 0);
    signal n_DWORD_ID_3094_3081_buffered : std_logic_vector(2 downto 0);
    signal pa_3102 : std_logic_vector(35 downto 0);
    signal r0_3127 : std_logic_vector(63 downto 0);
    signal r1_3139 : std_logic_vector(63 downto 0);
    signal r2_3151 : std_logic_vector(63 downto 0);
    signal r3_3163 : std_logic_vector(63 downto 0);
    signal r4_3175 : std_logic_vector(63 downto 0);
    signal r5_3187 : std_logic_vector(63 downto 0);
    signal r6_3199 : std_logic_vector(63 downto 0);
    signal r7_3211 : std_logic_vector(63 downto 0);
    signal rval_3112 : std_logic_vector(63 downto 0);
    signal s0_2928_delayed_8_0_3123 : std_logic_vector(0 downto 0);
    signal s0_3120 : std_logic_vector(0 downto 0);
    signal s1_2937_delayed_8_0_3135 : std_logic_vector(0 downto 0);
    signal s1_3132 : std_logic_vector(0 downto 0);
    signal s2_2946_delayed_8_0_3147 : std_logic_vector(0 downto 0);
    signal s2_3144 : std_logic_vector(0 downto 0);
    signal s3_2955_delayed_8_0_3159 : std_logic_vector(0 downto 0);
    signal s3_3156 : std_logic_vector(0 downto 0);
    signal s4_2964_delayed_8_0_3171 : std_logic_vector(0 downto 0);
    signal s4_3168 : std_logic_vector(0 downto 0);
    signal s5_2973_delayed_8_0_3183 : std_logic_vector(0 downto 0);
    signal s5_3180 : std_logic_vector(0 downto 0);
    signal s6_2982_delayed_8_0_3195 : std_logic_vector(0 downto 0);
    signal s6_3192 : std_logic_vector(0 downto 0);
    signal s7_2991_delayed_8_0_3207 : std_logic_vector(0 downto 0);
    signal s7_3204 : std_logic_vector(0 downto 0);
    signal type_cast_3083_wire_constant : std_logic_vector(2 downto 0);
    signal type_cast_3100_wire_constant : std_logic_vector(2 downto 0);
    signal type_cast_3104_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_3110_wire_constant : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    NOT_u8_u8_3107_wire_constant <= "11111111";
    konst_3087_wire_constant <= "111";
    konst_3092_wire_constant <= "001";
    konst_3118_wire_constant <= "000";
    konst_3130_wire_constant <= "001";
    konst_3142_wire_constant <= "010";
    konst_3154_wire_constant <= "011";
    konst_3166_wire_constant <= "100";
    konst_3178_wire_constant <= "101";
    konst_3190_wire_constant <= "110";
    konst_3202_wire_constant <= "111";
    type_cast_3083_wire_constant <= "000";
    type_cast_3100_wire_constant <= "000";
    type_cast_3104_wire_constant <= "1";
    type_cast_3110_wire_constant <= "0000000000000000000000000000000000000000000000000000000000000000";
    phi_stmt_3079: Block -- phi operator 
      signal idata: std_logic_vector(5 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= n_DWORD_ID_3094_3081_buffered & type_cast_3083_wire_constant;
      req <= phi_stmt_3079_req_0 & phi_stmt_3079_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3079",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 3) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3079_ack_0,
          idata => idata,
          odata => DWORD_ID_3079,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3079
    W_r0_3125_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= W_r0_3125_inst_req_0;
      W_r0_3125_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= W_r0_3125_inst_req_1;
      W_r0_3125_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  s0_2928_delayed_8_0_3123(0);
      W_r0_3125_inst_gI: SplitGuardInterface generic map(name => "W_r0_3125_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      W_r0_3125_inst : InterlockBuffer generic map ( -- 
        name => "W_r0_3125_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rval_3112,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => r0_3127,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_r1_3137_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= W_r1_3137_inst_req_0;
      W_r1_3137_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= W_r1_3137_inst_req_1;
      W_r1_3137_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  s1_2937_delayed_8_0_3135(0);
      W_r1_3137_inst_gI: SplitGuardInterface generic map(name => "W_r1_3137_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      W_r1_3137_inst : InterlockBuffer generic map ( -- 
        name => "W_r1_3137_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rval_3112,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => r1_3139,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_r2_3149_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= W_r2_3149_inst_req_0;
      W_r2_3149_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= W_r2_3149_inst_req_1;
      W_r2_3149_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  s2_2946_delayed_8_0_3147(0);
      W_r2_3149_inst_gI: SplitGuardInterface generic map(name => "W_r2_3149_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      W_r2_3149_inst : InterlockBuffer generic map ( -- 
        name => "W_r2_3149_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rval_3112,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => r2_3151,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_r3_3161_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= W_r3_3161_inst_req_0;
      W_r3_3161_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= W_r3_3161_inst_req_1;
      W_r3_3161_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  s3_2955_delayed_8_0_3159(0);
      W_r3_3161_inst_gI: SplitGuardInterface generic map(name => "W_r3_3161_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      W_r3_3161_inst : InterlockBuffer generic map ( -- 
        name => "W_r3_3161_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rval_3112,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => r3_3163,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_r4_3173_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= W_r4_3173_inst_req_0;
      W_r4_3173_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= W_r4_3173_inst_req_1;
      W_r4_3173_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  s4_2964_delayed_8_0_3171(0);
      W_r4_3173_inst_gI: SplitGuardInterface generic map(name => "W_r4_3173_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      W_r4_3173_inst : InterlockBuffer generic map ( -- 
        name => "W_r4_3173_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rval_3112,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => r4_3175,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_r5_3185_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= W_r5_3185_inst_req_0;
      W_r5_3185_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= W_r5_3185_inst_req_1;
      W_r5_3185_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  s5_2973_delayed_8_0_3183(0);
      W_r5_3185_inst_gI: SplitGuardInterface generic map(name => "W_r5_3185_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      W_r5_3185_inst : InterlockBuffer generic map ( -- 
        name => "W_r5_3185_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rval_3112,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => r5_3187,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_r6_3197_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= W_r6_3197_inst_req_0;
      W_r6_3197_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= W_r6_3197_inst_req_1;
      W_r6_3197_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  s6_2982_delayed_8_0_3195(0);
      W_r6_3197_inst_gI: SplitGuardInterface generic map(name => "W_r6_3197_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      W_r6_3197_inst : InterlockBuffer generic map ( -- 
        name => "W_r6_3197_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rval_3112,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => r6_3199,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_r7_3209_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      signal wreq_ug, wack_ug, rreq_ug, rack_ug: BooleanArray(0 downto 0); 
      signal guard_vector : std_logic_vector(0 downto 0); 
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      -- 
    begin -- 
      wreq_ug(0) <= W_r7_3209_inst_req_0;
      W_r7_3209_inst_ack_0<= wack_ug(0);
      rreq_ug(0) <= W_r7_3209_inst_req_1;
      W_r7_3209_inst_ack_1<= rack_ug(0);
      guard_vector(0) <=  s7_2991_delayed_8_0_3207(0);
      W_r7_3209_inst_gI: SplitGuardInterface generic map(name => "W_r7_3209_inst_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => wreq_ug,
        sr_out => wreq,
        sa_in => wack,
        sa_out => wack_ug,
        cr_in => rreq_ug,
        cr_out => rreq,
        ca_in => rack,
        ca_out => rack_ug,
        guards => guard_vector); -- 
      W_r7_3209_inst : InterlockBuffer generic map ( -- 
        name => "W_r7_3209_inst",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 64,
        out_data_width => 64,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => rval_3112,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => r7_3211,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_s0_2928_delayed_8_0_3121_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_s0_2928_delayed_8_0_3121_inst_req_0;
      W_s0_2928_delayed_8_0_3121_inst_ack_0<= wack(0);
      rreq(0) <= W_s0_2928_delayed_8_0_3121_inst_req_1;
      W_s0_2928_delayed_8_0_3121_inst_ack_1<= rack(0);
      W_s0_2928_delayed_8_0_3121_inst : InterlockBuffer generic map ( -- 
        name => "W_s0_2928_delayed_8_0_3121_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => s0_3120,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => s0_2928_delayed_8_0_3123,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_s1_2937_delayed_8_0_3133_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_s1_2937_delayed_8_0_3133_inst_req_0;
      W_s1_2937_delayed_8_0_3133_inst_ack_0<= wack(0);
      rreq(0) <= W_s1_2937_delayed_8_0_3133_inst_req_1;
      W_s1_2937_delayed_8_0_3133_inst_ack_1<= rack(0);
      W_s1_2937_delayed_8_0_3133_inst : InterlockBuffer generic map ( -- 
        name => "W_s1_2937_delayed_8_0_3133_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => s1_3132,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => s1_2937_delayed_8_0_3135,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_s2_2946_delayed_8_0_3145_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_s2_2946_delayed_8_0_3145_inst_req_0;
      W_s2_2946_delayed_8_0_3145_inst_ack_0<= wack(0);
      rreq(0) <= W_s2_2946_delayed_8_0_3145_inst_req_1;
      W_s2_2946_delayed_8_0_3145_inst_ack_1<= rack(0);
      W_s2_2946_delayed_8_0_3145_inst : InterlockBuffer generic map ( -- 
        name => "W_s2_2946_delayed_8_0_3145_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => s2_3144,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => s2_2946_delayed_8_0_3147,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_s3_2955_delayed_8_0_3157_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_s3_2955_delayed_8_0_3157_inst_req_0;
      W_s3_2955_delayed_8_0_3157_inst_ack_0<= wack(0);
      rreq(0) <= W_s3_2955_delayed_8_0_3157_inst_req_1;
      W_s3_2955_delayed_8_0_3157_inst_ack_1<= rack(0);
      W_s3_2955_delayed_8_0_3157_inst : InterlockBuffer generic map ( -- 
        name => "W_s3_2955_delayed_8_0_3157_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => s3_3156,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => s3_2955_delayed_8_0_3159,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_s4_2964_delayed_8_0_3169_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_s4_2964_delayed_8_0_3169_inst_req_0;
      W_s4_2964_delayed_8_0_3169_inst_ack_0<= wack(0);
      rreq(0) <= W_s4_2964_delayed_8_0_3169_inst_req_1;
      W_s4_2964_delayed_8_0_3169_inst_ack_1<= rack(0);
      W_s4_2964_delayed_8_0_3169_inst : InterlockBuffer generic map ( -- 
        name => "W_s4_2964_delayed_8_0_3169_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => s4_3168,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => s4_2964_delayed_8_0_3171,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_s5_2973_delayed_8_0_3181_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_s5_2973_delayed_8_0_3181_inst_req_0;
      W_s5_2973_delayed_8_0_3181_inst_ack_0<= wack(0);
      rreq(0) <= W_s5_2973_delayed_8_0_3181_inst_req_1;
      W_s5_2973_delayed_8_0_3181_inst_ack_1<= rack(0);
      W_s5_2973_delayed_8_0_3181_inst : InterlockBuffer generic map ( -- 
        name => "W_s5_2973_delayed_8_0_3181_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => s5_3180,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => s5_2973_delayed_8_0_3183,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_s6_2982_delayed_8_0_3193_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_s6_2982_delayed_8_0_3193_inst_req_0;
      W_s6_2982_delayed_8_0_3193_inst_ack_0<= wack(0);
      rreq(0) <= W_s6_2982_delayed_8_0_3193_inst_req_1;
      W_s6_2982_delayed_8_0_3193_inst_ack_1<= rack(0);
      W_s6_2982_delayed_8_0_3193_inst : InterlockBuffer generic map ( -- 
        name => "W_s6_2982_delayed_8_0_3193_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => s6_3192,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => s6_2982_delayed_8_0_3195,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    W_s7_2991_delayed_8_0_3205_inst_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= W_s7_2991_delayed_8_0_3205_inst_req_0;
      W_s7_2991_delayed_8_0_3205_inst_ack_0<= wack(0);
      rreq(0) <= W_s7_2991_delayed_8_0_3205_inst_req_1;
      W_s7_2991_delayed_8_0_3205_inst_ack_1<= rack(0);
      W_s7_2991_delayed_8_0_3205_inst : InterlockBuffer generic map ( -- 
        name => "W_s7_2991_delayed_8_0_3205_inst",
        buffer_size => 8,
        flow_through =>  false ,
        cut_through =>  true ,
        in_data_width => 1,
        out_data_width => 1,
        bypass_flag =>  true 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => s7_3204,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => s7_2991_delayed_8_0_3207,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    n_DWORD_ID_3094_3081_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= n_DWORD_ID_3094_3081_buf_req_0;
      n_DWORD_ID_3094_3081_buf_ack_0<= wack(0);
      rreq(0) <= n_DWORD_ID_3094_3081_buf_req_1;
      n_DWORD_ID_3094_3081_buf_ack_1<= rack(0);
      n_DWORD_ID_3094_3081_buf : InterlockBuffer generic map ( -- 
        name => "n_DWORD_ID_3094_3081_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 3,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => n_DWORD_ID_3094,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => n_DWORD_ID_3094_3081_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_3077_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= continue_flag_3089;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_3077_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_3077_branch_req_0,
          ack0 => do_while_stmt_3077_branch_ack_0,
          ack1 => do_while_stmt_3077_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator ADD_u3_u3_3093_inst
    process(DWORD_ID_3079) -- 
      variable tmp_var : std_logic_vector(2 downto 0); -- 
    begin -- 
      ApIntAdd_proc(DWORD_ID_3079, konst_3092_wire_constant, tmp_var);
      n_DWORD_ID_3094 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u128_u256_3222_inst
    process(CONCAT_u64_u128_3218_wire, CONCAT_u64_u128_3221_wire) -- 
      variable tmp_var : std_logic_vector(255 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u64_u128_3218_wire, CONCAT_u64_u128_3221_wire, tmp_var);
      CONCAT_u128_u256_3222_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u128_u256_3229_inst
    process(CONCAT_u64_u128_3225_wire, CONCAT_u64_u128_3228_wire) -- 
      variable tmp_var : std_logic_vector(255 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u64_u128_3225_wire, CONCAT_u64_u128_3228_wire, tmp_var);
      CONCAT_u128_u256_3229_wire <= tmp_var; --
    end process;
    -- shared split operator group (3) : CONCAT_u256_u512_3230_inst 
    ApConcat_group_3: Block -- 
      signal data_in: std_logic_vector(511 downto 0);
      signal data_out: std_logic_vector(511 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      data_in <= CONCAT_u128_u256_3222_wire & CONCAT_u128_u256_3229_wire;
      rline_buffer <= data_out(511 downto 0);
      guard_vector(0)  <=  '1';
      reqL_unguarded(0) <= CONCAT_u256_u512_3230_inst_req_0;
      CONCAT_u256_u512_3230_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= CONCAT_u256_u512_3230_inst_req_1;
      CONCAT_u256_u512_3230_inst_ack_1 <= ackR_unguarded(0);
      ApConcat_group_3_gI: SplitGuardInterface generic map(name => "ApConcat_group_3_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      UnsharedOperator: UnsharedOperatorWithBuffering -- 
        generic map ( -- 
          operator_id => "ApConcat",
          name => "ApConcat_group_3",
          input1_is_int => true, 
          input1_characteristic_width => 0, 
          input1_mantissa_width    => 0, 
          iwidth_1  => 256,
          input2_is_int => true, 
          input2_characteristic_width => 0, 
          input2_mantissa_width => 0, 
          iwidth_2      => 256, 
          num_inputs    => 2,
          output_is_int => true,
          output_characteristic_width  => 0, 
          output_mantissa_width => 0, 
          owidth => 512,
          constant_operand => "0",
          constant_width => 1,
          buffering  => 1,
          flow_through => false,
          full_rate  => false,
          use_constant  => false
          --
        ) 
        port map ( -- 
          reqL => reqL(0),
          ackL => ackL(0),
          reqR => reqR(0),
          ackR => ackR(0),
          dataL => data_in, 
          dataR => data_out,
          clk => clk,
          reset => reset); -- 
      -- 
    end Block; -- split operator group 3
    -- binary operator CONCAT_u30_u33_3098_inst
    process(line_address_buffer, DWORD_ID_3079) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(line_address_buffer, DWORD_ID_3079, tmp_var);
      CONCAT_u30_u33_3098_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u33_u36_3101_inst
    process(CONCAT_u30_u33_3098_wire) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u30_u33_3098_wire, type_cast_3100_wire_constant, tmp_var);
      pa_3102 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u64_u128_3218_inst
    process(r0_3127, r1_3139) -- 
      variable tmp_var : std_logic_vector(127 downto 0); -- 
    begin -- 
      ApConcat_proc(r0_3127, r1_3139, tmp_var);
      CONCAT_u64_u128_3218_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u64_u128_3221_inst
    process(r2_3151, r3_3163) -- 
      variable tmp_var : std_logic_vector(127 downto 0); -- 
    begin -- 
      ApConcat_proc(r2_3151, r3_3163, tmp_var);
      CONCAT_u64_u128_3221_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u64_u128_3225_inst
    process(r4_3175, r5_3187) -- 
      variable tmp_var : std_logic_vector(127 downto 0); -- 
    begin -- 
      ApConcat_proc(r4_3175, r5_3187, tmp_var);
      CONCAT_u64_u128_3225_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u64_u128_3228_inst
    process(r6_3199, r7_3211) -- 
      variable tmp_var : std_logic_vector(127 downto 0); -- 
    begin -- 
      ApConcat_proc(r6_3199, r7_3211, tmp_var);
      CONCAT_u64_u128_3228_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_3119_inst
    process(DWORD_ID_3079) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(DWORD_ID_3079, konst_3118_wire_constant, tmp_var);
      s0_3120 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_3131_inst
    process(DWORD_ID_3079) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(DWORD_ID_3079, konst_3130_wire_constant, tmp_var);
      s1_3132 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_3143_inst
    process(DWORD_ID_3079) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(DWORD_ID_3079, konst_3142_wire_constant, tmp_var);
      s2_3144 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_3155_inst
    process(DWORD_ID_3079) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(DWORD_ID_3079, konst_3154_wire_constant, tmp_var);
      s3_3156 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_3167_inst
    process(DWORD_ID_3079) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(DWORD_ID_3079, konst_3166_wire_constant, tmp_var);
      s4_3168 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_3179_inst
    process(DWORD_ID_3079) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(DWORD_ID_3079, konst_3178_wire_constant, tmp_var);
      s5_3180 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_3191_inst
    process(DWORD_ID_3079) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(DWORD_ID_3079, konst_3190_wire_constant, tmp_var);
      s6_3192 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_3203_inst
    process(DWORD_ID_3079) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(DWORD_ID_3079, konst_3202_wire_constant, tmp_var);
      s7_3204 <= tmp_var; --
    end process;
    -- binary operator ULT_u3_u1_3088_inst
    process(DWORD_ID_3079) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntUlt_proc(DWORD_ID_3079, konst_3087_wire_constant, tmp_var);
      continue_flag_3089 <= tmp_var; --
    end process;
    -- shared inport operator group (0) : RPIPE_sys_mem_lock_3074_inst 
    InportGroup_0: Block -- 
      signal data_out: std_logic_vector(0 downto 0);
      signal reqL, ackL, reqR, ackR : BooleanArray( 0 downto 0);
      signal reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      reqL_unguarded(0) <= RPIPE_sys_mem_lock_3074_inst_req_0;
      RPIPE_sys_mem_lock_3074_inst_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= RPIPE_sys_mem_lock_3074_inst_req_1;
      RPIPE_sys_mem_lock_3074_inst_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      acquired_lock_3075 <= data_out(0 downto 0);
      sys_mem_lock_read_0_gI: SplitGuardInterface generic map(name => "sys_mem_lock_read_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => true) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL,
        sa_in => ackL,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      sys_mem_lock_read_0: InputPortRevised -- 
        generic map ( name => "sys_mem_lock_read_0", data_width => 1,  num_reqs => 1,  output_buffering => outBUFs,   nonblocking_read_flag => False,  no_arbitration => false)
        port map (-- 
          sample_req => reqL , 
          sample_ack => ackL, 
          update_req => reqR, 
          update_ack => ackR, 
          data => data_out, 
          oreq => sys_mem_lock_pipe_read_req(0),
          oack => sys_mem_lock_pipe_read_ack(0),
          odata => sys_mem_lock_pipe_read_data(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      -- 
    end Block; -- inport group 0
    -- shared call operator group (0) : call_stmt_3112_call 
    accessSysMem_call_group_0: Block -- 
      signal data_in: std_logic_vector(108 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => false);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 8);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_3112_call_req_0;
      call_stmt_3112_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_3112_call_req_1;
      call_stmt_3112_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  '1';
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessSysMem_call_group_0_gI: SplitGuardInterface generic map(name => "accessSysMem_call_group_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_3104_wire_constant & NOT_u8_u8_3107_wire_constant & pa_3102 & type_cast_3110_wire_constant;
      rval_3112 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 109,
        owidth => 109,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessSysMem_call_reqs(0),
          ackR => accessSysMem_call_acks(0),
          dataR => accessSysMem_call_data(108 downto 0),
          tagR => accessSysMem_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessSysMem_return_acks(0), -- cross-over
          ackL => accessSysMem_return_reqs(0), -- cross-over
          dataL => accessSysMem_return_data(63 downto 0),
          tagL => accessSysMem_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 0
    -- 
  end Block; -- data_path
  -- 
end readMemoryFromL2_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library l2_cache_lib;
use l2_cache_lib.l2_cache_global_package.all;
entity setId_Volatile is -- 
  port ( -- 
    pa : in  std_logic_vector(35 downto 0);
    set_id : out  std_logic_vector(8 downto 0)-- 
  );
  -- 
end entity setId_Volatile;
architecture setId_Volatile_arch of setId_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(36-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal pa_buffer :  std_logic_vector(35 downto 0);
  -- output port buffer signals
  signal set_id_buffer :  std_logic_vector(8 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  pa_buffer <= pa;
  -- output handling  -------------------------------------------------------
  set_id <= set_id_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    -- 
  begin -- 
    -- flow-through slice operator slice_3057_inst
    set_id_buffer <= pa_buffer(14 downto 6);
    -- 
  end Block; -- data_path
  -- 
end setId_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library l2_cache_lib;
use l2_cache_lib.l2_cache_global_package.all;
entity updateDirtyWordMask_Volatile is -- 
  port ( -- 
    invalidate : in  std_logic_vector(0 downto 0);
    read_write_access : in  std_logic_vector(0 downto 0);
    is_hit : in  std_logic_vector(0 downto 0);
    rwbar : in  std_logic_vector(0 downto 0);
    dword_id : in  std_logic_vector(2 downto 0);
    current_dirty_mask : in  std_logic_vector(7 downto 0);
    updated_dirty_mask : out  std_logic_vector(7 downto 0)-- 
  );
  -- 
end entity updateDirtyWordMask_Volatile;
architecture updateDirtyWordMask_Volatile_arch of updateDirtyWordMask_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(15-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal invalidate_buffer :  std_logic_vector(0 downto 0);
  signal read_write_access_buffer :  std_logic_vector(0 downto 0);
  signal is_hit_buffer :  std_logic_vector(0 downto 0);
  signal rwbar_buffer :  std_logic_vector(0 downto 0);
  signal dword_id_buffer :  std_logic_vector(2 downto 0);
  signal current_dirty_mask_buffer :  std_logic_vector(7 downto 0);
  -- output port buffer signals
  signal updated_dirty_mask_buffer :  std_logic_vector(7 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  invalidate_buffer <= invalidate;
  read_write_access_buffer <= read_write_access;
  is_hit_buffer <= is_hit;
  rwbar_buffer <= rwbar;
  dword_id_buffer <= dword_id;
  current_dirty_mask_buffer <= current_dirty_mask;
  -- output handling  -------------------------------------------------------
  updated_dirty_mask <= updated_dirty_mask_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_1768_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_1821_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_1829_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_1838_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_1846_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_1856_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_1864_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_1873_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_1881_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_1894_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_1899_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_1905_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_1910_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_1917_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_1922_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_1928_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_1933_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u1_u2_1833_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_1850_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_1868_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_1885_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_1900_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_1911_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_1923_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_1934_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u2_u4_1851_wire : std_logic_vector(3 downto 0);
    signal CONCAT_u2_u4_1886_wire : std_logic_vector(3 downto 0);
    signal CONCAT_u2_u4_1912_wire : std_logic_vector(3 downto 0);
    signal CONCAT_u2_u4_1935_wire : std_logic_vector(3 downto 0);
    signal EQ_u3_u1_1820_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1828_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1837_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1845_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1855_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1863_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1872_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1880_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1892_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1897_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1903_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1908_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1915_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1920_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1926_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_1931_wire : std_logic_vector(0 downto 0);
    signal MUX_1824_wire : std_logic_vector(0 downto 0);
    signal MUX_1832_wire : std_logic_vector(0 downto 0);
    signal MUX_1841_wire : std_logic_vector(0 downto 0);
    signal MUX_1849_wire : std_logic_vector(0 downto 0);
    signal MUX_1859_wire : std_logic_vector(0 downto 0);
    signal MUX_1867_wire : std_logic_vector(0 downto 0);
    signal MUX_1876_wire : std_logic_vector(0 downto 0);
    signal MUX_1884_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1757_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1759_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1767_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1775_wire : std_logic_vector(0 downto 0);
    signal NOT_u1_u1_1781_wire : std_logic_vector(0 downto 0);
    signal OR_u1_u1_1769_wire : std_logic_vector(0 downto 0);
    signal bitval_1761 : std_logic_vector(0 downto 0);
    signal clear_bits_1777 : std_logic_vector(0 downto 0);
    signal d0_1787 : std_logic_vector(0 downto 0);
    signal d1_1791 : std_logic_vector(0 downto 0);
    signal d2_1795 : std_logic_vector(0 downto 0);
    signal d3_1799 : std_logic_vector(0 downto 0);
    signal d4_1803 : std_logic_vector(0 downto 0);
    signal d5_1807 : std_logic_vector(0 downto 0);
    signal d6_1811 : std_logic_vector(0 downto 0);
    signal d7_1815 : std_logic_vector(0 downto 0);
    signal konst_1819_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1827_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1836_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1844_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1854_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1862_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1871_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1879_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1891_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1896_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1902_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1907_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1914_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1919_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1925_wire_constant : std_logic_vector(2 downto 0);
    signal konst_1930_wire_constant : std_logic_vector(2 downto 0);
    signal modified_dirty_mask_1888 : std_logic_vector(7 downto 0);
    signal modify_1771 : std_logic_vector(0 downto 0);
    signal new_dirty_mask_1937 : std_logic_vector(7 downto 0);
    signal set_bit_in_new_mask_1783 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    konst_1819_wire_constant <= "000";
    konst_1827_wire_constant <= "001";
    konst_1836_wire_constant <= "010";
    konst_1844_wire_constant <= "011";
    konst_1854_wire_constant <= "100";
    konst_1862_wire_constant <= "101";
    konst_1871_wire_constant <= "110";
    konst_1879_wire_constant <= "111";
    konst_1891_wire_constant <= "000";
    konst_1896_wire_constant <= "001";
    konst_1902_wire_constant <= "010";
    konst_1907_wire_constant <= "011";
    konst_1914_wire_constant <= "100";
    konst_1919_wire_constant <= "101";
    konst_1925_wire_constant <= "110";
    konst_1930_wire_constant <= "111";
    -- flow-through select operator MUX_1824_inst
    MUX_1824_wire <= bitval_1761 when (AND_u1_u1_1821_wire(0) /=  '0') else d0_1787;
    -- flow-through select operator MUX_1832_inst
    MUX_1832_wire <= bitval_1761 when (AND_u1_u1_1829_wire(0) /=  '0') else d1_1791;
    -- flow-through select operator MUX_1841_inst
    MUX_1841_wire <= bitval_1761 when (AND_u1_u1_1838_wire(0) /=  '0') else d2_1795;
    -- flow-through select operator MUX_1849_inst
    MUX_1849_wire <= bitval_1761 when (AND_u1_u1_1846_wire(0) /=  '0') else d3_1799;
    -- flow-through select operator MUX_1859_inst
    MUX_1859_wire <= bitval_1761 when (AND_u1_u1_1856_wire(0) /=  '0') else d4_1803;
    -- flow-through select operator MUX_1867_inst
    MUX_1867_wire <= bitval_1761 when (AND_u1_u1_1864_wire(0) /=  '0') else d5_1807;
    -- flow-through select operator MUX_1876_inst
    MUX_1876_wire <= bitval_1761 when (AND_u1_u1_1873_wire(0) /=  '0') else d6_1811;
    -- flow-through select operator MUX_1884_inst
    MUX_1884_wire <= bitval_1761 when (AND_u1_u1_1881_wire(0) /=  '0') else d7_1815;
    -- flow-through select operator MUX_1942_inst
    updated_dirty_mask_buffer <= new_dirty_mask_1937 when (clear_bits_1777(0) /=  '0') else modified_dirty_mask_1888;
    -- flow-through slice operator slice_1786_inst
    d0_1787 <= current_dirty_mask_buffer(7 downto 7);
    -- flow-through slice operator slice_1790_inst
    d1_1791 <= current_dirty_mask_buffer(6 downto 6);
    -- flow-through slice operator slice_1794_inst
    d2_1795 <= current_dirty_mask_buffer(5 downto 5);
    -- flow-through slice operator slice_1798_inst
    d3_1799 <= current_dirty_mask_buffer(4 downto 4);
    -- flow-through slice operator slice_1802_inst
    d4_1803 <= current_dirty_mask_buffer(3 downto 3);
    -- flow-through slice operator slice_1806_inst
    d5_1807 <= current_dirty_mask_buffer(2 downto 2);
    -- flow-through slice operator slice_1810_inst
    d6_1811 <= current_dirty_mask_buffer(1 downto 1);
    -- flow-through slice operator slice_1814_inst
    d7_1815 <= current_dirty_mask_buffer(0 downto 0);
    -- binary operator AND_u1_u1_1760_inst
    process(NOT_u1_u1_1757_wire, NOT_u1_u1_1759_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(NOT_u1_u1_1757_wire, NOT_u1_u1_1759_wire, tmp_var);
      bitval_1761 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1768_inst
    process(read_write_access_buffer, NOT_u1_u1_1767_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(read_write_access_buffer, NOT_u1_u1_1767_wire, tmp_var);
      AND_u1_u1_1768_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1770_inst
    process(is_hit_buffer, OR_u1_u1_1769_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(is_hit_buffer, OR_u1_u1_1769_wire, tmp_var);
      modify_1771 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1776_inst
    process(read_write_access_buffer, NOT_u1_u1_1775_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(read_write_access_buffer, NOT_u1_u1_1775_wire, tmp_var);
      clear_bits_1777 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1782_inst
    process(clear_bits_1777, NOT_u1_u1_1781_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(clear_bits_1777, NOT_u1_u1_1781_wire, tmp_var);
      set_bit_in_new_mask_1783 <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1821_inst
    process(modify_1771, EQ_u3_u1_1820_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(modify_1771, EQ_u3_u1_1820_wire, tmp_var);
      AND_u1_u1_1821_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1829_inst
    process(modify_1771, EQ_u3_u1_1828_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(modify_1771, EQ_u3_u1_1828_wire, tmp_var);
      AND_u1_u1_1829_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1838_inst
    process(modify_1771, EQ_u3_u1_1837_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(modify_1771, EQ_u3_u1_1837_wire, tmp_var);
      AND_u1_u1_1838_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1846_inst
    process(modify_1771, EQ_u3_u1_1845_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(modify_1771, EQ_u3_u1_1845_wire, tmp_var);
      AND_u1_u1_1846_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1856_inst
    process(modify_1771, EQ_u3_u1_1855_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(modify_1771, EQ_u3_u1_1855_wire, tmp_var);
      AND_u1_u1_1856_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1864_inst
    process(modify_1771, EQ_u3_u1_1863_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(modify_1771, EQ_u3_u1_1863_wire, tmp_var);
      AND_u1_u1_1864_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1873_inst
    process(modify_1771, EQ_u3_u1_1872_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(modify_1771, EQ_u3_u1_1872_wire, tmp_var);
      AND_u1_u1_1873_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1881_inst
    process(modify_1771, EQ_u3_u1_1880_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(modify_1771, EQ_u3_u1_1880_wire, tmp_var);
      AND_u1_u1_1881_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1894_inst
    process(EQ_u3_u1_1892_wire, set_bit_in_new_mask_1783) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u3_u1_1892_wire, set_bit_in_new_mask_1783, tmp_var);
      AND_u1_u1_1894_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1899_inst
    process(EQ_u3_u1_1897_wire, set_bit_in_new_mask_1783) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u3_u1_1897_wire, set_bit_in_new_mask_1783, tmp_var);
      AND_u1_u1_1899_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1905_inst
    process(EQ_u3_u1_1903_wire, set_bit_in_new_mask_1783) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u3_u1_1903_wire, set_bit_in_new_mask_1783, tmp_var);
      AND_u1_u1_1905_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1910_inst
    process(EQ_u3_u1_1908_wire, set_bit_in_new_mask_1783) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u3_u1_1908_wire, set_bit_in_new_mask_1783, tmp_var);
      AND_u1_u1_1910_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1917_inst
    process(EQ_u3_u1_1915_wire, set_bit_in_new_mask_1783) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u3_u1_1915_wire, set_bit_in_new_mask_1783, tmp_var);
      AND_u1_u1_1917_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1922_inst
    process(EQ_u3_u1_1920_wire, set_bit_in_new_mask_1783) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u3_u1_1920_wire, set_bit_in_new_mask_1783, tmp_var);
      AND_u1_u1_1922_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1928_inst
    process(EQ_u3_u1_1926_wire, set_bit_in_new_mask_1783) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u3_u1_1926_wire, set_bit_in_new_mask_1783, tmp_var);
      AND_u1_u1_1928_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_1933_inst
    process(EQ_u3_u1_1931_wire, set_bit_in_new_mask_1783) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(EQ_u3_u1_1931_wire, set_bit_in_new_mask_1783, tmp_var);
      AND_u1_u1_1933_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_1833_inst
    process(MUX_1824_wire, MUX_1832_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_1824_wire, MUX_1832_wire, tmp_var);
      CONCAT_u1_u2_1833_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_1850_inst
    process(MUX_1841_wire, MUX_1849_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_1841_wire, MUX_1849_wire, tmp_var);
      CONCAT_u1_u2_1850_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_1868_inst
    process(MUX_1859_wire, MUX_1867_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_1859_wire, MUX_1867_wire, tmp_var);
      CONCAT_u1_u2_1868_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_1885_inst
    process(MUX_1876_wire, MUX_1884_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_1876_wire, MUX_1884_wire, tmp_var);
      CONCAT_u1_u2_1885_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_1900_inst
    process(AND_u1_u1_1894_wire, AND_u1_u1_1899_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(AND_u1_u1_1894_wire, AND_u1_u1_1899_wire, tmp_var);
      CONCAT_u1_u2_1900_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_1911_inst
    process(AND_u1_u1_1905_wire, AND_u1_u1_1910_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(AND_u1_u1_1905_wire, AND_u1_u1_1910_wire, tmp_var);
      CONCAT_u1_u2_1911_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_1923_inst
    process(AND_u1_u1_1917_wire, AND_u1_u1_1922_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(AND_u1_u1_1917_wire, AND_u1_u1_1922_wire, tmp_var);
      CONCAT_u1_u2_1923_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_1934_inst
    process(AND_u1_u1_1928_wire, AND_u1_u1_1933_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(AND_u1_u1_1928_wire, AND_u1_u1_1933_wire, tmp_var);
      CONCAT_u1_u2_1934_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u2_u4_1851_inst
    process(CONCAT_u1_u2_1833_wire, CONCAT_u1_u2_1850_wire) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_1833_wire, CONCAT_u1_u2_1850_wire, tmp_var);
      CONCAT_u2_u4_1851_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u2_u4_1886_inst
    process(CONCAT_u1_u2_1868_wire, CONCAT_u1_u2_1885_wire) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_1868_wire, CONCAT_u1_u2_1885_wire, tmp_var);
      CONCAT_u2_u4_1886_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u2_u4_1912_inst
    process(CONCAT_u1_u2_1900_wire, CONCAT_u1_u2_1911_wire) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_1900_wire, CONCAT_u1_u2_1911_wire, tmp_var);
      CONCAT_u2_u4_1912_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u2_u4_1935_inst
    process(CONCAT_u1_u2_1923_wire, CONCAT_u1_u2_1934_wire) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_1923_wire, CONCAT_u1_u2_1934_wire, tmp_var);
      CONCAT_u2_u4_1935_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u4_u8_1887_inst
    process(CONCAT_u2_u4_1851_wire, CONCAT_u2_u4_1886_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u2_u4_1851_wire, CONCAT_u2_u4_1886_wire, tmp_var);
      modified_dirty_mask_1888 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u4_u8_1936_inst
    process(CONCAT_u2_u4_1912_wire, CONCAT_u2_u4_1935_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u2_u4_1912_wire, CONCAT_u2_u4_1935_wire, tmp_var);
      new_dirty_mask_1937 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1820_inst
    process(dword_id_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dword_id_buffer, konst_1819_wire_constant, tmp_var);
      EQ_u3_u1_1820_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1828_inst
    process(dword_id_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dword_id_buffer, konst_1827_wire_constant, tmp_var);
      EQ_u3_u1_1828_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1837_inst
    process(dword_id_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dword_id_buffer, konst_1836_wire_constant, tmp_var);
      EQ_u3_u1_1837_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1845_inst
    process(dword_id_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dword_id_buffer, konst_1844_wire_constant, tmp_var);
      EQ_u3_u1_1845_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1855_inst
    process(dword_id_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dword_id_buffer, konst_1854_wire_constant, tmp_var);
      EQ_u3_u1_1855_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1863_inst
    process(dword_id_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dword_id_buffer, konst_1862_wire_constant, tmp_var);
      EQ_u3_u1_1863_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1872_inst
    process(dword_id_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dword_id_buffer, konst_1871_wire_constant, tmp_var);
      EQ_u3_u1_1872_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1880_inst
    process(dword_id_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dword_id_buffer, konst_1879_wire_constant, tmp_var);
      EQ_u3_u1_1880_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1892_inst
    process(dword_id_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dword_id_buffer, konst_1891_wire_constant, tmp_var);
      EQ_u3_u1_1892_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1897_inst
    process(dword_id_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dword_id_buffer, konst_1896_wire_constant, tmp_var);
      EQ_u3_u1_1897_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1903_inst
    process(dword_id_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dword_id_buffer, konst_1902_wire_constant, tmp_var);
      EQ_u3_u1_1903_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1908_inst
    process(dword_id_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dword_id_buffer, konst_1907_wire_constant, tmp_var);
      EQ_u3_u1_1908_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1915_inst
    process(dword_id_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dword_id_buffer, konst_1914_wire_constant, tmp_var);
      EQ_u3_u1_1915_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1920_inst
    process(dword_id_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dword_id_buffer, konst_1919_wire_constant, tmp_var);
      EQ_u3_u1_1920_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1926_inst
    process(dword_id_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dword_id_buffer, konst_1925_wire_constant, tmp_var);
      EQ_u3_u1_1926_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_1931_inst
    process(dword_id_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(dword_id_buffer, konst_1930_wire_constant, tmp_var);
      EQ_u3_u1_1931_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1757_inst
    process(rwbar_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", rwbar_buffer, tmp_var);
      NOT_u1_u1_1757_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1759_inst
    process(invalidate_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", invalidate_buffer, tmp_var);
      NOT_u1_u1_1759_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1767_inst
    process(rwbar_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", rwbar_buffer, tmp_var);
      NOT_u1_u1_1767_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1775_inst
    process(is_hit_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", is_hit_buffer, tmp_var);
      NOT_u1_u1_1775_wire <= tmp_var; -- 
    end process;
    -- unary operator NOT_u1_u1_1781_inst
    process(rwbar_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", rwbar_buffer, tmp_var);
      NOT_u1_u1_1781_wire <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_1769_inst
    process(invalidate_buffer, AND_u1_u1_1768_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(invalidate_buffer, AND_u1_u1_1768_wire, tmp_var);
      OR_u1_u1_1769_wire <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end updateDirtyWordMask_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library l2_cache_lib;
use l2_cache_lib.l2_cache_global_package.all;
entity updateSetTags_Volatile is -- 
  port ( -- 
    read_write_access : in  std_logic_vector(0 downto 0);
    access_index : in  std_logic_vector(2 downto 0);
    pa_tag : in  std_logic_vector(20 downto 0);
    set_tags : in  std_logic_vector(167 downto 0);
    updated_set_tags : out  std_logic_vector(167 downto 0)-- 
  );
  -- 
end entity updateSetTags_Volatile;
architecture updateSetTags_Volatile_arch of updateSetTags_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(193-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal read_write_access_buffer :  std_logic_vector(0 downto 0);
  signal access_index_buffer :  std_logic_vector(2 downto 0);
  signal pa_tag_buffer :  std_logic_vector(20 downto 0);
  signal set_tags_buffer :  std_logic_vector(167 downto 0);
  -- output port buffer signals
  signal updated_set_tags_buffer :  std_logic_vector(167 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  read_write_access_buffer <= read_write_access;
  access_index_buffer <= access_index;
  pa_tag_buffer <= pa_tag;
  set_tags_buffer <= set_tags;
  -- output handling  -------------------------------------------------------
  updated_set_tags <= updated_set_tags_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_2119_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_2127_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_2136_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_2144_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_2154_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_2162_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_2171_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_2179_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u21_u42_2131_wire : std_logic_vector(41 downto 0);
    signal CONCAT_u21_u42_2148_wire : std_logic_vector(41 downto 0);
    signal CONCAT_u21_u42_2166_wire : std_logic_vector(41 downto 0);
    signal CONCAT_u21_u42_2183_wire : std_logic_vector(41 downto 0);
    signal CONCAT_u42_u84_2149_wire : std_logic_vector(83 downto 0);
    signal CONCAT_u42_u84_2184_wire : std_logic_vector(83 downto 0);
    signal EQ_u3_u1_2118_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2126_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2135_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2143_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2153_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2161_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2170_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2178_wire : std_logic_vector(0 downto 0);
    signal MUX_2122_wire : std_logic_vector(20 downto 0);
    signal MUX_2130_wire : std_logic_vector(20 downto 0);
    signal MUX_2139_wire : std_logic_vector(20 downto 0);
    signal MUX_2147_wire : std_logic_vector(20 downto 0);
    signal MUX_2157_wire : std_logic_vector(20 downto 0);
    signal MUX_2165_wire : std_logic_vector(20 downto 0);
    signal MUX_2174_wire : std_logic_vector(20 downto 0);
    signal MUX_2182_wire : std_logic_vector(20 downto 0);
    signal insert_bit_2081 : std_logic_vector(0 downto 0);
    signal konst_2117_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2125_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2134_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2142_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2152_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2160_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2169_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2177_wire_constant : std_logic_vector(2 downto 0);
    signal modified_set_tags_2186 : std_logic_vector(167 downto 0);
    signal t0_2085 : std_logic_vector(20 downto 0);
    signal t1_2089 : std_logic_vector(20 downto 0);
    signal t2_2093 : std_logic_vector(20 downto 0);
    signal t3_2097 : std_logic_vector(20 downto 0);
    signal t4_2101 : std_logic_vector(20 downto 0);
    signal t5_2105 : std_logic_vector(20 downto 0);
    signal t6_2109 : std_logic_vector(20 downto 0);
    signal t7_2113 : std_logic_vector(20 downto 0);
    -- 
  begin -- 
    konst_2117_wire_constant <= "000";
    konst_2125_wire_constant <= "001";
    konst_2134_wire_constant <= "010";
    konst_2142_wire_constant <= "011";
    konst_2152_wire_constant <= "100";
    konst_2160_wire_constant <= "101";
    konst_2169_wire_constant <= "110";
    konst_2177_wire_constant <= "111";
    -- flow-through select operator MUX_2122_inst
    MUX_2122_wire <= pa_tag_buffer when (AND_u1_u1_2119_wire(0) /=  '0') else t0_2085;
    -- flow-through select operator MUX_2130_inst
    MUX_2130_wire <= pa_tag_buffer when (AND_u1_u1_2127_wire(0) /=  '0') else t1_2089;
    -- flow-through select operator MUX_2139_inst
    MUX_2139_wire <= pa_tag_buffer when (AND_u1_u1_2136_wire(0) /=  '0') else t2_2093;
    -- flow-through select operator MUX_2147_inst
    MUX_2147_wire <= pa_tag_buffer when (AND_u1_u1_2144_wire(0) /=  '0') else t3_2097;
    -- flow-through select operator MUX_2157_inst
    MUX_2157_wire <= pa_tag_buffer when (AND_u1_u1_2154_wire(0) /=  '0') else t4_2101;
    -- flow-through select operator MUX_2165_inst
    MUX_2165_wire <= pa_tag_buffer when (AND_u1_u1_2162_wire(0) /=  '0') else t5_2105;
    -- flow-through select operator MUX_2174_inst
    MUX_2174_wire <= pa_tag_buffer when (AND_u1_u1_2171_wire(0) /=  '0') else t6_2109;
    -- flow-through select operator MUX_2182_inst
    MUX_2182_wire <= pa_tag_buffer when (AND_u1_u1_2179_wire(0) /=  '0') else t7_2113;
    -- flow-through select operator MUX_2191_inst
    updated_set_tags_buffer <= modified_set_tags_2186 when (read_write_access_buffer(0) /=  '0') else set_tags_buffer;
    -- flow-through slice operator slice_2084_inst
    t0_2085 <= set_tags_buffer(167 downto 147);
    -- flow-through slice operator slice_2088_inst
    t1_2089 <= set_tags_buffer(146 downto 126);
    -- flow-through slice operator slice_2092_inst
    t2_2093 <= set_tags_buffer(125 downto 105);
    -- flow-through slice operator slice_2096_inst
    t3_2097 <= set_tags_buffer(104 downto 84);
    -- flow-through slice operator slice_2100_inst
    t4_2101 <= set_tags_buffer(83 downto 63);
    -- flow-through slice operator slice_2104_inst
    t5_2105 <= set_tags_buffer(62 downto 42);
    -- flow-through slice operator slice_2108_inst
    t6_2109 <= set_tags_buffer(41 downto 21);
    -- flow-through slice operator slice_2112_inst
    t7_2113 <= set_tags_buffer(20 downto 0);
    -- interlock W_insert_bit_2079_inst
    process(read_write_access_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 0 downto 0) := read_write_access_buffer(0 downto 0);
      insert_bit_2081 <= tmp_var; -- 
    end process;
    -- binary operator AND_u1_u1_2119_inst
    process(insert_bit_2081, EQ_u3_u1_2118_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(insert_bit_2081, EQ_u3_u1_2118_wire, tmp_var);
      AND_u1_u1_2119_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2127_inst
    process(insert_bit_2081, EQ_u3_u1_2126_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(insert_bit_2081, EQ_u3_u1_2126_wire, tmp_var);
      AND_u1_u1_2127_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2136_inst
    process(insert_bit_2081, EQ_u3_u1_2135_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(insert_bit_2081, EQ_u3_u1_2135_wire, tmp_var);
      AND_u1_u1_2136_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2144_inst
    process(insert_bit_2081, EQ_u3_u1_2143_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(insert_bit_2081, EQ_u3_u1_2143_wire, tmp_var);
      AND_u1_u1_2144_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2154_inst
    process(insert_bit_2081, EQ_u3_u1_2153_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(insert_bit_2081, EQ_u3_u1_2153_wire, tmp_var);
      AND_u1_u1_2154_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2162_inst
    process(insert_bit_2081, EQ_u3_u1_2161_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(insert_bit_2081, EQ_u3_u1_2161_wire, tmp_var);
      AND_u1_u1_2162_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2171_inst
    process(insert_bit_2081, EQ_u3_u1_2170_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(insert_bit_2081, EQ_u3_u1_2170_wire, tmp_var);
      AND_u1_u1_2171_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2179_inst
    process(insert_bit_2081, EQ_u3_u1_2178_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(insert_bit_2081, EQ_u3_u1_2178_wire, tmp_var);
      AND_u1_u1_2179_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u21_u42_2131_inst
    process(MUX_2122_wire, MUX_2130_wire) -- 
      variable tmp_var : std_logic_vector(41 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_2122_wire, MUX_2130_wire, tmp_var);
      CONCAT_u21_u42_2131_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u21_u42_2148_inst
    process(MUX_2139_wire, MUX_2147_wire) -- 
      variable tmp_var : std_logic_vector(41 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_2139_wire, MUX_2147_wire, tmp_var);
      CONCAT_u21_u42_2148_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u21_u42_2166_inst
    process(MUX_2157_wire, MUX_2165_wire) -- 
      variable tmp_var : std_logic_vector(41 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_2157_wire, MUX_2165_wire, tmp_var);
      CONCAT_u21_u42_2166_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u21_u42_2183_inst
    process(MUX_2174_wire, MUX_2182_wire) -- 
      variable tmp_var : std_logic_vector(41 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_2174_wire, MUX_2182_wire, tmp_var);
      CONCAT_u21_u42_2183_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u42_u84_2149_inst
    process(CONCAT_u21_u42_2131_wire, CONCAT_u21_u42_2148_wire) -- 
      variable tmp_var : std_logic_vector(83 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u21_u42_2131_wire, CONCAT_u21_u42_2148_wire, tmp_var);
      CONCAT_u42_u84_2149_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u42_u84_2184_inst
    process(CONCAT_u21_u42_2166_wire, CONCAT_u21_u42_2183_wire) -- 
      variable tmp_var : std_logic_vector(83 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u21_u42_2166_wire, CONCAT_u21_u42_2183_wire, tmp_var);
      CONCAT_u42_u84_2184_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u84_u168_2185_inst
    process(CONCAT_u42_u84_2149_wire, CONCAT_u42_u84_2184_wire) -- 
      variable tmp_var : std_logic_vector(167 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u42_u84_2149_wire, CONCAT_u42_u84_2184_wire, tmp_var);
      modified_set_tags_2186 <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_2118_inst
    process(access_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(access_index_buffer, konst_2117_wire_constant, tmp_var);
      EQ_u3_u1_2118_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_2126_inst
    process(access_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(access_index_buffer, konst_2125_wire_constant, tmp_var);
      EQ_u3_u1_2126_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_2135_inst
    process(access_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(access_index_buffer, konst_2134_wire_constant, tmp_var);
      EQ_u3_u1_2135_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_2143_inst
    process(access_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(access_index_buffer, konst_2142_wire_constant, tmp_var);
      EQ_u3_u1_2143_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_2153_inst
    process(access_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(access_index_buffer, konst_2152_wire_constant, tmp_var);
      EQ_u3_u1_2153_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_2161_inst
    process(access_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(access_index_buffer, konst_2160_wire_constant, tmp_var);
      EQ_u3_u1_2161_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_2170_inst
    process(access_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(access_index_buffer, konst_2169_wire_constant, tmp_var);
      EQ_u3_u1_2170_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_2178_inst
    process(access_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(access_index_buffer, konst_2177_wire_constant, tmp_var);
      EQ_u3_u1_2178_wire <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end updateSetTags_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library l2_cache_lib;
use l2_cache_lib.l2_cache_global_package.all;
entity updateSetValids_Volatile is -- 
  port ( -- 
    invalidate : in  std_logic_vector(0 downto 0);
    read_write_access : in  std_logic_vector(0 downto 0);
    set_valids : in  std_logic_vector(7 downto 0);
    access_index : in  std_logic_vector(2 downto 0);
    updated_set_valids : out  std_logic_vector(7 downto 0)-- 
  );
  -- 
end entity updateSetValids_Volatile;
architecture updateSetValids_Volatile_arch of updateSetValids_Volatile is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector(13-1 downto 0);
  signal default_zero_sig: std_logic;
  -- input port buffer signals
  signal invalidate_buffer :  std_logic_vector(0 downto 0);
  signal read_write_access_buffer :  std_logic_vector(0 downto 0);
  signal set_valids_buffer :  std_logic_vector(7 downto 0);
  signal access_index_buffer :  std_logic_vector(2 downto 0);
  -- output port buffer signals
  signal updated_set_valids_buffer :  std_logic_vector(7 downto 0);
  -- volatile/operator module components. 
  -- 
begin --  
  -- input handling ------------------------------------------------
  invalidate_buffer <= invalidate;
  read_write_access_buffer <= read_write_access;
  set_valids_buffer <= set_valids;
  access_index_buffer <= access_index;
  -- output handling  -------------------------------------------------------
  updated_set_valids <= updated_set_valids_buffer;
  -- the control path --------------------------------------------------
  default_zero_sig <= '0';
  -- volatile module, no control path
  -- the data path
  data_path: Block -- 
    signal AND_u1_u1_2002_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_2010_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_2019_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_2027_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_2037_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_2045_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_2054_wire : std_logic_vector(0 downto 0);
    signal AND_u1_u1_2062_wire : std_logic_vector(0 downto 0);
    signal CONCAT_u1_u2_2014_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_2031_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_2049_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u1_u2_2066_wire : std_logic_vector(1 downto 0);
    signal CONCAT_u2_u4_2032_wire : std_logic_vector(3 downto 0);
    signal CONCAT_u2_u4_2067_wire : std_logic_vector(3 downto 0);
    signal EQ_u3_u1_2001_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2009_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2018_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2026_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2036_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2044_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2053_wire : std_logic_vector(0 downto 0);
    signal EQ_u3_u1_2061_wire : std_logic_vector(0 downto 0);
    signal MUX_2005_wire : std_logic_vector(0 downto 0);
    signal MUX_2013_wire : std_logic_vector(0 downto 0);
    signal MUX_2022_wire : std_logic_vector(0 downto 0);
    signal MUX_2030_wire : std_logic_vector(0 downto 0);
    signal MUX_2040_wire : std_logic_vector(0 downto 0);
    signal MUX_2048_wire : std_logic_vector(0 downto 0);
    signal MUX_2057_wire : std_logic_vector(0 downto 0);
    signal MUX_2065_wire : std_logic_vector(0 downto 0);
    signal bitval_1959 : std_logic_vector(0 downto 0);
    signal insert_bit_1964 : std_logic_vector(0 downto 0);
    signal konst_2000_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2008_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2017_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2025_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2035_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2043_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2052_wire_constant : std_logic_vector(2 downto 0);
    signal konst_2060_wire_constant : std_logic_vector(2 downto 0);
    signal v0_1968 : std_logic_vector(0 downto 0);
    signal v1_1972 : std_logic_vector(0 downto 0);
    signal v2_1976 : std_logic_vector(0 downto 0);
    signal v3_1980 : std_logic_vector(0 downto 0);
    signal v4_1984 : std_logic_vector(0 downto 0);
    signal v5_1988 : std_logic_vector(0 downto 0);
    signal v6_1992 : std_logic_vector(0 downto 0);
    signal v7_1996 : std_logic_vector(0 downto 0);
    -- 
  begin -- 
    konst_2000_wire_constant <= "000";
    konst_2008_wire_constant <= "001";
    konst_2017_wire_constant <= "010";
    konst_2025_wire_constant <= "011";
    konst_2035_wire_constant <= "100";
    konst_2043_wire_constant <= "101";
    konst_2052_wire_constant <= "110";
    konst_2060_wire_constant <= "111";
    -- flow-through select operator MUX_2005_inst
    MUX_2005_wire <= bitval_1959 when (AND_u1_u1_2002_wire(0) /=  '0') else v0_1968;
    -- flow-through select operator MUX_2013_inst
    MUX_2013_wire <= bitval_1959 when (AND_u1_u1_2010_wire(0) /=  '0') else v1_1972;
    -- flow-through select operator MUX_2022_inst
    MUX_2022_wire <= bitval_1959 when (AND_u1_u1_2019_wire(0) /=  '0') else v2_1976;
    -- flow-through select operator MUX_2030_inst
    MUX_2030_wire <= bitval_1959 when (AND_u1_u1_2027_wire(0) /=  '0') else v3_1980;
    -- flow-through select operator MUX_2040_inst
    MUX_2040_wire <= bitval_1959 when (AND_u1_u1_2037_wire(0) /=  '0') else v4_1984;
    -- flow-through select operator MUX_2048_inst
    MUX_2048_wire <= bitval_1959 when (AND_u1_u1_2045_wire(0) /=  '0') else v5_1988;
    -- flow-through select operator MUX_2057_inst
    MUX_2057_wire <= bitval_1959 when (AND_u1_u1_2054_wire(0) /=  '0') else v6_1992;
    -- flow-through select operator MUX_2065_inst
    MUX_2065_wire <= bitval_1959 when (AND_u1_u1_2062_wire(0) /=  '0') else v7_1996;
    -- flow-through slice operator slice_1967_inst
    v0_1968 <= set_valids_buffer(7 downto 7);
    -- flow-through slice operator slice_1971_inst
    v1_1972 <= set_valids_buffer(6 downto 6);
    -- flow-through slice operator slice_1975_inst
    v2_1976 <= set_valids_buffer(5 downto 5);
    -- flow-through slice operator slice_1979_inst
    v3_1980 <= set_valids_buffer(4 downto 4);
    -- flow-through slice operator slice_1983_inst
    v4_1984 <= set_valids_buffer(3 downto 3);
    -- flow-through slice operator slice_1987_inst
    v5_1988 <= set_valids_buffer(2 downto 2);
    -- flow-through slice operator slice_1991_inst
    v6_1992 <= set_valids_buffer(1 downto 1);
    -- flow-through slice operator slice_1995_inst
    v7_1996 <= set_valids_buffer(0 downto 0);
    -- binary operator AND_u1_u1_2002_inst
    process(insert_bit_1964, EQ_u3_u1_2001_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(insert_bit_1964, EQ_u3_u1_2001_wire, tmp_var);
      AND_u1_u1_2002_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2010_inst
    process(insert_bit_1964, EQ_u3_u1_2009_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(insert_bit_1964, EQ_u3_u1_2009_wire, tmp_var);
      AND_u1_u1_2010_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2019_inst
    process(insert_bit_1964, EQ_u3_u1_2018_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(insert_bit_1964, EQ_u3_u1_2018_wire, tmp_var);
      AND_u1_u1_2019_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2027_inst
    process(insert_bit_1964, EQ_u3_u1_2026_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(insert_bit_1964, EQ_u3_u1_2026_wire, tmp_var);
      AND_u1_u1_2027_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2037_inst
    process(insert_bit_1964, EQ_u3_u1_2036_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(insert_bit_1964, EQ_u3_u1_2036_wire, tmp_var);
      AND_u1_u1_2037_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2045_inst
    process(insert_bit_1964, EQ_u3_u1_2044_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(insert_bit_1964, EQ_u3_u1_2044_wire, tmp_var);
      AND_u1_u1_2045_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2054_inst
    process(insert_bit_1964, EQ_u3_u1_2053_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(insert_bit_1964, EQ_u3_u1_2053_wire, tmp_var);
      AND_u1_u1_2054_wire <= tmp_var; --
    end process;
    -- binary operator AND_u1_u1_2062_inst
    process(insert_bit_1964, EQ_u3_u1_2061_wire) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntAnd_proc(insert_bit_1964, EQ_u3_u1_2061_wire, tmp_var);
      AND_u1_u1_2062_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_2014_inst
    process(MUX_2005_wire, MUX_2013_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_2005_wire, MUX_2013_wire, tmp_var);
      CONCAT_u1_u2_2014_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_2031_inst
    process(MUX_2022_wire, MUX_2030_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_2022_wire, MUX_2030_wire, tmp_var);
      CONCAT_u1_u2_2031_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_2049_inst
    process(MUX_2040_wire, MUX_2048_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_2040_wire, MUX_2048_wire, tmp_var);
      CONCAT_u1_u2_2049_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u1_u2_2066_inst
    process(MUX_2057_wire, MUX_2065_wire) -- 
      variable tmp_var : std_logic_vector(1 downto 0); -- 
    begin -- 
      ApConcat_proc(MUX_2057_wire, MUX_2065_wire, tmp_var);
      CONCAT_u1_u2_2066_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u2_u4_2032_inst
    process(CONCAT_u1_u2_2014_wire, CONCAT_u1_u2_2031_wire) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_2014_wire, CONCAT_u1_u2_2031_wire, tmp_var);
      CONCAT_u2_u4_2032_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u2_u4_2067_inst
    process(CONCAT_u1_u2_2049_wire, CONCAT_u1_u2_2066_wire) -- 
      variable tmp_var : std_logic_vector(3 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u1_u2_2049_wire, CONCAT_u1_u2_2066_wire, tmp_var);
      CONCAT_u2_u4_2067_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u4_u8_2068_inst
    process(CONCAT_u2_u4_2032_wire, CONCAT_u2_u4_2067_wire) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u2_u4_2032_wire, CONCAT_u2_u4_2067_wire, tmp_var);
      updated_set_valids_buffer <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_2001_inst
    process(access_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(access_index_buffer, konst_2000_wire_constant, tmp_var);
      EQ_u3_u1_2001_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_2009_inst
    process(access_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(access_index_buffer, konst_2008_wire_constant, tmp_var);
      EQ_u3_u1_2009_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_2018_inst
    process(access_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(access_index_buffer, konst_2017_wire_constant, tmp_var);
      EQ_u3_u1_2018_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_2026_inst
    process(access_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(access_index_buffer, konst_2025_wire_constant, tmp_var);
      EQ_u3_u1_2026_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_2036_inst
    process(access_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(access_index_buffer, konst_2035_wire_constant, tmp_var);
      EQ_u3_u1_2036_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_2044_inst
    process(access_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(access_index_buffer, konst_2043_wire_constant, tmp_var);
      EQ_u3_u1_2044_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_2053_inst
    process(access_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(access_index_buffer, konst_2052_wire_constant, tmp_var);
      EQ_u3_u1_2053_wire <= tmp_var; --
    end process;
    -- binary operator EQ_u3_u1_2061_inst
    process(access_index_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntEq_proc(access_index_buffer, konst_2060_wire_constant, tmp_var);
      EQ_u3_u1_2061_wire <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_1958_inst
    process(invalidate_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", invalidate_buffer, tmp_var);
      bitval_1959 <= tmp_var; -- 
    end process;
    -- binary operator OR_u1_u1_1963_inst
    process(invalidate_buffer, read_write_access_buffer) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      ApIntOr_proc(invalidate_buffer, read_write_access_buffer, tmp_var);
      insert_bit_1964 <= tmp_var; --
    end process;
    -- 
  end Block; -- data_path
  -- 
end updateSetValids_Volatile_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library l2_cache_lib;
use l2_cache_lib.l2_cache_global_package.all;
entity writeMemoryFromL2 is -- 
  generic (tag_length : integer); 
  port ( -- 
    release_lock : in  std_logic_vector(0 downto 0);
    do_write : in  std_logic_vector(0 downto 0);
    dirty_word_mask : in  std_logic_vector(7 downto 0);
    line_address : in  std_logic_vector(29 downto 0);
    wline : in  std_logic_vector(511 downto 0);
    sys_mem_lock_pipe_write_req : out  std_logic_vector(0 downto 0);
    sys_mem_lock_pipe_write_ack : in   std_logic_vector(0 downto 0);
    sys_mem_lock_pipe_write_data : out  std_logic_vector(0 downto 0);
    accessSysMem_call_reqs : out  std_logic_vector(0 downto 0);
    accessSysMem_call_acks : in   std_logic_vector(0 downto 0);
    accessSysMem_call_data : out  std_logic_vector(108 downto 0);
    accessSysMem_call_tag  :  out  std_logic_vector(0 downto 0);
    accessSysMem_return_reqs : out  std_logic_vector(0 downto 0);
    accessSysMem_return_acks : in   std_logic_vector(0 downto 0);
    accessSysMem_return_data : in   std_logic_vector(63 downto 0);
    accessSysMem_return_tag :  in   std_logic_vector(0 downto 0);
    tag_in: in std_logic_vector(tag_length-1 downto 0);
    tag_out: out std_logic_vector(tag_length-1 downto 0) ;
    clk : in std_logic;
    reset : in std_logic;
    start_req : in std_logic;
    start_ack : out std_logic;
    fin_req : in std_logic;
    fin_ack   : out std_logic-- 
  );
  -- 
end entity writeMemoryFromL2;
architecture writeMemoryFromL2_arch of writeMemoryFromL2 is -- 
  -- always true...
  signal always_true_symbol: Boolean;
  signal in_buffer_data_in, in_buffer_data_out: std_logic_vector((tag_length + 552)-1 downto 0);
  signal default_zero_sig: std_logic;
  signal in_buffer_write_req: std_logic;
  signal in_buffer_write_ack: std_logic;
  signal in_buffer_unload_req_symbol: Boolean;
  signal in_buffer_unload_ack_symbol: Boolean;
  signal out_buffer_data_in, out_buffer_data_out: std_logic_vector((tag_length + 0)-1 downto 0);
  signal out_buffer_read_req: std_logic;
  signal out_buffer_read_ack: std_logic;
  signal out_buffer_write_req_symbol: Boolean;
  signal out_buffer_write_ack_symbol: Boolean;
  signal tag_ub_out, tag_ilock_out: std_logic_vector(tag_length-1 downto 0);
  signal tag_push_req, tag_push_ack, tag_pop_req, tag_pop_ack: std_logic;
  signal tag_unload_req_symbol, tag_unload_ack_symbol, tag_write_req_symbol, tag_write_ack_symbol: Boolean;
  signal tag_ilock_write_req_symbol, tag_ilock_write_ack_symbol, tag_ilock_read_req_symbol, tag_ilock_read_ack_symbol: Boolean;
  signal start_req_sig, fin_req_sig, start_ack_sig, fin_ack_sig: std_logic; 
  signal input_sample_reenable_symbol: Boolean;
  -- input port buffer signals
  signal release_lock_buffer :  std_logic_vector(0 downto 0);
  signal release_lock_update_enable: Boolean;
  signal do_write_buffer :  std_logic_vector(0 downto 0);
  signal do_write_update_enable: Boolean;
  signal dirty_word_mask_buffer :  std_logic_vector(7 downto 0);
  signal dirty_word_mask_update_enable: Boolean;
  signal line_address_buffer :  std_logic_vector(29 downto 0);
  signal line_address_update_enable: Boolean;
  signal wline_buffer :  std_logic_vector(511 downto 0);
  signal wline_update_enable: Boolean;
  -- output port buffer signals
  signal writeMemoryFromL2_CP_3057_start: Boolean;
  signal writeMemoryFromL2_CP_3057_symbol: Boolean;
  -- volatile/operator module components. 
  component extractDword_Volatile is -- 
    port ( -- 
      dword_id : in  std_logic_vector(2 downto 0);
      cache_line : in  std_logic_vector(511 downto 0);
      dword : out  std_logic_vector(63 downto 0)-- 
    );
    -- 
  end component; 
  component accessSysMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      byte_mask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEM_TO_L2CACHE_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEM_TO_L2CACHE_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEM_TO_L2CACHE_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      L2CACHE_TO_MEM_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      L2CACHE_TO_MEM_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      L2CACHE_TO_MEM_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  component getNextDirtyOffset_Volatile is -- 
    port ( -- 
      first_time : in  std_logic_vector(0 downto 0);
      last_offset : in  std_logic_vector(2 downto 0);
      dirty_mask : in  std_logic_vector(7 downto 0);
      none_found : out  std_logic_vector(0 downto 0);
      current_offset : out  std_logic_vector(2 downto 0)-- 
    );
    -- 
  end component; 
  -- links between control-path and data-path
  signal WPIPE_sys_mem_lock_3325_inst_ack_1 : boolean;
  signal call_stmt_3311_call_ack_0 : boolean;
  signal offset_3285_3278_buf_req_0 : boolean;
  signal phi_stmt_3268_req_1 : boolean;
  signal if_stmt_3264_branch_req_0 : boolean;
  signal phi_stmt_3274_ack_0 : boolean;
  signal call_stmt_3311_call_ack_1 : boolean;
  signal WPIPE_sys_mem_lock_3325_inst_req_1 : boolean;
  signal if_stmt_3264_branch_ack_0 : boolean;
  signal phi_stmt_3268_ack_0 : boolean;
  signal call_stmt_3311_call_req_0 : boolean;
  signal if_stmt_3264_branch_ack_1 : boolean;
  signal phi_stmt_3268_req_0 : boolean;
  signal call_stmt_3311_call_req_1 : boolean;
  signal phi_stmt_3274_req_0 : boolean;
  signal offset_3285_3278_buf_ack_1 : boolean;
  signal phi_stmt_3274_req_1 : boolean;
  signal WPIPE_sys_mem_lock_3325_inst_ack_0 : boolean;
  signal offset_3285_3278_buf_req_1 : boolean;
  signal WPIPE_sys_mem_lock_3325_inst_req_0 : boolean;
  signal offset_3285_3278_buf_ack_0 : boolean;
  signal do_while_stmt_3266_branch_ack_1 : boolean;
  signal do_while_stmt_3266_branch_ack_0 : boolean;
  signal do_while_stmt_3266_branch_req_0 : boolean;
  -- 
begin --  
  -- input handling ------------------------------------------------
  in_buffer: UnloadBuffer -- 
    generic map(name => "writeMemoryFromL2_input_buffer", -- 
      buffer_size => 0,
      bypass_flag => true,
      data_width => tag_length + 552) -- 
    port map(write_req => in_buffer_write_req, -- 
      write_ack => in_buffer_write_ack, 
      write_data => in_buffer_data_in,
      unload_req => in_buffer_unload_req_symbol, 
      unload_ack => in_buffer_unload_ack_symbol, 
      read_data => in_buffer_data_out,
      clk => clk, reset => reset); -- 
  in_buffer_data_in(0 downto 0) <= release_lock;
  release_lock_buffer <= in_buffer_data_out(0 downto 0);
  in_buffer_data_in(1 downto 1) <= do_write;
  do_write_buffer <= in_buffer_data_out(1 downto 1);
  in_buffer_data_in(9 downto 2) <= dirty_word_mask;
  dirty_word_mask_buffer <= in_buffer_data_out(9 downto 2);
  in_buffer_data_in(39 downto 10) <= line_address;
  line_address_buffer <= in_buffer_data_out(39 downto 10);
  in_buffer_data_in(551 downto 40) <= wline;
  wline_buffer <= in_buffer_data_out(551 downto 40);
  in_buffer_data_in(tag_length + 551 downto 552) <= tag_in;
  tag_ub_out <= in_buffer_data_out(tag_length + 551 downto 552);
  in_buffer_write_req <= start_req;
  start_ack <= in_buffer_write_ack;
  in_buffer_unload_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 1,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 32) := "in_buffer_unload_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= in_buffer_unload_ack_symbol & input_sample_reenable_symbol;
    gj_in_buffer_unload_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => in_buffer_unload_req_symbol, clk => clk, reset => reset); --
  end block;
  -- join of all unload_ack_symbols.. used to trigger CP.
  writeMemoryFromL2_CP_3057_start <= in_buffer_unload_ack_symbol;
  -- output handling  -------------------------------------------------------
  out_buffer: ReceiveBuffer -- 
    generic map(name => "writeMemoryFromL2_out_buffer", -- 
      buffer_size => 0,
      full_rate => false,
      data_width => tag_length + 0) --
    port map(write_req => out_buffer_write_req_symbol, -- 
      write_ack => out_buffer_write_ack_symbol, 
      write_data => out_buffer_data_in,
      read_req => out_buffer_read_req, 
      read_ack => out_buffer_read_ack, 
      read_data => out_buffer_data_out,
      clk => clk, reset => reset); -- 
  out_buffer_data_in(tag_length-1 downto 0) <= tag_ilock_out;
  tag_out <= out_buffer_data_out(tag_length-1 downto 0);
  out_buffer_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 0);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 1,2 => 0);
    constant joinName: string(1 to 32) := "out_buffer_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeMemoryFromL2_CP_3057_symbol & out_buffer_write_ack_symbol & tag_ilock_read_ack_symbol;
    gj_out_buffer_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => out_buffer_write_req_symbol, clk => clk, reset => reset); --
  end block;
  -- write-to output-buffer produces  reenable input sampling
  input_sample_reenable_symbol <= out_buffer_write_ack_symbol;
  -- fin-req/ack level protocol..
  out_buffer_read_req <= fin_req;
  fin_ack <= out_buffer_read_ack;
  ----- tag-queue --------------------------------------------------
  -- interlock buffer for TAG.. to provide required buffering.
  tagIlock: InterlockBuffer -- 
    generic map(name => "tag-interlock-buffer", -- 
      buffer_size => 1,
      bypass_flag => false,
      in_data_width => tag_length,
      out_data_width => tag_length) -- 
    port map(write_req => tag_ilock_write_req_symbol, -- 
      write_ack => tag_ilock_write_ack_symbol, 
      write_data => tag_ub_out,
      read_req => tag_ilock_read_req_symbol, 
      read_ack => tag_ilock_read_ack_symbol, 
      read_data => tag_ilock_out, 
      clk => clk, reset => reset); -- 
  -- tag ilock-buffer control logic. 
  tag_ilock_write_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 1) := (0 => 1,1 => 1);
    constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
    constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
    constant joinName: string(1 to 31) := "tag_ilock_write_req_symbol_join"; 
    signal preds: BooleanArray(1 to 2); -- 
  begin -- 
    preds <= writeMemoryFromL2_CP_3057_start & tag_ilock_write_ack_symbol;
    gj_tag_ilock_write_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_write_req_symbol, clk => clk, reset => reset); --
  end block;
  tag_ilock_read_req_symbol_join: block -- 
    constant place_capacities: IntegerArray(0 to 2) := (0 => 1,1 => 1,2 => 1);
    constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 1,2 => 1);
    constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
    constant joinName: string(1 to 30) := "tag_ilock_read_req_symbol_join"; 
    signal preds: BooleanArray(1 to 3); -- 
  begin -- 
    preds <= writeMemoryFromL2_CP_3057_start & tag_ilock_read_ack_symbol & out_buffer_write_ack_symbol;
    gj_tag_ilock_read_req_symbol_join : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
      port map(preds => preds, symbol_out => tag_ilock_read_req_symbol, clk => clk, reset => reset); --
  end block;
  -- the control path --------------------------------------------------
  always_true_symbol <= true; 
  default_zero_sig <= '0';
  writeMemoryFromL2_CP_3057: Block -- control-path 
    signal writeMemoryFromL2_CP_3057_elements: BooleanArray(65 downto 0);
    -- 
  begin -- 
    writeMemoryFromL2_CP_3057_elements(0) <= writeMemoryFromL2_CP_3057_start;
    writeMemoryFromL2_CP_3057_symbol <= writeMemoryFromL2_CP_3057_elements(65);
    -- CP-element group 0:  branch  transition  place  output  bypass 
    -- CP-element group 0: predecessors 
    -- CP-element group 0: successors 
    -- CP-element group 0: 	2 
    -- CP-element group 0: 	3 
    -- CP-element group 0:  members (13) 
      -- CP-element group 0: 	 branch_block_stmt_3263/$entry
      -- CP-element group 0: 	 assign_stmt_3255_to_assign_stmt_3258/$exit
      -- CP-element group 0: 	 branch_block_stmt_3263/if_stmt_3264_eval_test/branch_req
      -- CP-element group 0: 	 branch_block_stmt_3263/if_stmt_3264_else_link/$entry
      -- CP-element group 0: 	 assign_stmt_3255_to_assign_stmt_3258/$entry
      -- CP-element group 0: 	 branch_block_stmt_3263/if_stmt_3264_if_link/$entry
      -- CP-element group 0: 	 $entry
      -- CP-element group 0: 	 branch_block_stmt_3263/R_do_write_3265_place
      -- CP-element group 0: 	 branch_block_stmt_3263/if_stmt_3264__entry__
      -- CP-element group 0: 	 branch_block_stmt_3263/if_stmt_3264_eval_test/$exit
      -- CP-element group 0: 	 branch_block_stmt_3263/if_stmt_3264_eval_test/$entry
      -- CP-element group 0: 	 branch_block_stmt_3263/if_stmt_3264_dead_link/$entry
      -- CP-element group 0: 	 branch_block_stmt_3263/branch_block_stmt_3263__entry__
      -- 
    branch_req_3077_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " branch_req_3077_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeMemoryFromL2_CP_3057_elements(0), ack => if_stmt_3264_branch_req_0); -- 
    -- CP-element group 1:  merge  transition  place  output  bypass 
    -- CP-element group 1: predecessors 
    -- CP-element group 1: 	3 
    -- CP-element group 1: 	4 
    -- CP-element group 1: successors 
    -- CP-element group 1: 	64 
    -- CP-element group 1:  members (7) 
      -- CP-element group 1: 	 assign_stmt_3328/$entry
      -- CP-element group 1: 	 branch_block_stmt_3263/$exit
      -- CP-element group 1: 	 assign_stmt_3328/WPIPE_sys_mem_lock_3325_Sample/req
      -- CP-element group 1: 	 assign_stmt_3328/WPIPE_sys_mem_lock_3325_Sample/$entry
      -- CP-element group 1: 	 branch_block_stmt_3263/if_stmt_3264__exit__
      -- CP-element group 1: 	 assign_stmt_3328/WPIPE_sys_mem_lock_3325_sample_start_
      -- CP-element group 1: 	 branch_block_stmt_3263/branch_block_stmt_3263__exit__
      -- 
    req_3222_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3222_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeMemoryFromL2_CP_3057_elements(1), ack => WPIPE_sys_mem_lock_3325_inst_req_0); -- 
    writeMemoryFromL2_CP_3057_elements(1) <= OrReduce(writeMemoryFromL2_CP_3057_elements(3) & writeMemoryFromL2_CP_3057_elements(4));
    -- CP-element group 2:  transition  place  input  bypass 
    -- CP-element group 2: predecessors 
    -- CP-element group 2: 	0 
    -- CP-element group 2: successors 
    -- CP-element group 2: 	5 
    -- CP-element group 2:  members (3) 
      -- CP-element group 2: 	 branch_block_stmt_3263/if_stmt_3264_if_link/$exit
      -- CP-element group 2: 	 branch_block_stmt_3263/if_stmt_3264_if_link/if_choice_transition
      -- CP-element group 2: 	 branch_block_stmt_3263/do_while_stmt_3266__entry__
      -- 
    if_choice_transition_3082_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 2_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3264_branch_ack_1, ack => writeMemoryFromL2_CP_3057_elements(2)); -- 
    -- CP-element group 3:  transition  input  bypass 
    -- CP-element group 3: predecessors 
    -- CP-element group 3: 	0 
    -- CP-element group 3: successors 
    -- CP-element group 3: 	1 
    -- CP-element group 3:  members (2) 
      -- CP-element group 3: 	 branch_block_stmt_3263/if_stmt_3264_else_link/else_choice_transition
      -- CP-element group 3: 	 branch_block_stmt_3263/if_stmt_3264_else_link/$exit
      -- 
    else_choice_transition_3086_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 3_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => if_stmt_3264_branch_ack_0, ack => writeMemoryFromL2_CP_3057_elements(3)); -- 
    -- CP-element group 4:  place  bypass 
    -- CP-element group 4: predecessors 
    -- CP-element group 4: 	63 
    -- CP-element group 4: successors 
    -- CP-element group 4: 	1 
    -- CP-element group 4:  members (1) 
      -- CP-element group 4: 	 branch_block_stmt_3263/do_while_stmt_3266__exit__
      -- 
    writeMemoryFromL2_CP_3057_elements(4) <= writeMemoryFromL2_CP_3057_elements(63);
    -- CP-element group 5:  transition  place  bypass  pipeline-parent 
    -- CP-element group 5: predecessors 
    -- CP-element group 5: 	2 
    -- CP-element group 5: successors 
    -- CP-element group 5: 	11 
    -- CP-element group 5:  members (2) 
      -- CP-element group 5: 	 branch_block_stmt_3263/do_while_stmt_3266/$entry
      -- CP-element group 5: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266__entry__
      -- 
    writeMemoryFromL2_CP_3057_elements(5) <= writeMemoryFromL2_CP_3057_elements(2);
    -- CP-element group 6:  merge  place  bypass  pipeline-parent 
    -- CP-element group 6: predecessors 
    -- CP-element group 6: successors 
    -- CP-element group 6: 	63 
    -- CP-element group 6:  members (1) 
      -- CP-element group 6: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266__exit__
      -- 
    -- Element group writeMemoryFromL2_CP_3057_elements(6) is bound as output of CP function.
    -- CP-element group 7:  merge  place  bypass  pipeline-parent 
    -- CP-element group 7: predecessors 
    -- CP-element group 7: successors 
    -- CP-element group 7: 	10 
    -- CP-element group 7:  members (1) 
      -- CP-element group 7: 	 branch_block_stmt_3263/do_while_stmt_3266/loop_back
      -- 
    -- Element group writeMemoryFromL2_CP_3057_elements(7) is bound as output of CP function.
    -- CP-element group 8:  branch  transition  place  bypass  pipeline-parent 
    -- CP-element group 8: predecessors 
    -- CP-element group 8: 	13 
    -- CP-element group 8: successors 
    -- CP-element group 8: 	61 
    -- CP-element group 8: 	62 
    -- CP-element group 8:  members (3) 
      -- CP-element group 8: 	 branch_block_stmt_3263/do_while_stmt_3266/condition_done
      -- CP-element group 8: 	 branch_block_stmt_3263/do_while_stmt_3266/loop_exit/$entry
      -- CP-element group 8: 	 branch_block_stmt_3263/do_while_stmt_3266/loop_taken/$entry
      -- 
    writeMemoryFromL2_CP_3057_elements(8) <= writeMemoryFromL2_CP_3057_elements(13);
    -- CP-element group 9:  branch  place  bypass  pipeline-parent 
    -- CP-element group 9: predecessors 
    -- CP-element group 9: 	60 
    -- CP-element group 9: successors 
    -- CP-element group 9:  members (1) 
      -- CP-element group 9: 	 branch_block_stmt_3263/do_while_stmt_3266/loop_body_done
      -- 
    writeMemoryFromL2_CP_3057_elements(9) <= writeMemoryFromL2_CP_3057_elements(60);
    -- CP-element group 10:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 10: predecessors 
    -- CP-element group 10: 	7 
    -- CP-element group 10: successors 
    -- CP-element group 10: 	23 
    -- CP-element group 10: 	42 
    -- CP-element group 10:  members (1) 
      -- CP-element group 10: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/back_edge_to_loop_body
      -- 
    writeMemoryFromL2_CP_3057_elements(10) <= writeMemoryFromL2_CP_3057_elements(7);
    -- CP-element group 11:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 11: predecessors 
    -- CP-element group 11: 	5 
    -- CP-element group 11: successors 
    -- CP-element group 11: 	25 
    -- CP-element group 11: 	44 
    -- CP-element group 11:  members (1) 
      -- CP-element group 11: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/first_time_through_loop_body
      -- 
    writeMemoryFromL2_CP_3057_elements(11) <= writeMemoryFromL2_CP_3057_elements(5);
    -- CP-element group 12:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 12: predecessors 
    -- CP-element group 12: successors 
    -- CP-element group 12: 	59 
    -- CP-element group 12: 	19 
    -- CP-element group 12: 	20 
    -- CP-element group 12: 	36 
    -- CP-element group 12: 	37 
    -- CP-element group 12:  members (2) 
      -- CP-element group 12: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/loop_body_start
      -- CP-element group 12: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/$entry
      -- 
    -- Element group writeMemoryFromL2_CP_3057_elements(12) is bound as output of CP function.
    -- CP-element group 13:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 13: predecessors 
    -- CP-element group 13: 	59 
    -- CP-element group 13: 	16 
    -- CP-element group 13: 	18 
    -- CP-element group 13: successors 
    -- CP-element group 13: 	8 
    -- CP-element group 13:  members (1) 
      -- CP-element group 13: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/condition_evaluated
      -- 
    condition_evaluated_3103_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " condition_evaluated_3103_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeMemoryFromL2_CP_3057_elements(13), ack => do_while_stmt_3266_branch_req_0); -- 
    writeMemoryFromL2_cp_element_group_13: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 15);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 0);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "writeMemoryFromL2_cp_element_group_13"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeMemoryFromL2_CP_3057_elements(59) & writeMemoryFromL2_CP_3057_elements(16) & writeMemoryFromL2_CP_3057_elements(18);
      gj_writeMemoryFromL2_cp_element_group_13 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeMemoryFromL2_CP_3057_elements(13), clk => clk, reset => reset); --
    end block;
    -- CP-element group 14:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 14: predecessors 
    -- CP-element group 14: 	19 
    -- CP-element group 14: 	36 
    -- CP-element group 14: marked-predecessors 
    -- CP-element group 14: 	18 
    -- CP-element group 14: successors 
    -- CP-element group 14: 	38 
    -- CP-element group 14:  members (2) 
      -- CP-element group 14: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/phi_stmt_3268_sample_start__ps
      -- CP-element group 14: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/aggregated_phi_sample_req
      -- 
    writeMemoryFromL2_cp_element_group_14: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 0);
      constant joinName: string(1 to 37) := "writeMemoryFromL2_cp_element_group_14"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeMemoryFromL2_CP_3057_elements(19) & writeMemoryFromL2_CP_3057_elements(36) & writeMemoryFromL2_CP_3057_elements(18);
      gj_writeMemoryFromL2_cp_element_group_14 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeMemoryFromL2_CP_3057_elements(14), clk => clk, reset => reset); --
    end block;
    -- CP-element group 15:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 15: predecessors 
    -- CP-element group 15: 	21 
    -- CP-element group 15: 	39 
    -- CP-element group 15: successors 
    -- CP-element group 15: 	60 
    -- CP-element group 15: 	16 
    -- CP-element group 15: marked-successors 
    -- CP-element group 15: 	19 
    -- CP-element group 15: 	36 
    -- CP-element group 15:  members (3) 
      -- CP-element group 15: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/phi_stmt_3274_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/phi_stmt_3268_sample_completed_
      -- CP-element group 15: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/aggregated_phi_sample_ack
      -- 
    writeMemoryFromL2_cp_element_group_15: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writeMemoryFromL2_cp_element_group_15"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeMemoryFromL2_CP_3057_elements(21) & writeMemoryFromL2_CP_3057_elements(39);
      gj_writeMemoryFromL2_cp_element_group_15 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeMemoryFromL2_CP_3057_elements(15), clk => clk, reset => reset); --
    end block;
    -- CP-element group 16:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 16: predecessors 
    -- CP-element group 16: 	15 
    -- CP-element group 16: successors 
    -- CP-element group 16: 	13 
    -- CP-element group 16:  members (1) 
      -- CP-element group 16: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/aggregated_phi_sample_ack_d
      -- 
    -- Element group writeMemoryFromL2_CP_3057_elements(16) is a control-delay.
    cp_element_16_delay: control_delay_element  generic map(name => " 16_delay", delay_value => 1)  port map(req => writeMemoryFromL2_CP_3057_elements(15), ack => writeMemoryFromL2_CP_3057_elements(16), clk => clk, reset =>reset);
    -- CP-element group 17:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 17: predecessors 
    -- CP-element group 17: 	20 
    -- CP-element group 17: 	37 
    -- CP-element group 17: successors 
    -- CP-element group 17: 	40 
    -- CP-element group 17:  members (2) 
      -- CP-element group 17: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/phi_stmt_3268_update_start__ps
      -- CP-element group 17: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/aggregated_phi_update_req
      -- 
    writeMemoryFromL2_cp_element_group_17: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writeMemoryFromL2_cp_element_group_17"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeMemoryFromL2_CP_3057_elements(20) & writeMemoryFromL2_CP_3057_elements(37);
      gj_writeMemoryFromL2_cp_element_group_17 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeMemoryFromL2_CP_3057_elements(17), clk => clk, reset => reset); --
    end block;
    -- CP-element group 18:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 18: predecessors 
    -- CP-element group 18: 	22 
    -- CP-element group 18: 	41 
    -- CP-element group 18: successors 
    -- CP-element group 18: 	13 
    -- CP-element group 18: marked-successors 
    -- CP-element group 18: 	14 
    -- CP-element group 18:  members (1) 
      -- CP-element group 18: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/aggregated_phi_update_ack
      -- 
    writeMemoryFromL2_cp_element_group_18: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writeMemoryFromL2_cp_element_group_18"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeMemoryFromL2_CP_3057_elements(22) & writeMemoryFromL2_CP_3057_elements(41);
      gj_writeMemoryFromL2_cp_element_group_18 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeMemoryFromL2_CP_3057_elements(18), clk => clk, reset => reset); --
    end block;
    -- CP-element group 19:  join  transition  bypass  pipeline-parent 
    -- CP-element group 19: predecessors 
    -- CP-element group 19: 	12 
    -- CP-element group 19: marked-predecessors 
    -- CP-element group 19: 	15 
    -- CP-element group 19: successors 
    -- CP-element group 19: 	14 
    -- CP-element group 19:  members (1) 
      -- CP-element group 19: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/phi_stmt_3268_sample_start_
      -- 
    writeMemoryFromL2_cp_element_group_19: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "writeMemoryFromL2_cp_element_group_19"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeMemoryFromL2_CP_3057_elements(12) & writeMemoryFromL2_CP_3057_elements(15);
      gj_writeMemoryFromL2_cp_element_group_19 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeMemoryFromL2_CP_3057_elements(19), clk => clk, reset => reset); --
    end block;
    -- CP-element group 20:  join  transition  bypass  pipeline-parent 
    -- CP-element group 20: predecessors 
    -- CP-element group 20: 	12 
    -- CP-element group 20: marked-predecessors 
    -- CP-element group 20: 	57 
    -- CP-element group 20: successors 
    -- CP-element group 20: 	17 
    -- CP-element group 20:  members (1) 
      -- CP-element group 20: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/phi_stmt_3268_update_start_
      -- 
    writeMemoryFromL2_cp_element_group_20: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writeMemoryFromL2_cp_element_group_20"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeMemoryFromL2_CP_3057_elements(12) & writeMemoryFromL2_CP_3057_elements(57);
      gj_writeMemoryFromL2_cp_element_group_20 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeMemoryFromL2_CP_3057_elements(20), clk => clk, reset => reset); --
    end block;
    -- CP-element group 21:  join  transition  bypass  pipeline-parent 
    -- CP-element group 21: predecessors 
    -- CP-element group 21: successors 
    -- CP-element group 21: 	15 
    -- CP-element group 21:  members (1) 
      -- CP-element group 21: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/phi_stmt_3268_sample_completed__ps
      -- 
    -- Element group writeMemoryFromL2_CP_3057_elements(21) is bound as output of CP function.
    -- CP-element group 22:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 22: predecessors 
    -- CP-element group 22: successors 
    -- CP-element group 22: 	55 
    -- CP-element group 22: 	18 
    -- CP-element group 22:  members (2) 
      -- CP-element group 22: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/phi_stmt_3268_update_completed__ps
      -- CP-element group 22: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/phi_stmt_3268_update_completed_
      -- 
    -- Element group writeMemoryFromL2_CP_3057_elements(22) is bound as output of CP function.
    -- CP-element group 23:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 23: predecessors 
    -- CP-element group 23: 	10 
    -- CP-element group 23: successors 
    -- CP-element group 23:  members (1) 
      -- CP-element group 23: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/phi_stmt_3268_loopback_trigger
      -- 
    writeMemoryFromL2_CP_3057_elements(23) <= writeMemoryFromL2_CP_3057_elements(10);
    -- CP-element group 24:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 24: predecessors 
    -- CP-element group 24: successors 
    -- CP-element group 24:  members (2) 
      -- CP-element group 24: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/phi_stmt_3268_loopback_sample_req
      -- CP-element group 24: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/phi_stmt_3268_loopback_sample_req_ps
      -- 
    phi_stmt_3268_loopback_sample_req_3119_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3268_loopback_sample_req_3119_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeMemoryFromL2_CP_3057_elements(24), ack => phi_stmt_3268_req_1); -- 
    -- Element group writeMemoryFromL2_CP_3057_elements(24) is bound as output of CP function.
    -- CP-element group 25:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 25: predecessors 
    -- CP-element group 25: 	11 
    -- CP-element group 25: successors 
    -- CP-element group 25:  members (1) 
      -- CP-element group 25: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/phi_stmt_3268_entry_trigger
      -- 
    writeMemoryFromL2_CP_3057_elements(25) <= writeMemoryFromL2_CP_3057_elements(11);
    -- CP-element group 26:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 26: predecessors 
    -- CP-element group 26: successors 
    -- CP-element group 26:  members (2) 
      -- CP-element group 26: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/phi_stmt_3268_entry_sample_req_ps
      -- CP-element group 26: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/phi_stmt_3268_entry_sample_req
      -- 
    phi_stmt_3268_entry_sample_req_3122_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3268_entry_sample_req_3122_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeMemoryFromL2_CP_3057_elements(26), ack => phi_stmt_3268_req_0); -- 
    -- Element group writeMemoryFromL2_CP_3057_elements(26) is bound as output of CP function.
    -- CP-element group 27:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 27: predecessors 
    -- CP-element group 27: successors 
    -- CP-element group 27:  members (2) 
      -- CP-element group 27: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/phi_stmt_3268_phi_mux_ack
      -- CP-element group 27: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/phi_stmt_3268_phi_mux_ack_ps
      -- 
    phi_stmt_3268_phi_mux_ack_3125_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 27_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3268_ack_0, ack => writeMemoryFromL2_CP_3057_elements(27)); -- 
    -- CP-element group 28:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 28: predecessors 
    -- CP-element group 28: successors 
    -- CP-element group 28:  members (4) 
      -- CP-element group 28: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/type_cast_3271_sample_completed__ps
      -- CP-element group 28: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/type_cast_3271_sample_start__ps
      -- CP-element group 28: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/type_cast_3271_sample_start_
      -- CP-element group 28: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/type_cast_3271_sample_completed_
      -- 
    -- Element group writeMemoryFromL2_CP_3057_elements(28) is bound as output of CP function.
    -- CP-element group 29:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 29: predecessors 
    -- CP-element group 29: successors 
    -- CP-element group 29: 	31 
    -- CP-element group 29:  members (2) 
      -- CP-element group 29: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/type_cast_3271_update_start__ps
      -- CP-element group 29: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/type_cast_3271_update_start_
      -- 
    -- Element group writeMemoryFromL2_CP_3057_elements(29) is bound as output of CP function.
    -- CP-element group 30:  join  transition  bypass  pipeline-parent 
    -- CP-element group 30: predecessors 
    -- CP-element group 30: 	31 
    -- CP-element group 30: successors 
    -- CP-element group 30:  members (1) 
      -- CP-element group 30: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/type_cast_3271_update_completed__ps
      -- 
    writeMemoryFromL2_CP_3057_elements(30) <= writeMemoryFromL2_CP_3057_elements(31);
    -- CP-element group 31:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 31: predecessors 
    -- CP-element group 31: 	29 
    -- CP-element group 31: successors 
    -- CP-element group 31: 	30 
    -- CP-element group 31:  members (1) 
      -- CP-element group 31: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/type_cast_3271_update_completed_
      -- 
    -- Element group writeMemoryFromL2_CP_3057_elements(31) is a control-delay.
    cp_element_31_delay: control_delay_element  generic map(name => " 31_delay", delay_value => 1)  port map(req => writeMemoryFromL2_CP_3057_elements(29), ack => writeMemoryFromL2_CP_3057_elements(31), clk => clk, reset =>reset);
    -- CP-element group 32:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 32: predecessors 
    -- CP-element group 32: successors 
    -- CP-element group 32:  members (4) 
      -- CP-element group 32: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/type_cast_3273_sample_completed__ps
      -- CP-element group 32: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/type_cast_3273_sample_start__ps
      -- CP-element group 32: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/type_cast_3273_sample_completed_
      -- CP-element group 32: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/type_cast_3273_sample_start_
      -- 
    -- Element group writeMemoryFromL2_CP_3057_elements(32) is bound as output of CP function.
    -- CP-element group 33:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 33: predecessors 
    -- CP-element group 33: successors 
    -- CP-element group 33: 	35 
    -- CP-element group 33:  members (2) 
      -- CP-element group 33: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/type_cast_3273_update_start__ps
      -- CP-element group 33: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/type_cast_3273_update_start_
      -- 
    -- Element group writeMemoryFromL2_CP_3057_elements(33) is bound as output of CP function.
    -- CP-element group 34:  join  transition  bypass  pipeline-parent 
    -- CP-element group 34: predecessors 
    -- CP-element group 34: 	35 
    -- CP-element group 34: successors 
    -- CP-element group 34:  members (1) 
      -- CP-element group 34: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/type_cast_3273_update_completed__ps
      -- 
    writeMemoryFromL2_CP_3057_elements(34) <= writeMemoryFromL2_CP_3057_elements(35);
    -- CP-element group 35:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 35: predecessors 
    -- CP-element group 35: 	33 
    -- CP-element group 35: successors 
    -- CP-element group 35: 	34 
    -- CP-element group 35:  members (1) 
      -- CP-element group 35: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/type_cast_3273_update_completed_
      -- 
    -- Element group writeMemoryFromL2_CP_3057_elements(35) is a control-delay.
    cp_element_35_delay: control_delay_element  generic map(name => " 35_delay", delay_value => 1)  port map(req => writeMemoryFromL2_CP_3057_elements(33), ack => writeMemoryFromL2_CP_3057_elements(35), clk => clk, reset =>reset);
    -- CP-element group 36:  join  transition  bypass  pipeline-parent 
    -- CP-element group 36: predecessors 
    -- CP-element group 36: 	12 
    -- CP-element group 36: marked-predecessors 
    -- CP-element group 36: 	15 
    -- CP-element group 36: successors 
    -- CP-element group 36: 	14 
    -- CP-element group 36:  members (1) 
      -- CP-element group 36: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/phi_stmt_3274_sample_start_
      -- 
    writeMemoryFromL2_cp_element_group_36: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 1);
      constant joinName: string(1 to 37) := "writeMemoryFromL2_cp_element_group_36"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeMemoryFromL2_CP_3057_elements(12) & writeMemoryFromL2_CP_3057_elements(15);
      gj_writeMemoryFromL2_cp_element_group_36 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeMemoryFromL2_CP_3057_elements(36), clk => clk, reset => reset); --
    end block;
    -- CP-element group 37:  join  transition  bypass  pipeline-parent 
    -- CP-element group 37: predecessors 
    -- CP-element group 37: 	12 
    -- CP-element group 37: marked-predecessors 
    -- CP-element group 37: 	57 
    -- CP-element group 37: successors 
    -- CP-element group 37: 	17 
    -- CP-element group 37:  members (1) 
      -- CP-element group 37: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/phi_stmt_3274_update_start_
      -- 
    writeMemoryFromL2_cp_element_group_37: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 1);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 1);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writeMemoryFromL2_cp_element_group_37"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeMemoryFromL2_CP_3057_elements(12) & writeMemoryFromL2_CP_3057_elements(57);
      gj_writeMemoryFromL2_cp_element_group_37 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeMemoryFromL2_CP_3057_elements(37), clk => clk, reset => reset); --
    end block;
    -- CP-element group 38:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 38: predecessors 
    -- CP-element group 38: 	14 
    -- CP-element group 38: successors 
    -- CP-element group 38:  members (1) 
      -- CP-element group 38: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/phi_stmt_3274_sample_start__ps
      -- 
    writeMemoryFromL2_CP_3057_elements(38) <= writeMemoryFromL2_CP_3057_elements(14);
    -- CP-element group 39:  join  transition  bypass  pipeline-parent 
    -- CP-element group 39: predecessors 
    -- CP-element group 39: successors 
    -- CP-element group 39: 	15 
    -- CP-element group 39:  members (1) 
      -- CP-element group 39: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/phi_stmt_3274_sample_completed__ps
      -- 
    -- Element group writeMemoryFromL2_CP_3057_elements(39) is bound as output of CP function.
    -- CP-element group 40:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 40: predecessors 
    -- CP-element group 40: 	17 
    -- CP-element group 40: successors 
    -- CP-element group 40:  members (1) 
      -- CP-element group 40: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/phi_stmt_3274_update_start__ps
      -- 
    writeMemoryFromL2_CP_3057_elements(40) <= writeMemoryFromL2_CP_3057_elements(17);
    -- CP-element group 41:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 41: predecessors 
    -- CP-element group 41: successors 
    -- CP-element group 41: 	55 
    -- CP-element group 41: 	18 
    -- CP-element group 41:  members (2) 
      -- CP-element group 41: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/phi_stmt_3274_update_completed__ps
      -- CP-element group 41: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/phi_stmt_3274_update_completed_
      -- 
    -- Element group writeMemoryFromL2_CP_3057_elements(41) is bound as output of CP function.
    -- CP-element group 42:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 42: predecessors 
    -- CP-element group 42: 	10 
    -- CP-element group 42: successors 
    -- CP-element group 42:  members (1) 
      -- CP-element group 42: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/phi_stmt_3274_loopback_trigger
      -- 
    writeMemoryFromL2_CP_3057_elements(42) <= writeMemoryFromL2_CP_3057_elements(10);
    -- CP-element group 43:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 43: predecessors 
    -- CP-element group 43: successors 
    -- CP-element group 43:  members (2) 
      -- CP-element group 43: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/phi_stmt_3274_loopback_sample_req_ps
      -- CP-element group 43: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/phi_stmt_3274_loopback_sample_req
      -- 
    phi_stmt_3274_loopback_sample_req_3153_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3274_loopback_sample_req_3153_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeMemoryFromL2_CP_3057_elements(43), ack => phi_stmt_3274_req_1); -- 
    -- Element group writeMemoryFromL2_CP_3057_elements(43) is bound as output of CP function.
    -- CP-element group 44:  fork  transition  bypass  pipeline-parent 
    -- CP-element group 44: predecessors 
    -- CP-element group 44: 	11 
    -- CP-element group 44: successors 
    -- CP-element group 44:  members (1) 
      -- CP-element group 44: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/phi_stmt_3274_entry_trigger
      -- 
    writeMemoryFromL2_CP_3057_elements(44) <= writeMemoryFromL2_CP_3057_elements(11);
    -- CP-element group 45:  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 45: predecessors 
    -- CP-element group 45: successors 
    -- CP-element group 45:  members (2) 
      -- CP-element group 45: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/phi_stmt_3274_entry_sample_req_ps
      -- CP-element group 45: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/phi_stmt_3274_entry_sample_req
      -- 
    phi_stmt_3274_entry_sample_req_3156_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " phi_stmt_3274_entry_sample_req_3156_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeMemoryFromL2_CP_3057_elements(45), ack => phi_stmt_3274_req_0); -- 
    -- Element group writeMemoryFromL2_CP_3057_elements(45) is bound as output of CP function.
    -- CP-element group 46:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 46: predecessors 
    -- CP-element group 46: successors 
    -- CP-element group 46:  members (2) 
      -- CP-element group 46: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/phi_stmt_3274_phi_mux_ack
      -- CP-element group 46: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/phi_stmt_3274_phi_mux_ack_ps
      -- 
    phi_stmt_3274_phi_mux_ack_3159_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 46_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => phi_stmt_3274_ack_0, ack => writeMemoryFromL2_CP_3057_elements(46)); -- 
    -- CP-element group 47:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 47: predecessors 
    -- CP-element group 47: successors 
    -- CP-element group 47:  members (4) 
      -- CP-element group 47: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/type_cast_3277_sample_completed__ps
      -- CP-element group 47: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/type_cast_3277_sample_start__ps
      -- CP-element group 47: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/type_cast_3277_sample_completed_
      -- CP-element group 47: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/type_cast_3277_sample_start_
      -- 
    -- Element group writeMemoryFromL2_CP_3057_elements(47) is bound as output of CP function.
    -- CP-element group 48:  join  fork  transition  bypass  pipeline-parent 
    -- CP-element group 48: predecessors 
    -- CP-element group 48: successors 
    -- CP-element group 48: 	50 
    -- CP-element group 48:  members (2) 
      -- CP-element group 48: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/type_cast_3277_update_start__ps
      -- CP-element group 48: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/type_cast_3277_update_start_
      -- 
    -- Element group writeMemoryFromL2_CP_3057_elements(48) is bound as output of CP function.
    -- CP-element group 49:  join  transition  bypass  pipeline-parent 
    -- CP-element group 49: predecessors 
    -- CP-element group 49: 	50 
    -- CP-element group 49: successors 
    -- CP-element group 49:  members (1) 
      -- CP-element group 49: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/type_cast_3277_update_completed__ps
      -- 
    writeMemoryFromL2_CP_3057_elements(49) <= writeMemoryFromL2_CP_3057_elements(50);
    -- CP-element group 50:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 50: predecessors 
    -- CP-element group 50: 	48 
    -- CP-element group 50: successors 
    -- CP-element group 50: 	49 
    -- CP-element group 50:  members (1) 
      -- CP-element group 50: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/type_cast_3277_update_completed_
      -- 
    -- Element group writeMemoryFromL2_CP_3057_elements(50) is a control-delay.
    cp_element_50_delay: control_delay_element  generic map(name => " 50_delay", delay_value => 1)  port map(req => writeMemoryFromL2_CP_3057_elements(48), ack => writeMemoryFromL2_CP_3057_elements(50), clk => clk, reset =>reset);
    -- CP-element group 51:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 51: predecessors 
    -- CP-element group 51: successors 
    -- CP-element group 51: 	53 
    -- CP-element group 51:  members (4) 
      -- CP-element group 51: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/R_offset_3278_Sample/req
      -- CP-element group 51: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/R_offset_3278_Sample/$entry
      -- CP-element group 51: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/R_offset_3278_sample_start_
      -- CP-element group 51: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/R_offset_3278_sample_start__ps
      -- 
    req_3180_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3180_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeMemoryFromL2_CP_3057_elements(51), ack => offset_3285_3278_buf_req_0); -- 
    -- Element group writeMemoryFromL2_CP_3057_elements(51) is bound as output of CP function.
    -- CP-element group 52:  join  fork  transition  output  bypass  pipeline-parent 
    -- CP-element group 52: predecessors 
    -- CP-element group 52: successors 
    -- CP-element group 52: 	54 
    -- CP-element group 52:  members (4) 
      -- CP-element group 52: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/R_offset_3278_Update/req
      -- CP-element group 52: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/R_offset_3278_Update/$entry
      -- CP-element group 52: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/R_offset_3278_update_start_
      -- CP-element group 52: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/R_offset_3278_update_start__ps
      -- 
    req_3185_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3185_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeMemoryFromL2_CP_3057_elements(52), ack => offset_3285_3278_buf_req_1); -- 
    -- Element group writeMemoryFromL2_CP_3057_elements(52) is bound as output of CP function.
    -- CP-element group 53:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 53: predecessors 
    -- CP-element group 53: 	51 
    -- CP-element group 53: successors 
    -- CP-element group 53:  members (4) 
      -- CP-element group 53: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/R_offset_3278_Sample/ack
      -- CP-element group 53: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/R_offset_3278_Sample/$exit
      -- CP-element group 53: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/R_offset_3278_sample_completed_
      -- CP-element group 53: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/R_offset_3278_sample_completed__ps
      -- 
    ack_3181_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 53_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => offset_3285_3278_buf_ack_0, ack => writeMemoryFromL2_CP_3057_elements(53)); -- 
    -- CP-element group 54:  join  transition  input  bypass  pipeline-parent 
    -- CP-element group 54: predecessors 
    -- CP-element group 54: 	52 
    -- CP-element group 54: successors 
    -- CP-element group 54:  members (4) 
      -- CP-element group 54: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/R_offset_3278_Update/ack
      -- CP-element group 54: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/R_offset_3278_Update/$exit
      -- CP-element group 54: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/R_offset_3278_update_completed_
      -- CP-element group 54: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/R_offset_3278_update_completed__ps
      -- 
    ack_3186_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 54_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => offset_3285_3278_buf_ack_1, ack => writeMemoryFromL2_CP_3057_elements(54)); -- 
    -- CP-element group 55:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 55: predecessors 
    -- CP-element group 55: 	22 
    -- CP-element group 55: 	41 
    -- CP-element group 55: marked-predecessors 
    -- CP-element group 55: 	57 
    -- CP-element group 55: successors 
    -- CP-element group 55: 	57 
    -- CP-element group 55:  members (3) 
      -- CP-element group 55: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/call_stmt_3311_Sample/crr
      -- CP-element group 55: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/call_stmt_3311_Sample/$entry
      -- CP-element group 55: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/call_stmt_3311_sample_start_
      -- 
    crr_3195_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " crr_3195_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeMemoryFromL2_CP_3057_elements(55), ack => call_stmt_3311_call_req_0); -- 
    writeMemoryFromL2_cp_element_group_55: block -- 
      constant place_capacities: IntegerArray(0 to 2) := (0 => 15,1 => 15,2 => 1);
      constant place_markings: IntegerArray(0 to 2)  := (0 => 0,1 => 0,2 => 1);
      constant place_delays: IntegerArray(0 to 2) := (0 => 0,1 => 0,2 => 1);
      constant joinName: string(1 to 37) := "writeMemoryFromL2_cp_element_group_55"; 
      signal preds: BooleanArray(1 to 3); -- 
    begin -- 
      preds <= writeMemoryFromL2_CP_3057_elements(22) & writeMemoryFromL2_CP_3057_elements(41) & writeMemoryFromL2_CP_3057_elements(57);
      gj_writeMemoryFromL2_cp_element_group_55 : generic_join generic map(name => joinName, number_of_predecessors => 3, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeMemoryFromL2_CP_3057_elements(55), clk => clk, reset => reset); --
    end block;
    -- CP-element group 56:  join  transition  output  bypass  pipeline-parent 
    -- CP-element group 56: predecessors 
    -- CP-element group 56: marked-predecessors 
    -- CP-element group 56: 	58 
    -- CP-element group 56: successors 
    -- CP-element group 56: 	58 
    -- CP-element group 56:  members (3) 
      -- CP-element group 56: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/call_stmt_3311_update_start_
      -- CP-element group 56: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/call_stmt_3311_Update/ccr
      -- CP-element group 56: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/call_stmt_3311_Update/$entry
      -- 
    ccr_3200_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " ccr_3200_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeMemoryFromL2_CP_3057_elements(56), ack => call_stmt_3311_call_req_1); -- 
    writeMemoryFromL2_cp_element_group_56: block -- 
      constant place_capacities: IntegerArray(0 to 0) := (0 => 1);
      constant place_markings: IntegerArray(0 to 0)  := (0 => 1);
      constant place_delays: IntegerArray(0 to 0) := (0 => 0);
      constant joinName: string(1 to 37) := "writeMemoryFromL2_cp_element_group_56"; 
      signal preds: BooleanArray(1 to 1); -- 
    begin -- 
      preds(1) <= writeMemoryFromL2_CP_3057_elements(58);
      gj_writeMemoryFromL2_cp_element_group_56 : generic_join generic map(name => joinName, number_of_predecessors => 1, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeMemoryFromL2_CP_3057_elements(56), clk => clk, reset => reset); --
    end block;
    -- CP-element group 57:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 57: predecessors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: successors 
    -- CP-element group 57: marked-successors 
    -- CP-element group 57: 	55 
    -- CP-element group 57: 	20 
    -- CP-element group 57: 	37 
    -- CP-element group 57:  members (3) 
      -- CP-element group 57: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/call_stmt_3311_Sample/$exit
      -- CP-element group 57: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/call_stmt_3311_Sample/cra
      -- CP-element group 57: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/call_stmt_3311_sample_completed_
      -- 
    cra_3196_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 57_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_3311_call_ack_0, ack => writeMemoryFromL2_CP_3057_elements(57)); -- 
    -- CP-element group 58:  fork  transition  input  bypass  pipeline-parent 
    -- CP-element group 58: predecessors 
    -- CP-element group 58: 	56 
    -- CP-element group 58: successors 
    -- CP-element group 58: 	60 
    -- CP-element group 58: marked-successors 
    -- CP-element group 58: 	56 
    -- CP-element group 58:  members (3) 
      -- CP-element group 58: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/call_stmt_3311_Update/cca
      -- CP-element group 58: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/call_stmt_3311_update_completed_
      -- CP-element group 58: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/call_stmt_3311_Update/$exit
      -- 
    cca_3201_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 58_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => call_stmt_3311_call_ack_1, ack => writeMemoryFromL2_CP_3057_elements(58)); -- 
    -- CP-element group 59:  transition  delay-element  bypass  pipeline-parent 
    -- CP-element group 59: predecessors 
    -- CP-element group 59: 	12 
    -- CP-element group 59: successors 
    -- CP-element group 59: 	13 
    -- CP-element group 59:  members (1) 
      -- CP-element group 59: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/loop_body_delay_to_condition_start
      -- 
    -- Element group writeMemoryFromL2_CP_3057_elements(59) is a control-delay.
    cp_element_59_delay: control_delay_element  generic map(name => " 59_delay", delay_value => 1)  port map(req => writeMemoryFromL2_CP_3057_elements(12), ack => writeMemoryFromL2_CP_3057_elements(59), clk => clk, reset =>reset);
    -- CP-element group 60:  join  transition  bypass  pipeline-parent 
    -- CP-element group 60: predecessors 
    -- CP-element group 60: 	58 
    -- CP-element group 60: 	15 
    -- CP-element group 60: successors 
    -- CP-element group 60: 	9 
    -- CP-element group 60:  members (1) 
      -- CP-element group 60: 	 branch_block_stmt_3263/do_while_stmt_3266/do_while_stmt_3266_loop_body/$exit
      -- 
    writeMemoryFromL2_cp_element_group_60: block -- 
      constant place_capacities: IntegerArray(0 to 1) := (0 => 15,1 => 15);
      constant place_markings: IntegerArray(0 to 1)  := (0 => 0,1 => 0);
      constant place_delays: IntegerArray(0 to 1) := (0 => 0,1 => 0);
      constant joinName: string(1 to 37) := "writeMemoryFromL2_cp_element_group_60"; 
      signal preds: BooleanArray(1 to 2); -- 
    begin -- 
      preds <= writeMemoryFromL2_CP_3057_elements(58) & writeMemoryFromL2_CP_3057_elements(15);
      gj_writeMemoryFromL2_cp_element_group_60 : generic_join generic map(name => joinName, number_of_predecessors => 2, place_capacities => place_capacities, place_markings => place_markings, place_delays => place_delays) -- 
        port map(preds => preds, symbol_out => writeMemoryFromL2_CP_3057_elements(60), clk => clk, reset => reset); --
    end block;
    -- CP-element group 61:  transition  input  bypass  pipeline-parent 
    -- CP-element group 61: predecessors 
    -- CP-element group 61: 	8 
    -- CP-element group 61: successors 
    -- CP-element group 61:  members (2) 
      -- CP-element group 61: 	 branch_block_stmt_3263/do_while_stmt_3266/loop_exit/$exit
      -- CP-element group 61: 	 branch_block_stmt_3263/do_while_stmt_3266/loop_exit/ack
      -- 
    ack_3206_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 61_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_3266_branch_ack_0, ack => writeMemoryFromL2_CP_3057_elements(61)); -- 
    -- CP-element group 62:  transition  input  bypass  pipeline-parent 
    -- CP-element group 62: predecessors 
    -- CP-element group 62: 	8 
    -- CP-element group 62: successors 
    -- CP-element group 62:  members (2) 
      -- CP-element group 62: 	 branch_block_stmt_3263/do_while_stmt_3266/loop_taken/ack
      -- CP-element group 62: 	 branch_block_stmt_3263/do_while_stmt_3266/loop_taken/$exit
      -- 
    ack_3210_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 62_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => do_while_stmt_3266_branch_ack_1, ack => writeMemoryFromL2_CP_3057_elements(62)); -- 
    -- CP-element group 63:  transition  bypass  pipeline-parent 
    -- CP-element group 63: predecessors 
    -- CP-element group 63: 	6 
    -- CP-element group 63: successors 
    -- CP-element group 63: 	4 
    -- CP-element group 63:  members (1) 
      -- CP-element group 63: 	 branch_block_stmt_3263/do_while_stmt_3266/$exit
      -- 
    writeMemoryFromL2_CP_3057_elements(63) <= writeMemoryFromL2_CP_3057_elements(6);
    -- CP-element group 64:  transition  input  output  bypass 
    -- CP-element group 64: predecessors 
    -- CP-element group 64: 	1 
    -- CP-element group 64: successors 
    -- CP-element group 64: 	65 
    -- CP-element group 64:  members (6) 
      -- CP-element group 64: 	 assign_stmt_3328/WPIPE_sys_mem_lock_3325_Update/req
      -- CP-element group 64: 	 assign_stmt_3328/WPIPE_sys_mem_lock_3325_Update/$entry
      -- CP-element group 64: 	 assign_stmt_3328/WPIPE_sys_mem_lock_3325_Sample/ack
      -- CP-element group 64: 	 assign_stmt_3328/WPIPE_sys_mem_lock_3325_Sample/$exit
      -- CP-element group 64: 	 assign_stmt_3328/WPIPE_sys_mem_lock_3325_update_start_
      -- CP-element group 64: 	 assign_stmt_3328/WPIPE_sys_mem_lock_3325_sample_completed_
      -- 
    ack_3223_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 64_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_sys_mem_lock_3325_inst_ack_0, ack => writeMemoryFromL2_CP_3057_elements(64)); -- 
    req_3227_symbol_link_to_dp: control_delay_element -- 
      generic map(name => " req_3227_symbol_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => writeMemoryFromL2_CP_3057_elements(64), ack => WPIPE_sys_mem_lock_3325_inst_req_1); -- 
    -- CP-element group 65:  transition  input  bypass 
    -- CP-element group 65: predecessors 
    -- CP-element group 65: 	64 
    -- CP-element group 65: successors 
    -- CP-element group 65:  members (5) 
      -- CP-element group 65: 	 assign_stmt_3328/$exit
      -- CP-element group 65: 	 assign_stmt_3328/WPIPE_sys_mem_lock_3325_Update/ack
      -- CP-element group 65: 	 $exit
      -- CP-element group 65: 	 assign_stmt_3328/WPIPE_sys_mem_lock_3325_Update/$exit
      -- CP-element group 65: 	 assign_stmt_3328/WPIPE_sys_mem_lock_3325_update_completed_
      -- 
    ack_3228_symbol_link_from_dp: control_delay_element -- 
      generic map(name => " 65_delay",delay_value => 0)
      port map(clk => clk, reset => reset, req => WPIPE_sys_mem_lock_3325_inst_ack_1, ack => writeMemoryFromL2_CP_3057_elements(65)); -- 
    writeMemoryFromL2_do_while_stmt_3266_terminator_3211: loop_terminator -- 
      generic map (name => " writeMemoryFromL2_do_while_stmt_3266_terminator_3211", max_iterations_in_flight =>15) 
      port map(loop_body_exit => writeMemoryFromL2_CP_3057_elements(9),loop_continue => writeMemoryFromL2_CP_3057_elements(62),loop_terminate => writeMemoryFromL2_CP_3057_elements(61),loop_back => writeMemoryFromL2_CP_3057_elements(7),loop_exit => writeMemoryFromL2_CP_3057_elements(6),clk => clk, reset => reset); -- 
    phi_stmt_3268_phi_seq_3143_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= writeMemoryFromL2_CP_3057_elements(25);
      writeMemoryFromL2_CP_3057_elements(28)<= src_sample_reqs(0);
      src_sample_acks(0)  <= writeMemoryFromL2_CP_3057_elements(28);
      writeMemoryFromL2_CP_3057_elements(29)<= src_update_reqs(0);
      src_update_acks(0)  <= writeMemoryFromL2_CP_3057_elements(30);
      writeMemoryFromL2_CP_3057_elements(26) <= phi_mux_reqs(0);
      triggers(1)  <= writeMemoryFromL2_CP_3057_elements(23);
      writeMemoryFromL2_CP_3057_elements(32)<= src_sample_reqs(1);
      src_sample_acks(1)  <= writeMemoryFromL2_CP_3057_elements(32);
      writeMemoryFromL2_CP_3057_elements(33)<= src_update_reqs(1);
      src_update_acks(1)  <= writeMemoryFromL2_CP_3057_elements(34);
      writeMemoryFromL2_CP_3057_elements(24) <= phi_mux_reqs(1);
      phi_stmt_3268_phi_seq_3143 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_3268_phi_seq_3143") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => writeMemoryFromL2_CP_3057_elements(14), 
          phi_sample_ack => writeMemoryFromL2_CP_3057_elements(21), 
          phi_update_req => writeMemoryFromL2_CP_3057_elements(17), 
          phi_update_ack => writeMemoryFromL2_CP_3057_elements(22), 
          phi_mux_ack => writeMemoryFromL2_CP_3057_elements(27), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    phi_stmt_3274_phi_seq_3187_block : block -- 
      signal triggers, src_sample_reqs, src_sample_acks, src_update_reqs, src_update_acks : BooleanArray(0 to 1);
      signal phi_mux_reqs : BooleanArray(0 to 1); -- 
    begin -- 
      triggers(0)  <= writeMemoryFromL2_CP_3057_elements(44);
      writeMemoryFromL2_CP_3057_elements(47)<= src_sample_reqs(0);
      src_sample_acks(0)  <= writeMemoryFromL2_CP_3057_elements(47);
      writeMemoryFromL2_CP_3057_elements(48)<= src_update_reqs(0);
      src_update_acks(0)  <= writeMemoryFromL2_CP_3057_elements(49);
      writeMemoryFromL2_CP_3057_elements(45) <= phi_mux_reqs(0);
      triggers(1)  <= writeMemoryFromL2_CP_3057_elements(42);
      writeMemoryFromL2_CP_3057_elements(51)<= src_sample_reqs(1);
      src_sample_acks(1)  <= writeMemoryFromL2_CP_3057_elements(53);
      writeMemoryFromL2_CP_3057_elements(52)<= src_update_reqs(1);
      src_update_acks(1)  <= writeMemoryFromL2_CP_3057_elements(54);
      writeMemoryFromL2_CP_3057_elements(43) <= phi_mux_reqs(1);
      phi_stmt_3274_phi_seq_3187 : phi_sequencer_v2-- 
        generic map (place_capacity => 15, ntriggers => 2, name => "phi_stmt_3274_phi_seq_3187") 
        port map ( -- 
          triggers => triggers, src_sample_starts => src_sample_reqs, 
          src_sample_completes => src_sample_acks, src_update_starts => src_update_reqs, 
          src_update_completes => src_update_acks,
          phi_mux_select_reqs => phi_mux_reqs, 
          phi_sample_req => writeMemoryFromL2_CP_3057_elements(38), 
          phi_sample_ack => writeMemoryFromL2_CP_3057_elements(39), 
          phi_update_req => writeMemoryFromL2_CP_3057_elements(40), 
          phi_update_ack => writeMemoryFromL2_CP_3057_elements(41), 
          phi_mux_ack => writeMemoryFromL2_CP_3057_elements(46), 
          clk => clk, reset => reset -- 
        );
        -- 
    end block;
    entry_tmerge_3104_block : block -- 
      signal preds : BooleanArray(0 to 1);
      begin -- 
        preds(0)  <= writeMemoryFromL2_CP_3057_elements(10);
        preds(1)  <= writeMemoryFromL2_CP_3057_elements(11);
        entry_tmerge_3104 : transition_merge -- 
          generic map(name => " entry_tmerge_3104")
          port map (preds => preds, symbol_out => writeMemoryFromL2_CP_3057_elements(12));
          -- 
    end block;
    --  hookup: inputs to control-path 
    -- hookup: output from control-path 
    -- 
  end Block; -- control-path
  -- the data path
  data_path: Block -- 
    signal CONCAT_u30_u33_3297_wire : std_logic_vector(32 downto 0);
    signal NOT_u8_u8_3307_wire_constant : std_logic_vector(7 downto 0);
    signal continue_flag_3289 : std_logic_vector(0 downto 0);
    signal dirty_word_mask_qualified_3258 : std_logic_vector(7 downto 0);
    signal first_time_3268 : std_logic_vector(0 downto 0);
    signal last_offset_3274 : std_logic_vector(2 downto 0);
    signal none_found_3285 : std_logic_vector(0 downto 0);
    signal offset_3285 : std_logic_vector(2 downto 0);
    signal offset_3285_3278_buffered : std_logic_vector(2 downto 0);
    signal pa_3301 : std_logic_vector(35 downto 0);
    signal pa_base_3255 : std_logic_vector(35 downto 0);
    signal rval_3311 : std_logic_vector(63 downto 0);
    signal type_cast_3253_wire_constant : std_logic_vector(5 downto 0);
    signal type_cast_3271_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_3273_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_3277_wire_constant : std_logic_vector(2 downto 0);
    signal type_cast_3299_wire_constant : std_logic_vector(2 downto 0);
    signal type_cast_3304_wire_constant : std_logic_vector(0 downto 0);
    signal type_cast_3327_wire_constant : std_logic_vector(0 downto 0);
    signal wdata_3293 : std_logic_vector(63 downto 0);
    -- 
  begin -- 
    NOT_u8_u8_3307_wire_constant <= "11111111";
    type_cast_3253_wire_constant <= "000000";
    type_cast_3271_wire_constant <= "1";
    type_cast_3273_wire_constant <= "0";
    type_cast_3277_wire_constant <= "000";
    type_cast_3299_wire_constant <= "000";
    type_cast_3304_wire_constant <= "0";
    type_cast_3327_wire_constant <= "1";
    phi_stmt_3268: Block -- phi operator 
      signal idata: std_logic_vector(1 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3271_wire_constant & type_cast_3273_wire_constant;
      req <= phi_stmt_3268_req_0 & phi_stmt_3268_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3268",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 1) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3268_ack_0,
          idata => idata,
          odata => first_time_3268,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3268
    phi_stmt_3274: Block -- phi operator 
      signal idata: std_logic_vector(5 downto 0);
      signal req: BooleanArray(1 downto 0);
      --
    begin -- 
      idata <= type_cast_3277_wire_constant & offset_3285_3278_buffered;
      req <= phi_stmt_3274_req_0 & phi_stmt_3274_req_1;
      phi: PhiBase -- 
        generic map( -- 
          name => "phi_stmt_3274",
          num_reqs => 2,
          bypass_flag => true,
          data_width => 3) -- 
        port map( -- 
          req => req, 
          ack => phi_stmt_3274_ack_0,
          idata => idata,
          odata => last_offset_3274,
          clk => clk,
          reset => reset ); -- 
      -- 
    end Block; -- phi operator phi_stmt_3274
    -- interlock W_dirty_word_mask_qualified_3256_inst
    process(dirty_word_mask_buffer) -- 
      variable tmp_var : std_logic_vector(7 downto 0); -- 
    begin -- 
      tmp_var := (others => '0'); 
      tmp_var( 7 downto 0) := dirty_word_mask_buffer(7 downto 0);
      dirty_word_mask_qualified_3258 <= tmp_var; -- 
    end process;
    offset_3285_3278_buf_block: block -- 
      signal wreq, wack, rreq, rack: BooleanArray(0 downto 0); 
      -- 
    begin -- 
      wreq(0) <= offset_3285_3278_buf_req_0;
      offset_3285_3278_buf_ack_0<= wack(0);
      rreq(0) <= offset_3285_3278_buf_req_1;
      offset_3285_3278_buf_ack_1<= rack(0);
      offset_3285_3278_buf : InterlockBuffer generic map ( -- 
        name => "offset_3285_3278_buf",
        buffer_size => 1,
        flow_through =>  false ,
        cut_through =>  false ,
        in_data_width => 3,
        out_data_width => 3,
        bypass_flag =>  false 
        -- 
      )port map ( -- 
        write_req => wreq(0), 
        write_ack => wack(0), 
        write_data => offset_3285,
        read_req => rreq(0),  
        read_ack => rack(0), 
        read_data => offset_3285_3278_buffered,
        clk => clk, reset => reset
        -- 
      );
      end block; -- 
    do_while_stmt_3266_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= continue_flag_3289;
      branch_instance: BranchBase -- 
        generic map( name => "do_while_stmt_3266_branch", condition_width => 1,  bypass_flag => true)
        port map( -- 
          condition => condition_sig,
          req => do_while_stmt_3266_branch_req_0,
          ack0 => do_while_stmt_3266_branch_ack_0,
          ack1 => do_while_stmt_3266_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    if_stmt_3264_branch: Block -- 
      -- branch-block
      signal condition_sig : std_logic_vector(0 downto 0);
      begin 
      condition_sig <= do_write_buffer;
      branch_instance: BranchBase -- 
        generic map( name => "if_stmt_3264_branch", condition_width => 1,  bypass_flag => false)
        port map( -- 
          condition => condition_sig,
          req => if_stmt_3264_branch_req_0,
          ack0 => if_stmt_3264_branch_ack_0,
          ack1 => if_stmt_3264_branch_ack_1,
          clk => clk,
          reset => reset); -- 
      --
    end Block; -- branch-block
    -- binary operator CONCAT_u30_u33_3297_inst
    process(line_address_buffer, offset_3285) -- 
      variable tmp_var : std_logic_vector(32 downto 0); -- 
    begin -- 
      ApConcat_proc(line_address_buffer, offset_3285, tmp_var);
      CONCAT_u30_u33_3297_wire <= tmp_var; --
    end process;
    -- binary operator CONCAT_u30_u36_3254_inst
    process(line_address_buffer) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(line_address_buffer, type_cast_3253_wire_constant, tmp_var);
      pa_base_3255 <= tmp_var; --
    end process;
    -- binary operator CONCAT_u33_u36_3300_inst
    process(CONCAT_u30_u33_3297_wire) -- 
      variable tmp_var : std_logic_vector(35 downto 0); -- 
    begin -- 
      ApConcat_proc(CONCAT_u30_u33_3297_wire, type_cast_3299_wire_constant, tmp_var);
      pa_3301 <= tmp_var; --
    end process;
    -- unary operator NOT_u1_u1_3288_inst
    process(none_found_3285) -- 
      variable tmp_var : std_logic_vector(0 downto 0); -- 
    begin -- 
      SingleInputOperation("ApIntNot", none_found_3285, tmp_var);
      continue_flag_3289 <= tmp_var; -- 
    end process;
    -- shared outport operator group (0) : WPIPE_sys_mem_lock_3325_inst 
    OutportGroup_0: Block -- 
      signal data_in: std_logic_vector(0 downto 0);
      signal sample_req, sample_ack : BooleanArray( 0 downto 0);
      signal update_req, update_ack : BooleanArray( 0 downto 0);
      signal sample_req_unguarded, sample_ack_unguarded : BooleanArray( 0 downto 0);
      signal update_req_unguarded, update_ack_unguarded : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 0);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 2);
      -- 
    begin -- 
      sample_req_unguarded(0) <= WPIPE_sys_mem_lock_3325_inst_req_0;
      WPIPE_sys_mem_lock_3325_inst_ack_0 <= sample_ack_unguarded(0);
      update_req_unguarded(0) <= WPIPE_sys_mem_lock_3325_inst_req_1;
      WPIPE_sys_mem_lock_3325_inst_ack_1 <= update_ack_unguarded(0);
      guard_vector(0)  <= release_lock_buffer(0);
      data_in <= type_cast_3327_wire_constant;
      sys_mem_lock_write_0_gI: SplitGuardInterface generic map(name => "sys_mem_lock_write_0_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => true,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => sample_req_unguarded,
        sr_out => sample_req,
        sa_in => sample_ack,
        sa_out => sample_ack_unguarded,
        cr_in => update_req_unguarded,
        cr_out => update_req,
        ca_in => update_ack,
        ca_out => update_ack_unguarded,
        guards => guard_vector); -- 
      sys_mem_lock_write_0: OutputPortRevised -- 
        generic map ( name => "sys_mem_lock", data_width => 1, num_reqs => 1, input_buffering => inBUFs, full_rate => false,
        no_arbitration => false)
        port map (--
          sample_req => sample_req , 
          sample_ack => sample_ack , 
          update_req => update_req , 
          update_ack => update_ack , 
          data => data_in, 
          oreq => sys_mem_lock_pipe_write_req(0),
          oack => sys_mem_lock_pipe_write_ack(0),
          odata => sys_mem_lock_pipe_write_data(0 downto 0),
          clk => clk, reset => reset -- 
        );-- 
      -- 
    end Block; -- outport group 0
    volatile_operator_getNextDirtyOffset_6078: getNextDirtyOffset_Volatile port map(first_time => first_time_3268, last_offset => last_offset_3274, dirty_mask => dirty_word_mask_qualified_3258, none_found => none_found_3285, current_offset => offset_3285); 
    volatile_operator_extractDword_6080: extractDword_Volatile port map(dword_id => offset_3285, cache_line => wline_buffer, dword => wdata_3293); 
    -- shared call operator group (2) : call_stmt_3311_call 
    accessSysMem_call_group_2: Block -- 
      signal data_in: std_logic_vector(108 downto 0);
      signal data_out: std_logic_vector(63 downto 0);
      signal reqR, ackR, reqL, ackL : BooleanArray( 0 downto 0);
      signal reqR_unguarded, ackR_unguarded, reqL_unguarded, ackL_unguarded : BooleanArray( 0 downto 0);
      signal reqL_unregulated, ackL_unregulated : BooleanArray( 0 downto 0);
      signal guard_vector : std_logic_vector( 0 downto 0);
      constant inBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant outBUFs : IntegerArray(0 downto 0) := (0 => 1);
      constant guardFlags : BooleanArray(0 downto 0) := (0 => true);
      constant guardBuffering: IntegerArray(0 downto 0)  := (0 => 8);
      -- 
    begin -- 
      reqL_unguarded(0) <= call_stmt_3311_call_req_0;
      call_stmt_3311_call_ack_0 <= ackL_unguarded(0);
      reqR_unguarded(0) <= call_stmt_3311_call_req_1;
      call_stmt_3311_call_ack_1 <= ackR_unguarded(0);
      guard_vector(0)  <=  not none_found_3285(0);
      reqL <= reqL_unregulated;
      ackL_unregulated <= ackL;
      accessSysMem_call_group_2_gI: SplitGuardInterface generic map(name => "accessSysMem_call_group_2_gI", nreqs => 1, buffering => guardBuffering, use_guards => guardFlags,  sample_only => false,  update_only => false) -- 
        port map(clk => clk, reset => reset,
        sr_in => reqL_unguarded,
        sr_out => reqL_unregulated,
        sa_in => ackL_unregulated,
        sa_out => ackL_unguarded,
        cr_in => reqR_unguarded,
        cr_out => reqR,
        ca_in => ackR,
        ca_out => ackR_unguarded,
        guards => guard_vector); -- 
      data_in <= type_cast_3304_wire_constant & NOT_u8_u8_3307_wire_constant & pa_3301 & wdata_3293;
      rval_3311 <= data_out(63 downto 0);
      CallReq: InputMuxWithBuffering -- 
        generic map (name => "InputMuxWithBuffering",
        iwidth => 109,
        owidth => 109,
        buffering => inBUFs,
        full_rate =>  true,
        twidth => 1,
        nreqs => 1,
        registered_output => false,
        no_arbitration => false)
        port map ( -- 
          reqL => reqL , 
          ackL => ackL , 
          dataL => data_in, 
          reqR => accessSysMem_call_reqs(0),
          ackR => accessSysMem_call_acks(0),
          dataR => accessSysMem_call_data(108 downto 0),
          tagR => accessSysMem_call_tag(0 downto 0),
          clk => clk, reset => reset -- 
        ); -- 
      CallComplete: OutputDemuxBaseWithBuffering -- 
        generic map ( -- 
          iwidth => 64,
          owidth => 64,
          detailed_buffering_per_output => outBUFs, 
          full_rate => true, 
          twidth => 1,
          name => "OutputDemuxBaseWithBuffering",
          nreqs => 1) -- 
        port map ( -- 
          reqR => reqR , 
          ackR => ackR , 
          dataR => data_out, 
          reqL => accessSysMem_return_acks(0), -- cross-over
          ackL => accessSysMem_return_reqs(0), -- cross-over
          dataL => accessSysMem_return_data(63 downto 0),
          tagL => accessSysMem_return_tag(0 downto 0),
          clk => clk,
          reset => reset -- 
        ); -- 
      -- 
    end Block; -- call group 2
    -- 
  end Block; -- data_path
  -- 
end writeMemoryFromL2_arch;
library std;
use std.standard.all;
library ieee;
use ieee.std_logic_1164.all;
library aHiR_ieee_proposed;
use aHiR_ieee_proposed.math_utility_pkg.all;
use aHiR_ieee_proposed.fixed_pkg.all;
use aHiR_ieee_proposed.float_pkg.all;
library ahir;
use ahir.memory_subsystem_package.all;
use ahir.types.all;
use ahir.subprograms.all;
use ahir.components.all;
use ahir.basecomponents.all;
use ahir.operatorpackage.all;
use ahir.floatoperatorpackage.all;
use ahir.utilities.all;
use ahir.functionLibraryComponents.all;
library AjitCustom;
use AjitCustom.AjitCustomComponents.all;
library l2_cache_lib;
use l2_cache_lib.l2_cache_global_package.all;
entity l2_cache is  -- system 
  port (-- 
    clk : in std_logic;
    reset : in std_logic;
    L2CACHE_TO_MEM_REQUEST_pipe_read_data: out std_logic_vector(109 downto 0);
    L2CACHE_TO_MEM_REQUEST_pipe_read_req : in std_logic_vector(0 downto 0);
    L2CACHE_TO_MEM_REQUEST_pipe_read_ack : out std_logic_vector(0 downto 0);
    L2_RESPONSE_pipe_read_data: out std_logic_vector(64 downto 0);
    L2_RESPONSE_pipe_read_req : in std_logic_vector(0 downto 0);
    L2_RESPONSE_pipe_read_ack : out std_logic_vector(0 downto 0);
    L2_TO_L1_INVALIDATE_pipe_read_data: out std_logic_vector(29 downto 0);
    L2_TO_L1_INVALIDATE_pipe_read_req : in std_logic_vector(0 downto 0);
    L2_TO_L1_INVALIDATE_pipe_read_ack : out std_logic_vector(0 downto 0);
    MEM_TO_L2CACHE_RESPONSE_pipe_write_data: in std_logic_vector(64 downto 0);
    MEM_TO_L2CACHE_RESPONSE_pipe_write_req : in std_logic_vector(0 downto 0);
    MEM_TO_L2CACHE_RESPONSE_pipe_write_ack : out std_logic_vector(0 downto 0);
    NOBLOCK_L2_INVALIDATE_pipe_write_data: in std_logic_vector(30 downto 0);
    NOBLOCK_L2_INVALIDATE_pipe_write_req : in std_logic_vector(0 downto 0);
    NOBLOCK_L2_INVALIDATE_pipe_write_ack : out std_logic_vector(0 downto 0);
    NOBLOCK_L2_REQUEST_pipe_write_data: in std_logic_vector(110 downto 0);
    NOBLOCK_L2_REQUEST_pipe_write_req : in std_logic_vector(0 downto 0);
    NOBLOCK_L2_REQUEST_pipe_write_ack : out std_logic_vector(0 downto 0)); -- 
  -- 
end entity; 
architecture l2_cache_arch  of l2_cache is -- system-architecture 
  -- interface signals to connect to memory space memory_space_1
  -- declarations related to module accessL2DataMemX4096X512
  -- declarations related to module accessL2TagMemX4096X8
  -- declarations related to module accessL2TagsDaemon
  component accessL2TagsDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      NOBLOCK_L2_TAGS_REQUEST_pipe_read_req : out  std_logic_vector(0 downto 0);
      NOBLOCK_L2_TAGS_REQUEST_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NOBLOCK_L2_TAGS_REQUEST_pipe_read_data : in   std_logic_vector(44 downto 0);
      L2_TAGS_RESPONSE_pipe_write_req : out  std_logic_vector(0 downto 0);
      L2_TAGS_RESPONSE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      L2_TAGS_RESPONSE_pipe_write_data : out  std_logic_vector(33 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module accessL2TagsDaemon
  signal accessL2TagsDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal accessL2TagsDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal accessL2TagsDaemon_start_req : std_logic;
  signal accessL2TagsDaemon_start_ack : std_logic;
  signal accessL2TagsDaemon_fin_req   : std_logic;
  signal accessL2TagsDaemon_fin_ack : std_logic;
  -- declarations related to module accessSysMem
  component accessSysMem is -- 
    generic (tag_length : integer); 
    port ( -- 
      rwbar : in  std_logic_vector(0 downto 0);
      byte_mask : in  std_logic_vector(7 downto 0);
      addr : in  std_logic_vector(35 downto 0);
      wdata : in  std_logic_vector(63 downto 0);
      rdata : out  std_logic_vector(63 downto 0);
      MEM_TO_L2CACHE_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      MEM_TO_L2CACHE_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      MEM_TO_L2CACHE_RESPONSE_pipe_read_data : in   std_logic_vector(64 downto 0);
      L2CACHE_TO_MEM_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      L2CACHE_TO_MEM_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      L2CACHE_TO_MEM_REQUEST_pipe_write_data : out  std_logic_vector(109 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module accessSysMem
  signal accessSysMem_rwbar :  std_logic_vector(0 downto 0);
  signal accessSysMem_byte_mask :  std_logic_vector(7 downto 0);
  signal accessSysMem_addr :  std_logic_vector(35 downto 0);
  signal accessSysMem_wdata :  std_logic_vector(63 downto 0);
  signal accessSysMem_rdata :  std_logic_vector(63 downto 0);
  signal accessSysMem_in_args    : std_logic_vector(108 downto 0);
  signal accessSysMem_out_args   : std_logic_vector(63 downto 0);
  signal accessSysMem_tag_in    : std_logic_vector(2 downto 0) := (others => '0');
  signal accessSysMem_tag_out   : std_logic_vector(2 downto 0);
  signal accessSysMem_start_req : std_logic;
  signal accessSysMem_start_ack : std_logic;
  signal accessSysMem_fin_req   : std_logic;
  signal accessSysMem_fin_ack : std_logic;
  -- caller side aggregated signals for module accessSysMem
  signal accessSysMem_call_reqs: std_logic_vector(1 downto 0);
  signal accessSysMem_call_acks: std_logic_vector(1 downto 0);
  signal accessSysMem_return_reqs: std_logic_vector(1 downto 0);
  signal accessSysMem_return_acks: std_logic_vector(1 downto 0);
  signal accessSysMem_call_data: std_logic_vector(217 downto 0);
  signal accessSysMem_call_tag: std_logic_vector(1 downto 0);
  signal accessSysMem_return_data: std_logic_vector(127 downto 0);
  signal accessSysMem_return_tag: std_logic_vector(1 downto 0);
  -- declarations related to module calculateHits
  -- declarations related to module dwordId
  -- declarations related to module extractDword
  -- declarations related to module getNextDirtyOffset
  -- declarations related to module insBytes
  -- declarations related to module insertIntoSetDirtyDwordMasks
  -- declarations related to module l2CacheDaemon
  component l2CacheDaemon is -- 
    generic (tag_length : integer); 
    port ( -- 
      NOBLOCK_L2_REQUEST_pipe_read_req : out  std_logic_vector(0 downto 0);
      NOBLOCK_L2_REQUEST_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NOBLOCK_L2_REQUEST_pipe_read_data : in   std_logic_vector(110 downto 0);
      L2_TAGS_RESPONSE_pipe_read_req : out  std_logic_vector(0 downto 0);
      L2_TAGS_RESPONSE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      L2_TAGS_RESPONSE_pipe_read_data : in   std_logic_vector(33 downto 0);
      NOBLOCK_L2_INVALIDATE_pipe_read_req : out  std_logic_vector(0 downto 0);
      NOBLOCK_L2_INVALIDATE_pipe_read_ack : in   std_logic_vector(0 downto 0);
      NOBLOCK_L2_INVALIDATE_pipe_read_data : in   std_logic_vector(30 downto 0);
      NOBLOCK_L2_TAGS_REQUEST_pipe_write_req : out  std_logic_vector(0 downto 0);
      NOBLOCK_L2_TAGS_REQUEST_pipe_write_ack : in   std_logic_vector(0 downto 0);
      NOBLOCK_L2_TAGS_REQUEST_pipe_write_data : out  std_logic_vector(44 downto 0);
      L2_RESPONSE_pipe_write_req : out  std_logic_vector(0 downto 0);
      L2_RESPONSE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      L2_RESPONSE_pipe_write_data : out  std_logic_vector(64 downto 0);
      L2_TO_L1_INVALIDATE_pipe_write_req : out  std_logic_vector(0 downto 0);
      L2_TO_L1_INVALIDATE_pipe_write_ack : in   std_logic_vector(0 downto 0);
      L2_TO_L1_INVALIDATE_pipe_write_data : out  std_logic_vector(29 downto 0);
      sys_mem_lock_pipe_write_req : out  std_logic_vector(0 downto 0);
      sys_mem_lock_pipe_write_ack : in   std_logic_vector(0 downto 0);
      sys_mem_lock_pipe_write_data : out  std_logic_vector(0 downto 0);
      readMemoryFromL2_call_reqs : out  std_logic_vector(0 downto 0);
      readMemoryFromL2_call_acks : in   std_logic_vector(0 downto 0);
      readMemoryFromL2_call_data : out  std_logic_vector(29 downto 0);
      readMemoryFromL2_call_tag  :  out  std_logic_vector(0 downto 0);
      readMemoryFromL2_return_reqs : out  std_logic_vector(0 downto 0);
      readMemoryFromL2_return_acks : in   std_logic_vector(0 downto 0);
      readMemoryFromL2_return_data : in   std_logic_vector(511 downto 0);
      readMemoryFromL2_return_tag :  in   std_logic_vector(0 downto 0);
      writeMemoryFromL2_call_reqs : out  std_logic_vector(0 downto 0);
      writeMemoryFromL2_call_acks : in   std_logic_vector(0 downto 0);
      writeMemoryFromL2_call_data : out  std_logic_vector(551 downto 0);
      writeMemoryFromL2_call_tag  :  out  std_logic_vector(0 downto 0);
      writeMemoryFromL2_return_reqs : out  std_logic_vector(0 downto 0);
      writeMemoryFromL2_return_acks : in   std_logic_vector(0 downto 0);
      writeMemoryFromL2_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module l2CacheDaemon
  signal l2CacheDaemon_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal l2CacheDaemon_tag_out   : std_logic_vector(1 downto 0);
  signal l2CacheDaemon_start_req : std_logic;
  signal l2CacheDaemon_start_ack : std_logic;
  signal l2CacheDaemon_fin_req   : std_logic;
  signal l2CacheDaemon_fin_ack : std_logic;
  -- declarations related to module lineAddress
  -- declarations related to module nextFreeIndex
  -- declarations related to module paTag
  -- declarations related to module readMemoryFromL2
  component readMemoryFromL2 is -- 
    generic (tag_length : integer); 
    port ( -- 
      line_address : in  std_logic_vector(29 downto 0);
      rline : out  std_logic_vector(511 downto 0);
      sys_mem_lock_pipe_read_req : out  std_logic_vector(0 downto 0);
      sys_mem_lock_pipe_read_ack : in   std_logic_vector(0 downto 0);
      sys_mem_lock_pipe_read_data : in   std_logic_vector(0 downto 0);
      accessSysMem_call_reqs : out  std_logic_vector(0 downto 0);
      accessSysMem_call_acks : in   std_logic_vector(0 downto 0);
      accessSysMem_call_data : out  std_logic_vector(108 downto 0);
      accessSysMem_call_tag  :  out  std_logic_vector(0 downto 0);
      accessSysMem_return_reqs : out  std_logic_vector(0 downto 0);
      accessSysMem_return_acks : in   std_logic_vector(0 downto 0);
      accessSysMem_return_data : in   std_logic_vector(63 downto 0);
      accessSysMem_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module readMemoryFromL2
  signal readMemoryFromL2_line_address :  std_logic_vector(29 downto 0);
  signal readMemoryFromL2_rline :  std_logic_vector(511 downto 0);
  signal readMemoryFromL2_in_args    : std_logic_vector(29 downto 0);
  signal readMemoryFromL2_out_args   : std_logic_vector(511 downto 0);
  signal readMemoryFromL2_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal readMemoryFromL2_tag_out   : std_logic_vector(1 downto 0);
  signal readMemoryFromL2_start_req : std_logic;
  signal readMemoryFromL2_start_ack : std_logic;
  signal readMemoryFromL2_fin_req   : std_logic;
  signal readMemoryFromL2_fin_ack : std_logic;
  -- caller side aggregated signals for module readMemoryFromL2
  signal readMemoryFromL2_call_reqs: std_logic_vector(0 downto 0);
  signal readMemoryFromL2_call_acks: std_logic_vector(0 downto 0);
  signal readMemoryFromL2_return_reqs: std_logic_vector(0 downto 0);
  signal readMemoryFromL2_return_acks: std_logic_vector(0 downto 0);
  signal readMemoryFromL2_call_data: std_logic_vector(29 downto 0);
  signal readMemoryFromL2_call_tag: std_logic_vector(0 downto 0);
  signal readMemoryFromL2_return_data: std_logic_vector(511 downto 0);
  signal readMemoryFromL2_return_tag: std_logic_vector(0 downto 0);
  -- declarations related to module setId
  -- declarations related to module updateDirtyWordMask
  -- declarations related to module updateSetTags
  -- declarations related to module updateSetValids
  -- declarations related to module writeMemoryFromL2
  component writeMemoryFromL2 is -- 
    generic (tag_length : integer); 
    port ( -- 
      release_lock : in  std_logic_vector(0 downto 0);
      do_write : in  std_logic_vector(0 downto 0);
      dirty_word_mask : in  std_logic_vector(7 downto 0);
      line_address : in  std_logic_vector(29 downto 0);
      wline : in  std_logic_vector(511 downto 0);
      sys_mem_lock_pipe_write_req : out  std_logic_vector(0 downto 0);
      sys_mem_lock_pipe_write_ack : in   std_logic_vector(0 downto 0);
      sys_mem_lock_pipe_write_data : out  std_logic_vector(0 downto 0);
      accessSysMem_call_reqs : out  std_logic_vector(0 downto 0);
      accessSysMem_call_acks : in   std_logic_vector(0 downto 0);
      accessSysMem_call_data : out  std_logic_vector(108 downto 0);
      accessSysMem_call_tag  :  out  std_logic_vector(0 downto 0);
      accessSysMem_return_reqs : out  std_logic_vector(0 downto 0);
      accessSysMem_return_acks : in   std_logic_vector(0 downto 0);
      accessSysMem_return_data : in   std_logic_vector(63 downto 0);
      accessSysMem_return_tag :  in   std_logic_vector(0 downto 0);
      tag_in: in std_logic_vector(tag_length-1 downto 0);
      tag_out: out std_logic_vector(tag_length-1 downto 0) ;
      clk : in std_logic;
      reset : in std_logic;
      start_req : in std_logic;
      start_ack : out std_logic;
      fin_req : in std_logic;
      fin_ack   : out std_logic-- 
    );
    -- 
  end component;
  -- argument signals for module writeMemoryFromL2
  signal writeMemoryFromL2_release_lock :  std_logic_vector(0 downto 0);
  signal writeMemoryFromL2_do_write :  std_logic_vector(0 downto 0);
  signal writeMemoryFromL2_dirty_word_mask :  std_logic_vector(7 downto 0);
  signal writeMemoryFromL2_line_address :  std_logic_vector(29 downto 0);
  signal writeMemoryFromL2_wline :  std_logic_vector(511 downto 0);
  signal writeMemoryFromL2_in_args    : std_logic_vector(551 downto 0);
  signal writeMemoryFromL2_tag_in    : std_logic_vector(1 downto 0) := (others => '0');
  signal writeMemoryFromL2_tag_out   : std_logic_vector(1 downto 0);
  signal writeMemoryFromL2_start_req : std_logic;
  signal writeMemoryFromL2_start_ack : std_logic;
  signal writeMemoryFromL2_fin_req   : std_logic;
  signal writeMemoryFromL2_fin_ack : std_logic;
  -- caller side aggregated signals for module writeMemoryFromL2
  signal writeMemoryFromL2_call_reqs: std_logic_vector(0 downto 0);
  signal writeMemoryFromL2_call_acks: std_logic_vector(0 downto 0);
  signal writeMemoryFromL2_return_reqs: std_logic_vector(0 downto 0);
  signal writeMemoryFromL2_return_acks: std_logic_vector(0 downto 0);
  signal writeMemoryFromL2_call_data: std_logic_vector(551 downto 0);
  signal writeMemoryFromL2_call_tag: std_logic_vector(0 downto 0);
  signal writeMemoryFromL2_return_tag: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe L2CACHE_TO_MEM_REQUEST
  signal L2CACHE_TO_MEM_REQUEST_pipe_write_data: std_logic_vector(109 downto 0);
  signal L2CACHE_TO_MEM_REQUEST_pipe_write_req: std_logic_vector(0 downto 0);
  signal L2CACHE_TO_MEM_REQUEST_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe L2_RESPONSE
  signal L2_RESPONSE_pipe_write_data: std_logic_vector(64 downto 0);
  signal L2_RESPONSE_pipe_write_req: std_logic_vector(0 downto 0);
  signal L2_RESPONSE_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe L2_TAGS_RESPONSE
  signal L2_TAGS_RESPONSE_pipe_write_data: std_logic_vector(33 downto 0);
  signal L2_TAGS_RESPONSE_pipe_write_req: std_logic_vector(0 downto 0);
  signal L2_TAGS_RESPONSE_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe L2_TAGS_RESPONSE
  signal L2_TAGS_RESPONSE_pipe_read_data: std_logic_vector(33 downto 0);
  signal L2_TAGS_RESPONSE_pipe_read_req: std_logic_vector(0 downto 0);
  signal L2_TAGS_RESPONSE_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe L2_TO_L1_INVALIDATE
  signal L2_TO_L1_INVALIDATE_pipe_write_data: std_logic_vector(29 downto 0);
  signal L2_TO_L1_INVALIDATE_pipe_write_req: std_logic_vector(0 downto 0);
  signal L2_TO_L1_INVALIDATE_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe MEM_TO_L2CACHE_RESPONSE
  signal MEM_TO_L2CACHE_RESPONSE_pipe_read_data: std_logic_vector(64 downto 0);
  signal MEM_TO_L2CACHE_RESPONSE_pipe_read_req: std_logic_vector(0 downto 0);
  signal MEM_TO_L2CACHE_RESPONSE_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe NOBLOCK_L2_INVALIDATE
  signal NOBLOCK_L2_INVALIDATE_pipe_read_data: std_logic_vector(30 downto 0);
  signal NOBLOCK_L2_INVALIDATE_pipe_read_req: std_logic_vector(0 downto 0);
  signal NOBLOCK_L2_INVALIDATE_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe NOBLOCK_L2_REQUEST
  signal NOBLOCK_L2_REQUEST_pipe_read_data: std_logic_vector(110 downto 0);
  signal NOBLOCK_L2_REQUEST_pipe_read_req: std_logic_vector(0 downto 0);
  signal NOBLOCK_L2_REQUEST_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe NOBLOCK_L2_TAGS_REQUEST
  signal NOBLOCK_L2_TAGS_REQUEST_pipe_write_data: std_logic_vector(44 downto 0);
  signal NOBLOCK_L2_TAGS_REQUEST_pipe_write_req: std_logic_vector(0 downto 0);
  signal NOBLOCK_L2_TAGS_REQUEST_pipe_write_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for read from pipe NOBLOCK_L2_TAGS_REQUEST
  signal NOBLOCK_L2_TAGS_REQUEST_pipe_read_data: std_logic_vector(44 downto 0);
  signal NOBLOCK_L2_TAGS_REQUEST_pipe_read_req: std_logic_vector(0 downto 0);
  signal NOBLOCK_L2_TAGS_REQUEST_pipe_read_ack: std_logic_vector(0 downto 0);
  -- aggregate signals for write to pipe sys_mem_lock
  signal sys_mem_lock_pipe_write_data: std_logic_vector(1 downto 0);
  signal sys_mem_lock_pipe_write_req: std_logic_vector(1 downto 0);
  signal sys_mem_lock_pipe_write_ack: std_logic_vector(1 downto 0);
  -- aggregate signals for read from pipe sys_mem_lock
  signal sys_mem_lock_pipe_read_data: std_logic_vector(0 downto 0);
  signal sys_mem_lock_pipe_read_req: std_logic_vector(0 downto 0);
  signal sys_mem_lock_pipe_read_ack: std_logic_vector(0 downto 0);
  -- gated clock signal declarations.
  -- 
begin -- 
  -- module accessL2TagsDaemon
  accessL2TagsDaemon_instance:accessL2TagsDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => accessL2TagsDaemon_start_req,
      start_ack => accessL2TagsDaemon_start_ack,
      fin_req => accessL2TagsDaemon_fin_req,
      fin_ack => accessL2TagsDaemon_fin_ack,
      clk => clk,
      reset => reset,
      NOBLOCK_L2_TAGS_REQUEST_pipe_read_req => NOBLOCK_L2_TAGS_REQUEST_pipe_read_req(0 downto 0),
      NOBLOCK_L2_TAGS_REQUEST_pipe_read_ack => NOBLOCK_L2_TAGS_REQUEST_pipe_read_ack(0 downto 0),
      NOBLOCK_L2_TAGS_REQUEST_pipe_read_data => NOBLOCK_L2_TAGS_REQUEST_pipe_read_data(44 downto 0),
      L2_TAGS_RESPONSE_pipe_write_req => L2_TAGS_RESPONSE_pipe_write_req(0 downto 0),
      L2_TAGS_RESPONSE_pipe_write_ack => L2_TAGS_RESPONSE_pipe_write_ack(0 downto 0),
      L2_TAGS_RESPONSE_pipe_write_data => L2_TAGS_RESPONSE_pipe_write_data(33 downto 0),
      tag_in => accessL2TagsDaemon_tag_in,
      tag_out => accessL2TagsDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  accessL2TagsDaemon_tag_in <= (others => '0');
  accessL2TagsDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => accessL2TagsDaemon_start_req, start_ack => accessL2TagsDaemon_start_ack,  fin_req => accessL2TagsDaemon_fin_req,  fin_ack => accessL2TagsDaemon_fin_ack);
  -- module accessSysMem
  accessSysMem_rwbar <= accessSysMem_in_args(108 downto 108);
  accessSysMem_byte_mask <= accessSysMem_in_args(107 downto 100);
  accessSysMem_addr <= accessSysMem_in_args(99 downto 64);
  accessSysMem_wdata <= accessSysMem_in_args(63 downto 0);
  accessSysMem_out_args <= accessSysMem_rdata ;
  -- call arbiter for module accessSysMem
  accessSysMem_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 2,
      call_data_width => 109,
      return_data_width => 64,
      callee_tag_length => 2,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => accessSysMem_call_reqs,
      call_acks => accessSysMem_call_acks,
      return_reqs => accessSysMem_return_reqs,
      return_acks => accessSysMem_return_acks,
      call_data  => accessSysMem_call_data,
      call_tag  => accessSysMem_call_tag,
      return_tag  => accessSysMem_return_tag,
      call_mtag => accessSysMem_tag_in,
      return_mtag => accessSysMem_tag_out,
      return_data =>accessSysMem_return_data,
      call_mreq => accessSysMem_start_req,
      call_mack => accessSysMem_start_ack,
      return_mreq => accessSysMem_fin_req,
      return_mack => accessSysMem_fin_ack,
      call_mdata => accessSysMem_in_args,
      return_mdata => accessSysMem_out_args,
      clk => clk, 
      reset => reset --
    ); --
  accessSysMem_instance:accessSysMem-- 
    generic map(tag_length => 3)
    port map(-- 
      rwbar => accessSysMem_rwbar,
      byte_mask => accessSysMem_byte_mask,
      addr => accessSysMem_addr,
      wdata => accessSysMem_wdata,
      rdata => accessSysMem_rdata,
      start_req => accessSysMem_start_req,
      start_ack => accessSysMem_start_ack,
      fin_req => accessSysMem_fin_req,
      fin_ack => accessSysMem_fin_ack,
      clk => clk,
      reset => reset,
      MEM_TO_L2CACHE_RESPONSE_pipe_read_req => MEM_TO_L2CACHE_RESPONSE_pipe_read_req(0 downto 0),
      MEM_TO_L2CACHE_RESPONSE_pipe_read_ack => MEM_TO_L2CACHE_RESPONSE_pipe_read_ack(0 downto 0),
      MEM_TO_L2CACHE_RESPONSE_pipe_read_data => MEM_TO_L2CACHE_RESPONSE_pipe_read_data(64 downto 0),
      L2CACHE_TO_MEM_REQUEST_pipe_write_req => L2CACHE_TO_MEM_REQUEST_pipe_write_req(0 downto 0),
      L2CACHE_TO_MEM_REQUEST_pipe_write_ack => L2CACHE_TO_MEM_REQUEST_pipe_write_ack(0 downto 0),
      L2CACHE_TO_MEM_REQUEST_pipe_write_data => L2CACHE_TO_MEM_REQUEST_pipe_write_data(109 downto 0),
      tag_in => accessSysMem_tag_in,
      tag_out => accessSysMem_tag_out-- 
    ); -- 
  -- module l2CacheDaemon
  l2CacheDaemon_instance:l2CacheDaemon-- 
    generic map(tag_length => 2)
    port map(-- 
      start_req => l2CacheDaemon_start_req,
      start_ack => l2CacheDaemon_start_ack,
      fin_req => l2CacheDaemon_fin_req,
      fin_ack => l2CacheDaemon_fin_ack,
      clk => clk,
      reset => reset,
      NOBLOCK_L2_REQUEST_pipe_read_req => NOBLOCK_L2_REQUEST_pipe_read_req(0 downto 0),
      NOBLOCK_L2_REQUEST_pipe_read_ack => NOBLOCK_L2_REQUEST_pipe_read_ack(0 downto 0),
      NOBLOCK_L2_REQUEST_pipe_read_data => NOBLOCK_L2_REQUEST_pipe_read_data(110 downto 0),
      L2_TAGS_RESPONSE_pipe_read_req => L2_TAGS_RESPONSE_pipe_read_req(0 downto 0),
      L2_TAGS_RESPONSE_pipe_read_ack => L2_TAGS_RESPONSE_pipe_read_ack(0 downto 0),
      L2_TAGS_RESPONSE_pipe_read_data => L2_TAGS_RESPONSE_pipe_read_data(33 downto 0),
      NOBLOCK_L2_INVALIDATE_pipe_read_req => NOBLOCK_L2_INVALIDATE_pipe_read_req(0 downto 0),
      NOBLOCK_L2_INVALIDATE_pipe_read_ack => NOBLOCK_L2_INVALIDATE_pipe_read_ack(0 downto 0),
      NOBLOCK_L2_INVALIDATE_pipe_read_data => NOBLOCK_L2_INVALIDATE_pipe_read_data(30 downto 0),
      NOBLOCK_L2_TAGS_REQUEST_pipe_write_req => NOBLOCK_L2_TAGS_REQUEST_pipe_write_req(0 downto 0),
      NOBLOCK_L2_TAGS_REQUEST_pipe_write_ack => NOBLOCK_L2_TAGS_REQUEST_pipe_write_ack(0 downto 0),
      NOBLOCK_L2_TAGS_REQUEST_pipe_write_data => NOBLOCK_L2_TAGS_REQUEST_pipe_write_data(44 downto 0),
      L2_RESPONSE_pipe_write_req => L2_RESPONSE_pipe_write_req(0 downto 0),
      L2_RESPONSE_pipe_write_ack => L2_RESPONSE_pipe_write_ack(0 downto 0),
      L2_RESPONSE_pipe_write_data => L2_RESPONSE_pipe_write_data(64 downto 0),
      L2_TO_L1_INVALIDATE_pipe_write_req => L2_TO_L1_INVALIDATE_pipe_write_req(0 downto 0),
      L2_TO_L1_INVALIDATE_pipe_write_ack => L2_TO_L1_INVALIDATE_pipe_write_ack(0 downto 0),
      L2_TO_L1_INVALIDATE_pipe_write_data => L2_TO_L1_INVALIDATE_pipe_write_data(29 downto 0),
      sys_mem_lock_pipe_write_req => sys_mem_lock_pipe_write_req(1 downto 1),
      sys_mem_lock_pipe_write_ack => sys_mem_lock_pipe_write_ack(1 downto 1),
      sys_mem_lock_pipe_write_data => sys_mem_lock_pipe_write_data(1 downto 1),
      readMemoryFromL2_call_reqs => readMemoryFromL2_call_reqs(0 downto 0),
      readMemoryFromL2_call_acks => readMemoryFromL2_call_acks(0 downto 0),
      readMemoryFromL2_call_data => readMemoryFromL2_call_data(29 downto 0),
      readMemoryFromL2_call_tag => readMemoryFromL2_call_tag(0 downto 0),
      readMemoryFromL2_return_reqs => readMemoryFromL2_return_reqs(0 downto 0),
      readMemoryFromL2_return_acks => readMemoryFromL2_return_acks(0 downto 0),
      readMemoryFromL2_return_data => readMemoryFromL2_return_data(511 downto 0),
      readMemoryFromL2_return_tag => readMemoryFromL2_return_tag(0 downto 0),
      writeMemoryFromL2_call_reqs => writeMemoryFromL2_call_reqs(0 downto 0),
      writeMemoryFromL2_call_acks => writeMemoryFromL2_call_acks(0 downto 0),
      writeMemoryFromL2_call_data => writeMemoryFromL2_call_data(551 downto 0),
      writeMemoryFromL2_call_tag => writeMemoryFromL2_call_tag(0 downto 0),
      writeMemoryFromL2_return_reqs => writeMemoryFromL2_return_reqs(0 downto 0),
      writeMemoryFromL2_return_acks => writeMemoryFromL2_return_acks(0 downto 0),
      writeMemoryFromL2_return_tag => writeMemoryFromL2_return_tag(0 downto 0),
      tag_in => l2CacheDaemon_tag_in,
      tag_out => l2CacheDaemon_tag_out-- 
    ); -- 
  -- module will be run forever 
  l2CacheDaemon_tag_in <= (others => '0');
  l2CacheDaemon_auto_run: auto_run generic map(use_delay => true)  port map(clk => clk, reset => reset, start_req => l2CacheDaemon_start_req, start_ack => l2CacheDaemon_start_ack,  fin_req => l2CacheDaemon_fin_req,  fin_ack => l2CacheDaemon_fin_ack);
  -- module readMemoryFromL2
  readMemoryFromL2_line_address <= readMemoryFromL2_in_args(29 downto 0);
  readMemoryFromL2_out_args <= readMemoryFromL2_rline ;
  -- call arbiter for module readMemoryFromL2
  readMemoryFromL2_arbiter: SplitCallArbiter -- 
    generic map( --
      name => "SplitCallArbiter", num_reqs => 1,
      call_data_width => 30,
      return_data_width => 512,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => readMemoryFromL2_call_reqs,
      call_acks => readMemoryFromL2_call_acks,
      return_reqs => readMemoryFromL2_return_reqs,
      return_acks => readMemoryFromL2_return_acks,
      call_data  => readMemoryFromL2_call_data,
      call_tag  => readMemoryFromL2_call_tag,
      return_tag  => readMemoryFromL2_return_tag,
      call_mtag => readMemoryFromL2_tag_in,
      return_mtag => readMemoryFromL2_tag_out,
      return_data =>readMemoryFromL2_return_data,
      call_mreq => readMemoryFromL2_start_req,
      call_mack => readMemoryFromL2_start_ack,
      return_mreq => readMemoryFromL2_fin_req,
      return_mack => readMemoryFromL2_fin_ack,
      call_mdata => readMemoryFromL2_in_args,
      return_mdata => readMemoryFromL2_out_args,
      clk => clk, 
      reset => reset --
    ); --
  readMemoryFromL2_instance:readMemoryFromL2-- 
    generic map(tag_length => 2)
    port map(-- 
      line_address => readMemoryFromL2_line_address,
      rline => readMemoryFromL2_rline,
      start_req => readMemoryFromL2_start_req,
      start_ack => readMemoryFromL2_start_ack,
      fin_req => readMemoryFromL2_fin_req,
      fin_ack => readMemoryFromL2_fin_ack,
      clk => clk,
      reset => reset,
      sys_mem_lock_pipe_read_req => sys_mem_lock_pipe_read_req(0 downto 0),
      sys_mem_lock_pipe_read_ack => sys_mem_lock_pipe_read_ack(0 downto 0),
      sys_mem_lock_pipe_read_data => sys_mem_lock_pipe_read_data(0 downto 0),
      accessSysMem_call_reqs => accessSysMem_call_reqs(1 downto 1),
      accessSysMem_call_acks => accessSysMem_call_acks(1 downto 1),
      accessSysMem_call_data => accessSysMem_call_data(217 downto 109),
      accessSysMem_call_tag => accessSysMem_call_tag(1 downto 1),
      accessSysMem_return_reqs => accessSysMem_return_reqs(1 downto 1),
      accessSysMem_return_acks => accessSysMem_return_acks(1 downto 1),
      accessSysMem_return_data => accessSysMem_return_data(127 downto 64),
      accessSysMem_return_tag => accessSysMem_return_tag(1 downto 1),
      tag_in => readMemoryFromL2_tag_in,
      tag_out => readMemoryFromL2_tag_out-- 
    ); -- 
  -- module writeMemoryFromL2
  writeMemoryFromL2_release_lock <= writeMemoryFromL2_in_args(551 downto 551);
  writeMemoryFromL2_do_write <= writeMemoryFromL2_in_args(550 downto 550);
  writeMemoryFromL2_dirty_word_mask <= writeMemoryFromL2_in_args(549 downto 542);
  writeMemoryFromL2_line_address <= writeMemoryFromL2_in_args(541 downto 512);
  writeMemoryFromL2_wline <= writeMemoryFromL2_in_args(511 downto 0);
  -- call arbiter for module writeMemoryFromL2
  writeMemoryFromL2_arbiter: SplitCallArbiterNoOutargs -- 
    generic map( --
      name => "SplitCallArbiterNoOutargs", num_reqs => 1,
      call_data_width => 552,
      callee_tag_length => 1,
      caller_tag_length => 1--
    )
    port map(-- 
      call_reqs => writeMemoryFromL2_call_reqs,
      call_acks => writeMemoryFromL2_call_acks,
      return_reqs => writeMemoryFromL2_return_reqs,
      return_acks => writeMemoryFromL2_return_acks,
      call_data  => writeMemoryFromL2_call_data,
      call_tag  => writeMemoryFromL2_call_tag,
      return_tag  => writeMemoryFromL2_return_tag,
      call_mtag => writeMemoryFromL2_tag_in,
      return_mtag => writeMemoryFromL2_tag_out,
      call_mreq => writeMemoryFromL2_start_req,
      call_mack => writeMemoryFromL2_start_ack,
      return_mreq => writeMemoryFromL2_fin_req,
      return_mack => writeMemoryFromL2_fin_ack,
      call_mdata => writeMemoryFromL2_in_args,
      clk => clk, 
      reset => reset --
    ); --
  writeMemoryFromL2_instance:writeMemoryFromL2-- 
    generic map(tag_length => 2)
    port map(-- 
      release_lock => writeMemoryFromL2_release_lock,
      do_write => writeMemoryFromL2_do_write,
      dirty_word_mask => writeMemoryFromL2_dirty_word_mask,
      line_address => writeMemoryFromL2_line_address,
      wline => writeMemoryFromL2_wline,
      start_req => writeMemoryFromL2_start_req,
      start_ack => writeMemoryFromL2_start_ack,
      fin_req => writeMemoryFromL2_fin_req,
      fin_ack => writeMemoryFromL2_fin_ack,
      clk => clk,
      reset => reset,
      sys_mem_lock_pipe_write_req => sys_mem_lock_pipe_write_req(0 downto 0),
      sys_mem_lock_pipe_write_ack => sys_mem_lock_pipe_write_ack(0 downto 0),
      sys_mem_lock_pipe_write_data => sys_mem_lock_pipe_write_data(0 downto 0),
      accessSysMem_call_reqs => accessSysMem_call_reqs(0 downto 0),
      accessSysMem_call_acks => accessSysMem_call_acks(0 downto 0),
      accessSysMem_call_data => accessSysMem_call_data(108 downto 0),
      accessSysMem_call_tag => accessSysMem_call_tag(0 downto 0),
      accessSysMem_return_reqs => accessSysMem_return_reqs(0 downto 0),
      accessSysMem_return_acks => accessSysMem_return_acks(0 downto 0),
      accessSysMem_return_data => accessSysMem_return_data(63 downto 0),
      accessSysMem_return_tag => accessSysMem_return_tag(0 downto 0),
      tag_in => writeMemoryFromL2_tag_in,
      tag_out => writeMemoryFromL2_tag_out-- 
    ); -- 
  L2CACHE_TO_MEM_REQUEST_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe L2CACHE_TO_MEM_REQUEST",
      num_reads => 1,
      num_writes => 1,
      data_width => 110,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => L2CACHE_TO_MEM_REQUEST_pipe_read_req,
      read_ack => L2CACHE_TO_MEM_REQUEST_pipe_read_ack,
      read_data => L2CACHE_TO_MEM_REQUEST_pipe_read_data,
      write_req => L2CACHE_TO_MEM_REQUEST_pipe_write_req,
      write_ack => L2CACHE_TO_MEM_REQUEST_pipe_write_ack,
      write_data => L2CACHE_TO_MEM_REQUEST_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  L2_RESPONSE_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe L2_RESPONSE",
      num_reads => 1,
      num_writes => 1,
      data_width => 65,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => L2_RESPONSE_pipe_read_req,
      read_ack => L2_RESPONSE_pipe_read_ack,
      read_data => L2_RESPONSE_pipe_read_data,
      write_req => L2_RESPONSE_pipe_write_req,
      write_ack => L2_RESPONSE_pipe_write_ack,
      write_data => L2_RESPONSE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  L2_TAGS_RESPONSE_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe L2_TAGS_RESPONSE",
      num_reads => 1,
      num_writes => 1,
      data_width => 34,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => true,
      depth => 0 --
    )
    port map( -- 
      read_req => L2_TAGS_RESPONSE_pipe_read_req,
      read_ack => L2_TAGS_RESPONSE_pipe_read_ack,
      read_data => L2_TAGS_RESPONSE_pipe_read_data,
      write_req => L2_TAGS_RESPONSE_pipe_write_req,
      write_ack => L2_TAGS_RESPONSE_pipe_write_ack,
      write_data => L2_TAGS_RESPONSE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  L2_TO_L1_INVALIDATE_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe L2_TO_L1_INVALIDATE",
      num_reads => 1,
      num_writes => 1,
      data_width => 30,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => L2_TO_L1_INVALIDATE_pipe_read_req,
      read_ack => L2_TO_L1_INVALIDATE_pipe_read_ack,
      read_data => L2_TO_L1_INVALIDATE_pipe_read_data,
      write_req => L2_TO_L1_INVALIDATE_pipe_write_req,
      write_ack => L2_TO_L1_INVALIDATE_pipe_write_ack,
      write_data => L2_TO_L1_INVALIDATE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  MEM_TO_L2CACHE_RESPONSE_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe MEM_TO_L2CACHE_RESPONSE",
      num_reads => 1,
      num_writes => 1,
      data_width => 65,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => MEM_TO_L2CACHE_RESPONSE_pipe_read_req,
      read_ack => MEM_TO_L2CACHE_RESPONSE_pipe_read_ack,
      read_data => MEM_TO_L2CACHE_RESPONSE_pipe_read_data,
      write_req => MEM_TO_L2CACHE_RESPONSE_pipe_write_req,
      write_ack => MEM_TO_L2CACHE_RESPONSE_pipe_write_ack,
      write_data => MEM_TO_L2CACHE_RESPONSE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  NOBLOCK_L2_INVALIDATE_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe NOBLOCK_L2_INVALIDATE",
      num_reads => 1,
      num_writes => 1,
      data_width => 31,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => NOBLOCK_L2_INVALIDATE_pipe_read_req,
      read_ack => NOBLOCK_L2_INVALIDATE_pipe_read_ack,
      read_data => NOBLOCK_L2_INVALIDATE_pipe_read_data,
      write_req => NOBLOCK_L2_INVALIDATE_pipe_write_req,
      write_ack => NOBLOCK_L2_INVALIDATE_pipe_write_ack,
      write_data => NOBLOCK_L2_INVALIDATE_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  NOBLOCK_L2_REQUEST_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe NOBLOCK_L2_REQUEST",
      num_reads => 1,
      num_writes => 1,
      data_width => 111,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 0 --
    )
    port map( -- 
      read_req => NOBLOCK_L2_REQUEST_pipe_read_req,
      read_ack => NOBLOCK_L2_REQUEST_pipe_read_ack,
      read_data => NOBLOCK_L2_REQUEST_pipe_read_data,
      write_req => NOBLOCK_L2_REQUEST_pipe_write_req,
      write_ack => NOBLOCK_L2_REQUEST_pipe_write_ack,
      write_data => NOBLOCK_L2_REQUEST_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- non-blocking pipe... Input-ports must have non-blocking-flag => true
  NOBLOCK_L2_TAGS_REQUEST_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe NOBLOCK_L2_TAGS_REQUEST",
      num_reads => 1,
      num_writes => 1,
      data_width => 45,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => true,
      depth => 0 --
    )
    port map( -- 
      read_req => NOBLOCK_L2_TAGS_REQUEST_pipe_read_req,
      read_ack => NOBLOCK_L2_TAGS_REQUEST_pipe_read_ack,
      read_data => NOBLOCK_L2_TAGS_REQUEST_pipe_read_data,
      write_req => NOBLOCK_L2_TAGS_REQUEST_pipe_write_req,
      write_ack => NOBLOCK_L2_TAGS_REQUEST_pipe_write_ack,
      write_data => NOBLOCK_L2_TAGS_REQUEST_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  sys_mem_lock_Pipe: PipeBase -- 
    generic map( -- 
      name => "pipe sys_mem_lock",
      num_reads => 1,
      num_writes => 2,
      data_width => 1,
      lifo_mode => false,
      full_rate => false,
      shift_register_mode => false,
      bypass => false,
      depth => 1 --
    )
    port map( -- 
      read_req => sys_mem_lock_pipe_read_req,
      read_ack => sys_mem_lock_pipe_read_ack,
      read_data => sys_mem_lock_pipe_read_data,
      write_req => sys_mem_lock_pipe_write_req,
      write_ack => sys_mem_lock_pipe_write_ack,
      write_data => sys_mem_lock_pipe_write_data,
      clk => clk,reset => reset -- 
    ); -- 
  -- gated clock generators 
  -- 
end l2_cache_arch;
